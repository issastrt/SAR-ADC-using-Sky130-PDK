magic
tech sky130A
magscale 1 2
timestamp 1757042133
<< nwell >>
rect 0 -882 8762 928
<< pwell >>
rect 0 978 8762 1782
rect 0 -1736 8762 -932
<< metal1 >>
rect -97 1831 -33 1837
rect -97 1779 -91 1831
rect -39 1828 -33 1831
rect -39 1782 8762 1828
rect -39 1779 -33 1782
rect -97 1773 -33 1779
rect 349 985 395 1204
rect 340 979 404 985
rect 340 927 346 979
rect 398 927 404 979
rect 340 921 404 927
rect 1698 979 1762 985
rect 1698 927 1704 979
rect 1756 927 1762 979
rect 1698 921 1762 927
rect 2535 979 2599 985
rect 2535 927 2541 979
rect 2593 927 2599 979
rect 2535 921 2599 927
rect 3670 979 3734 985
rect 3670 927 3676 979
rect 3728 927 3734 979
rect 3670 921 3734 927
rect 6609 979 6673 985
rect 6609 927 6615 979
rect 6667 927 6673 979
rect 6609 921 6673 927
rect 7744 979 7808 985
rect 7744 927 7750 979
rect 7802 927 7808 979
rect 7744 921 7808 927
rect 349 672 395 921
rect 3056 859 3120 865
rect 3056 807 3062 859
rect 3114 807 3120 859
rect 3056 801 3120 807
rect 7130 859 7194 865
rect 7130 807 7136 859
rect 7188 807 7194 859
rect 7130 801 7194 807
rect 4507 721 4571 727
rect 4507 669 4513 721
rect 4565 669 4571 721
rect 4507 663 4571 669
rect 5772 721 5836 727
rect 5772 669 5778 721
rect 5830 669 5836 721
rect 5772 663 5836 669
rect 4385 401 4449 407
rect 441 395 505 401
rect 441 343 447 395
rect 499 343 505 395
rect 4385 349 4391 401
rect 4443 349 4449 401
rect 4385 343 4449 349
rect 8459 401 8523 407
rect 8459 349 8465 401
rect 8517 349 8523 401
rect 8459 343 8523 349
rect 441 337 505 343
rect 1120 305 1184 311
rect 1120 253 1126 305
rect 1178 253 1184 305
rect 1120 247 1184 253
rect 2312 305 2376 311
rect 2312 253 2318 305
rect 2370 253 2376 305
rect 2312 247 2376 253
rect 4248 305 4312 311
rect 4248 253 4254 305
rect 4306 253 4312 305
rect 4248 247 4312 253
rect 6386 305 6450 311
rect 6386 253 6392 305
rect 6444 253 6450 305
rect 6386 247 6450 253
rect 8322 305 8386 311
rect 8322 253 8328 305
rect 8380 253 8386 305
rect 8322 247 8386 253
rect 0 0 8762 46
rect 1120 -207 1184 -201
rect 1120 -259 1126 -207
rect 1178 -259 1184 -207
rect 1120 -265 1184 -259
rect 2312 -207 2376 -201
rect 2312 -259 2318 -207
rect 2370 -259 2376 -207
rect 2312 -265 2376 -259
rect 4248 -207 4312 -201
rect 4248 -259 4254 -207
rect 4306 -259 4312 -207
rect 4248 -265 4312 -259
rect 6386 -207 6450 -201
rect 6386 -259 6392 -207
rect 6444 -259 6450 -207
rect 6386 -265 6450 -259
rect 8322 -207 8386 -201
rect 8322 -259 8328 -207
rect 8380 -259 8386 -207
rect 8322 -265 8386 -259
rect 4385 -304 4449 -298
rect 4385 -356 4391 -304
rect 4443 -356 4449 -304
rect 4385 -362 4449 -356
rect 8459 -304 8523 -298
rect 8459 -356 8465 -304
rect 8517 -356 8523 -304
rect 8459 -362 8523 -356
rect 4507 -623 4571 -617
rect 4507 -675 4513 -623
rect 4565 -675 4571 -623
rect 4507 -681 4571 -675
rect 5772 -623 5836 -617
rect 5772 -675 5778 -623
rect 5830 -675 5836 -623
rect 5772 -681 5836 -675
rect 3056 -761 3120 -755
rect 3056 -813 3062 -761
rect 3114 -813 3120 -761
rect 3056 -819 3120 -813
rect 7130 -761 7194 -755
rect 7130 -813 7136 -761
rect 7188 -813 7194 -761
rect 7130 -819 7194 -813
rect 1698 -881 1762 -875
rect 1698 -933 1704 -881
rect 1756 -933 1762 -881
rect 1698 -939 1762 -933
rect 2535 -881 2599 -875
rect 2535 -933 2541 -881
rect 2593 -933 2599 -881
rect 2535 -939 2599 -933
rect 3670 -881 3734 -875
rect 3670 -933 3676 -881
rect 3728 -933 3734 -881
rect 3670 -939 3734 -933
rect 5251 -881 5315 -875
rect 5251 -933 5257 -881
rect 5309 -933 5315 -881
rect 5251 -939 5315 -933
rect 6386 -881 6450 -875
rect 6386 -933 6392 -881
rect 6444 -933 6450 -881
rect 6386 -939 6450 -933
rect 6609 -881 6673 -875
rect 6609 -933 6615 -881
rect 6667 -933 6673 -881
rect 6609 -939 6673 -933
rect 7744 -881 7808 -875
rect 7744 -933 7750 -881
rect 7802 -933 7808 -881
rect 7744 -939 7808 -933
rect 2312 -1109 2376 -1103
rect 2312 -1161 2318 -1109
rect 2370 -1161 2376 -1109
rect 2312 -1167 2376 -1161
rect 5028 -1109 5092 -1103
rect 5028 -1161 5034 -1109
rect 5086 -1161 5092 -1109
rect 5028 -1167 5092 -1161
rect -97 -1733 -33 -1727
rect -97 -1785 -91 -1733
rect -39 -1736 -33 -1733
rect -39 -1782 8762 -1736
rect -39 -1785 -33 -1782
rect -97 -1791 -33 -1785
<< via1 >>
rect -91 1779 -39 1831
rect 346 927 398 979
rect 1704 927 1756 979
rect 2541 927 2593 979
rect 3676 927 3728 979
rect 6615 927 6667 979
rect 7750 927 7802 979
rect 3062 807 3114 859
rect 7136 807 7188 859
rect 4513 669 4565 721
rect 5778 669 5830 721
rect 447 343 499 395
rect 4391 349 4443 401
rect 8465 349 8517 401
rect 1126 253 1178 305
rect 2318 253 2370 305
rect 4254 253 4306 305
rect 6392 253 6444 305
rect 8328 253 8380 305
rect 1126 -259 1178 -207
rect 2318 -259 2370 -207
rect 4254 -259 4306 -207
rect 6392 -259 6444 -207
rect 8328 -259 8380 -207
rect 4391 -356 4443 -304
rect 8465 -356 8517 -304
rect 4513 -675 4565 -623
rect 5778 -675 5830 -623
rect 3062 -813 3114 -761
rect 7136 -813 7188 -761
rect 1704 -933 1756 -881
rect 2541 -933 2593 -881
rect 3676 -933 3728 -881
rect 5257 -933 5309 -881
rect 6392 -933 6444 -881
rect 6615 -933 6667 -881
rect 7750 -933 7802 -881
rect 2318 -1161 2370 -1109
rect 5034 -1161 5086 -1109
rect -91 -1785 -39 -1733
<< metal2 >>
rect -102 1833 -28 1842
rect -102 1777 -93 1833
rect -37 1777 -28 1833
rect -102 1768 -28 1777
rect 340 979 404 985
rect 340 927 346 979
rect 398 976 404 979
rect 1698 979 1762 985
rect 1698 976 1704 979
rect 398 930 1704 976
rect 398 927 404 930
rect 340 921 404 927
rect 1698 927 1704 930
rect 1756 927 1762 979
rect 1698 921 1762 927
rect 2535 979 2599 985
rect 2535 927 2541 979
rect 2593 976 2599 979
rect 3670 979 3734 985
rect 3670 976 3676 979
rect 2593 930 3676 976
rect 2593 927 2599 930
rect 2535 921 2599 927
rect 3670 927 3676 930
rect 3728 927 3734 979
rect 3670 921 3734 927
rect 6609 979 6673 985
rect 6609 927 6615 979
rect 6667 976 6673 979
rect 7744 979 7808 985
rect 7744 976 7750 979
rect 6667 930 7750 976
rect 6667 927 6673 930
rect 6609 921 6673 927
rect 7744 927 7750 930
rect 7802 927 7808 979
rect 7744 921 7808 927
rect 1250 861 1324 870
rect 1250 805 1259 861
rect 1315 856 1324 861
rect 3056 859 3120 865
rect 3056 856 3062 859
rect 1315 810 3062 856
rect 1315 805 1324 810
rect 1250 796 1324 805
rect 3056 807 3062 810
rect 3114 856 3120 859
rect 7130 859 7194 865
rect 7130 856 7136 859
rect 3114 810 7136 856
rect 3114 807 3120 810
rect 3056 801 3120 807
rect 7130 807 7136 810
rect 7188 807 7194 859
rect 7130 801 7194 807
rect 4507 721 4571 727
rect 4507 669 4513 721
rect 4565 718 4571 721
rect 5772 721 5836 727
rect 5772 718 5778 721
rect 4565 672 5778 718
rect 4565 669 4571 672
rect 4507 663 4571 669
rect 5772 669 5778 672
rect 5830 669 5836 721
rect 5772 663 5836 669
rect 441 395 505 401
rect 441 343 447 395
rect 499 392 505 395
rect 565 397 639 406
rect 565 392 574 397
rect 499 346 574 392
rect 499 343 505 346
rect 441 337 505 343
rect 565 341 574 346
rect 630 341 639 397
rect 565 332 639 341
rect 4380 403 4454 412
rect 4380 347 4389 403
rect 4445 347 4454 403
rect 4380 338 4454 347
rect 8454 403 8528 412
rect 8454 347 8463 403
rect 8519 347 8528 403
rect 8454 338 8528 347
rect 1120 305 1184 311
rect 1120 253 1126 305
rect 1178 302 1184 305
rect 1399 307 1473 316
rect 1399 302 1408 307
rect 1178 256 1408 302
rect 1178 253 1184 256
rect 1120 247 1184 253
rect 1399 251 1408 256
rect 1464 251 1473 307
rect 1399 242 1473 251
rect 2307 307 2381 316
rect 2307 251 2316 307
rect 2372 251 2381 307
rect 2307 242 2381 251
rect 4243 307 4317 316
rect 4243 251 4252 307
rect 4308 251 4317 307
rect 4243 242 4317 251
rect 6381 307 6455 316
rect 6381 251 6390 307
rect 6446 251 6455 307
rect 6381 242 6455 251
rect 8317 307 8391 316
rect 8317 251 8326 307
rect 8382 251 8391 307
rect 8317 242 8391 251
rect 1120 -207 1184 -201
rect 1120 -210 1126 -207
rect 1118 -256 1126 -210
rect 1120 -259 1126 -256
rect 1178 -210 1184 -207
rect 1250 -205 1324 -196
rect 1250 -210 1259 -205
rect 1178 -256 1259 -210
rect 1178 -259 1184 -256
rect 1120 -265 1184 -259
rect 1250 -261 1259 -256
rect 1315 -261 1324 -205
rect 1250 -270 1324 -261
rect 2307 -205 2381 -196
rect 2307 -261 2316 -205
rect 2372 -261 2381 -205
rect 2307 -270 2381 -261
rect 4248 -207 4312 -201
rect 4248 -259 4254 -207
rect 4306 -210 4312 -207
rect 4380 -205 4454 -196
rect 4380 -210 4389 -205
rect 4306 -256 4389 -210
rect 4306 -259 4312 -256
rect 4248 -265 4312 -259
rect 4380 -261 4389 -256
rect 4445 -261 4454 -205
rect 4380 -270 4454 -261
rect 6381 -205 6455 -196
rect 6381 -261 6390 -205
rect 6446 -261 6455 -205
rect 6381 -270 6455 -261
rect 8322 -207 8386 -201
rect 8322 -259 8328 -207
rect 8380 -210 8386 -207
rect 8454 -205 8528 -196
rect 8454 -210 8463 -205
rect 8380 -256 8463 -210
rect 8380 -259 8386 -256
rect 8322 -265 8386 -259
rect 8454 -261 8463 -256
rect 8519 -261 8528 -205
rect 8454 -270 8528 -261
rect 4243 -302 4317 -293
rect 4243 -358 4252 -302
rect 4308 -307 4317 -302
rect 4385 -304 4449 -298
rect 4385 -307 4391 -304
rect 4308 -353 4391 -307
rect 4308 -358 4317 -353
rect 4243 -367 4317 -358
rect 4385 -356 4391 -353
rect 4443 -356 4449 -304
rect 4385 -362 4449 -356
rect 8317 -302 8391 -293
rect 8317 -358 8326 -302
rect 8382 -307 8391 -302
rect 8459 -304 8523 -298
rect 8459 -307 8465 -304
rect 8382 -353 8465 -307
rect 8382 -358 8391 -353
rect 8317 -367 8391 -358
rect 8459 -356 8465 -353
rect 8517 -356 8523 -304
rect 8459 -362 8523 -356
rect 4507 -623 4571 -617
rect 4507 -675 4513 -623
rect 4565 -626 4571 -623
rect 5772 -623 5836 -617
rect 5772 -626 5778 -623
rect 4565 -672 5778 -626
rect 4565 -675 4571 -672
rect 4507 -681 4571 -675
rect 5772 -675 5778 -672
rect 5830 -675 5836 -623
rect 5772 -681 5836 -675
rect 1399 -759 1473 -750
rect 1399 -815 1408 -759
rect 1464 -764 1473 -759
rect 3056 -761 3120 -755
rect 3056 -764 3062 -761
rect 1464 -810 3062 -764
rect 1464 -815 1473 -810
rect 1399 -824 1473 -815
rect 3056 -813 3062 -810
rect 3114 -764 3120 -761
rect 7130 -761 7194 -755
rect 7130 -764 7136 -761
rect 3114 -810 7136 -764
rect 3114 -813 3120 -810
rect 3056 -819 3120 -813
rect 7130 -813 7136 -810
rect 7188 -813 7194 -761
rect 7130 -819 7194 -813
rect 565 -879 639 -870
rect 565 -935 574 -879
rect 630 -884 639 -879
rect 1698 -881 1762 -875
rect 1698 -884 1704 -881
rect 630 -930 1704 -884
rect 630 -935 639 -930
rect 565 -944 639 -935
rect 1698 -933 1704 -930
rect 1756 -933 1762 -881
rect 1698 -939 1762 -933
rect 2535 -881 2599 -875
rect 2535 -933 2541 -881
rect 2593 -884 2599 -881
rect 3670 -881 3734 -875
rect 3670 -884 3676 -881
rect 2593 -930 3676 -884
rect 2593 -933 2599 -930
rect 2535 -939 2599 -933
rect 3670 -933 3676 -930
rect 3728 -933 3734 -881
rect 3670 -939 3734 -933
rect 5251 -881 5315 -875
rect 5251 -933 5257 -881
rect 5309 -884 5315 -881
rect 6386 -881 6450 -875
rect 6386 -884 6392 -881
rect 5309 -930 6392 -884
rect 5309 -933 5315 -930
rect 5251 -939 5315 -933
rect 6386 -933 6392 -930
rect 6444 -933 6450 -881
rect 6386 -939 6450 -933
rect 6609 -881 6673 -875
rect 6609 -933 6615 -881
rect 6667 -884 6673 -881
rect 7744 -881 7808 -875
rect 7744 -884 7750 -881
rect 6667 -930 7750 -884
rect 6667 -933 6673 -930
rect 6609 -939 6673 -933
rect 7744 -933 7750 -930
rect 7802 -933 7808 -881
rect 7744 -939 7808 -933
rect 2312 -1109 2376 -1103
rect 2312 -1161 2318 -1109
rect 2370 -1112 2376 -1109
rect 5028 -1109 5092 -1103
rect 5028 -1112 5034 -1109
rect 2370 -1158 5034 -1112
rect 2370 -1161 2376 -1158
rect 2312 -1167 2376 -1161
rect 5028 -1161 5034 -1158
rect 5086 -1161 5092 -1109
rect 5028 -1167 5092 -1161
rect -102 -1731 -28 -1722
rect -102 -1787 -93 -1731
rect -37 -1787 -28 -1731
rect -102 -1796 -28 -1787
<< via2 >>
rect -93 1831 -37 1833
rect -93 1779 -91 1831
rect -91 1779 -39 1831
rect -39 1779 -37 1831
rect -93 1777 -37 1779
rect 1259 805 1315 861
rect 574 341 630 397
rect 4389 401 4445 403
rect 4389 349 4391 401
rect 4391 349 4443 401
rect 4443 349 4445 401
rect 4389 347 4445 349
rect 8463 401 8519 403
rect 8463 349 8465 401
rect 8465 349 8517 401
rect 8517 349 8519 401
rect 8463 347 8519 349
rect 1408 251 1464 307
rect 2316 305 2372 307
rect 2316 253 2318 305
rect 2318 253 2370 305
rect 2370 253 2372 305
rect 2316 251 2372 253
rect 4252 305 4308 307
rect 4252 253 4254 305
rect 4254 253 4306 305
rect 4306 253 4308 305
rect 4252 251 4308 253
rect 6390 305 6446 307
rect 6390 253 6392 305
rect 6392 253 6444 305
rect 6444 253 6446 305
rect 6390 251 6446 253
rect 8326 305 8382 307
rect 8326 253 8328 305
rect 8328 253 8380 305
rect 8380 253 8382 305
rect 8326 251 8382 253
rect 1259 -261 1315 -205
rect 2316 -207 2372 -205
rect 2316 -259 2318 -207
rect 2318 -259 2370 -207
rect 2370 -259 2372 -207
rect 2316 -261 2372 -259
rect 4389 -261 4445 -205
rect 6390 -207 6446 -205
rect 6390 -259 6392 -207
rect 6392 -259 6444 -207
rect 6444 -259 6446 -207
rect 6390 -261 6446 -259
rect 8463 -261 8519 -205
rect 4252 -358 4308 -302
rect 8326 -358 8382 -302
rect 1408 -815 1464 -759
rect 574 -935 630 -879
rect -93 -1733 -37 -1731
rect -93 -1785 -91 -1733
rect -91 -1785 -39 -1733
rect -39 -1785 -37 -1733
rect -93 -1787 -37 -1785
<< metal3 >>
rect -98 1833 -32 1838
rect -98 1777 -93 1833
rect -37 1777 -32 1833
rect -98 1772 -32 1777
rect -95 -1726 -35 1772
rect 1254 861 1320 866
rect 1254 805 1259 861
rect 1315 805 1320 861
rect 1254 800 1320 805
rect 569 397 635 402
rect 569 341 574 397
rect 630 341 635 397
rect 569 336 635 341
rect 572 -874 632 336
rect 1257 -200 1317 800
rect 4384 403 4450 408
rect 4384 347 4389 403
rect 4445 347 4450 403
rect 4384 342 4450 347
rect 8458 403 8524 408
rect 8458 347 8463 403
rect 8519 347 8524 403
rect 8458 342 8524 347
rect 1403 307 1469 312
rect 1403 251 1408 307
rect 1464 251 1469 307
rect 1403 246 1469 251
rect 2311 307 2377 312
rect 2311 251 2316 307
rect 2372 251 2377 307
rect 2311 246 2377 251
rect 4247 307 4313 312
rect 4247 251 4252 307
rect 4308 251 4313 307
rect 4247 246 4313 251
rect 1254 -205 1320 -200
rect 1254 -261 1259 -205
rect 1315 -261 1320 -205
rect 1254 -266 1320 -261
rect 1406 -754 1466 246
rect 2314 -200 2374 246
rect 2311 -205 2377 -200
rect 2311 -261 2316 -205
rect 2372 -261 2377 -205
rect 2311 -266 2377 -261
rect 4250 -297 4310 246
rect 4387 -200 4447 342
rect 6385 307 6451 312
rect 6385 251 6390 307
rect 6446 251 6451 307
rect 6385 246 6451 251
rect 8321 307 8387 312
rect 8321 251 8326 307
rect 8382 251 8387 307
rect 8321 246 8387 251
rect 6388 -200 6448 246
rect 4384 -205 4450 -200
rect 4384 -261 4389 -205
rect 4445 -261 4450 -205
rect 4384 -266 4450 -261
rect 6385 -205 6451 -200
rect 6385 -261 6390 -205
rect 6446 -261 6451 -205
rect 6385 -266 6451 -261
rect 8324 -297 8384 246
rect 8461 -200 8521 342
rect 8458 -205 8524 -200
rect 8458 -261 8463 -205
rect 8519 -261 8524 -205
rect 8458 -266 8524 -261
rect 4247 -302 4313 -297
rect 4247 -358 4252 -302
rect 4308 -358 4313 -302
rect 4247 -363 4313 -358
rect 8321 -302 8387 -297
rect 8321 -358 8326 -302
rect 8382 -358 8387 -302
rect 8321 -363 8387 -358
rect 1403 -759 1469 -754
rect 1403 -815 1408 -759
rect 1464 -815 1469 -759
rect 1403 -820 1469 -815
rect 569 -879 635 -874
rect 569 -935 574 -879
rect 630 -935 635 -879
rect 569 -940 635 -935
rect -98 -1731 -32 -1726
rect -98 -1787 -93 -1731
rect -37 -1787 -32 -1731
rect -98 -1792 -32 -1787
use 3-input-nand  3-input-nand_0
timestamp 1756481424
transform 1 0 -1279 0 -1 400
box 2023 -1428 3995 400
use 3-input-nand  3-input-nand_1
timestamp 1756481424
transform 1 0 -1279 0 1 -354
box 2023 -1428 3995 400
use 3-input-nand  3-input-nand_2
timestamp 1756481424
transform 1 0 693 0 -1 400
box 2023 -1428 3995 400
use 3-input-nand  3-input-nand_3
timestamp 1756481424
transform 1 0 693 0 1 -354
box 2023 -1428 3995 400
use 3-input-nand  3-input-nand_4
timestamp 1756481424
transform 1 0 4767 0 -1 400
box 2023 -1428 3995 400
use 3-input-nand  3-input-nand_5
timestamp 1756481424
transform 1 0 4767 0 1 -354
box 2023 -1428 3995 400
use Inverter  Inverter_0
timestamp 1756481424
transform 1 0 -1366 0 -1 942
box 1366 -886 2110 942
use Inverter  Inverter_1
timestamp 1756481424
transform 1 0 3322 0 1 -896
box 1366 -886 2110 942
use Nand_Gate  Nand_Gate_0
timestamp 1756481424
transform 1 0 3526 0 -1 1298
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_1
timestamp 1756481424
transform 1 0 3526 0 1 -1252
box 1906 -530 3264 1298
<< labels >>
flabel metal1 349 672 395 1204 0 FreeSans 160 0 0 0 D
port 1 nsew
flabel metal3 2314 -205 2374 251 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 1257 -205 1317 805 0 FreeSans 160 90 0 0 nPRE
port 4 nsew
flabel metal3 1406 -759 1466 251 0 FreeSans 160 90 0 0 nCLR
port 3 nsew
flabel metal3 8461 -205 8521 347 0 FreeSans 160 0 0 0 Q
port 6 nsew
flabel metal1 0 0 8762 46 0 FreeSans 160 0 0 0 VDD
port 7 nsew
flabel metal1 -42 1782 8762 1828 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal3 8324 -302 8384 251 0 FreeSans 160 0 0 0 Qbar
port 5 nsew
<< end >>
