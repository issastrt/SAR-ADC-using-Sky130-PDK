* NGSPICE file created from SAR-ADC-using-Sky130-PDK.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_CY7YBN a_n130_n144# a_72_n144# w_n330_n441# a_n72_n241#
X0 a_72_n144# a_n72_n241# a_n130_n144# w_n330_n441# sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P a_n202_n144# a_n144_n232# a_144_n144#
+ VSUBS
X0 a_144_n144# a_n144_n232# a_n202_n144# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
.ends

.subckt Inverter GND VDD Vout Vin
XXM1 VDD Vout VDD Vin sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM2 GND Vin Vout GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
.ends

.subckt Nand_Gate GND A B Vout VDD
XXM1 VDD Vout VDD B sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM2 Vout VDD VDD A sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM3 m1_2428_n226# B Vout GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
XXM4 GND A m1_2428_n226# GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
.ends

.subckt And_Gate VDD B Vout A GND
XInverter_0 GND VDD Vout Inverter_0/Vin Inverter
XNand_Gate_0 GND A B Inverter_0/Vin VDD Nand_Gate
.ends

.subckt x3-input-nand GND A B Vout C VDD
XXM1 VDD Vout VDD C sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM2 Vout VDD VDD B sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM3 VDD Vout VDD A sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM4 m1_3159_n1124# C Vout GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
XXM5 m1_2545_n1124# B m1_3159_n1124# GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
XXM6 GND A m1_2545_n1124# GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
.ends

.subckt D_FlipFlop CLK nCLR nPRE Qbar Q D VDD GND
XInverter_1 GND VDD Nand_Gate_1/B CLK Inverter
XInverter_0 GND VDD Inverter_0/Vout D Inverter
X3-input-nand_0 GND nCLR D 3-input-nand_2/B CLK VDD x3-input-nand
X3-input-nand_1 GND nPRE Inverter_0/Vout 3-input-nand_3/B CLK VDD x3-input-nand
X3-input-nand_3 GND nCLR 3-input-nand_3/B Nand_Gate_1/A Nand_Gate_0/A VDD x3-input-nand
X3-input-nand_2 GND nPRE 3-input-nand_2/B Nand_Gate_0/A Nand_Gate_1/A VDD x3-input-nand
X3-input-nand_4 GND nPRE Nand_Gate_0/Vout Q Qbar VDD x3-input-nand
X3-input-nand_5 GND nCLR Nand_Gate_1/Vout Qbar Q VDD x3-input-nand
XNand_Gate_0 GND Nand_Gate_0/A Nand_Gate_1/B Nand_Gate_0/Vout VDD Nand_Gate
XNand_Gate_1 GND Nand_Gate_1/A Nand_Gate_1/B Nand_Gate_1/Vout VDD Nand_Gate
.ends

.subckt switch GND VDD Z A B Vref
XXM1 B Z VDD m1_1636_n741# sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM2 Z Vref B GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
XXM3 Z A VDD Vref sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM4 A m1_1636_n741# Z GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
XXM5 VDD m1_1636_n741# VDD Vref sky130_fd_pr__pfet_g5v0d10v5_CY7YBN
XXM6 GND Vref m1_1636_n741# GND sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_XAJUMH m4_n2619_n280# c2_n2539_n200#
X0 c2_n2539_n200# m4_n2619_n280# sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
.ends

.subckt CDAC8 GND VDD OUT b1 b4 b7 b6 b0 b5 b3 b2
Xswitch_0 GND VDD switch_0/Z GND VDD b2 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_28 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_39 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_17 switch_2/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_193 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_182 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_171 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_160 switch_0/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_1 GND VDD switch_1/Z GND VDD b0 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_29 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_18 switch_0/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_194 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_183 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_150 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_161 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_172 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_2 GND VDD switch_2/Z GND VDD b1 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_19 switch_0/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_195 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_184 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_140 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_162 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_173 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_196 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_185 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_130 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_141 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_152 switch_0/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_163 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_174 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_120 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_197 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_186 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_131 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_142 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_164 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_153 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_175 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_5 GND VDD switch_5/Z GND VDD b3 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_121 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_198 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_187 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_110 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_132 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_143 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_165 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_154 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_176 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_6 GND VDD switch_6/Z GND VDD b6 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_122 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_199 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_188 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_177 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_133 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_100 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_144 switch_2/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_166 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_155 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_111 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_7 GND VDD switch_7/Z GND VDD b7 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_123 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_189 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_178 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_134 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_145 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_101 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_112 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_167 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_156 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_8 GND VDD switch_8/Z GND VDD b4 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_124 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_113 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_179 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_135 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_102 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_146 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_168 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_157 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xswitch_9 GND VDD switch_9/Z GND VDD b5 switch
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_0 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_125 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_114 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_169 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_103 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_147 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_158 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_1 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_126 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_115 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_104 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_137 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_148 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_159 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_2 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_127 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_116 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_105 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_138 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_149 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_3 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_128 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_117 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_106 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_139 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_4 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_118 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_129 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_107 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_5 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_119 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_108 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_6 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_109 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_7 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_8 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_9 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_250 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_251 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_240 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_252 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_241 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_230 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_253 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_242 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_231 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_220 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_90 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_254 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_243 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_232 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_221 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_210 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_80 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_91 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_255 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_244 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_233 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_222 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_211 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_200 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_70 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_81 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_92 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_256 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_245 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_234 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_223 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_212 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_201 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_71 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_82 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_93 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_60 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_246 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_235 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_224 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_213 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_202 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_50 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_72 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_83 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_94 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_61 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_247 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_225 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_236 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_214 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_203 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_51 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_73 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_40 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_84 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_95 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_62 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_248 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_226 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_237 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_215 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_204 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_30 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_52 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_74 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_41 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_96 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_85 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_63 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_249 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_227 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_238 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_216 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_205 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_20 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_31 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_53 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_75 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_42 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_64 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_86 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_97 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_228 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_239 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_217 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_206 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_32 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_54 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_43 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_10 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_76 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_65 switch_1/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_98 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_87 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_21 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_229 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_218 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_207 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_44 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_11 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_55 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_77 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_22 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_99 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_66 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_33 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_88 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_219 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_208 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_45 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_12 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_78 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_23 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_56 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_67 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_34 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_89 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_209 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_46 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_13 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_79 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_24 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_57 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_68 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_35 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_47 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_14 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_69 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_25 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_58 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_36 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_190 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_15 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_48 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_26 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_59 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_37 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_191 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_180 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_49 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_27 switch_8/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_38 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_16 switch_9/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_192 switch_5/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_181 switch_6/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
Xsky130_fd_pr__cap_mim_m3_2_XAJUMH_170 switch_7/Z OUT sky130_fd_pr__cap_mim_m3_2_XAJUMH
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DTGLBV a_100_n2000# a_n100_n2088# a_n292_n2222#
+ a_n158_n2000#
X0 a_100_n2000# a_n100_n2088# a_n158_n2000# a_n292_n2222# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_AZGBXE m4_n884_n280# c2_n804_n200#
X0 c2_n804_n200# m4_n884_n280# sky130_fd_pr__cap_mim_m3_2 l=2 w=5.35
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q a_100_n5000# w_n358_n5297# a_n158_n5000#
+ a_n100_n5097#
X0 a_100_n5000# a_n100_n5097# a_n158_n5000# w_n358_n5297# sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_Q3M7H8 a_n100_n1088# a_n292_n1222# a_n158_n1000#
+ a_100_n1000#
X0 a_100_n1000# a_n100_n1088# a_n158_n1000# a_n292_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_94KJBV a_100_n1500# a_n100_n1588# a_n292_n1722#
+ a_n158_n1500#
X0 a_100_n1500# a_n100_n1588# a_n158_n1500# a_n292_n1722# sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_UX3D7Q a_n100_n6097# a_100_n6000# w_n358_n6297#
+ a_n158_n6000#
X0 a_100_n6000# a_n100_n6097# a_n158_n6000# w_n358_n6297# sky130_fd_pr__pfet_g5v0d10v5 ad=17.4 pd=120.58 as=17.4 ps=120.58 w=60 l=1
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_2WP2GG a_n703_n15546# a_n573_14984# a_n573_n15416#
X0 a_n573_14984# a_n573_n15416# a_n703_n15546# sky130_fd_pr__res_xhigh_po_5p73 l=150
.ends

.subckt Comparator VDD Vinm Vinp Vout VSS
Xsky130_fd_pr__nfet_g5v0d10v5_DTGLBV_2 VSS m1_25981_n1645# VSS m1_25981_n1645# sky130_fd_pr__nfet_g5v0d10v5_DTGLBV
Xsky130_fd_pr__cap_mim_m3_2_AZGBXE_0 VSS Vout sky130_fd_pr__cap_mim_m3_2_AZGBXE
XXM3 VDD VDD m1_27718_12003# m1_27718_12003# sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q
Xsky130_fd_pr__cap_mim_m3_2_AZGBXE_1 Vout m1_28569_18903# sky130_fd_pr__cap_mim_m3_2_AZGBXE
XXM4 m1_28569_18903# VDD VDD m1_27718_12003# sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q
XXM6 m1_25981_n1645# VSS VSS Vout sky130_fd_pr__nfet_g5v0d10v5_Q3M7H8
Xsky130_fd_pr__nfet_g5v0d10v5_94KJBV_0 m1_27975_9075# Vinm VSS m1_27718_12003# sky130_fd_pr__nfet_g5v0d10v5_94KJBV
Xsky130_fd_pr__nfet_g5v0d10v5_94KJBV_1 m1_28569_18903# Vinp VSS m1_27975_9075# sky130_fd_pr__nfet_g5v0d10v5_94KJBV
XXM9 m1_28569_18903# Vout VDD VDD sky130_fd_pr__pfet_g5v0d10v5_UX3D7Q
Xsky130_fd_pr__res_xhigh_po_5p73_2WP2GG_0 VSS VDD m1_25981_n1645# sky130_fd_pr__res_xhigh_po_5p73_2WP2GG
Xsky130_fd_pr__nfet_g5v0d10v5_DTGLBV_1 VSS m1_25981_n1645# VSS m1_27975_9075# sky130_fd_pr__nfet_g5v0d10v5_DTGLBV
.ends

.subckt RingCounter Q0 Q1 Q2 Q3 Q4 Q5 Q6 Q7 Q8 Q9 Q10 Q11 Q12 Q13 Q14 Q15 VDD CLK
+ EN GND
XD_FlipFlop_10 CLK VDD EN D_FlipFlop_10/Qbar Q8 Q7 VDD GND D_FlipFlop
XD_FlipFlop_11 CLK VDD EN D_FlipFlop_11/Qbar Q10 Q9 VDD GND D_FlipFlop
XD_FlipFlop_12 CLK VDD EN D_FlipFlop_12/Qbar Q11 Q10 VDD GND D_FlipFlop
XD_FlipFlop_13 CLK VDD EN D_FlipFlop_13/Qbar Q12 Q11 VDD GND D_FlipFlop
XD_FlipFlop_14 CLK VDD EN D_FlipFlop_14/Qbar Q13 Q12 VDD GND D_FlipFlop
XD_FlipFlop_15 CLK VDD EN D_FlipFlop_15/Qbar Q14 Q13 VDD GND D_FlipFlop
XD_FlipFlop_16 CLK VDD EN D_FlipFlop_16/Qbar D_FlipFlop_17/D Q15 VDD GND D_FlipFlop
XD_FlipFlop_17 CLK EN VDD D_FlipFlop_17/Qbar Q0 D_FlipFlop_17/D VDD GND D_FlipFlop
XD_FlipFlop_1 CLK VDD EN D_FlipFlop_1/Qbar Q1 Q0 VDD GND D_FlipFlop
XD_FlipFlop_3 CLK VDD EN D_FlipFlop_3/Qbar Q3 Q2 VDD GND D_FlipFlop
XD_FlipFlop_2 CLK VDD EN D_FlipFlop_2/Qbar Q2 Q1 VDD GND D_FlipFlop
XD_FlipFlop_4 CLK VDD EN D_FlipFlop_4/Qbar Q4 Q3 VDD GND D_FlipFlop
XD_FlipFlop_5 CLK VDD EN D_FlipFlop_5/Qbar Q5 Q4 VDD GND D_FlipFlop
XD_FlipFlop_6 CLK VDD EN D_FlipFlop_6/Qbar Q7 Q6 VDD GND D_FlipFlop
XD_FlipFlop_7 CLK VDD EN D_FlipFlop_7/Qbar Q6 Q5 VDD GND D_FlipFlop
XD_FlipFlop_8 CLK VDD EN D_FlipFlop_8/Qbar Q15 Q14 VDD GND D_FlipFlop
XD_FlipFlop_9 CLK VDD EN D_FlipFlop_9/Qbar Q9 Q8 VDD GND D_FlipFlop
.ends

.subckt SAR-ADC-using-Sky130-PDK CLK Q0 Q1 Q2 Q3 Q4 Q6 Q5 Q7 VDD EN GND Vbias Vin
XAnd_Gate_0 VDD And_Gate_0/B And_Gate_0/Vout CLK GND And_Gate
XAnd_Gate_1 VDD And_Gate_1/B And_Gate_1/Vout CLK GND And_Gate
XAnd_Gate_3 VDD And_Gate_3/B And_Gate_3/Vout CLK GND And_Gate
XAnd_Gate_2 VDD And_Gate_2/B And_Gate_2/Vout CLK GND And_Gate
XAnd_Gate_4 VDD CLK And_Gate_4/Vout And_Gate_4/A GND And_Gate
XAnd_Gate_5 VDD CLK And_Gate_5/Vout And_Gate_5/A GND And_Gate
XAnd_Gate_6 VDD CLK And_Gate_6/Vout And_Gate_6/A GND And_Gate
XAnd_Gate_7 VDD CLK And_Gate_7/Vout And_Gate_7/A GND And_Gate
XD_FlipFlop_0 And_Gate_7/Vout FFCLR Nand_Gate_5/A D_FlipFlop_0/Qbar Q4 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XD_FlipFlop_1 And_Gate_5/Vout EN FFCLR D_FlipFlop_1/Qbar Q7 D_FlipFlop_7/D VDD GND
+ D_FlipFlop
XCDAC8_0 GND VDD CDAC8_0/OUT Q1 Q4 Q7 Q6 Q0 Q5 Q3 Q2 CDAC8
XD_FlipFlop_2 And_Gate_4/Vout FFCLR Nand_Gate_0/A D_FlipFlop_2/Qbar Q6 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XD_FlipFlop_3 And_Gate_6/Vout FFCLR Nand_Gate_2/A D_FlipFlop_3/Qbar Q5 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XD_FlipFlop_4 And_Gate_3/Vout FFCLR Nand_Gate_1/B D_FlipFlop_4/Qbar Q3 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XComparator_0 VDD CDAC8_0/OUT Vin D_FlipFlop_7/D Vbias Comparator
XD_FlipFlop_5 And_Gate_2/Vout FFCLR Nand_Gate_6/B D_FlipFlop_5/Qbar Q2 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XD_FlipFlop_6 And_Gate_0/Vout FFCLR Nand_Gate_7/B D_FlipFlop_6/Qbar Q1 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XD_FlipFlop_7 And_Gate_1/Vout FFCLR Nand_Gate_4/B D_FlipFlop_7/Qbar Q0 D_FlipFlop_7/D
+ VDD GND D_FlipFlop
XNand_Gate_0 GND Nand_Gate_0/A Nand_Gate_0/B And_Gate_4/A VDD Nand_Gate
XNand_Gate_1 GND Nand_Gate_1/A Nand_Gate_1/B And_Gate_3/B VDD Nand_Gate
XNand_Gate_2 GND Nand_Gate_2/A Nand_Gate_2/B And_Gate_6/A VDD Nand_Gate
XNand_Gate_4 GND Nand_Gate_4/A Nand_Gate_4/B And_Gate_1/B VDD Nand_Gate
XNand_Gate_3 GND FFCLR Nand_Gate_3/B And_Gate_5/A VDD Nand_Gate
XNand_Gate_5 GND Nand_Gate_5/A Nand_Gate_5/B And_Gate_7/A VDD Nand_Gate
XNand_Gate_6 GND Nand_Gate_6/A Nand_Gate_6/B And_Gate_2/B VDD Nand_Gate
XRingCounter_0 FFCLR Nand_Gate_3/B Nand_Gate_0/A Nand_Gate_0/B Nand_Gate_2/A Nand_Gate_2/B
+ Nand_Gate_5/A Nand_Gate_5/B Nand_Gate_1/B Nand_Gate_1/A Nand_Gate_6/B Nand_Gate_6/A
+ Nand_Gate_7/B Nand_Gate_7/A Nand_Gate_4/B Nand_Gate_4/A VDD CLK EN GND RingCounter
XNand_Gate_7 GND Nand_Gate_7/A Nand_Gate_7/B And_Gate_0/B VDD Nand_Gate
.ends

