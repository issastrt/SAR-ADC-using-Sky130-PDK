magic
tech sky130A
magscale 1 2
timestamp 1755260286
<< pwell >>
rect -739 -15582 739 15582
<< psubdiff >>
rect -703 15512 -607 15546
rect 607 15512 703 15546
rect -703 15450 -669 15512
rect 669 15450 703 15512
rect -703 -15512 -669 -15450
rect 669 -15512 703 -15450
rect -703 -15546 -607 -15512
rect 607 -15546 703 -15512
<< psubdiffcont >>
rect -607 15512 607 15546
rect -703 -15450 -669 15450
rect 669 -15450 703 15450
rect -607 -15546 607 -15512
<< xpolycontact >>
rect -573 14984 573 15416
rect -573 -15416 573 -14984
<< xpolyres >>
rect -573 -14984 573 14984
<< locali >>
rect -703 15512 -607 15546
rect 607 15512 703 15546
rect -703 15450 -669 15512
rect 669 15450 703 15512
rect -703 -15512 -669 -15450
rect 669 -15512 703 -15450
rect -703 -15546 -607 -15512
rect 607 -15546 703 -15512
<< viali >>
rect -557 15001 557 15398
rect -557 -15398 557 -15001
<< metal1 >>
rect -569 15398 569 15404
rect -569 15001 -557 15398
rect 557 15001 569 15398
rect -569 14995 569 15001
rect -569 -15001 569 -14995
rect -569 -15398 -557 -15001
rect 557 -15398 569 -15001
rect -569 -15404 569 -15398
<< properties >>
string FIXED_BBOX -686 -15529 686 15529
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 150.0 m 1 nx 1 wmin 5.730 lmin 0.50 class resistor rho 2000 val 52.421k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0 mult 1
<< end >>
