* NGSPICE file created from SAR-ADC-using-Sky130-PDK.ext - technology: sky130A

.subckt SAR-ADC-using-Sky130-PDK CLK Q0 Q1 Q2 Q3 Q4 Q6 Q5 Q7 VDD EN GND Vbias Vin
X0 Comparator_0.Vinm CDAC8_0.switch_7.Z.t131 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1 a_64511_52572# EN.t0 GND.t581 GND.t580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X2 a_45761_13083# CLK.t0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 GND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X3 GND.t577 EN.t1 a_29289_15797# GND.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X4 VDD.t943 Nand_Gate_4.A.t4 RingCounter_0.D_FlipFlop_8.Qbar VDD.t626 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X5 D_FlipFlop_6.3-input-nand_2.C.t0 D_FlipFlop_6.3-input-nand_1.Vout VDD.t225 VDD.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X6 a_51499_49858# EN.t2 GND.t573 GND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X7 GND.t579 EN.t3 a_46375_13083# GND.t578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 VDD.t762 VDD.t763 VDD.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X9 a_100961_13083# CLK.t1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 GND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X10 Comparator_0.Vinm CDAC8_0.switch_7.Z.t130 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X11 Comparator_0.Vinm CDAC8_0.switch_8.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X12 D_FlipFlop_7.Qbar D_FlipFlop_7.Nand_Gate_1.Vout VDD.t803 VDD.t652 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X13 a_124399_52572# RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_123785_52572# GND.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X14 a_68585_52572# EN.t4 GND.t575 GND.t574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X15 a_51369_13083# RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 a_50755_13083# GND.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X16 Comparator_0.Vinm CDAC8_0.switch_6.Z.t67 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X17 VDD.t966 D_FlipFlop_1.3-input-nand_2.Vout.t4 D_FlipFlop_1.3-input-nand_2.C.t0 VDD.t778 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X18 GND.t571 EN.t5 a_101575_13083# GND.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X19 a_65125_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_64511_52572# GND.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X20 Comparator_0.Vinm CDAC8_0.switch_6.Z.t66 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X21 Comparator_0.Vinm CDAC8_0.switch_6.Z.t65 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X22 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_7.D.t3 VDD.t807 VDD.t806 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X23 VDD.t1100 CLK.t2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 VDD.t1048 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X24 Nand_Gate_0.A.t1 RingCounter_0.D_FlipFlop_2.Qbar a_69199_52572# GND.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X25 Comparator_0.Vinm CDAC8_0.switch_6.Z.t64 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X26 VDD.t539 EN.t6 D_FlipFlop_1.3-input-nand_2.C.t2 VDD.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X27 a_52113_49858# RingCounter_0.D_FlipFlop_1.3-input-nand_1.B a_51499_49858# GND.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X28 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 a_56187_49858# GND.t714 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X29 VDD.t795 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 VDD.t794 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X30 VDD.t34 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_2.A.t0 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X31 a_48565_16975# CLK.t3 GND.t79 GND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X32 a_134283_17072# And_Gate_1.Vout.t2 D_FlipFlop_7.3-input-nand_1.Vout GND.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X33 VDD.t780 Nand_Gate_2.B.t4 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X34 VDD.t1103 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 VDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X35 a_123785_52572# EN.t7 GND.t569 GND.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X36 VDD.t766 And_Gate_4.Vout.t2 D_FlipFlop_2.3-input-nand_1.Vout VDD.t657 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X37 D_FlipFlop_0.CLK.t1 And_Gate_7.Nand_Gate_0.Vout GND.t645 GND.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X38 a_134283_27764# And_Gate_3.Vout.t2 D_FlipFlop_4.3-input-nand_1.Vout GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X39 a_71017_47663# Nand_Gate_0.A.t4 GND.t747 GND.t746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X40 a_74807_15797# RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout GND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X41 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_2.3-input-nand_2.C.t4 VDD.t909 VDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X42 Comparator_0.Vinm CDAC8_0.switch_9.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X43 Nand_Gate_5.B.t1 RingCounter_0.D_FlipFlop_6.Qbar a_124399_52572# GND.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X44 GND.t103 VDD.t1108 a_51369_13083# GND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X45 Comparator_0.Vinm CDAC8_0.switch_7.Z.t129 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X46 a_79495_15797# Nand_Gate_6.A.t4 a_78881_15797# GND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X47 Nand_Gate_6.A.t0 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t161 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X48 GND.t275 FFCLR.t4 a_132925_37007# GND.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X49 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 a_111387_49858# GND.t729 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X50 a_107927_13083# RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 GND.t882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X51 a_56187_49858# RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 GND.t812 GND.t811 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X52 Comparator_0.Vinm CDAC8_0.switch_7.Z.t128 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X53 Comparator_0.Vinm CDAC8_0.switch_9.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X54 GND.t105 VDD.t1109 a_57415_15797# GND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X55 a_134897_43285# D_FlipFlop_7.D.t4 a_134283_43285# GND.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X56 Nand_Gate_2.A.t2 RingCounter_0.D_FlipFlop_4.Qbar VDD.t313 VDD.t312 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X57 a_108671_52572# EN.t8 GND.t567 GND.t566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X58 VDD.t30 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X59 Comparator_0.Vinm CDAC8_0.switch_8.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X60 VDD.t537 EN.t9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 VDD.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X61 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 a_109285_52572# GND.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X62 Comparator_0.Vinm CDAC8_0.switch_7.Z.t127 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X63 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 VDD.t760 VDD.t761 VDD.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X64 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 EN.t10 VDD.t535 VDD.t534 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X65 D_FlipFlop_1.3-input-nand_2.Vout.t0 D_FlipFlop_1.3-input-nand_0.Vout VDD.t413 VDD.t412 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X66 VDD.t661 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 VDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X67 a_76909_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 GND.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X68 Comparator_0.Vinm CDAC8_0.switch_6.Z.t63 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X69 VDD.t533 EN.t11 Nand_Gate_6.A.t1 VDD.t532 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X70 GND.t107 VDD.t1110 a_112615_15797# GND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X71 D_FlipFlop_0.3-input-nand_2.Vout.t0 D_FlipFlop_0.3-input-nand_0.Vout VDD.t76 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X72 a_110029_13083# RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 GND.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X73 VDD.t216 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 VDD.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X74 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 CLK.t4 GND.t12 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X75 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 VDD.t136 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X76 GND.t873 D_FlipFlop_5.3-input-nand_2.C.t4 a_130209_24200# GND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X77 a_75898_39392# Q6.t4 GND.t702 GND.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X78 Comparator_0.Vinm CDAC8_0.switch_7.Z.t126 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X79 CDAC8_0.switch_2.Z.t0 a_75898_21528# VDD.t569 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X80 Comparator_0.Vinm CDAC8_0.switch_8.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X81 VDD.t993 Q3.t4 CDAC8_0.switch_5.Z.t2 GND.t876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X82 Nand_Gate_5.Vout.t1 Nand_Gate_5.B.t4 a_115177_47663# GND.t874 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X83 a_109285_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_108671_52572# GND.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X84 GND.t680 Nand_Gate_6.B.t4 a_134897_24200# GND.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X85 VDD.t244 FFCLR.t5 D_FlipFlop_5.3-input-nand_0.Vout VDD.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X86 VDD.t1099 CLK.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 VDD.t1045 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X87 GND.t14 CLK.t6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 GND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X88 VDD.t321 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_5.Qbar VDD.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X89 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B Nand_Gate_2.A.t4 GND.t722 GND.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X90 RingCounter_0.D_FlipFlop_17.Qbar EN.t12 VDD.t531 VDD.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X91 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t758 VDD.t759 VDD.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X92 VDD.t995 Q3.t5 D_FlipFlop_4.Qbar VDD.t994 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X93 VDD.t860 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 VDD.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X94 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 CLK.t7 GND.t16 GND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X95 VDD.t967 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 VDD.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X96 a_86591_49858# VDD.t1111 GND.t109 GND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X97 RingCounter_0.D_FlipFlop_17.Qbar FFCLR.t6 VDD.t246 VDD.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X98 VDD.t1098 CLK.t8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 VDD.t1042 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X99 CDAC8_0.switch_5.Z.t1 a_75898_28676# GND.t97 GND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X100 a_115177_47663# Nand_Gate_5.A.t4 GND.t847 GND.t846 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X101 a_118967_15797# RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout GND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X102 RingCounter_0.D_FlipFlop_5.Qbar VDD.t756 VDD.t757 VDD.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X103 a_138533_35417.t2 D_FlipFlop_7.D.t0 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X104 Nand_Gate_4.B.t3 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t861 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X105 Comparator_0.Vinm CDAC8_0.switch_9.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X106 a_132311_40571# D_FlipFlop_3.3-input-nand_2.Vout.t4 D_FlipFlop_3.3-input-nand_2.C.t2 GND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X107 Comparator_0.Vinm CDAC8_0.switch_7.Z.t125 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X108 GND.t698 D_FlipFlop_7.D.t5 D_FlipFlop_5.3-input-nand_1.B GND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X109 VDD.t613 D_FlipFlop_3.3-input-nand_2.C.t4 D_FlipFlop_3.3-input-nand_2.Vout.t2 VDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X110 GND.t247 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 a_85847_13083# GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X111 VDD.t248 FFCLR.t7 D_FlipFlop_2.3-input-nand_0.Vout VDD.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X112 RingCounter_0.D_FlipFlop_5.Qbar Nand_Gate_2.B.t5 VDD.t918 VDD.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X113 Comparator_0.Vinm CDAC8_0.switch_7.Z.t124 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X114 a_128237_39721# D_FlipFlop_2.Qbar Q6.t3 GND.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X115 D_FlipFlop_4.Qbar D_FlipFlop_4.Nand_Gate_1.Vout VDD.t826 VDD.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X116 VDD.t842 Nand_Gate_2.A.t5 D_FlipFlop_3.3-input-nand_2.Vout.t0 VDD.t384 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X117 VDD.t234 D_FlipFlop_0.3-input-nand_2.Vout.t4 D_FlipFlop_0.3-input-nand_2.C.t2 VDD.t233 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X118 VDD.t323 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout VDD.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X119 VDD.t407 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout VDD.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X120 a_87205_49858# RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 a_86591_49858# GND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X121 GND.t723 Nand_Gate_2.A.t6 a_128851_43285# GND.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X122 GND.t616 D_FlipFlop_6.3-input-nand_2.C.t4 a_130209_20636# GND.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X123 VDD.t250 FFCLR.t8 D_FlipFlop_0.3-input-nand_2.C.t3 VDD.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X124 VDD.t529 EN.t13 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 VDD.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X125 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 CLK.t9 a_41073_52572# GND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X126 VDD.t527 EN.t14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 VDD.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X127 Comparator_0.Vinm CDAC8_0.switch_8.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X128 a_43789_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 GND.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X129 GND.t271 Nand_Gate_7.B.t4 a_134897_20636# GND.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X130 VDD.t251 FFCLR.t9 D_FlipFlop_6.3-input-nand_0.Vout VDD.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X131 a_128237_23350# D_FlipFlop_6.Qbar Q1.t3 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X132 CDAC8_0.switch_6.Z.t0 a_75898_39392# VDD.t132 VDD.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X133 VDD.t525 EN.t15 Nand_Gate_4.B.t2 VDD.t524 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X134 Comparator_0.Vinm CDAC8_0.switch_7.Z.t123 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X135 Comparator_0.Vinm CDAC8_0.switch_6.Z.t62 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X136 a_132925_40571# D_FlipFlop_3.3-input-nand_1.Vout a_132311_40571# GND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X137 VDD.t81 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X138 Comparator_0.Vinm CDAC8_0.switch_7.Z.t122 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X139 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 VDD.t325 VDD.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X140 CDAC8_0.switch_1.Z.t0 a_75898_18814# VDD.t22 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X141 a_75898_28676# Q3.t6 VDD.t997 VDD.t996 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X142 a_134897_19786# D_FlipFlop_7.D.t6 a_134283_19786# GND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X143 VDD.t260 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 VDD.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X144 a_103765_47663# Nand_Gate_2.Vout.t3 GND.t744 GND.t743 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X145 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B Nand_Gate_3.B.t4 GND.t407 GND.t406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X146 GND.t19 CLK.t10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 GND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X147 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t754 VDD.t755 VDD.t463 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X148 VDD.t268 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X149 And_Gate_3.Vout.t0 And_Gate_3.Nand_Gate_0.Vout VDD.t302 VDD.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X150 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 CLK.t11 VDD.t1097 VDD.t1096 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X151 Comparator_0.Vinm CDAC8_0.switch_6.Z.t61 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X152 VDD.t523 EN.t16 Nand_Gate_1.B.t1 VDD.t522 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X153 VDD.t563 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 VDD.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X154 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 CLK.t12 a_96273_49858# GND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X155 GND.t283 Q7.t4 CDAC8_0.switch_7.Z.t0 VDD.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X156 VDD.t119 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X157 GND.t228 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 a_52727_13083# GND.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X158 VDD.t275 And_Gate_5.Vout.t2 D_FlipFlop_1.3-input-nand_1.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X159 Comparator_0.Vinm CDAC8_0.switch_7.Z.t121 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X160 VDD.t369 Nand_Gate_3.B.t5 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X161 Comparator_0.Vinm CDAC8_0.switch_7.Z.t120 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X162 D_FlipFlop_1.Nand_Gate_1.Vout D_FlipFlop_1.3-input-nand_2.C.t4 VDD.t777 VDD.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X163 a_57545_49858# VDD.t1112 GND.t111 GND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X164 Comparator_0.Vinm CDAC8_0.switch_7.Z.t119 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X165 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 VDD.t553 VDD.t552 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X166 Comparator_0.Vinm CDAC8_0.switch_9.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X167 a_75898_42964# Q5.t4 VDD.t855 VDD.t854 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X168 a_130209_33443# D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout GND.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X169 VDD.t180 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout VDD.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X170 VDD.t163 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X171 VDD.t990 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_0.Vout VDD.t988 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X172 a_112745_49858# VDD.t1113 GND.t113 GND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X173 VDD.t949 D_FlipFlop_7.3-input-nand_2.C.t4 D_FlipFlop_7.3-input-nand_2.Vout.t2 VDD.t948 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X174 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 VDD.t381 VDD.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X175 GND.t790 D_FlipFlop_2.3-input-nand_2.C.t5 a_130209_37007# GND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X176 Nand_Gate_1.Vout.t0 Nand_Gate_1.B.t4 VDD.t277 VDD.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X177 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 VDD.t218 VDD.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X178 GND.t748 Nand_Gate_0.A.t5 a_134897_37007# GND.t542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X179 Comparator_0.Vinm CDAC8_0.switch_7.Z.t118 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X180 a_69199_52572# RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_68585_52572# GND.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X181 Comparator_0.Vinm CDAC8_0.switch_7.Z.t117 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X182 GND.t1 Nand_Gate_7.A.t4 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B GND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X183 VDD.t561 Nand_Gate_4.B.t4 D_FlipFlop_7.3-input-nand_2.Vout.t3 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X184 Comparator_0.Vinm CDAC8_0.switch_7.Z.t116 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X185 Comparator_0.Vinm CDAC8_0.switch_9.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X186 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B Nand_Gate_2.B.t6 GND.t799 GND.t798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X187 GND.t192 Nand_Gate_4.B.t5 a_128851_19786# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X188 a_132311_26914# D_FlipFlop_5.3-input-nand_2.C.t5 D_FlipFlop_5.3-input-nand_2.Vout.t0 GND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X189 a_72835_13083# Nand_Gate_7.B.t5 RingCounter_0.D_FlipFlop_13.Qbar GND.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X190 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t752 VDD.t753 VDD.t457 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X191 a_77523_13083# RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 a_76909_13083# GND.t733 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X192 Comparator_0.Vinm CDAC8_0.switch_6.Z.t60 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X193 a_73579_52572# VDD.t1114 GND.t115 GND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X194 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK.t13 VDD.t1095 VDD.t1030 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X195 GND.t336 Nand_Gate_1.B.t5 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B GND.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X196 VDD.t210 FFCLR.t10 D_FlipFlop_6.Qbar VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X197 GND.t430 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 a_63767_15797# GND.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X198 GND.t250 And_Gate_2.Vout.t2 D_FlipFlop_5.Inverter_1.Vout GND.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X199 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 CLK.t14 a_63153_49858# GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X200 Comparator_0.Vinm CDAC8_0.switch_6.Z.t59 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X201 VDD.t1094 CLK.t15 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 VDD.t1050 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X202 VDD.t209 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X203 Comparator_0.Vinm CDAC8_0.switch_7.Z.t115 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X204 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 CLK.t16 VDD.t1093 VDD.t1060 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X205 Comparator_0.Vinm CDAC8_0.switch_6.Z.t58 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X206 a_132925_26914# D_FlipFlop_5.3-input-nand_0.Vout a_132311_26914# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X207 VDD.t977 And_Gate_4.A.t3 And_Gate_4.Nand_Gate_0.Vout VDD.t976 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X208 Comparator_0.Vinm CDAC8_0.switch_6.Z.t57 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X209 VDD.t154 Nand_Gate_4.B.t6 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B VDD.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X210 GND.t117 VDD.t1115 a_77523_13083# GND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X211 Comparator_0.Vinm CDAC8_0.switch_7.Z.t114 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X212 Comparator_0.Vinm CDAC8_0.switch_7.Z.t113 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X213 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 EN.t17 VDD.t521 VDD.t520 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X214 a_84489_15797# RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_83875_15797# GND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X215 Comparator_0.Vinm CDAC8_0.switch_9.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X216 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 a_78267_52572# GND.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X217 a_75898_25104# Q2.t4 VDD.t409 VDD.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X218 VDD.t843 Nand_Gate_2.A.t7 D_FlipFlop_3.3-input-nand_1.Vout VDD.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X219 a_128237_36157# D_FlipFlop_1.Qbar Q7.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X220 a_117609_13083# RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 a_116995_13083# GND.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X221 RingCounter_0.D_FlipFlop_11.Qbar RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 VDD.t870 VDD.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X222 VDD.t519 EN.t18 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 VDD.t518 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X223 VDD.t66 Nand_Gate_1.A.t4 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X224 VDD.t813 Q6.t5 CDAC8_0.switch_6.Z.t3 GND.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X225 a_128237_46849# D_FlipFlop_0.Qbar Q4.t0 GND.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X226 Comparator_0.Vinm CDAC8_0.switch_7.Z.t112 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X227 GND.t750 Nand_Gate_0.A.t6 a_132925_39721# GND.t749 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X228 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 VDD.t83 VDD.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X229 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_7.D.t7 VDD.t600 VDD.t599 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X230 a_83875_15797# RingCounter_0.D_FlipFlop_12.Qbar Nand_Gate_6.A.t2 GND.t627 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X231 VDD.t42 And_Gate_6.Vout.t2 D_FlipFlop_3.3-input-nand_0.Vout VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X232 a_88563_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 a_87949_15797# GND.t617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X233 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.3-input-nand_2.Vout.t5 VDD.t165 VDD.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X234 Comparator_0.Vinm CDAC8_0.switch_7.Z.t111 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X235 VDD.t1092 CLK.t17 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 VDD.t1091 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X236 Comparator_0.Vinm CDAC8_0.switch_7.Z.t110 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X237 GND.t565 EN.t19 a_84489_15797# GND.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X238 VDD.t789 Nand_Gate_6.B.t5 RingCounter_0.D_FlipFlop_11.Qbar VDD.t788 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X239 GND.t884 And_Gate_0.Vout.t2 D_FlipFlop_6.Inverter_1.Vout GND.t883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X240 VDD.t556 D_FlipFlop_0.CLK.t2 D_FlipFlop_0.3-input-nand_1.Vout VDD.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X241 VDD.t411 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Qbar VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X242 a_128237_30478# D_FlipFlop_4.Qbar Q3.t2 GND.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X243 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_0.3-input-nand_2.C.t4 VDD.t273 VDD.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X244 a_44403_13083# RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 a_43789_13083# GND.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X245 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 VDD.t134 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X246 CDAC8_0.switch_6.Z.t1 a_75898_39392# GND.t101 GND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X247 GND.t274 Nand_Gate_7.B.t6 a_132925_23350# GND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X248 And_Gate_7.Nand_Gate_0.Vout CLK.t18 VDD.t1090 VDD.t1089 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X249 And_Gate_5.A.t2 Nand_Gate_3.B.t6 VDD.t371 VDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X250 a_40459_52572# EN.t20 GND.t563 GND.t562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X251 GND.t119 VDD.t1116 a_117609_13083# GND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X252 VDD.t751 VDD.t750 RingCounter_0.D_FlipFlop_11.Qbar VDD.t473 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X253 a_134283_24200# And_Gate_2.Vout.t3 D_FlipFlop_5.3-input-nand_1.Vout GND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X254 VDD.t749 VDD.t748 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 VDD.t461 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X255 a_130209_44135# D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X256 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 Nand_Gate_7.A.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X257 a_132311_17072# D_FlipFlop_7.3-input-nand_2.Vout.t4 D_FlipFlop_7.3-input-nand_2.C.t2 GND.t858 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X258 VDD.t212 FFCLR.t11 Q7.t2 VDD.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X259 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 EN.t21 VDD.t517 VDD.t516 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X260 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_7.D.t8 VDD.t602 VDD.t601 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X261 a_134897_40571# D_FlipFlop_3.3-input-nand_1.B a_134283_40571# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X262 GND.t561 EN.t22 a_88563_15797# GND.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X263 Comparator_0.Vinm CDAC8_0.switch_8.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X264 a_132311_27764# D_FlipFlop_4.3-input-nand_2.Vout.t4 D_FlipFlop_4.3-input-nand_2.C.t2 GND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X265 VDD.t770 D_FlipFlop_4.3-input-nand_2.C.t4 D_FlipFlop_4.3-input-nand_2.Vout.t2 VDD.t769 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X266 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 VDD.t309 VDD.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X267 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 CLK.t19 VDD.t1088 VDD.t1056 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X268 a_29289_13083# RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 a_28675_13083# GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X269 Comparator_0.Vinm CDAC8_0.switch_7.Z.t109 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X270 VDD.t959 Nand_Gate_5.A.t5 Q4.t3 VDD.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X271 Comparator_0.Vinm CDAC8_0.switch_7.Z.t108 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X272 Comparator_0.Vinm CDAC8_0.switch_0.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X273 VDD.t375 RingCounter_0.D_FlipFlop_13.Qbar Nand_Gate_7.B.t1 VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X274 a_128851_43285# D_FlipFlop_3.Nand_Gate_0.Vout a_128237_43285# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X275 Comparator_0.Vinm CDAC8_0.switch_6.Z.t56 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X276 GND.t121 VDD.t1117 a_44403_13083# GND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X277 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 Nand_Gate_1.B.t6 VDD.t416 VDD.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X278 VDD.t417 Nand_Gate_1.B.t7 D_FlipFlop_4.3-input-nand_2.Vout.t1 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X279 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 VDD.t329 VDD.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X280 Comparator_0.Vinm CDAC8_0.switch_6.Z.t55 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X281 a_41073_52572# RingCounter_0.D_FlipFlop_16.Q.t4 a_40459_52572# GND.t676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X282 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_7.D.t9 VDD.t604 VDD.t603 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X283 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 a_76165_49858# GND.t768 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X284 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 a_45147_52572# GND.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X285 VDD.t286 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 VDD.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X286 a_132925_17072# D_FlipFlop_7.3-input-nand_1.Vout a_132311_17072# GND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X287 VDD.t414 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 VDD.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X288 VDD.t515 EN.t23 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 VDD.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X289 a_28675_13083# RingCounter_0.D_FlipFlop_16.Q.t5 RingCounter_0.D_FlipFlop_16.Qbar GND.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X290 a_122427_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 GND.t65 GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X291 GND.t877 Q3.t7 CDAC8_0.switch_5.Z.t3 VDD.t998 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X292 a_95659_49858# EN.t24 GND.t559 GND.t558 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X293 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 VDD.t828 VDD.t827 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X294 a_132925_27764# D_FlipFlop_4.3-input-nand_1.Vout a_132311_27764# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X295 GND.t123 VDD.t1118 a_29289_13083# GND.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X296 a_82057_16975# Nand_Gate_6.A.t5 GND.t82 GND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X297 Comparator_0.Vinm CDAC8_0.switch_7.Z.t107 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X298 a_50755_15797# RingCounter_0.D_FlipFlop_15.Qbar Nand_Gate_4.B.t1 GND.t349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X299 a_134283_20636# And_Gate_0.Vout.t3 D_FlipFlop_6.3-input-nand_1.Vout GND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X300 Comparator_0.Vinm CDAC8_0.switch_7.Z.t106 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X301 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 a_100347_52572# GND.t413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X302 Nand_Gate_0.A.t3 EN.t25 VDD.t507 VDD.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X303 a_55443_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 a_54829_15797# GND.t408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X304 Vbias.t8 a_138485_16882.t3 D_FlipFlop_7.D.t2 Vbias.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X305 VDD.t117 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X306 VDD.t3 Nand_Gate_7.A.t6 RingCounter_0.D_FlipFlop_14.Qbar VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X307 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 VDD.t851 VDD.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X308 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 VDD.t894 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X309 VDD.t156 Nand_Gate_4.B.t7 D_FlipFlop_7.3-input-nand_1.Vout VDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X310 a_107313_52572# Nand_Gate_2.B.t7 a_106699_52572# GND.t800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X311 Comparator_0.Vinm CDAC8_0.switch_6.Z.t54 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X312 VDD.t747 VDD.t746 RingCounter_0.D_FlipFlop_14.Qbar VDD.t469 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X313 Comparator_0.Vinm CDAC8_0.switch_7.Z.t105 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X314 a_96273_49858# RingCounter_0.D_FlipFlop_5.3-input-nand_1.B a_95659_49858# GND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X315 Comparator_0.Vinm CDAC8_0.switch_9.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X316 VDD.t290 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 VDD.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X317 Nand_Gate_5.B.t3 EN.t26 VDD.t513 VDD.t512 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X318 a_110643_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 a_110029_15797# GND.t756 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X319 CDAC8_0.switch_7.Z.t3 a_75898_35820# VDD.t885 VDD.t884 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X320 GND.t658 And_Gate_4.Vout.t3 D_FlipFlop_2.Inverter_1.Vout GND.t657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X321 Comparator_0.Vinm CDAC8_0.switch_9.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X322 VDD.t912 And_Gate_1.Vout.t3 D_FlipFlop_7.3-input-nand_0.Vout VDD.t911 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X323 a_90665_52572# EN.t27 GND.t557 GND.t556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X324 Comparator_0.Vinm CDAC8_0.switch_6.Z.t53 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X325 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 VDD.t150 VDD.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X326 GND.t555 EN.t28 a_55443_15797# GND.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X327 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.3-input-nand_2.Vout.t5 VDD.t971 VDD.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X328 GND.t236 FFCLR.t12 a_128851_40571# GND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X329 Nand_Gate_2.A.t1 RingCounter_0.D_FlipFlop_4.Qbar a_91279_52572# GND.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X330 VDD.t547 RingCounter_0.D_FlipFlop_10.Qbar Nand_Gate_1.B.t3 VDD.t546 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X331 Comparator_0.Vinm CDAC8_0.switch_7.Z.t104 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X332 GND.t203 Q5.t5 CDAC8_0.switch_9.Z.t0 VDD.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X333 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK.t20 a_107313_52572# GND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X334 And_Gate_1.Vout.t1 And_Gate_1.Nand_Gate_0.Vout GND.t807 GND.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X335 a_74807_13083# RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 GND.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X336 a_70645_16975# CLK.t21 GND.t70 GND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X337 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 EN.t29 VDD.t511 VDD.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X338 Comparator_0.Vinm CDAC8_0.switch_8.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X339 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 a_43045_49858# GND.t878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X340 a_79495_13083# RingCounter_0.D_FlipFlop_13.3-input-nand_1.B a_78881_13083# GND.t755 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X341 GND.t553 EN.t30 a_110643_15797# GND.t552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X342 a_120325_49858# RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 a_119711_49858# GND.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X343 a_75551_52572# EN.t31 GND.t551 GND.t550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X344 VDD.t901 Q1.t4 D_FlipFlop_6.Qbar VDD.t856 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X345 RingCounter_0.D_FlipFlop_9.Qbar RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 VDD.t635 VDD.t634 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X346 VDD.t774 Nand_Gate_1.A.t5 Nand_Gate_1.Vout.t2 VDD.t773 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X347 VDD.t92 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X348 a_62539_49858# EN.t32 GND.t549 GND.t548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X349 GND.t547 EN.t33 a_57415_13083# GND.t546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X350 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 VDD.t744 VDD.t745 VDD.t475 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X351 a_128851_19786# D_FlipFlop_7.Nand_Gate_0.Vout a_128237_19786# GND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X352 D_FlipFlop_5.3-input-nand_2.C.t3 D_FlipFlop_5.3-input-nand_1.Vout VDD.t979 VDD.t567 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X353 a_134897_26914# D_FlipFlop_7.D.t10 a_134283_26914# GND.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X354 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 VDD.t281 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X355 a_76909_13083# RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 GND.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X356 Comparator_0.Vinm CDAC8_0.switch_7.Z.t103 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X357 GND.t238 FFCLR.t13 a_132925_36157# GND.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X358 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 VDD.t111 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X359 a_89307_49858# RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 GND.t233 GND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X360 GND.t545 EN.t34 a_112615_13083# GND.t544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X361 VDD.t509 EN.t35 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 VDD.t508 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X362 a_134283_37007# And_Gate_4.Vout.t4 D_FlipFlop_2.3-input-nand_1.Vout GND.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X363 a_76165_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_75551_52572# GND.t866 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X364 D_FlipFlop_6.Qbar D_FlipFlop_6.Nand_Gate_1.Vout VDD.t404 VDD.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X365 VDD.t743 VDD.t742 RingCounter_0.D_FlipFlop_9.Qbar VDD.t467 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X366 VDD.t236 RingCounter_0.D_FlipFlop_16.Qbar RingCounter_0.D_FlipFlop_16.Q.t1 VDD.t235 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X367 GND.t394 Nand_Gate_5.A.t6 a_132925_46849# GND.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X368 Comparator_0.Vinm CDAC8_0.switch_6.Z.t52 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X369 a_63153_49858# RingCounter_0.D_FlipFlop_2.3-input-nand_1.B a_62539_49858# GND.t864 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X370 And_Gate_3.Nand_Gate_0.Vout Nand_Gate_1.Vout.t3 a_114805_16975# GND.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X371 And_Gate_1.B.t0 Nand_Gate_4.B.t8 a_37897_16975# GND.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X372 VDD.t18 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X373 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 a_67227_49858# GND.t587 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X374 Comparator_0.Vinm CDAC8_0.switch_7.Z.t102 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X375 GND.t367 D_FlipFlop_2.3-input-nand_2.Vout.t4 a_130209_39721# GND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X376 Comparator_0.Vinm CDAC8_0.switch_9.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X377 VDD.t200 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X378 GND.t240 FFCLR.t14 a_134897_39721# GND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X379 Comparator_0.Vinm CDAC8_0.switch_6.Z.t51 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X380 a_85847_15797# RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout GND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X381 VDD.t606 D_FlipFlop_7.D.t11 D_FlipFlop_3.3-input-nand_1.B VDD.t605 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X382 GND.t468 Nand_Gate_1.B.t8 a_132925_30478# GND.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X383 Comparator_0.Vinm CDAC8_0.switch_7.Z.t101 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X384 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 a_122427_49858# GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X385 a_118967_13083# RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 GND.t879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X386 GND.t463 Q2.t5 CDAC8_0.switch_0.Z.t3 VDD.t410 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X387 GND.t608 D_FlipFlop_6.3-input-nand_2.Vout.t4 a_130209_23350# GND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X388 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.3-input-nand_1.B VDD.t121 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X389 Comparator_0.Vinm CDAC8_0.switch_8.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X390 GND.t242 FFCLR.t15 a_134897_23350# GND.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X391 GND.t125 VDD.t1119 a_68455_15797# GND.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X392 a_42431_52572# VDD.t1120 GND.t127 GND.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X393 VDD.t419 Nand_Gate_1.B.t9 D_FlipFlop_4.3-input-nand_1.Vout VDD.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X394 Comparator_0.Vinm CDAC8_0.switch_9.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X395 VDD.t169 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X396 VDD.t115 D_FlipFlop_1.Qbar Q7.t0 VDD.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X397 VDD.t505 EN.t36 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 VDD.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X398 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 VDD.t740 VDD.t741 VDD.t471 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X399 a_87949_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 GND.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X400 VDD.t363 D_FlipFlop_0.Qbar Q4.t1 VDD.t362 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X401 VDD.t5 And_Gate_3.Vout.t3 D_FlipFlop_4.3-input-nand_0.Vout VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X402 GND.t129 VDD.t1121 a_123655_15797# GND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X403 a_43789_13083# RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 GND.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X404 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.3-input-nand_2.Vout.t5 VDD.t928 VDD.t771 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X405 VDD.t96 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 VDD.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X406 Comparator_0.Vinm CDAC8_0.switch_7.Z.t100 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X407 GND.t681 Nand_Gate_6.B.t6 a_128851_26914# GND.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X408 VDD.t214 FFCLR.t16 And_Gate_5.A.t0 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X409 a_102319_52572# RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_101705_52572# GND.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X410 Comparator_0.Vinm CDAC8_0.switch_0.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X411 Comparator_0.Vinm CDAC8_0.switch_7.Z.t99 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X412 a_43045_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 a_42431_52572# GND.t760 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X413 VDD.t1087 CLK.t22 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 VDD.t1018 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X414 a_91279_49858# RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 a_90665_49858# GND.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X415 VDD.t850 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_7.Qbar VDD.t431 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X416 FFCLR.t2 RingCounter_0.D_FlipFlop_17.Qbar a_47119_52572# GND.t708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X417 Q7.t3 D_FlipFlop_1.Nand_Gate_0.Vout VDD.t615 VDD.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X418 a_134897_17072# D_FlipFlop_7.3-input-nand_1.B a_134283_17072# GND.t865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X419 VDD.t739 VDD.t738 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 VDD.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X420 VDD.t978 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X421 a_97631_49858# VDD.t1122 GND.t131 GND.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X422 RingCounter_0.D_FlipFlop_1.Qbar Nand_Gate_3.B.t7 VDD.t372 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X423 VDD.t197 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 VDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X424 Q4.t2 D_FlipFlop_0.Nand_Gate_0.Vout VDD.t398 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X425 a_134897_27764# D_FlipFlop_4.3-input-nand_1.B a_134283_27764# GND.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X426 And_Gate_6.Vout.t1 And_Gate_6.Nand_Gate_0.Vout GND.t758 GND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X427 VDD.t1086 CLK.t23 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 VDD.t1016 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X428 a_52727_15797# RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout GND.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X429 Comparator_0.Vinm CDAC8_0.switch_7.Z.t98 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X430 Nand_Gate_2.B.t0 RingCounter_0.D_FlipFlop_5.Qbar a_102319_52572# GND.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X431 a_57415_15797# Nand_Gate_7.A.t7 a_56801_15797# GND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X432 Comparator_0.Vinm CDAC8_0.switch_9.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X433 a_128237_33443# Q7.t5 D_FlipFlop_1.Qbar GND.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X434 Nand_Gate_7.A.t3 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t1101 VDD.t892 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X435 Comparator_0.Vinm CDAC8_0.switch_7.Z.t97 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X436 a_75898_42964# Q5.t6 GND.t205 GND.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X437 RingCounter_0.D_FlipFlop_7.Qbar Nand_Gate_5.A.t7 VDD.t350 VDD.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X438 GND.t264 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 a_30647_15797# GND.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X439 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B VDD.t586 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X440 a_75898_46095# Q4.t4 GND.t374 GND.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X441 GND.t133 VDD.t1123 a_35335_15797# GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X442 CDAC8_0.switch_5.Z.t0 a_75898_28676# VDD.t123 VDD.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X443 VDD.t945 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 VDD.t944 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X444 And_Gate_2.Nand_Gate_0.Vout Nand_Gate_6.Vout.t3 VDD.t400 VDD.t399 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X445 a_98245_49858# RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 a_97631_49858# GND.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X446 a_112615_15797# Nand_Gate_1.B.t10 a_112001_15797# GND.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X447 a_67227_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 GND.t312 GND.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X448 Comparator_0.Vinm CDAC8_0.switch_6.Z.t50 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X449 VDD.t503 EN.t37 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 VDD.t502 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X450 Comparator_0.Vinm CDAC8_0.switch_9.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X451 VDD.t501 EN.t38 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 VDD.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X452 a_54829_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 GND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X453 VDD.t608 D_FlipFlop_7.D.t12 D_FlipFlop_7.3-input-nand_1.B VDD.t607 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X454 Comparator_0.Vinm CDAC8_0.switch_7.Z.t96 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X455 VDD.t159 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X456 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B VDD.t573 VDD.t572 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X457 Comparator_0.Vinm CDAC8_0.switch_7.Z.t95 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X458 Comparator_0.Vinm CDAC8_0.switch_5.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X459 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.3-input-nand_1.B VDD.t981 VDD.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X460 a_106699_52572# VDD.t1124 GND.t135 GND.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X461 Comparator_0.Vinm CDAC8_0.switch_7.Z.t94 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X462 VDD.t387 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 VDD.t386 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X463 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B Nand_Gate_2.B.t8 VDD.t920 VDD.t919 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X464 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 VDD.t946 VDD.t632 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X465 VDD.t499 EN.t39 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 VDD.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X466 D_FlipFlop_2.3-input-nand_2.C.t2 D_FlipFlop_2.3-input-nand_1.Vout VDD.t430 VDD.t429 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X467 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 EN.t40 VDD.t497 VDD.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X468 Comparator_0.Vinm CDAC8_0.switch_2.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X469 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B Nand_Gate_0.A.t7 GND.t752 GND.t751 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X470 GND.t225 CLK.t24 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 GND.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X471 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t736 VDD.t737 VDD.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X472 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 VDD.t565 VDD.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X473 VDD.t105 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X474 Comparator_0.Vinm CDAC8_0.switch_6.Z.t49 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X475 VDD.t891 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X476 GND.t421 FFCLR.t17 a_128851_17072# GND.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X477 a_132311_24200# D_FlipFlop_5.3-input-nand_2.Vout.t4 D_FlipFlop_5.3-input-nand_2.C.t0 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X478 a_64511_49858# VDD.t1125 GND.t137 GND.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X479 VDD.t991 D_FlipFlop_5.3-input-nand_2.C.t6 D_FlipFlop_5.3-input-nand_2.Vout.t1 VDD.t597 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X480 a_128851_40571# D_FlipFlop_3.Nand_Gate_1.Vout a_128237_40571# GND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X481 Comparator_0.Vinm CDAC8_0.switch_6.Z.t48 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X482 Comparator_0.Vinm CDAC8_0.switch_7.Z.t93 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X483 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 CLK.t25 VDD.t1085 VDD.t1084 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X484 GND.t84 Nand_Gate_6.A.t6 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X485 CDAC8_0.switch_9.Z.t2 a_75898_42964# VDD.t986 VDD.t985 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X486 VDD.t566 a_138485_16882.t0 Vbias.t2 sky130_fd_pr__res_xhigh_po_5p73 l=150
X487 VDD.t790 Nand_Gate_6.B.t7 D_FlipFlop_5.3-input-nand_2.Vout.t3 VDD.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X488 GND.t423 FFCLR.t18 a_128851_27764# GND.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X489 Comparator_0.Vinm CDAC8_0.switch_7.Z.t92 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X490 GND.t853 D_FlipFlop_1.3-input-nand_2.Vout.t5 a_130209_36157# GND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X491 Comparator_0.Vinm CDAC8_0.switch_9.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X492 GND.t543 EN.t41 a_134897_36157# GND.t542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X493 GND.t683 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 a_63767_13083# GND.t682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X494 Comparator_0.Vinm CDAC8_0.switch_7.Z.t91 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X495 VDD.t44 And_Gate_6.Vout.t3 D_FlipFlop_3.Inverter_1.Vout VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X496 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B VDD.t152 VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X497 a_75898_25104# Q2.t6 GND.t48 GND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X498 VDD.t872 Nand_Gate_0.A.t8 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t871 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X499 GND.t266 D_FlipFlop_0.3-input-nand_2.Vout.t5 a_130209_46849# GND.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X500 a_124399_49858# RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 a_123785_49858# GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X501 VDD.t1083 CLK.t26 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 VDD.t1082 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X502 a_68585_49858# VDD.t1126 GND.t139 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X503 GND.t425 FFCLR.t19 a_134897_46849# GND.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X504 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 VDD.t238 VDD.t237 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X505 a_116995_15797# RingCounter_0.D_FlipFlop_10.Qbar Nand_Gate_1.B.t2 GND.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X506 a_132925_24200# D_FlipFlop_5.3-input-nand_1.Vout a_132311_24200# GND.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X507 a_65125_49858# RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 a_64511_49858# GND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X508 VDD.t910 D_FlipFlop_2.3-input-nand_2.C.t6 D_FlipFlop_2.3-input-nand_2.Vout.t1 VDD.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X509 Comparator_0.Vinm CDAC8_0.switch_7.Z.t90 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X510 RingCounter_0.D_FlipFlop_2.Qbar Nand_Gate_0.A.t9 a_69199_49858# GND.t753 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X511 a_75898_18814# Q0.t4 GND.t695 GND.t694 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X512 And_Gate_4.Vout.t0 And_Gate_4.Nand_Gate_0.Vout VDD.t171 VDD.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X513 a_84489_13083# RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 a_83875_13083# GND.t775 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X514 VDD.t873 Nand_Gate_0.A.t10 D_FlipFlop_2.3-input-nand_2.Vout.t2 VDD.t642 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X515 GND.t804 D_FlipFlop_4.3-input-nand_2.Vout.t6 a_130209_30478# GND.t674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X516 Comparator_0.Vinm CDAC8_0.switch_7.Z.t89 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X517 Comparator_0.Vinm CDAC8_0.switch_7.Z.t88 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X518 a_123785_49858# VDD.t1127 GND.t141 GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X519 GND.t426 FFCLR.t20 a_134897_30478# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X520 Comparator_0.Vinm CDAC8_0.switch_9.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X521 VDD.t232 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 VDD.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X522 Comparator_0.Vinm CDAC8_0.switch_5.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X523 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 VDD.t98 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X524 a_132311_20636# D_FlipFlop_6.3-input-nand_2.Vout.t5 D_FlipFlop_6.3-input-nand_2.C.t2 GND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X525 VDD.t579 D_FlipFlop_6.3-input-nand_2.C.t5 D_FlipFlop_6.3-input-nand_2.Vout.t1 VDD.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X526 a_80239_52572# RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_79625_52572# GND.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X527 RingCounter_0.D_FlipFlop_6.Qbar Nand_Gate_5.B.t5 a_124399_49858# GND.t875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X528 a_128237_44135# Q4.t5 D_FlipFlop_0.Qbar GND.t375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X529 VDD.t240 Nand_Gate_7.B.t7 D_FlipFlop_6.3-input-nand_2.Vout.t3 VDD.t239 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X530 a_83875_13083# Nand_Gate_6.A.t7 RingCounter_0.D_FlipFlop_12.Qbar GND.t686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X531 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 EN.t42 VDD.t495 VDD.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X532 a_88563_13083# RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 a_87949_13083# GND.t710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X533 a_139804_27676.t1 Vin.t0 a_138533_35417.t0 Vbias.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X534 a_108671_49858# VDD.t1128 GND.t143 GND.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X535 GND.t145 VDD.t1129 a_84489_13083# GND.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X536 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK.t27 VDD.t1081 VDD.t1004 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X537 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 CLK.t28 VDD.t1080 VDD.t1079 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X538 a_89921_15797# CLK.t29 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 GND.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X539 Comparator_0.Vinm CDAC8_0.switch_7.Z.t87 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X540 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 a_109285_49858# GND.t405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X541 a_132925_20636# D_FlipFlop_6.3-input-nand_1.Vout a_132311_20636# GND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X542 CDAC8_0.switch_0.Z.t0 a_75898_25104# VDD.t138 VDD.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X543 VDD.t610 D_FlipFlop_7.D.t13 D_FlipFlop_4.3-input-nand_1.B VDD.t609 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X544 VDD.t376 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X545 VDD.t383 FFCLR.t21 D_FlipFlop_5.Qbar VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X546 a_134283_39721# And_Gate_4.Vout.t5 D_FlipFlop_2.3-input-nand_0.Vout GND.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X547 And_Gate_4.A.t1 Nand_Gate_0.B.t4 VDD.t129 VDD.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X548 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 CLK.t30 VDD.t1078 VDD.t1032 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X549 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.3-input-nand_1.B VDD.t982 VDD.t806 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X550 VDD.t887 RingCounter_0.D_FlipFlop_16.Q.t6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 VDD.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X551 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 CLK.t31 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X552 VDD.t125 Nand_Gate_7.A.t8 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B VDD.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X553 GND.t147 VDD.t1130 a_88563_13083# GND.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X554 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 VDD.t295 VDD.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X555 a_109285_49858# RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 a_108671_49858# GND.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X556 a_95529_15797# RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_94915_15797# GND.t582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X557 Comparator_0.Vinm CDAC8_0.switch_7.Z.t86 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X558 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 CLK.t32 GND.t260 GND.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X559 a_134283_23350# And_Gate_0.Vout.t4 D_FlipFlop_6.3-input-nand_0.Vout GND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X560 Comparator_0.Vinm CDAC8_0.switch_9.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X561 GND.t541 EN.t43 a_132925_33443# GND.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X562 D_FlipFlop_0.CLK.t0 And_Gate_7.Nand_Gate_0.Vout VDD.t630 VDD.t629 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X563 Comparator_0.Vinm CDAC8_0.switch_7.Z.t85 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X564 a_130209_43285# D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X565 VDD.t1075 CLK.t33 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 VDD.t1074 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X566 VDD.t304 Nand_Gate_1.B.t11 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B VDD.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X567 a_128851_26914# D_FlipFlop_5.Nand_Gate_0.Vout a_128237_26914# GND.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X568 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 VDD.t379 VDD.t378 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X569 Comparator_0.Vinm CDAC8_0.switch_7.Z.t84 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X570 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 VDD.t389 VDD.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X571 VDD.t914 And_Gate_1.Vout.t4 D_FlipFlop_7.Inverter_1.Vout VDD.t913 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X572 RingCounter_0.D_FlipFlop_3.Qbar VDD.t734 VDD.t735 VDD.t459 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X573 Comparator_0.Vinm CDAC8_0.switch_9.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X574 VDD.t348 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout VDD.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X575 a_47119_52572# RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 a_46505_52572# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X576 Comparator_0.Vinm CDAC8_0.switch_6.Z.t47 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X577 a_50755_13083# Nand_Gate_4.B.t9 RingCounter_0.D_FlipFlop_15.Qbar GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X578 Comparator_0.Vinm CDAC8_0.switch_8.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X579 GND.t540 EN.t44 a_95529_15797# GND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X580 VDD.t264 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_1.Qbar VDD.t263 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X581 a_132311_37007# D_FlipFlop_2.3-input-nand_2.Vout.t5 D_FlipFlop_2.3-input-nand_2.C.t1 GND.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X582 a_55443_13083# RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 a_54829_13083# GND.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X583 Comparator_0.Vinm CDAC8_0.switch_7.Z.t83 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X584 And_Gate_5.Nand_Gate_0.Vout CLK.t34 VDD.t1073 VDD.t1072 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X585 Comparator_0.Vinm CDAC8_0.switch_6.Z.t46 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X586 Comparator_0.Vinm CDAC8_0.switch_6.Z.t45 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X587 D_FlipFlop_1.3-input-nand_2.C.t3 D_FlipFlop_1.3-input-nand_1.Vout VDD.t550 VDD.t412 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X588 Comparator_0.Vinm CDAC8_0.switch_6.Z.t44 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X589 VDD.t733 VDD.t732 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 VDD.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X590 a_56801_15797# CLK.t35 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 GND.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X591 VDD.t426 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 VDD.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X592 Nand_Gate_2.A.t3 EN.t45 VDD.t493 VDD.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X593 VDD.t177 Q5.t7 CDAC8_0.switch_9.Z.t1 GND.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X594 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK.t36 a_41073_49858# GND.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X595 VDD.t1071 CLK.t37 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 VDD.t1022 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X596 a_110643_13083# RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 a_110029_13083# GND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X597 Comparator_0.Vinm CDAC8_0.switch_7.Z.t82 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X598 VDD.t781 Q4.t6 CDAC8_0.switch_8.Z.t2 GND.t678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X599 Nand_Gate_5.Vout.t2 Nand_Gate_5.B.t6 VDD.t647 VDD.t646 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X600 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 CLK.t38 VDD.t1070 VDD.t1028 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X601 VDD.t591 RingCounter_0.D_FlipFlop_12.Qbar Nand_Gate_6.A.t3 VDD.t590 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X602 VDD.t1069 CLK.t39 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 VDD.t1068 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X603 a_112001_15797# CLK.t40 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 GND.t414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X604 a_132925_37007# D_FlipFlop_2.3-input-nand_1.Vout a_132311_37007# GND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X605 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK.t41 a_74193_52572# GND.t415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X606 GND.t149 VDD.t1131 a_55443_13083# GND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X607 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 VDD.t582 VDD.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X608 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 EN.t46 VDD.t491 VDD.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X609 a_62409_15797# RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_61795_15797# GND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X610 CDAC8_0.switch_9.Z.t3 a_75898_42964# GND.t869 GND.t868 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X611 VDD.t1067 CLK.t42 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 VDD.t1020 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X612 VDD.t924 And_Gate_2.Vout.t4 D_FlipFlop_5.3-input-nand_0.Vout VDD.t923 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X613 CDAC8_0.switch_8.Z.t1 a_75898_46095# GND.t231 GND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X614 And_Gate_5.Nand_Gate_0.Vout CLK.t43 a_59605_47663# GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X615 RingCounter_0.D_FlipFlop_13.Qbar RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 VDD.t40 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X616 VDD.t489 EN.t47 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 VDD.t488 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X617 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.3-input-nand_2.Vout.t5 VDD.t596 VDD.t595 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X618 Comparator_0.Vinm CDAC8_0.switch_9.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X619 Comparator_0.Vinm CDAC8_0.switch_7.Z.t81 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X620 GND.t151 VDD.t1132 a_110643_13083# GND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X621 And_Gate_0.Vout.t1 And_Gate_0.Nand_Gate_0.Vout GND.t216 GND.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X622 Comparator_0.Vinm CDAC8_0.switch_7.Z.t80 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X623 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 VDD.t570 VDD.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X624 VDD.t167 D_FlipFlop_3.3-input-nand_2.Vout.t6 D_FlipFlop_3.3-input-nand_2.C.t1 VDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X625 a_66483_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 a_65869_15797# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X626 VDD.t385 FFCLR.t22 D_FlipFlop_3.3-input-nand_2.C.t0 VDD.t384 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X627 Comparator_0.Vinm CDAC8_0.switch_6.Z.t43 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X628 VDD.t1106 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 VDD.t848 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X629 VDD.t983 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 VDD.t794 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X630 GND.t538 EN.t48 a_62409_15797# GND.t537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X631 a_128851_17072# D_FlipFlop_7.Nand_Gate_1.Vout a_128237_17072# GND.t687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X632 Comparator_0.Vinm CDAC8_0.switch_5.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X633 a_134897_24200# D_FlipFlop_5.3-input-nand_1.B a_134283_24200# GND.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X634 a_118353_52572# Nand_Gate_5.A.t8 a_117739_52572# GND.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X635 VDD.t658 And_Gate_4.Vout.t6 D_FlipFlop_2.3-input-nand_0.Vout VDD.t657 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X636 And_Gate_6.Nand_Gate_0.Vout CLK.t44 VDD.t1066 VDD.t1065 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X637 VDD.t731 VDD.t730 RingCounter_0.D_FlipFlop_13.Qbar VDD.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X638 VDD.t242 Nand_Gate_7.B.t8 D_FlipFlop_6.3-input-nand_1.Vout VDD.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X639 a_130209_19786# D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X640 a_128851_27764# D_FlipFlop_4.Nand_Gate_1.Vout a_128237_27764# GND.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X641 Comparator_0.Vinm CDAC8_0.switch_7.Z.t79 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X642 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t173 VDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X643 Comparator_0.Vinm CDAC8_0.switch_6.Z.t42 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X644 Comparator_0.Vinm CDAC8_0.switch_6.Z.t41 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X645 a_121683_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 a_121069_15797# GND.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X646 Comparator_0.Vinm CDAC8_0.switch_6.Z.t40 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X647 Comparator_0.Vinm CDAC8_0.switch_7.Z.t78 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X648 GND.t428 FFCLR.t23 a_132925_44135# GND.t427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X649 a_75898_46095# Q4.t7 VDD.t783 VDD.t782 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X650 VDD.t1064 CLK.t45 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 VDD.t1014 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X651 VDD.t53 Q2.t7 CDAC8_0.switch_0.Z.t2 GND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X652 VDD.t831 And_Gate_0.Vout.t5 D_FlipFlop_6.3-input-nand_0.Vout VDD.t830 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X653 Comparator_0.Vinm CDAC8_0.switch_6.Z.t39 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X654 Comparator_0.Vinm CDAC8_0.switch_7.Z.t77 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X655 VDD.t127 Nand_Gate_7.A.t9 And_Gate_0.B.t0 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X656 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.3-input-nand_2.Vout.t6 VDD.t636 VDD.t580 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X657 VDD.t7 And_Gate_3.Vout.t4 D_FlipFlop_4.Inverter_1.Vout VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X658 VDD.t293 RingCounter_0.D_FlipFlop_15.Qbar Nand_Gate_4.B.t0 VDD.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X659 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK.t46 a_118353_52572# GND.t417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X660 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 VDD.t374 VDD.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X661 a_69199_49858# RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 a_68585_49858# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X662 And_Gate_0.B.t2 Nand_Gate_7.B.t9 a_59977_16975# GND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X663 a_85847_13083# RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 GND.t637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X664 VDD.t10 FFCLR.t24 D_FlipFlop_2.Qbar VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X665 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 VDD.t728 VDD.t729 VDD.t534 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X666 a_106569_15797# RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_105955_15797# GND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X667 VDD.t805 Q0.t5 CDAC8_0.switch_1.Z.t3 GND.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X668 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 EN.t49 VDD.t487 VDD.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X669 a_134283_36157# And_Gate_5.Vout.t3 D_FlipFlop_1.3-input-nand_0.Vout GND.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X670 D_FlipFlop_3.3-input-nand_2.Vout.t1 D_FlipFlop_3.3-input-nand_0.Vout VDD.t221 VDD.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X671 CDAC8_0.switch_0.Z.t1 a_75898_25104# GND.t186 GND.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X672 RingCounter_0.D_FlipFlop_10.Qbar RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 VDD.t194 VDD.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X673 RingCounter_0.D_FlipFlop_8.Qbar RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 VDD.t327 VDD.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X674 VDD.t485 EN.t50 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 VDD.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X675 a_100347_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 GND.t411 GND.t410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X676 a_134283_46849# D_FlipFlop_0.CLK.t3 D_FlipFlop_0.3-input-nand_0.Vout GND.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X677 D_FlipFlop_0.3-input-nand_2.C.t0 D_FlipFlop_0.3-input-nand_1.Vout VDD.t108 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X678 VDD.t144 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X679 a_73579_49858# EN.t51 GND.t536 GND.t535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X680 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 a_87205_52572# GND.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X681 GND.t534 EN.t52 a_68455_13083# GND.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X682 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 VDD.t877 VDD.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X683 And_Gate_3.Vout.t1 And_Gate_3.Nand_Gate_0.Vout GND.t356 GND.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X684 a_134897_20636# D_FlipFlop_6.3-input-nand_1.B a_134283_20636# GND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X685 Comparator_0.Vinm CDAC8_0.switch_7.Z.t76 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X686 VDD.t55 Q2.t8 D_FlipFlop_5.Qbar VDD.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X687 CDAC8_0.switch_1.Z.t1 a_75898_18814# GND.t22 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X688 VDD.t587 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_2.B.t3 VDD.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X689 Comparator_0.Vinm CDAC8_0.switch_9.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X690 GND.t736 D_FlipFlop_7.D.t14 D_FlipFlop_2.3-input-nand_1.B GND.t735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X691 FFCLR.t1 VDD.t726 VDD.t727 VDD.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X692 a_33363_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_32749_15797# GND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X693 a_139663_37417.t1 a_139663_37417.t0 VDD.t90 VDD.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X694 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 VDD.t377 VDD.t314 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X695 GND.t153 VDD.t1133 a_90535_15797# GND.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X696 a_87949_13083# RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 GND.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X697 VDD.t203 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 VDD.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X698 GND.t532 EN.t53 a_106569_15797# GND.t531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X699 a_134283_30478# And_Gate_3.Vout.t5 D_FlipFlop_4.3-input-nand_0.Vout GND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X700 FFCLR.t3 RingCounter_0.D_FlipFlop_17.Qbar VDD.t819 VDD.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X701 VDD.t723 VDD.t722 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 VDD.t449 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X702 GND.t530 EN.t54 a_123655_13083# GND.t529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X703 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 VDD.t822 VDD.t821 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X704 VDD.t179 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout VDD.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X705 Nand_Gate_2.Vout.t1 Nand_Gate_2.B.t9 a_93097_47663# GND.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X706 GND.t314 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 a_96887_15797# GND.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X707 VDD.t725 VDD.t724 RingCounter_0.D_FlipFlop_8.Qbar VDD.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X708 GND.t6 FFCLR.t25 a_128851_24200# GND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X709 GND.t675 D_FlipFlop_1.3-input-nand_2.C.t5 a_130209_33443# GND.t674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X710 VDD.t656 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_3.Qbar VDD.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X711 VDD.t627 RingCounter_0.D_FlipFlop_8.Qbar Nand_Gate_4.A.t3 VDD.t626 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X712 GND.t738 D_FlipFlop_7.D.t15 D_FlipFlop_6.3-input-nand_1.B GND.t737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X713 Nand_Gate_2.B.t2 EN.t55 VDD.t483 VDD.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X714 GND.t8 FFCLR.t26 a_134897_33443# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X715 VDD.t481 EN.t56 D_FlipFlop_1.3-input-nand_0.Vout VDD.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X716 VDD.t972 D_FlipFlop_7.3-input-nand_2.Vout.t6 D_FlipFlop_7.3-input-nand_2.C.t3 VDD.t948 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X717 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 a_78267_49858# GND.t848 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X718 Comparator_0.Vinm CDAC8_0.switch_7.Z.t75 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X719 D_FlipFlop_5.Qbar D_FlipFlop_5.Nand_Gate_1.Vout VDD.t936 VDD.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X720 VDD.t620 Nand_Gate_0.A.t11 And_Gate_4.A.t2 VDD.t619 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X721 Comparator_0.Vinm CDAC8_0.switch_7.Z.t74 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X722 Comparator_0.Vinm CDAC8_0.switch_7.Z.t73 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X723 Nand_Gate_2.B.t1 RingCounter_0.D_FlipFlop_5.Qbar VDD.t306 VDD.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X724 Comparator_0.Vinm CDAC8_0.switch_7.Z.t72 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X725 VDD.t12 FFCLR.t27 D_FlipFlop_0.3-input-nand_0.Vout VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X726 GND.t528 EN.t57 a_33363_15797# GND.t527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X727 VDD.t14 FFCLR.t28 D_FlipFlop_7.3-input-nand_2.C.t1 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X728 RingCounter_0.D_FlipFlop_16.Qbar RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 VDD.t862 VDD.t427 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X729 a_96887_15797# RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout GND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X730 VDD.t973 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 VDD.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X731 Comparator_0.Vinm CDAC8_0.switch_6.Z.t38 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X732 Nand_Gate_1.Vout.t1 Nand_Gate_1.B.t12 a_104137_16975# GND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X733 a_52727_13083# RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 GND.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X734 And_Gate_1.Nand_Gate_0.Vout And_Gate_1.B.t3 VDD.t955 VDD.t954 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X735 RingCounter_0.D_FlipFlop_3.Qbar Nand_Gate_0.B.t5 VDD.t130 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X736 a_57415_13083# RingCounter_0.D_FlipFlop_15.3-input-nand_1.B a_56801_13083# GND.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X737 Comparator_0.Vinm CDAC8_0.switch_5.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X738 a_53471_52572# EN.t58 GND.t526 GND.t525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X739 GND.t278 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 a_30647_13083# GND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X740 VDD.t345 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X741 a_40459_49858# VDD.t1134 GND.t155 GND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X742 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 a_54085_52572# GND.t369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X743 GND.t524 EN.t59 a_35335_13083# GND.t523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X744 VDD.t1063 CLK.t47 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 VDD.t1062 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X745 Comparator_0.Vinm CDAC8_0.switch_6.Z.t37 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X746 And_Gate_4.Nand_Gate_0.Vout CLK.t48 a_81685_47663# GND.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X747 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 VDD.t720 VDD.t721 VDD.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X748 VDD.t719 VDD.t718 RingCounter_0.D_FlipFlop_16.Qbar VDD.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X749 Comparator_0.Vinm CDAC8_0.switch_6.Z.t36 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X750 a_112615_13083# RingCounter_0.D_FlipFlop_9.3-input-nand_1.B a_112001_13083# GND.t867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X751 GND.t10 FFCLR.t29 a_128851_20636# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X752 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B VDD.t859 VDD.t858 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X753 Comparator_0.Vinm CDAC8_0.switch_7.Z.t71 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X754 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t820 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X755 a_54829_13083# RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X756 Comparator_0.Vinm CDAC8_0.switch_9.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X757 a_134897_37007# D_FlipFlop_2.3-input-nand_1.B a_134283_37007# GND.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X758 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B Nand_Gate_0.A.t12 VDD.t622 VDD.t621 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X759 a_113359_52572# RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_112745_52572# GND.t474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X760 D_FlipFlop_7.3-input-nand_2.Vout.t0 D_FlipFlop_7.3-input-nand_0.Vout VDD.t288 VDD.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X761 a_54085_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_53471_52572# GND.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X762 Comparator_0.Vinm CDAC8_0.switch_7.Z.t70 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X763 a_81685_47663# And_Gate_4.A.t4 GND.t863 GND.t862 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X764 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 EN.t60 VDD.t479 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X765 Nand_Gate_3.B.t0 RingCounter_0.D_FlipFlop_1.Qbar a_58159_52572# GND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X766 VDD.t332 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_6.Qbar VDD.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X767 a_41073_49858# RingCounter_0.D_FlipFlop_17.3-input-nand_1.B a_40459_49858# GND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X768 VDD.t864 D_FlipFlop_7.D.t16 D_FlipFlop_5.3-input-nand_1.B VDD.t863 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X769 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 VDD.t85 VDD.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X770 Comparator_0.Vinm CDAC8_0.switch_7.Z.t69 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X771 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 VDD.t905 VDD.t593 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X772 VDD.t717 VDD.t716 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 VDD.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X773 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 a_45147_49858# GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X774 And_Gate_2.Vout.t0 And_Gate_2.Nand_Gate_0.Vout VDD.t584 VDD.t583 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X775 VDD.t352 Nand_Gate_5.A.t9 Nand_Gate_5.Vout.t0 VDD.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X776 RingCounter_0.D_FlipFlop_2.Qbar Nand_Gate_0.A.t13 VDD.t623 VDD.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X777 a_122427_49858# RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 GND.t347 GND.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X778 VDD.t45 And_Gate_6.Vout.t4 D_FlipFlop_3.3-input-nand_1.Vout VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X779 Comparator_0.Vinm CDAC8_0.switch_7.Z.t68 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X780 a_74193_52572# Nand_Gate_0.A.t14 a_73579_52572# GND.t638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X781 a_63767_15797# RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout GND.t391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X782 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_3.3-input-nand_2.C.t5 VDD.t614 VDD.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X783 VDD.t219 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 VDD.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X784 Nand_Gate_5.A.t2 RingCounter_0.D_FlipFlop_7.Qbar a_113359_52572# GND.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X785 a_68455_15797# Nand_Gate_7.B.t10 a_67841_15797# GND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X786 a_132311_39721# D_FlipFlop_2.3-input-nand_2.C.t7 D_FlipFlop_2.3-input-nand_2.Vout.t0 GND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X787 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 a_100347_49858# GND.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X788 a_130209_40571# D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X789 VDD.t62 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X790 RingCounter_0.D_FlipFlop_6.Qbar Nand_Gate_5.B.t7 VDD.t648 VDD.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X791 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B VDD.t876 VDD.t800 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X792 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 VDD.t551 VDD.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X793 VDD.t866 D_FlipFlop_7.D.t17 D_FlipFlop_2.3-input-nand_1.B VDD.t865 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X794 VDD.t989 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout VDD.t988 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X795 a_107313_49858# RingCounter_0.D_FlipFlop_7.3-input-nand_1.B a_106699_49858# GND.t433 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X796 VDD.t559 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X797 a_123655_15797# Nand_Gate_5.B.t8 a_123041_15797# GND.t654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X798 VDD.t477 EN.t61 D_FlipFlop_1.Qbar VDD.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X799 GND.t320 D_FlipFlop_0.3-input-nand_2.C.t5 a_130209_44135# GND.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X800 a_78267_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 GND.t788 GND.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X801 a_132311_23350# D_FlipFlop_6.3-input-nand_2.C.t6 D_FlipFlop_6.3-input-nand_2.Vout.t0 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X802 And_Gate_7.Nand_Gate_0.Vout CLK.t49 a_125845_47663# GND.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X803 And_Gate_5.A.t1 Nand_Gate_3.B.t8 a_48937_47663# GND.t795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X804 GND.t396 Nand_Gate_5.A.t10 a_134897_44135# GND.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X805 a_65869_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 GND.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X806 a_116995_13083# Nand_Gate_1.B.t13 RingCounter_0.D_FlipFlop_10.Qbar GND.t359 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X807 VDD.t929 D_FlipFlop_4.3-input-nand_2.Vout.t7 D_FlipFlop_4.3-input-nand_2.C.t3 VDD.t769 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X808 VDD.t868 D_FlipFlop_7.D.t18 D_FlipFlop_6.3-input-nand_1.B VDD.t867 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X809 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 VDD.t227 VDD.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X810 a_90665_49858# VDD.t1135 GND.t157 GND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X811 a_132925_39721# D_FlipFlop_2.3-input-nand_0.Vout a_132311_39721# GND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X812 VDD.t592 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X813 VDD.t16 FFCLR.t30 D_FlipFlop_4.3-input-nand_2.C.t1 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X814 a_117739_52572# VDD.t1136 GND.t159 GND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X815 Nand_Gate_6.Vout.t2 Nand_Gate_6.B.t8 VDD.t792 VDD.t791 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X816 VDD.t809 Q6.t6 D_FlipFlop_2.Qbar VDD.t808 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X817 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B Nand_Gate_5.A.t11 VDD.t575 VDD.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X818 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.3-input-nand_1.B VDD.t852 VDD.t603 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X819 RingCounter_0.D_FlipFlop_4.Qbar Nand_Gate_2.A.t8 a_91279_49858# GND.t724 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X820 VDD.t715 VDD.t714 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 VDD.t441 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X821 GND.t785 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 a_107927_15797# GND.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X822 GND.t385 FFCLR.t31 a_128851_37007# GND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X823 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 CLK.t50 a_107313_49858# GND.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X824 a_121069_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 GND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X825 GND.t740 D_FlipFlop_7.D.t19 D_FlipFlop_1.3-input-nand_1.B GND.t739 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X826 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B Nand_Gate_0.B.t6 GND.t24 GND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X827 Comparator_0.Vinm CDAC8_0.switch_7.Z.t67 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X828 GND.t679 Q4.t8 CDAC8_0.switch_8.Z.t3 VDD.t784 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X829 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 VDD.t107 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X830 VDD.t713 VDD.t712 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X831 a_132925_23350# D_FlipFlop_6.3-input-nand_0.Vout a_132311_23350# GND.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X832 Comparator_0.Vinm CDAC8_0.switch_7.Z.t66 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X833 GND.t742 D_FlipFlop_7.D.t20 D_FlipFlop_0.3-input-nand_1.B GND.t741 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X834 VDD.t78 Nand_Gate_5.Vout.t3 And_Gate_7.Nand_Gate_0.Vout VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X835 VDD.t282 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X836 Comparator_0.Vinm CDAC8_0.switch_7.Z.t65 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X837 a_75551_49858# VDD.t1137 GND.t161 GND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X838 Comparator_0.Vinm CDAC8_0.switch_7.Z.t64 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X839 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK.t51 VDD.t1061 VDD.t1060 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X840 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 CLK.t52 VDD.t1059 VDD.t1058 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X841 a_30647_15797# RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout GND.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X842 VDD.t201 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X843 D_FlipFlop_2.Qbar D_FlipFlop_2.Nand_Gate_1.Vout VDD.t319 VDD.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X844 a_35335_15797# Nand_Gate_4.A.t5 a_34721_15797# GND.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X845 a_89921_13083# CLK.t53 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 GND.t381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X846 Comparator_0.Vinm CDAC8_0.switch_6.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X847 GND.t436 D_FlipFlop_7.D.t21 D_FlipFlop_4.3-input-nand_1.B GND.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X848 GND.t332 And_Gate_5.Vout.t4 D_FlipFlop_1.Inverter_1.Vout GND.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X849 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B VDD.t935 VDD.t934 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X850 a_128237_43285# D_FlipFlop_3.Qbar Q5.t2 GND.t375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X851 Comparator_0.Vinm CDAC8_0.switch_7.Z.t63 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X852 Comparator_0.Vinm CDAC8_0.switch_8.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X853 Comparator_0.Vinm CDAC8_0.switch_9.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X854 D_FlipFlop_4.3-input-nand_2.Vout.t0 D_FlipFlop_4.3-input-nand_0.Vout VDD.t392 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X855 Comparator_0.Vinm CDAC8_0.switch_6.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X856 And_Gate_0.Nand_Gate_0.Vout And_Gate_0.B.t3 VDD.t421 VDD.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X857 a_76165_49858# RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 a_75551_49858# GND.t685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X858 Comparator_0.Vinm CDAC8_0.switch_6.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X859 a_45147_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 GND.t860 GND.t859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X860 VDD.t915 And_Gate_1.Vout.t5 D_FlipFlop_7.3-input-nand_1.Vout VDD.t911 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X861 a_32749_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 GND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X862 D_FlipFlop_7.Nand_Gate_1.Vout D_FlipFlop_7.3-input-nand_2.C.t5 VDD.t223 VDD.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X863 a_95529_13083# RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 a_94915_13083# GND.t745 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X864 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B VDD.t397 VDD.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X865 VDD.t797 Nand_Gate_6.A.t8 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B VDD.t796 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X866 VDD.t38 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 FFCLR.t0 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X867 Comparator_0.Vinm CDAC8_0.switch_8.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X868 VDD.t1104 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 VDD.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X869 VDD.t50 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X870 a_128851_24200# D_FlipFlop_5.Nand_Gate_1.Vout a_128237_24200# GND.t725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X871 Comparator_0.Vinm CDAC8_0.switch_6.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X872 VDD.t711 VDD.t710 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 VDD.t437 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X873 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B FFCLR.t32 GND.t387 GND.t386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X874 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_7.D.t22 VDD.t394 VDD.t393 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X875 Comparator_0.Vinm CDAC8_0.switch_6.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X876 a_130209_26914# D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout GND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X877 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t708 VDD.t709 VDD.t516 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X878 Comparator_0.Vinm CDAC8_0.switch_7.Z.t62 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X879 VDD.t844 Nand_Gate_2.A.t9 Q5.t1 VDD.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X880 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_7.D.t23 VDD.t395 VDD.t333 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X881 a_42431_49858# EN.t62 GND.t522 GND.t521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X882 GND.t163 VDD.t1138 a_95529_13083# GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X883 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK.t54 VDD.t1057 VDD.t1056 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X884 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 CLK.t55 VDD.t1055 VDD.t1054 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X885 VDD.t340 FFCLR.t33 D_FlipFlop_0.Qbar VDD.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X886 a_39715_15797# RingCounter_0.D_FlipFlop_8.Qbar Nand_Gate_4.A.t2 GND.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X887 a_134283_33443# And_Gate_5.Vout.t5 D_FlipFlop_1.3-input-nand_1.Vout GND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X888 a_56801_13083# CLK.t56 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 GND.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X889 VDD.t229 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X890 Comparator_0.Vinm CDAC8_0.switch_6.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X891 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 CLK.t57 VDD.t1053 VDD.t1052 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X892 VDD.t342 FFCLR.t34 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X893 a_102319_49858# RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 a_101705_49858# GND.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X894 VDD.t765 Nand_Gate_7.B.t11 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B VDD.t764 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X895 Comparator_0.Vinm CDAC8_0.switch_7.Z.t61 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X896 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 VDD.t829 VDD.t827 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X897 Comparator_0.Vinm CDAC8_0.switch_8.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X898 Comparator_0.Vinm CDAC8_0.switch_9.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X899 And_Gate_1.B.t1 Nand_Gate_4.B.t10 VDD.t969 VDD.t968 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X900 a_43045_49858# RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_42431_49858# GND.t732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X901 a_132311_36157# D_FlipFlop_1.3-input-nand_2.C.t6 D_FlipFlop_1.3-input-nand_2.Vout.t1 GND.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X902 RingCounter_0.D_FlipFlop_17.Qbar FFCLR.t35 a_47119_49858# GND.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X903 a_112001_13083# CLK.t58 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 GND.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X904 a_128851_20636# D_FlipFlop_6.Nand_Gate_1.Vout a_128237_20636# GND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X905 Comparator_0.Vinm CDAC8_0.switch_7.Z.t60 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X906 VDD.t775 Nand_Gate_1.A.t6 RingCounter_0.D_FlipFlop_9.Qbar VDD.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X907 And_Gate_5.Vout.t0 And_Gate_5.Nand_Gate_0.Vout VDD.t847 VDD.t846 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X908 a_62409_13083# RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 a_61795_13083# GND.t769 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X909 a_79625_52572# EN.t63 GND.t520 GND.t519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X910 a_132311_46849# D_FlipFlop_0.3-input-nand_2.C.t6 D_FlipFlop_0.3-input-nand_2.Vout.t2 GND.t861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X911 VDD.t650 Nand_Gate_5.B.t9 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B VDD.t649 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X912 VDD.t1051 CLK.t59 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 VDD.t1050 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X913 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 VDD.t331 VDD.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X914 Comparator_0.Vinm CDAC8_0.switch_8.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X915 a_128237_19786# D_FlipFlop_7.Qbar Q0.t2 GND.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X916 a_58159_52572# RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_57545_52572# GND.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X917 RingCounter_0.D_FlipFlop_5.Qbar Nand_Gate_2.B.t10 a_102319_49858# GND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X918 VDD.t833 And_Gate_0.Vout.t6 D_FlipFlop_6.Inverter_1.Vout VDD.t832 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X919 VDD.t576 Nand_Gate_5.A.t12 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X920 Comparator_0.Vinm CDAC8_0.switch_7.Z.t59 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X921 Comparator_0.Vinm CDAC8_0.switch_6.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X922 a_132311_30478# D_FlipFlop_4.3-input-nand_2.C.t5 D_FlipFlop_4.3-input-nand_2.Vout.t3 GND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X923 a_132925_36157# D_FlipFlop_1.3-input-nand_0.Vout a_132311_36157# GND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X924 GND.t595 D_FlipFlop_0.CLK.t4 D_FlipFlop_0.Inverter_1.Vout GND.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X925 VDD.t110 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_2.Qbar VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X926 Comparator_0.Vinm CDAC8_0.switch_6.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X927 VDD.t269 Q7.t6 D_FlipFlop_1.Qbar VDD.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X928 a_66483_13083# RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 a_65869_13083# GND.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X929 GND.t165 VDD.t1139 a_62409_13083# GND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X930 a_132925_46849# D_FlipFlop_0.3-input-nand_0.Vout a_132311_46849# GND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X931 Nand_Gate_6.B.t1 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t542 VDD.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X932 a_67841_15797# CLK.t60 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 GND.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X933 a_37897_16975# Nand_Gate_4.A.t6 GND.t290 GND.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X934 a_114805_16975# CLK.t61 GND.t325 GND.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X935 VDD.t8 And_Gate_3.Vout.t6 D_FlipFlop_4.3-input-nand_1.Vout VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X936 a_67227_49858# RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 GND.t309 GND.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X937 VDD.t904 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 VDD.t835 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X938 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_4.3-input-nand_2.C.t6 VDD.t772 VDD.t771 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X939 a_130209_17072# D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X940 a_134897_39721# D_FlipFlop_7.D.t24 a_134283_39721# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X941 a_119711_52572# EN.t64 GND.t518 GND.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X942 VDD.t1049 CLK.t62 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 VDD.t1048 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X943 a_121683_13083# RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 a_121069_13083# GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X944 a_132925_30478# D_FlipFlop_4.3-input-nand_0.Vout a_132311_30478# GND.t434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X945 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 CLK.t63 VDD.t1047 VDD.t1002 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X946 a_130209_27764# D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout GND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X947 VDD.t817 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_0.Vout VDD.t815 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X948 a_106699_49858# EN.t65 GND.t516 GND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X949 Comparator_0.Vinm CDAC8_0.switch_6.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X950 VDD.t897 RingCounter_0.D_FlipFlop_11.Qbar Nand_Gate_6.B.t3 VDD.t788 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X951 VDD.t942 Nand_Gate_4.A.t7 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B VDD.t941 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X952 VDD.t970 Nand_Gate_4.B.t11 Q0.t1 VDD.t639 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X953 D_FlipFlop_1.Qbar D_FlipFlop_1.Nand_Gate_1.Vout VDD.t361 VDD.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X954 Comparator_0.Vinm CDAC8_0.switch_6.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X955 a_123041_15797# CLK.t64 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 GND.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X956 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK.t65 a_85233_52572# GND.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X957 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 VDD.t300 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X958 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 EN.t66 VDD.t476 VDD.t475 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X959 VDD.t474 EN.t67 Nand_Gate_6.B.t0 VDD.t473 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X960 a_73449_15797# RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_72835_15797# GND.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X961 a_134897_23350# D_FlipFlop_7.D.t25 a_134283_23350# GND.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X962 Comparator_0.Vinm CDAC8_0.switch_7.Z.t58 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X963 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 CLK.t66 GND.t329 GND.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X964 Comparator_0.Vinm CDAC8_0.switch_7.Z.t57 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X965 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 VDD.t585 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X966 a_46505_52572# VDD.t1140 GND.t167 GND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X967 a_106569_13083# RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 a_105955_13083# GND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X968 Comparator_0.Vinm CDAC8_0.switch_9.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X969 Comparator_0.Vinm CDAC8_0.switch_7.Z.t56 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X970 RingCounter_0.D_FlipFlop_12.Qbar RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 VDD.t899 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X971 VDD.t799 Nand_Gate_6.A.t9 Nand_Gate_6.Vout.t0 VDD.t798 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X972 Comparator_0.Vinm CDAC8_0.switch_7.Z.t55 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X973 GND.t841 CLK.t67 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 GND.t840 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X974 a_128851_37007# D_FlipFlop_2.Nand_Gate_1.Vout a_128237_37007# GND.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X975 GND.t716 Nand_Gate_2.A.t10 a_132925_43285# GND.t427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X976 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 VDD.t1105 VDD.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X977 RingCounter_0.D_FlipFlop_1.Qbar VDD.t704 VDD.t705 VDD.t435 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X978 a_134283_44135# D_FlipFlop_0.CLK.t5 D_FlipFlop_0.3-input-nand_1.Vout GND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X979 CDAC8_0.switch_8.Z.t0 a_75898_46095# VDD.t207 VDD.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X980 VDD.t999 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X981 VDD.t274 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X982 a_101705_52572# EN.t68 GND.t512 GND.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X983 GND.t514 EN.t69 a_73449_15797# GND.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X984 a_33363_13083# RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 a_32749_13083# GND.t759 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X985 GND.t510 EN.t70 a_90535_13083# GND.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X986 Comparator_0.Vinm CDAC8_0.switch_7.Z.t54 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X987 GND.t169 VDD.t1141 a_106569_13083# GND.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X988 RingCounter_0.D_FlipFlop_7.Qbar VDD.t706 VDD.t707 VDD.t433 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X989 VDD.t703 VDD.t702 RingCounter_0.D_FlipFlop_12.Qbar VDD.t532 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X990 Comparator_0.Vinm CDAC8_0.switch_1.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X991 a_34721_15797# CLK.t68 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout GND.t842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X992 GND.t282 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 a_96887_13083# GND.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X993 And_Gate_2.Nand_Gate_0.Vout Nand_Gate_6.Vout.t4 a_92725_16975# GND.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X994 VDD.t793 Nand_Gate_6.B.t9 D_FlipFlop_5.3-input-nand_1.Vout VDD.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X995 VDD.t1046 CLK.t69 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 VDD.t1045 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X996 GND.t639 Nand_Gate_0.A.t15 a_128851_39721# GND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X997 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK.t70 VDD.t1044 VDD.t1000 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X998 VDD.t900 RingCounter_0.D_FlipFlop_14.Qbar Nand_Gate_7.A.t2 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X999 a_59605_47663# And_Gate_5.A.t3 GND.t334 GND.t333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1000 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK.t71 a_52113_52572# GND.t843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1001 GND.t171 VDD.t1142 a_33363_13083# GND.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1002 Comparator_0.Vinm CDAC8_0.switch_6.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1003 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 VDD.t32 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1004 a_80239_49858# RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 a_79625_49858# GND.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1005 a_96887_13083# RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 GND.t808 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1006 VDD.t560 D_FlipFlop_3.Qbar Q5.t3 VDD.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1007 Comparator_0.Vinm CDAC8_0.switch_7.Z.t53 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1008 Comparator_0.Vinm CDAC8_0.switch_6.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1009 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 EN.t71 VDD.t472 VDD.t471 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1010 VDD.t470 EN.t72 Nand_Gate_7.A.t0 VDD.t469 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1011 a_40329_15797# RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_39715_15797# GND.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1012 VDD.t1043 CLK.t72 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 VDD.t1042 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1013 Comparator_0.Vinm CDAC8_0.switch_7.Z.t52 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1014 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 CLK.t73 GND.t845 GND.t844 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1015 VDD.t785 Q4.t9 D_FlipFlop_0.Qbar VDD.t362 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1016 GND.t663 Nand_Gate_7.B.t12 a_128851_23350# GND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1017 VDD.t1041 CLK.t74 And_Gate_2.Nand_Gate_0.Vout VDD.t1040 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1018 RingCounter_0.D_FlipFlop_15.Qbar RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 VDD.t100 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1019 Comparator_0.Vinm CDAC8_0.switch_7.Z.t51 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1020 a_111387_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 GND.t257 GND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1021 Comparator_0.Vinm CDAC8_0.switch_9.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1022 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 VDD.t571 VDD.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1023 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 a_98245_52572# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1024 VDD.t432 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_5.A.t0 VDD.t431 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1025 Q5.t0 D_FlipFlop_3.Nand_Gate_0.Vout VDD.t64 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1026 VDD.t188 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1027 GND.t508 EN.t73 a_40329_15797# GND.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1028 Comparator_0.Vinm CDAC8_0.switch_7.Z.t50 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1029 Comparator_0.Vinm CDAC8_0.switch_7.Z.t49 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1030 VDD.t701 VDD.t700 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 VDD.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1031 Comparator_0.Vinm CDAC8_0.switch_6.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1032 Nand_Gate_3.B.t1 RingCounter_0.D_FlipFlop_1.Qbar VDD.t142 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1033 VDD.t895 Nand_Gate_1.B.t14 Q3.t1 VDD.t644 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1034 D_FlipFlop_0.Qbar D_FlipFlop_0.Nand_Gate_1.Vout VDD.t336 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1035 VDD.t699 VDD.t698 RingCounter_0.D_FlipFlop_15.Qbar VDD.t524 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1036 Nand_Gate_1.A.t3 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t818 VDD.t634 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1037 GND.t506 EN.t74 a_121683_15797# GND.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1038 Comparator_0.Vinm CDAC8_0.switch_7.Z.t48 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1039 VDD.t195 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_4.Qbar VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1040 VDD.t391 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1041 GND.t854 Nand_Gate_4.B.t12 a_132925_19786# GND.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1042 a_128237_40571# Q5.t8 D_FlipFlop_3.Qbar GND.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1043 Nand_Gate_5.A.t3 RingCounter_0.D_FlipFlop_7.Qbar VDD.t930 VDD.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1044 VDD.t637 D_FlipFlop_6.3-input-nand_2.Vout.t7 D_FlipFlop_6.3-input-nand_2.C.t3 VDD.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1045 D_FlipFlop_5.3-input-nand_2.Vout.t2 D_FlipFlop_5.3-input-nand_0.Vout VDD.t568 VDD.t567 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1046 And_Gate_4.Vout.t1 And_Gate_4.Nand_Gate_0.Vout GND.t202 GND.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1047 VDD.t987 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD.t944 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1048 Nand_Gate_0.B.t0 RingCounter_0.D_FlipFlop_3.Qbar a_80239_52572# GND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1049 VDD.t940 Nand_Gate_4.A.t8 And_Gate_1.B.t2 VDD.t939 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1050 VDD.t343 FFCLR.t36 D_FlipFlop_6.3-input-nand_2.C.t1 VDD.t239 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1051 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t52 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1052 a_47119_49858# RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_46505_49858# GND.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1053 VDD.t697 VDD.t696 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 VDD.t508 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1054 a_63767_13083# RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 GND.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1055 a_134897_36157# D_FlipFlop_7.D.t26 a_134283_36157# GND.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1056 VDD.t468 EN.t75 Nand_Gate_1.A.t0 VDD.t467 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1057 RingCounter_0.D_FlipFlop_4.Qbar Nand_Gate_2.A.t11 VDD.t837 VDD.t312 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1058 a_68455_13083# RingCounter_0.D_FlipFlop_14.3-input-nand_1.B a_67841_13083# GND.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1059 Comparator_0.Vinm CDAC8_0.switch_7.Z.t47 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1060 VDD.t906 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 VDD.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1061 VDD.t695 VDD.t694 RingCounter_0.D_FlipFlop_10.Qbar VDD.t522 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1062 a_134897_46849# D_FlipFlop_7.D.t27 a_134283_46849# GND.t439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1063 Comparator_0.Vinm CDAC8_0.switch_7.Z.t46 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1064 GND.t665 Nand_Gate_7.B.t13 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B GND.t664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1065 VDD.t367 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 VDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1066 VDD.t767 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1067 a_90535_15797# Nand_Gate_6.B.t10 a_89921_15797# GND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1068 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 a_65125_52572# GND.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1069 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B Nand_Gate_5.A.t13 GND.t613 GND.t612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1070 VDD.t1039 CLK.t75 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 VDD.t1038 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1071 D_FlipFlop_2.3-input-nand_2.Vout.t3 D_FlipFlop_2.3-input-nand_0.Vout VDD.t824 VDD.t429 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1072 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t692 VDD.t693 VDD.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1073 a_123655_13083# RingCounter_0.D_FlipFlop_10.3-input-nand_1.B a_123041_13083# GND.t611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1074 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 VDD.t908 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1075 a_134897_30478# D_FlipFlop_7.D.t28 a_134283_30478# GND.t648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1076 VDD.t874 D_FlipFlop_7.Qbar Q0.t3 VDD.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1077 a_84619_52572# VDD.t1143 GND.t173 GND.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1078 a_65869_13083# RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 GND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1079 Comparator_0.Vinm CDAC8_0.switch_9.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1080 GND.t656 Nand_Gate_5.B.t10 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B GND.t655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1081 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B Nand_Gate_0.B.t7 VDD.t24 VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1082 Comparator_0.Vinm CDAC8_0.switch_7.Z.t45 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1083 Comparator_0.Vinm CDAC8_0.switch_7.Z.t44 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1084 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 a_120325_52572# GND.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1085 Comparator_0.Vinm CDAC8_0.switch_9.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1086 And_Gate_4.A.t0 Nand_Gate_0.B.t8 a_71017_47663# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1087 GND.t630 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 a_74807_15797# GND.t629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1088 Comparator_0.Vinm CDAC8_0.switch_6.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1089 D_FlipFlop_6.3-input-nand_2.Vout.t2 D_FlipFlop_6.3-input-nand_0.Vout VDD.t823 VDD.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1090 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 CLK.t76 a_74193_49858# GND.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1091 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 EN.t76 VDD.t466 VDD.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1092 GND.t602 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 a_107927_13083# GND.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1093 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 VDD.t589 VDD.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1094 VDD.t691 VDD.t690 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 VDD.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1095 a_121069_13083# RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 GND.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1096 GND.t597 D_FlipFlop_3.3-input-nand_2.Vout.t7 a_130209_43285# GND.t319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1097 Comparator_0.Vinm CDAC8_0.switch_6.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1098 Comparator_0.Vinm CDAC8_0.switch_8.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1099 GND.t390 FFCLR.t37 a_134897_43285# GND.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1100 Q0.t0 D_FlipFlop_7.Nand_Gate_0.Vout VDD.t653 VDD.t652 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1101 a_85233_52572# Nand_Gate_0.B.t9 a_84619_52572# GND.t692 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1102 Comparator_0.Vinm CDAC8_0.switch_0.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1103 VDD.t1037 CLK.t77 And_Gate_1.Nand_Gate_0.Vout VDD.t1036 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1104 a_132311_33443# D_FlipFlop_1.3-input-nand_2.Vout.t6 D_FlipFlop_1.3-input-nand_2.C.t1 GND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1105 VDD.t779 D_FlipFlop_1.3-input-nand_2.C.t7 D_FlipFlop_1.3-input-nand_2.Vout.t2 VDD.t778 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1106 Comparator_0.Vinm CDAC8_0.switch_8.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1107 VDD.t255 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 VDD.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1108 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 a_89307_52572# GND.t586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1109 VDD.t624 Nand_Gate_0.A.t16 D_FlipFlop_2.3-input-nand_1.Vout VDD.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1110 a_30647_13083# RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 GND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1111 Comparator_0.Vinm CDAC8_0.switch_6.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1112 VDD.t880 FFCLR.t38 D_FlipFlop_1.3-input-nand_2.Vout.t3 VDD.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1113 VDD.t975 D_FlipFlop_0.3-input-nand_2.C.t7 D_FlipFlop_0.3-input-nand_2.Vout.t3 VDD.t233 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1114 Comparator_0.Vinm CDAC8_0.switch_6.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1115 a_35335_13083# RingCounter_0.D_FlipFlop_16.3-input-nand_1.B a_34721_13083# GND.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1116 GND.t761 FFCLR.t39 a_128851_36157# GND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1117 VDD.t577 Nand_Gate_5.A.t14 D_FlipFlop_0.3-input-nand_2.Vout.t1 VDD.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1118 a_118353_49858# RingCounter_0.D_FlipFlop_6.3-input-nand_1.B a_117739_49858# GND.t345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1119 a_94915_15797# RingCounter_0.D_FlipFlop_11.Qbar Nand_Gate_6.B.t2 GND.t773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1120 GND.t92 Nand_Gate_4.A.t9 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B GND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1121 VDD.t198 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1122 GND.t615 Nand_Gate_5.A.t15 a_128851_46849# GND.t614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1123 Comparator_0.Vinm CDAC8_0.switch_7.Z.t43 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1124 a_99603_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 a_98989_15797# GND.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1125 VDD.t1035 CLK.t78 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 VDD.t1034 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1126 a_132925_33443# D_FlipFlop_1.3-input-nand_1.Vout a_132311_33443# GND.t434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1127 a_128237_26914# D_FlipFlop_5.Qbar Q2.t1 GND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1128 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 VDD.t974 VDD.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1129 a_51499_52572# VDD.t1144 GND.t175 GND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1130 a_32749_13083# RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 GND.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1131 GND.t771 Nand_Gate_1.B.t15 a_128851_30478# GND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1132 VDD.t898 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 VDD.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1133 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B FFCLR.t40 VDD.t882 VDD.t881 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1134 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 Nand_Gate_7.B.t14 VDD.t68 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1135 GND.t667 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 a_118967_15797# GND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1136 GND.t445 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 a_41687_15797# GND.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1137 VDD.t689 VDD.t688 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 VDD.t518 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1138 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 CLK.t79 a_118353_49858# GND.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1139 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 EN.t77 VDD.t464 VDD.t463 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1140 VDD.t146 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 VDD.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1141 GND.t504 EN.t78 a_99603_15797# GND.t503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1142 Comparator_0.Vinm CDAC8_0.switch_7.Z.t42 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1143 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 VDD.t588 VDD.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1144 VDD.t687 VDD.t686 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 VDD.t502 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1145 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.3-input-nand_1.B VDD.t875 VDD.t599 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1146 And_Gate_0.Vout.t0 And_Gate_0.Nand_Gate_0.Vout VDD.t190 VDD.t189 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1147 a_128851_39721# D_FlipFlop_2.Nand_Gate_0.Vout a_128237_39721# GND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1148 a_130209_24200# D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout GND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1149 VDD.t158 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1150 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK.t80 VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1151 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 Nand_Gate_5.B.t11 VDD.t651 VDD.t572 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1152 a_100347_49858# RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 GND.t34 GND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1153 Comparator_0.Vinm CDAC8_0.switch_6.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1154 a_52113_52572# FFCLR.t41 a_51499_52572# GND.t762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1155 a_41687_15797# RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1156 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 a_87205_49858# GND.t688 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1157 VDD.t617 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 VDD.t386 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1158 a_75898_21528# Q1.t5 GND.t778 GND.t777 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1159 VDD.t291 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 VDD.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1160 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 a_56187_52572# GND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1161 a_46375_15797# Nand_Gate_4.B.t13 a_45761_15797# GND.t855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1162 Comparator_0.Vinm CDAC8_0.switch_7.Z.t41 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1163 Comparator_0.Vinm CDAC8_0.switch_8.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1164 VDD.t685 VDD.t684 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 VDD.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1165 VDD.t980 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 VDD.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1166 a_39715_13083# Nand_Gate_4.A.t10 RingCounter_0.D_FlipFlop_8.Qbar GND.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1167 VDD.t1107 D_FlipFlop_4.Qbar Q3.t3 VDD.t994 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1168 VDD.t462 EN.t79 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 VDD.t461 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1169 a_128851_23350# D_FlipFlop_6.Nand_Gate_0.Vout a_128237_23350# GND.t725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1170 Comparator_0.Vinm CDAC8_0.switch_6.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1171 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B VDD.t230 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1172 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 VDD.t554 VDD.t552 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1173 GND.t763 FFCLR.t42 a_132925_40571# GND.t749 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1174 Comparator_0.Vinm CDAC8_0.switch_6.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1175 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 VDD.t907 VDD.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1176 Comparator_0.Vinm CDAC8_0.switch_7.Z.t40 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1177 GND.t341 D_FlipFlop_7.3-input-nand_2.Vout.t7 a_130209_19786# GND.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1178 VDD.t36 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1179 a_61795_15797# RingCounter_0.D_FlipFlop_14.Qbar Nand_Gate_7.A.t1 GND.t776 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1180 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B RingCounter_0.D_FlipFlop_16.Q.t7 VDD.t889 VDD.t888 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1181 VDD.t612 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1182 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 a_111387_52572# GND.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1183 a_101575_15797# Nand_Gate_1.A.t7 a_100961_15797# GND.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1184 Nand_Gate_0.B.t3 EN.t80 VDD.t460 VDD.t459 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1185 a_56187_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 GND.t871 GND.t870 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1186 GND.t764 FFCLR.t43 a_134897_19786# GND.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1187 VDD.t347 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout VDD.t346 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1188 And_Gate_6.Nand_Gate_0.Vout CLK.t81 a_103765_47663# GND.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1189 VDD.t70 Nand_Gate_7.B.t15 RingCounter_0.D_FlipFlop_13.Qbar VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1190 VDD.t834 And_Gate_0.Vout.t7 D_FlipFlop_6.3-input-nand_1.Vout VDD.t830 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1191 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B VDD.t984 VDD.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1192 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 VDD.t382 VDD.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1193 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 VDD.t1102 VDD.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1194 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_6.3-input-nand_2.C.t7 VDD.t581 VDD.t580 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1195 GND.t296 CLK.t82 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 GND.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1196 Comparator_0.Vinm CDAC8_0.switch_0.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1197 VDD.t26 Nand_Gate_6.B.t11 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1198 VDD.t424 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout Nand_Gate_3.B.t2 VDD.t263 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1199 Q3.t0 D_FlipFlop_4.Nand_Gate_0.Vout VDD.t299 VDD.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1200 And_Gate_0.B.t1 Nand_Gate_7.B.t16 VDD.t72 VDD.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1201 a_132311_44135# D_FlipFlop_0.3-input-nand_2.Vout.t6 D_FlipFlop_0.3-input-nand_2.C.t1 GND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1202 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout Nand_Gate_4.A.t11 VDD.t938 VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1203 a_130209_20636# D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1204 VDD.t406 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout VDD.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1205 D_FlipFlop_3.3-input-nand_2.C.t3 D_FlipFlop_3.3-input-nand_1.Vout VDD.t853 VDD.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1206 VDD.t683 VDD.t682 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 VDD.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1207 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 EN.t81 VDD.t458 VDD.t457 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1208 VDD.t804 Nand_Gate_0.B.t10 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1209 a_128237_17072# Q0.t6 D_FlipFlop_7.Qbar GND.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1210 Comparator_0.Vinm CDAC8_0.switch_7.Z.t39 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1211 GND.t478 EN.t82 a_66483_15797# GND.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1212 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 CLK.t83 VDD.t1031 VDD.t1030 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1213 Comparator_0.Vinm CDAC8_0.switch_9.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1214 VDD.t958 Nand_Gate_2.Vout.t4 And_Gate_6.Nand_Gate_0.Vout VDD.t957 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1215 Comparator_0.Vinm CDAC8_0.switch_7.Z.t38 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1216 Comparator_0.Vinm CDAC8_0.switch_7.Z.t37 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1217 a_128237_27764# Q3.t8 D_FlipFlop_4.Qbar GND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1218 a_53471_49858# VDD.t1145 GND.t177 GND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1219 Comparator_0.Vinm CDAC8_0.switch_9.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1220 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK.t84 VDD.t1029 VDD.t1028 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1221 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 a_54085_49858# GND.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1222 VDD.t283 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 VDD.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1223 a_132925_44135# D_FlipFlop_0.3-input-nand_1.Vout a_132311_44135# GND.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1224 a_86591_52572# EN.t83 GND.t480 GND.t479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1225 a_67841_13083# CLK.t85 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 GND.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1226 Nand_Gate_2.Vout.t2 Nand_Gate_2.B.t11 VDD.t922 VDD.t921 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1227 VDD.t402 a_138533_35417.t3 D_FlipFlop_7.D.t1 VDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=17.4 pd=120.58 as=17.4 ps=120.58 w=60 l=1
X1228 a_113359_49858# RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 a_112745_49858# GND.t730 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1229 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 VDD.t680 VDD.t681 VDD.t520 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1230 VDD.t883 FFCLR.t44 D_FlipFlop_1.3-input-nand_1.Vout VDD.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1231 a_105955_15797# RingCounter_0.D_FlipFlop_9.Qbar Nand_Gate_1.A.t1 GND.t585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1232 a_54085_49858# RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 a_53471_49858# GND.t712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1233 RingCounter_0.D_FlipFlop_1.Qbar Nand_Gate_3.B.t9 a_58159_49858# GND.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1234 a_123041_13083# CLK.t86 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 GND.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1235 VDD.t896 Nand_Gate_1.B.t16 RingCounter_0.D_FlipFlop_10.Qbar VDD.t546 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1236 a_73449_13083# RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 a_72835_13083# GND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1237 a_87205_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_86591_52572# GND.t321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1238 VDD.t102 And_Gate_5.Vout.t6 D_FlipFlop_1.3-input-nand_0.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1239 VDD.t28 Nand_Gate_6.B.t12 Q2.t3 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1240 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.3-input-nand_2.Vout.t7 VDD.t192 VDD.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1241 Comparator_0.Vinm CDAC8_0.switch_2.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1242 a_74193_49858# RingCounter_0.D_FlipFlop_3.3-input-nand_1.B a_73579_49858# GND.t767 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1243 Comparator_0.Vinm CDAC8_0.switch_7.Z.t36 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1244 RingCounter_0.D_FlipFlop_7.Qbar Nand_Gate_5.A.t16 a_113359_49858# GND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1245 VDD.t557 D_FlipFlop_0.CLK.t6 D_FlipFlop_0.3-input-nand_0.Vout VDD.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1246 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.3-input-nand_2.Vout.t7 VDD.t205 VDD.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1247 VDD.t616 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1248 a_93097_47663# Nand_Gate_2.A.t12 GND.t718 GND.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1249 a_130209_37007# D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout GND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1250 VDD.t926 And_Gate_2.Vout.t5 D_FlipFlop_5.Inverter_1.Vout VDD.t925 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1251 GND.t28 Nand_Gate_6.B.t13 a_132925_26914# GND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1252 And_Gate_1.Nand_Gate_0.Vout And_Gate_1.B.t4 a_48565_16975# GND.t838 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1253 And_Gate_4.Nand_Gate_0.Vout CLK.t87 VDD.t1027 VDD.t1026 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1254 GND.t179 VDD.t1146 a_73449_13083# GND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1255 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 CLK.t88 VDD.t1025 VDD.t1024 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1256 a_134897_33443# D_FlipFlop_1.3-input-nand_1.B a_134283_33443# GND.t648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1257 a_78881_15797# CLK.t89 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 GND.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1258 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.3-input-nand_1.B VDD.t631 VDD.t601 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1259 a_78267_49858# RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 GND.t184 GND.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1260 VDD.t625 Nand_Gate_0.A.t17 Q6.t0 VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1261 Comparator_0.Vinm CDAC8_0.switch_7.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1262 a_34721_13083# CLK.t90 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 GND.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1263 GND.t181 VDD.t1147 a_79495_15797# GND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1264 Comparator_0.Vinm CDAC8_0.switch_7.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1265 D_FlipFlop_7.3-input-nand_2.C.t0 D_FlipFlop_7.3-input-nand_1.Vout VDD.t113 VDD.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1266 a_128851_36157# D_FlipFlop_1.Nand_Gate_0.Vout a_128237_36157# GND.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1267 Comparator_0.Vinm CDAC8_0.switch_7.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1268 Comparator_0.Vinm CDAC8_0.switch_7.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1269 VDD.t890 RingCounter_0.D_FlipFlop_16.Q.t8 RingCounter_0.D_FlipFlop_16.Qbar VDD.t235 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1270 a_134283_43285# And_Gate_6.Vout.t5 D_FlipFlop_3.3-input-nand_0.Vout GND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1271 Comparator_0.Vinm CDAC8_0.switch_9.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1272 a_117739_49858# EN.t84 GND.t502 GND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1273 Comparator_0.Vinm CDAC8_0.switch_7.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1274 a_128851_46849# D_FlipFlop_0.Nand_Gate_0.Vout a_128237_46849# GND.t442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1275 a_104137_16975# Nand_Gate_1.A.t8 GND.t672 GND.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1276 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK.t91 a_96273_52572# GND.t301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1277 a_98989_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 GND.t673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1278 VDD.t74 Nand_Gate_7.B.t17 Q1.t1 VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1279 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 CLK.t92 GND.t303 GND.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1280 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 VDD.t315 VDD.t314 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1281 a_57545_52572# EN.t85 GND.t500 GND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1282 a_40329_13083# RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 a_39715_13083# GND.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1283 Comparator_0.Vinm CDAC8_0.switch_5.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1284 Comparator_0.Vinm CDAC8_0.switch_6.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1285 a_128851_30478# D_FlipFlop_4.Nand_Gate_0.Vout a_128237_30478# GND.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1286 Comparator_0.Vinm CDAC8_0.switch_7.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1287 VDD.t1023 CLK.t93 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 VDD.t1022 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1288 GND.t447 CLK.t94 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 GND.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1289 And_Gate_2.Vout.t1 And_Gate_2.Nand_Gate_0.Vout GND.t619 GND.t618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1290 RingCounter_0.D_FlipFlop_2.Qbar VDD.t678 VDD.t679 VDD.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1291 VDD.t61 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1292 VDD.t869 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1293 VDD.t254 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout Nand_Gate_0.B.t2 VDD.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1294 Comparator_0.Vinm CDAC8_0.switch_7.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1295 GND.t636 D_FlipFlop_3.3-input-nand_2.C.t6 a_130209_40571# GND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1296 VDD.t326 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 VDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1297 a_112745_52572# EN.t86 GND.t498 GND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1298 GND.t719 Nand_Gate_2.A.t13 a_134897_40571# GND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1299 VDD.t354 FFCLR.t45 D_FlipFlop_3.3-input-nand_0.Vout VDD.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1300 VDD.t1021 CLK.t95 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 VDD.t1020 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1301 a_75898_35820# Q7.t7 GND.t317 GND.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1302 GND.t814 VDD.t1148 a_40329_13083# GND.t813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1303 RingCounter_0.D_FlipFlop_6.Qbar VDD.t676 VDD.t677 VDD.t512 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1304 VDD.t79 Nand_Gate_5.A.t17 D_FlipFlop_0.3-input-nand_1.Vout VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1305 Nand_Gate_7.B.t3 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t628 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1306 VDD.t902 Q1.t6 CDAC8_0.switch_2.Z.t2 GND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1307 a_45761_15797# CLK.t96 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 GND.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1308 a_45147_49858# RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 GND.t371 GND.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1309 GND.t496 EN.t87 a_128851_33443# GND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1310 GND.t816 VDD.t1149 a_121683_13083# GND.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1311 GND.t818 VDD.t1150 a_46375_15797# GND.t817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1312 Nand_Gate_0.B.t1 RingCounter_0.D_FlipFlop_3.Qbar VDD.t47 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1313 VDD.t1019 CLK.t97 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 VDD.t1018 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1314 GND.t398 FFCLR.t46 a_132925_17072# GND.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1315 Comparator_0.Vinm CDAC8_0.switch_7.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1316 Comparator_0.Vinm CDAC8_0.switch_7.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1317 VDD.t849 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t848 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1318 Comparator_0.Vinm CDAC8_0.switch_7.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1319 Comparator_0.Vinm CDAC8_0.switch_9.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1320 VDD.t456 EN.t88 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 VDD.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1321 CDAC8_0.switch_2.Z.t1 a_75898_21528# GND.t606 GND.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1322 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 VDD.t674 VDD.t675 VDD.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1323 a_100961_15797# CLK.t98 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 GND.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1324 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK.t99 a_63153_52572# GND.t450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1325 GND.t399 FFCLR.t47 a_132925_27764# GND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1326 Nand_Gate_6.Vout.t1 Nand_Gate_6.B.t14 a_82057_16975# GND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1327 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 EN.t89 VDD.t454 VDD.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1328 a_51369_15797# RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_50755_15797# GND.t734 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1329 VDD.t452 EN.t90 Nand_Gate_7.B.t2 VDD.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1330 GND.t820 VDD.t1151 a_101575_15797# GND.t819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1331 VDD.t1017 CLK.t100 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 VDD.t1016 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1332 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 CLK.t101 GND.t452 GND.t451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1333 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 VDD.t148 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1334 Comparator_0.Vinm CDAC8_0.switch_6.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1335 RingCounter_0.D_FlipFlop_14.Qbar RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 VDD.t893 VDD.t892 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1336 Comparator_0.Vinm CDAC8_0.switch_6.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1337 a_125845_47663# Nand_Gate_5.Vout.t4 GND.t59 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1338 a_48937_47663# FFCLR.t48 GND.t401 GND.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1339 Comparator_0.Vinm CDAC8_0.switch_5.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1340 VDD.t1015 CLK.t102 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t1014 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1341 GND.t454 CLK.t103 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 GND.t453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1342 a_134283_19786# And_Gate_1.Vout.t6 D_FlipFlop_7.3-input-nand_0.Vout GND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1343 a_134897_44135# D_FlipFlop_0.3-input-nand_1.B a_134283_44135# GND.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1344 Comparator_0.Vinm CDAC8_0.switch_7.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1345 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t672 VDD.t673 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1346 a_90535_13083# RingCounter_0.D_FlipFlop_12.3-input-nand_1.B a_89921_13083# GND.t731 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1347 Comparator_0.Vinm CDAC8_0.switch_8.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1348 VDD.t182 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_5.B.t0 VDD.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1349 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 CLK.t104 GND.t456 GND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1350 D_FlipFlop_4.3-input-nand_2.C.t0 D_FlipFlop_4.3-input-nand_1.Vout VDD.t94 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1351 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 VDD.t947 VDD.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1352 GND.t494 EN.t91 a_51369_15797# GND.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1353 GND.t31 Nand_Gate_6.B.t15 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1354 VDD.t787 a_139663_37417.t3 a_138533_35417.t1 VDD.t786 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X1355 VDD.t671 VDD.t670 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 VDD.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1356 Nand_Gate_0.A.t2 RingCounter_0.D_FlipFlop_2.Qbar VDD.t365 VDD.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1357 a_107927_15797# RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout GND.t728 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1358 a_75898_21528# Q1.t7 VDD.t903 VDD.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1359 Nand_Gate_1.B.t0 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t307 VDD.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1360 Nand_Gate_4.A.t0 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t297 VDD.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1361 GND.t783 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 a_74807_13083# GND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1362 VDD.t660 And_Gate_4.Vout.t7 D_FlipFlop_2.Inverter_1.Vout VDD.t659 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1363 VDD.t49 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1364 Comparator_0.Vinm CDAC8_0.switch_7.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1365 VDD.t265 D_FlipFlop_5.Qbar Q2.t0 VDD.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1366 VDD.t962 D_FlipFlop_7.D.t29 D_FlipFlop_1.3-input-nand_1.B VDD.t961 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1367 VDD.t839 Nand_Gate_2.A.t14 Nand_Gate_2.Vout.t0 VDD.t838 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1368 Comparator_0.Vinm CDAC8_0.switch_6.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1369 a_79625_49858# VDD.t1152 GND.t822 GND.t821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1370 Nand_Gate_5.B.t2 RingCounter_0.D_FlipFlop_6.Qbar VDD.t184 VDD.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1371 Comparator_0.Vinm CDAC8_0.switch_7.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1372 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 VDD.t140 VDD.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1373 Comparator_0.Vinm CDAC8_0.switch_6.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1374 VDD.t355 FFCLR.t49 D_FlipFlop_7.3-input-nand_0.Vout VDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1375 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.3-input-nand_1.B VDD.t638 VDD.t393 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1376 VDD.t964 D_FlipFlop_7.D.t30 D_FlipFlop_0.3-input-nand_1.B VDD.t963 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1377 Comparator_0.Vinm CDAC8_0.switch_7.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1378 VDD.t450 EN.t92 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 VDD.t449 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1379 a_110029_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 GND.t603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1380 VDD.t598 D_FlipFlop_5.3-input-nand_2.Vout.t6 D_FlipFlop_5.3-input-nand_2.C.t2 VDD.t597 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1381 a_58159_49858# RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 a_57545_49858# GND.t691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1382 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 VDD.t956 VDD.t821 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1383 VDD.t357 FFCLR.t50 D_FlipFlop_3.Qbar VDD.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1384 GND.t632 D_FlipFlop_5.3-input-nand_2.Vout.t7 a_130209_26914# GND.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1385 Comparator_0.Vinm CDAC8_0.switch_7.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1386 VDD.t448 EN.t93 Nand_Gate_4.A.t1 VDD.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1387 Comparator_0.Vinm CDAC8_0.switch_9.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1388 VDD.t359 FFCLR.t51 D_FlipFlop_5.3-input-nand_2.C.t1 VDD.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1389 GND.t650 FFCLR.t52 a_134897_26914# GND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1390 And_Gate_1.Vout.t0 And_Gate_1.Nand_Gate_0.Vout VDD.t932 VDD.t931 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1391 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 VDD.t287 VDD.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1392 VDD.t1013 CLK.t105 And_Gate_0.Nand_Gate_0.Vout VDD.t1012 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1393 Q2.t2 D_FlipFlop_5.Nand_Gate_0.Vout VDD.t423 VDD.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1394 Comparator_0.Vinm CDAC8_0.switch_6.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1395 VDD.t825 D_FlipFlop_2.Qbar Q6.t2 VDD.t808 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1396 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 a_76165_52572# GND.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1397 GND.t458 CLK.t106 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 GND.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1398 GND.t460 CLK.t107 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 GND.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1399 VDD.t1011 CLK.t108 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 VDD.t1010 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1400 a_94915_13083# Nand_Gate_6.B.t16 RingCounter_0.D_FlipFlop_11.Qbar GND.t810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1401 RingCounter_0.D_FlipFlop_16.Q.t2 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t428 VDD.t427 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1402 GND.t652 FFCLR.t53 a_128851_44135# GND.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1403 a_99603_13083# RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 a_98989_13083# GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1404 Comparator_0.Vinm CDAC8_0.switch_7.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1405 a_75898_39392# Q6.t7 VDD.t811 VDD.t810 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1406 GND.t850 D_FlipFlop_7.D.t31 D_FlipFlop_3.3-input-nand_1.B GND.t849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1407 a_138485_16882.t2 a_138485_16882.t1 Vbias.t6 Vbias.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X1408 Comparator_0.Vinm CDAC8_0.switch_5.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1409 a_119711_49858# VDD.t1153 GND.t824 GND.t823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1410 a_95659_52572# VDD.t1154 GND.t826 GND.t825 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1411 a_128237_24200# Q2.t9 D_FlipFlop_5.Qbar GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1412 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B Nand_Gate_2.A.t15 VDD.t841 VDD.t840 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1413 Comparator_0.Vinm CDAC8_0.switch_7.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1414 VDD.t857 D_FlipFlop_6.Qbar Q1.t2 VDD.t856 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1415 a_75898_18814# Q0.t7 VDD.t87 VDD.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1416 GND.t245 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 a_85847_15797# GND.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1417 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 CLK.t109 a_85233_49858# GND.t461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1418 Q6.t1 D_FlipFlop_2.Nand_Gate_0.Vout VDD.t540 VDD.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1419 GND.t363 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 a_41687_13083# GND.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1420 GND.t40 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 a_118967_13083# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1421 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 VDD.t776 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1422 VDD.t446 EN.t94 RingCounter_0.D_FlipFlop_16.Q.t3 VDD.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1423 a_46505_49858# EN.t95 GND.t492 GND.t491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1424 GND.t828 VDD.t1155 a_99603_13083# GND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1425 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 Nand_Gate_6.B.t17 VDD.t937 VDD.t858 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1426 GND.t621 And_Gate_6.Vout.t6 D_FlipFlop_3.Inverter_1.Vout GND.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1427 Comparator_0.Vinm CDAC8_0.switch_7.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1428 And_Gate_5.Vout.t1 And_Gate_5.Nand_Gate_0.Vout GND.t727 GND.t726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1429 Comparator_0.Vinm CDAC8_0.switch_6.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1430 And_Gate_3.Nand_Gate_0.Vout Nand_Gate_1.Vout.t4 VDD.t951 VDD.t950 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1431 a_96273_52572# Nand_Gate_2.A.t16 a_95659_52572# GND.t720 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1432 Comparator_0.Vinm CDAC8_0.switch_7.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1433 Comparator_0.Vinm CDAC8_0.switch_6.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1434 Q1.t0 D_FlipFlop_6.Nand_Gate_0.Vout VDD.t845 VDD.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1435 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B RingCounter_0.D_FlipFlop_16.Q.t9 GND.t642 GND.t641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1436 a_41687_13083# RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1437 a_130209_39721# D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1438 a_46375_13083# RingCounter_0.D_FlipFlop_8.3-input-nand_1.B a_45761_13083# GND.t809 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1439 a_101705_49858# VDD.t1156 GND.t830 GND.t829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1440 Comparator_0.Vinm CDAC8_0.switch_7.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1441 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 VDD.t594 VDD.t593 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1442 VDD.t1009 CLK.t110 And_Gate_3.Nand_Gate_0.Vout VDD.t1008 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1443 Comparator_0.Vinm CDAC8_0.switch_9.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1444 GND.t857 Nand_Gate_4.B.t14 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B GND.t856 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1445 a_128237_20636# Q1.t8 D_FlipFlop_6.Qbar GND.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1446 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 a_43045_52572# GND.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1447 VDD.t1007 CLK.t111 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 VDD.t1006 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1448 Comparator_0.Vinm CDAC8_0.switch_6.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1449 GND.t253 D_FlipFlop_7.3-input-nand_2.C.t6 a_130209_17072# GND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1450 a_61795_13083# Nand_Gate_7.A.t10 RingCounter_0.D_FlipFlop_14.Qbar GND.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1451 a_130209_23350# D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout GND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1452 a_101575_13083# RingCounter_0.D_FlipFlop_11.3-input-nand_1.B a_100961_13083# GND.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1453 VDD.t816 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout VDD.t815 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1454 a_120325_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_119711_52572# GND.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1455 GND.t837 Nand_Gate_4.B.t15 a_134897_17072# GND.t836 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1456 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_7.D.t32 VDD.t965 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1457 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 VDD.t633 VDD.t632 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1458 Comparator_0.Vinm CDAC8_0.switch_7.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1459 VDD.t640 FFCLR.t54 D_FlipFlop_7.Qbar VDD.t639 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1460 GND.t669 D_FlipFlop_4.3-input-nand_2.C.t7 a_130209_27764# GND.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1461 a_62539_52572# VDD.t1157 GND.t832 GND.t831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1462 VDD.t270 Q7.t8 CDAC8_0.switch_7.Z.t1 GND.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1463 GND.t705 Nand_Gate_1.A.t9 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B GND.t704 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1464 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B Nand_Gate_3.B.t10 VDD.t917 VDD.t916 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1465 GND.t772 Nand_Gate_1.B.t17 a_134897_27764# GND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1466 VDD.t641 FFCLR.t55 D_FlipFlop_4.3-input-nand_0.Vout VDD.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1467 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_0.3-input-nand_1.B VDD.t334 VDD.t333 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1468 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 Nand_Gate_6.A.t10 VDD.t801 VDD.t800 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1469 GND.t625 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 a_52727_15797# GND.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1470 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 CLK.t112 a_52113_49858# GND.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1471 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 EN.t96 VDD.t444 VDD.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1472 a_128851_33443# D_FlipFlop_1.Nand_Gate_1.Vout a_128237_33443# GND.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1473 VDD.t258 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 VDD.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1474 a_134283_40571# And_Gate_6.Vout.t7 D_FlipFlop_3.3-input-nand_1.Vout GND.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1475 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 VDD.t618 VDD.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1476 D_FlipFlop_7.D.t33 Vbias.t0 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X1477 a_89307_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 GND.t690 GND.t689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1478 CDAC8_0.switch_7.Z.t2 a_75898_35820# GND.t766 GND.t765 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1479 GND.t834 VDD.t1158 a_66483_13083# GND.t833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1480 GND.t852 D_FlipFlop_7.D.t34 D_FlipFlop_7.3-input-nand_1.B GND.t851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1481 a_111387_49858# RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 GND.t344 GND.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1482 a_63153_52572# Nand_Gate_3.B.t11 a_62539_52572# GND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1483 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 a_98245_49858# GND.t412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1484 VDD.t20 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1485 a_139663_37417.t2 Comparator_0.Vinm a_139804_27676.t2 Vbias.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X1486 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 a_67227_52572# GND.t588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1487 VDD.t104 And_Gate_5.Vout.t7 D_FlipFlop_1.Inverter_1.Vout VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1488 Comparator_0.Vinm CDAC8_0.switch_7.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1489 And_Gate_6.Vout.t0 And_Gate_6.Nand_Gate_0.Vout VDD.t879 VDD.t878 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1490 VDD.t442 EN.t97 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 VDD.t441 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1491 a_132311_43285# D_FlipFlop_3.3-input-nand_2.C.t7 D_FlipFlop_3.3-input-nand_2.Vout.t3 GND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1492 VDD.t886 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 VDD.t871 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1493 VDD.t440 EN.t98 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 VDD.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1494 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 VDD.t960 VDD.t237 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1495 VDD.t175 D_FlipFlop_2.3-input-nand_2.Vout.t7 D_FlipFlop_2.3-input-nand_2.C.t0 VDD.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1496 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 VDD.t768 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1497 a_72835_15797# RingCounter_0.D_FlipFlop_13.Qbar Nand_Gate_7.B.t0 GND.t409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1498 a_139804_27676.t0 a_138485_16882.t4 Vbias.t4 Vbias.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X1499 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 a_122427_52572# GND.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1500 a_77523_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 a_76909_15797# GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1501 VDD.t643 FFCLR.t56 D_FlipFlop_2.3-input-nand_2.C.t3 VDD.t642 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1502 a_105955_13083# Nand_Gate_1.A.t10 RingCounter_0.D_FlipFlop_9.Qbar GND.t706 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1503 VDD.t802 Nand_Gate_6.A.t11 RingCounter_0.D_FlipFlop_12.Qbar VDD.t590 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1504 Comparator_0.Vinm CDAC8_0.switch_7.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1505 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 VDD.t267 VDD.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1506 Comparator_0.Vinm CDAC8_0.switch_7.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1507 VDD.t252 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout Nand_Gate_0.A.t0 VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1508 Comparator_0.Vinm CDAC8_0.switch_7.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1509 a_132925_43285# D_FlipFlop_3.3-input-nand_0.Vout a_132311_43285# GND.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1510 a_128237_37007# Q6.t8 D_FlipFlop_2.Qbar GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1511 VDD.t655 And_Gate_5.A.t4 And_Gate_5.Nand_Gate_0.Vout VDD.t654 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1512 Comparator_0.Vinm CDAC8_0.switch_7.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1513 GND.t786 Q1.t9 CDAC8_0.switch_2.Z.t3 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1514 a_75898_28676# Q3.t9 GND.t590 GND.t589 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1515 VDD.t279 Q5.t9 D_FlipFlop_3.Qbar VDD.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1516 Comparator_0.Vinm CDAC8_0.switch_7.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1517 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 Nand_Gate_4.B.t16 VDD.t952 VDD.t934 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1518 VDD.t927 And_Gate_2.Vout.t6 D_FlipFlop_5.3-input-nand_1.Vout VDD.t923 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1519 RingCounter_0.D_FlipFlop_3.Qbar Nand_Gate_0.B.t11 a_80239_49858# GND.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1520 VDD.t669 VDD.t668 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 VDD.t488 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1521 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_5.3-input-nand_2.C.t7 VDD.t992 VDD.t595 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1522 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD.t666 VDD.t667 VDD.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1523 VDD.t836 Nand_Gate_2.A.t17 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t835 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1524 GND.t482 EN.t99 a_77523_15797# GND.t481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1525 Comparator_0.Vinm CDAC8_0.switch_6.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1526 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 VDD.t285 VDD.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1527 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 CLK.t113 VDD.t1005 VDD.t1004 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1528 Comparator_0.Vinm CDAC8_0.switch_9.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1529 Comparator_0.Vinm CDAC8_0.switch_7.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1530 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK.t114 VDD.t1003 VDD.t1002 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1531 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 Nand_Gate_1.A.t11 VDD.t814 VDD.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1532 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.D.t35 VDD.t338 VDD.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1533 a_91279_52572# RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_90665_52572# GND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1534 a_92725_16975# CLK.t115 GND.t306 GND.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1535 a_117609_15797# RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_116995_15797# GND.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1536 GND.t653 FFCLR.t57 a_132925_24200# GND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1537 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 a_65125_49858# GND.t709 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1538 Comparator_0.Vinm CDAC8_0.switch_7.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1539 VDD.t311 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 VDD.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1540 Comparator_0.Vinm CDAC8_0.switch_6.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1541 D_FlipFlop_3.Qbar D_FlipFlop_3.Nand_Gate_1.Vout VDD.t294 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1542 VDD.t317 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1543 a_78881_13083# CLK.t116 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 GND.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1544 a_97631_52572# EN.t100 GND.t490 GND.t489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1545 VDD.t438 EN.t101 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 VDD.t437 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1546 VDD.t186 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1547 Comparator_0.Vinm CDAC8_0.switch_7.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1548 Comparator_0.Vinm CDAC8_0.switch_5.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1549 VDD.t645 FFCLR.t58 D_FlipFlop_4.Qbar VDD.t644 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1550 And_Gate_0.Nand_Gate_0.Vout And_Gate_0.B.t4 a_70645_16975# GND.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1551 a_84619_49858# EN.t102 GND.t488 GND.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1552 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 VDD.t57 VDD.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1553 GND.t486 EN.t103 a_79495_13083# GND.t485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1554 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 a_120325_49858# GND.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1555 a_44403_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 a_43789_15797# GND.t839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1556 Nand_Gate_3.B.t3 EN.t104 VDD.t436 VDD.t435 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1557 a_130209_36157# D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout GND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1558 a_128851_44135# D_FlipFlop_0.Nand_Gate_1.Vout a_128237_44135# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1559 a_98989_13083# RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 GND.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1560 GND.t700 Q6.t9 CDAC8_0.switch_6.Z.t2 VDD.t812 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1561 GND.t484 EN.t105 a_117609_15797# GND.t483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1562 VDD.t953 Nand_Gate_4.B.t17 RingCounter_0.D_FlipFlop_15.Qbar VDD.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1563 a_134283_26914# And_Gate_2.Vout.t7 D_FlipFlop_5.3-input-nand_0.Vout GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1564 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 VDD.t543 VDD.t378 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1565 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 VDD.t611 VDD.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1566 a_130209_46849# D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_0.Vout GND.t872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1567 a_98245_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_97631_52572# GND.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1568 a_132311_19786# D_FlipFlop_7.3-input-nand_2.C.t7 D_FlipFlop_7.3-input-nand_2.Vout.t1 GND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1569 GND.t73 Q0.t8 CDAC8_0.switch_1.Z.t2 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1570 Comparator_0.Vinm CDAC8_0.switch_7.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1571 a_85233_49858# RingCounter_0.D_FlipFlop_4.3-input-nand_1.B a_84619_49858# GND.t472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1572 Nand_Gate_5.A.t1 EN.t106 VDD.t434 VDD.t433 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1573 VDD.t59 D_FlipFlop_0.CLK.t7 D_FlipFlop_0.Inverter_1.Vout VDD.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1574 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 a_89307_49858# GND.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1575 VDD.t665 VDD.t664 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 VDD.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1576 a_29289_15797# RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_28675_15797# GND.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1577 VDD.t933 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1578 GND.t339 FFCLR.t59 a_132925_20636# GND.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1579 a_130209_30478# D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_0.Vout GND.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1580 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 VDD.t262 VDD.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1581 GND.t476 EN.t107 a_44403_15797# GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1582 GND.t794 And_Gate_1.Vout.t7 D_FlipFlop_7.Inverter_1.Vout GND.t793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1583 VDD.t549 RingCounter_0.D_FlipFlop_9.Qbar Nand_Gate_1.A.t2 VDD.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1584 Comparator_0.Vinm CDAC8_0.switch_6.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1585 RingCounter_0.D_FlipFlop_4.Qbar VDD.t662 VDD.t663 VDD.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1586 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 CLK.t117 VDD.t1001 VDD.t1000 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1587 a_132925_19786# D_FlipFlop_7.3-input-nand_0.Vout a_132311_19786# GND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1588 Comparator_0.Vinm CDAC8_0.switch_7.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1589 a_59977_16975# Nand_Gate_7.A.t11 GND.t432 GND.t431 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1590 GND.t4 And_Gate_3.Vout.t7 D_FlipFlop_4.Inverter_1.Vout GND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1591 a_75898_35820# Q7.t9 VDD.t272 VDD.t271 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1592 a_28675_15797# RingCounter_0.D_FlipFlop_16.Qbar RingCounter_0.D_FlipFlop_16.Q.t0 GND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1593 VDD.t545 Q0.t9 D_FlipFlop_7.Qbar VDD.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
R0 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.t0 168.609
R1 CDAC8_0.switch_7.Z CDAC8_0.switch_7.Z.t3 168.565
R2 CDAC8_0.switch_7.Z.n0 CDAC8_0.switch_7.Z.t2 60.321
R3 CDAC8_0.switch_7.Z.n0 CDAC8_0.switch_7.Z.t1 60.321
R4 CDAC8_0.switch_7.Z.n237 CDAC8_0.switch_7.Z.n236 40.463
R5 CDAC8_0.switch_7.Z.n296 CDAC8_0.switch_7.Z.n2 20.4699
R6 CDAC8_0.switch_7.Z.n296 CDAC8_0.switch_7.Z.n295 19.9889
R7 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.n296 11.6479
R8 CDAC8_0.switch_7.Z.n48 CDAC8_0.switch_7.Z.n47 4.61363
R9 CDAC8_0.switch_7.Z.n46 CDAC8_0.switch_7.Z.n36 4.61363
R10 CDAC8_0.switch_7.Z.n53 CDAC8_0.switch_7.Z.n52 4.61363
R11 CDAC8_0.switch_7.Z.n34 CDAC8_0.switch_7.Z.n26 4.61363
R12 CDAC8_0.switch_7.Z.n56 CDAC8_0.switch_7.Z.n55 4.61363
R13 CDAC8_0.switch_7.Z.n32 CDAC8_0.switch_7.Z.n24 4.61363
R14 CDAC8_0.switch_7.Z.n61 CDAC8_0.switch_7.Z.n60 4.61363
R15 CDAC8_0.switch_7.Z.n30 CDAC8_0.switch_7.Z.n22 4.61363
R16 CDAC8_0.switch_7.Z.n65 CDAC8_0.switch_7.Z.n64 4.61363
R17 CDAC8_0.switch_7.Z.n28 CDAC8_0.switch_7.Z.n20 4.61363
R18 CDAC8_0.switch_7.Z.n69 CDAC8_0.switch_7.Z.n18 4.61363
R19 CDAC8_0.switch_7.Z.n70 CDAC8_0.switch_7.Z.n13 4.61363
R20 CDAC8_0.switch_7.Z.n74 CDAC8_0.switch_7.Z.n3 4.61363
R21 CDAC8_0.switch_7.Z.n75 CDAC8_0.switch_7.Z.n74 4.61363
R22 CDAC8_0.switch_7.Z.n15 CDAC8_0.switch_7.Z.n5 4.61363
R23 CDAC8_0.switch_7.Z.n293 CDAC8_0.switch_7.Z.n292 4.61363
R24 CDAC8_0.switch_7.Z.n287 CDAC8_0.switch_7.Z.n9 4.61363
R25 CDAC8_0.switch_7.Z.n288 CDAC8_0.switch_7.Z.n8 4.61363
R26 CDAC8_0.switch_7.Z.n283 CDAC8_0.switch_7.Z.n282 4.61363
R27 CDAC8_0.switch_7.Z.n239 CDAC8_0.switch_7.Z.n80 4.61363
R28 CDAC8_0.switch_7.Z.n280 CDAC8_0.switch_7.Z.n279 4.61363
R29 CDAC8_0.switch_7.Z.n241 CDAC8_0.switch_7.Z.n83 4.61363
R30 CDAC8_0.switch_7.Z.n275 CDAC8_0.switch_7.Z.n274 4.61363
R31 CDAC8_0.switch_7.Z.n243 CDAC8_0.switch_7.Z.n85 4.61363
R32 CDAC8_0.switch_7.Z.n272 CDAC8_0.switch_7.Z.n271 4.61363
R33 CDAC8_0.switch_7.Z.n245 CDAC8_0.switch_7.Z.n87 4.61363
R34 CDAC8_0.switch_7.Z.n247 CDAC8_0.switch_7.Z.n89 4.61363
R35 CDAC8_0.switch_7.Z.n267 CDAC8_0.switch_7.Z.n266 4.61363
R36 CDAC8_0.switch_7.Z.n264 CDAC8_0.switch_7.Z.n263 4.61363
R37 CDAC8_0.switch_7.Z.n261 CDAC8_0.switch_7.Z.n249 4.61363
R38 CDAC8_0.switch_7.Z.n221 CDAC8_0.switch_7.Z.n220 4.61363
R39 CDAC8_0.switch_7.Z.n159 CDAC8_0.switch_7.Z.n158 4.61363
R40 CDAC8_0.switch_7.Z.n156 CDAC8_0.switch_7.Z.n144 4.61363
R41 CDAC8_0.switch_7.Z.n162 CDAC8_0.switch_7.Z.n161 4.61363
R42 CDAC8_0.switch_7.Z.n142 CDAC8_0.switch_7.Z.n132 4.61363
R43 CDAC8_0.switch_7.Z.n167 CDAC8_0.switch_7.Z.n166 4.61363
R44 CDAC8_0.switch_7.Z.n140 CDAC8_0.switch_7.Z.n130 4.61363
R45 CDAC8_0.switch_7.Z.n170 CDAC8_0.switch_7.Z.n169 4.61363
R46 CDAC8_0.switch_7.Z.n138 CDAC8_0.switch_7.Z.n128 4.61363
R47 CDAC8_0.switch_7.Z.n175 CDAC8_0.switch_7.Z.n174 4.61363
R48 CDAC8_0.switch_7.Z.n136 CDAC8_0.switch_7.Z.n126 4.61363
R49 CDAC8_0.switch_7.Z.n179 CDAC8_0.switch_7.Z.n178 4.61363
R50 CDAC8_0.switch_7.Z.n134 CDAC8_0.switch_7.Z.n124 4.61363
R51 CDAC8_0.switch_7.Z.n183 CDAC8_0.switch_7.Z.n122 4.61363
R52 CDAC8_0.switch_7.Z.n184 CDAC8_0.switch_7.Z.n121 4.61363
R53 CDAC8_0.switch_7.Z.n192 CDAC8_0.switch_7.Z.n191 4.61363
R54 CDAC8_0.switch_7.Z.n188 CDAC8_0.switch_7.Z.n118 4.61363
R55 CDAC8_0.switch_7.Z.n196 CDAC8_0.switch_7.Z.n90 4.61363
R56 CDAC8_0.switch_7.Z.n197 CDAC8_0.switch_7.Z.n115 4.61363
R57 CDAC8_0.switch_7.Z.n234 CDAC8_0.switch_7.Z.n233 4.61363
R58 CDAC8_0.switch_7.Z.n113 CDAC8_0.switch_7.Z.n92 4.61363
R59 CDAC8_0.switch_7.Z.n229 CDAC8_0.switch_7.Z.n228 4.61363
R60 CDAC8_0.switch_7.Z.n111 CDAC8_0.switch_7.Z.n95 4.61363
R61 CDAC8_0.switch_7.Z.n226 CDAC8_0.switch_7.Z.n225 4.61363
R62 CDAC8_0.switch_7.Z.n109 CDAC8_0.switch_7.Z.n97 4.61363
R63 CDAC8_0.switch_7.Z.n107 CDAC8_0.switch_7.Z.n99 4.61363
R64 CDAC8_0.switch_7.Z.n218 CDAC8_0.switch_7.Z.n217 4.61363
R65 CDAC8_0.switch_7.Z.n105 CDAC8_0.switch_7.Z.n101 4.61363
R66 CDAC8_0.switch_7.Z.n211 CDAC8_0.switch_7.Z.n102 4.61363
R67 CDAC8_0.switch_7.Z.n213 CDAC8_0.switch_7.Z.n212 4.61363
R68 CDAC8_0.switch_7.Z.n48 CDAC8_0.switch_7.Z.n46 4.23363
R69 CDAC8_0.switch_7.Z.n52 CDAC8_0.switch_7.Z.n26 4.23363
R70 CDAC8_0.switch_7.Z.n56 CDAC8_0.switch_7.Z.n24 4.23363
R71 CDAC8_0.switch_7.Z.n60 CDAC8_0.switch_7.Z.n22 4.23363
R72 CDAC8_0.switch_7.Z.n65 CDAC8_0.switch_7.Z.n20 4.23363
R73 CDAC8_0.switch_7.Z.n70 CDAC8_0.switch_7.Z.n69 4.23363
R74 CDAC8_0.switch_7.Z.n292 CDAC8_0.switch_7.Z.n5 4.23363
R75 CDAC8_0.switch_7.Z.n288 CDAC8_0.switch_7.Z.n287 4.23363
R76 CDAC8_0.switch_7.Z.n283 CDAC8_0.switch_7.Z.n80 4.23363
R77 CDAC8_0.switch_7.Z.n279 CDAC8_0.switch_7.Z.n83 4.23363
R78 CDAC8_0.switch_7.Z.n275 CDAC8_0.switch_7.Z.n85 4.23363
R79 CDAC8_0.switch_7.Z.n271 CDAC8_0.switch_7.Z.n87 4.23363
R80 CDAC8_0.switch_7.Z.n267 CDAC8_0.switch_7.Z.n89 4.23363
R81 CDAC8_0.switch_7.Z.n263 CDAC8_0.switch_7.Z.n261 4.23363
R82 CDAC8_0.switch_7.Z.n158 CDAC8_0.switch_7.Z.n156 4.23363
R83 CDAC8_0.switch_7.Z.n162 CDAC8_0.switch_7.Z.n132 4.23363
R84 CDAC8_0.switch_7.Z.n166 CDAC8_0.switch_7.Z.n130 4.23363
R85 CDAC8_0.switch_7.Z.n170 CDAC8_0.switch_7.Z.n128 4.23363
R86 CDAC8_0.switch_7.Z.n174 CDAC8_0.switch_7.Z.n126 4.23363
R87 CDAC8_0.switch_7.Z.n179 CDAC8_0.switch_7.Z.n124 4.23363
R88 CDAC8_0.switch_7.Z.n184 CDAC8_0.switch_7.Z.n183 4.23363
R89 CDAC8_0.switch_7.Z.n192 CDAC8_0.switch_7.Z.n188 4.23363
R90 CDAC8_0.switch_7.Z.n197 CDAC8_0.switch_7.Z.n196 4.23363
R91 CDAC8_0.switch_7.Z.n233 CDAC8_0.switch_7.Z.n92 4.23363
R92 CDAC8_0.switch_7.Z.n229 CDAC8_0.switch_7.Z.n95 4.23363
R93 CDAC8_0.switch_7.Z.n225 CDAC8_0.switch_7.Z.n97 4.23363
R94 CDAC8_0.switch_7.Z.n221 CDAC8_0.switch_7.Z.n99 4.23363
R95 CDAC8_0.switch_7.Z.n217 CDAC8_0.switch_7.Z.n101 4.23363
R96 CDAC8_0.switch_7.Z.n213 CDAC8_0.switch_7.Z.n211 4.23363
R97 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.n1 1.60376
R98 CDAC8_0.switch_7.Z.n262 CDAC8_0.switch_7.Z.t127 0.726216
R99 CDAC8_0.switch_7.Z.n260 CDAC8_0.switch_7.Z.t43 0.726216
R100 CDAC8_0.switch_7.Z.n264 CDAC8_0.switch_7.Z.t9 0.726216
R101 CDAC8_0.switch_7.Z.n249 CDAC8_0.switch_7.Z.t105 0.726216
R102 CDAC8_0.switch_7.Z.n210 CDAC8_0.switch_7.Z.t80 0.726216
R103 CDAC8_0.switch_7.Z.n214 CDAC8_0.switch_7.Z.t40 0.726216
R104 CDAC8_0.switch_7.Z.n102 CDAC8_0.switch_7.Z.t19 0.726216
R105 CDAC8_0.switch_7.Z.n212 CDAC8_0.switch_7.Z.t101 0.726216
R106 CDAC8_0.switch_7.Z.n159 CDAC8_0.switch_7.Z.t90 0.658247
R107 CDAC8_0.switch_7.Z.n36 CDAC8_0.switch_7.Z.t98 0.658247
R108 CDAC8_0.switch_7.Z.n47 CDAC8_0.switch_7.Z.t129 0.658247
R109 CDAC8_0.switch_7.Z.n45 CDAC8_0.switch_7.Z.t36 0.658247
R110 CDAC8_0.switch_7.Z.n49 CDAC8_0.switch_7.Z.t117 0.658247
R111 CDAC8_0.switch_7.Z.n144 CDAC8_0.switch_7.Z.t8 0.658247
R112 CDAC8_0.switch_7.Z.n157 CDAC8_0.switch_7.Z.t30 0.658247
R113 CDAC8_0.switch_7.Z.n155 CDAC8_0.switch_7.Z.t70 0.658247
R114 CDAC8_0.switch_7.Z.n160 CDAC8_0.switch_7.Z.t86 0.611304
R115 CDAC8_0.switch_7.Z.n129 CDAC8_0.switch_7.Z.t112 0.611304
R116 CDAC8_0.switch_7.Z.n168 CDAC8_0.switch_7.Z.t107 0.611304
R117 CDAC8_0.switch_7.Z.n125 CDAC8_0.switch_7.Z.t32 0.611304
R118 CDAC8_0.switch_7.Z.n176 CDAC8_0.switch_7.Z.t49 0.611304
R119 CDAC8_0.switch_7.Z.n177 CDAC8_0.switch_7.Z.t44 0.611304
R120 CDAC8_0.switch_7.Z.n189 CDAC8_0.switch_7.Z.t69 0.611304
R121 CDAC8_0.switch_7.Z.n190 CDAC8_0.switch_7.Z.t65 0.611304
R122 CDAC8_0.switch_7.Z.n35 CDAC8_0.switch_7.Z.t92 0.611304
R123 CDAC8_0.switch_7.Z.n33 CDAC8_0.switch_7.Z.t120 0.611304
R124 CDAC8_0.switch_7.Z.n31 CDAC8_0.switch_7.Z.t113 0.611304
R125 CDAC8_0.switch_7.Z.n29 CDAC8_0.switch_7.Z.t39 0.611304
R126 CDAC8_0.switch_7.Z.n27 CDAC8_0.switch_7.Z.t58 0.611304
R127 CDAC8_0.switch_7.Z.n12 CDAC8_0.switch_7.Z.t51 0.611304
R128 CDAC8_0.switch_7.Z.n294 CDAC8_0.switch_7.Z.t76 0.611304
R129 CDAC8_0.switch_7.Z.n4 CDAC8_0.switch_7.Z.t71 0.611304
R130 CDAC8_0.switch_7.Z.n238 CDAC8_0.switch_7.Z.t128 0.611304
R131 CDAC8_0.switch_7.Z.n240 CDAC8_0.switch_7.Z.t21 0.611304
R132 CDAC8_0.switch_7.Z.n242 CDAC8_0.switch_7.Z.t16 0.611304
R133 CDAC8_0.switch_7.Z.n244 CDAC8_0.switch_7.Z.t38 0.611304
R134 CDAC8_0.switch_7.Z.n246 CDAC8_0.switch_7.Z.t89 0.611304
R135 CDAC8_0.switch_7.Z.n248 CDAC8_0.switch_7.Z.t84 0.611304
R136 CDAC8_0.switch_7.Z.n25 CDAC8_0.switch_7.Z.t125 0.611304
R137 CDAC8_0.switch_7.Z.n54 CDAC8_0.switch_7.Z.t23 0.611304
R138 CDAC8_0.switch_7.Z.n21 CDAC8_0.switch_7.Z.t17 0.611304
R139 CDAC8_0.switch_7.Z.n62 CDAC8_0.switch_7.Z.t66 0.611304
R140 CDAC8_0.switch_7.Z.n63 CDAC8_0.switch_7.Z.t85 0.611304
R141 CDAC8_0.switch_7.Z.n17 CDAC8_0.switch_7.Z.t81 0.611304
R142 CDAC8_0.switch_7.Z.n16 CDAC8_0.switch_7.Z.t106 0.611304
R143 CDAC8_0.switch_7.Z.n14 CDAC8_0.switch_7.Z.t103 0.611304
R144 CDAC8_0.switch_7.Z.n81 CDAC8_0.switch_7.Z.t35 0.611304
R145 CDAC8_0.switch_7.Z.n281 CDAC8_0.switch_7.Z.t52 0.611304
R146 CDAC8_0.switch_7.Z.n82 CDAC8_0.switch_7.Z.t46 0.611304
R147 CDAC8_0.switch_7.Z.n273 CDAC8_0.switch_7.Z.t64 0.611304
R148 CDAC8_0.switch_7.Z.n86 CDAC8_0.switch_7.Z.t122 0.611304
R149 CDAC8_0.switch_7.Z.n44 CDAC8_0.switch_7.Z.t29 0.611304
R150 CDAC8_0.switch_7.Z.n42 CDAC8_0.switch_7.Z.t54 0.611304
R151 CDAC8_0.switch_7.Z.n40 CDAC8_0.switch_7.Z.t48 0.611304
R152 CDAC8_0.switch_7.Z.n38 CDAC8_0.switch_7.Z.t100 0.611304
R153 CDAC8_0.switch_7.Z.n11 CDAC8_0.switch_7.Z.t121 0.611304
R154 CDAC8_0.switch_7.Z.n72 CDAC8_0.switch_7.Z.t114 0.611304
R155 CDAC8_0.switch_7.Z.n6 CDAC8_0.switch_7.Z.t14 0.611304
R156 CDAC8_0.switch_7.Z.n290 CDAC8_0.switch_7.Z.t6 0.611304
R157 CDAC8_0.switch_7.Z.n7 CDAC8_0.switch_7.Z.t62 0.611304
R158 CDAC8_0.switch_7.Z.n251 CDAC8_0.switch_7.Z.t82 0.611304
R159 CDAC8_0.switch_7.Z.n253 CDAC8_0.switch_7.Z.t77 0.611304
R160 CDAC8_0.switch_7.Z.n255 CDAC8_0.switch_7.Z.t99 0.611304
R161 CDAC8_0.switch_7.Z.n50 CDAC8_0.switch_7.Z.t111 0.611304
R162 CDAC8_0.switch_7.Z.n23 CDAC8_0.switch_7.Z.t12 0.611304
R163 CDAC8_0.switch_7.Z.n58 CDAC8_0.switch_7.Z.t5 0.611304
R164 CDAC8_0.switch_7.Z.n19 CDAC8_0.switch_7.Z.t57 0.611304
R165 CDAC8_0.switch_7.Z.n67 CDAC8_0.switch_7.Z.t74 0.611304
R166 CDAC8_0.switch_7.Z.n10 CDAC8_0.switch_7.Z.t68 0.611304
R167 CDAC8_0.switch_7.Z.n76 CDAC8_0.switch_7.Z.t97 0.611304
R168 CDAC8_0.switch_7.Z.n78 CDAC8_0.switch_7.Z.t91 0.611304
R169 CDAC8_0.switch_7.Z.n285 CDAC8_0.switch_7.Z.t20 0.611304
R170 CDAC8_0.switch_7.Z.n79 CDAC8_0.switch_7.Z.t42 0.611304
R171 CDAC8_0.switch_7.Z.n277 CDAC8_0.switch_7.Z.t37 0.611304
R172 CDAC8_0.switch_7.Z.n84 CDAC8_0.switch_7.Z.t55 0.611304
R173 CDAC8_0.switch_7.Z.n269 CDAC8_0.switch_7.Z.t109 0.611304
R174 CDAC8_0.switch_7.Z.n88 CDAC8_0.switch_7.Z.t104 0.611304
R175 CDAC8_0.switch_7.Z.n257 CDAC8_0.switch_7.Z.t28 0.611304
R176 CDAC8_0.switch_7.Z.n259 CDAC8_0.switch_7.Z.t22 0.611304
R177 CDAC8_0.switch_7.Z.n265 CDAC8_0.switch_7.Z.t118 0.611304
R178 CDAC8_0.switch_7.Z.n235 CDAC8_0.switch_7.Z.t123 0.611304
R179 CDAC8_0.switch_7.Z.n91 CDAC8_0.switch_7.Z.t15 0.611304
R180 CDAC8_0.switch_7.Z.n227 CDAC8_0.switch_7.Z.t10 0.611304
R181 CDAC8_0.switch_7.Z.n96 CDAC8_0.switch_7.Z.t31 0.611304
R182 CDAC8_0.switch_7.Z.n219 CDAC8_0.switch_7.Z.t83 0.611304
R183 CDAC8_0.switch_7.Z.n100 CDAC8_0.switch_7.Z.t79 0.611304
R184 CDAC8_0.switch_7.Z.n143 CDAC8_0.switch_7.Z.t4 0.611304
R185 CDAC8_0.switch_7.Z.n141 CDAC8_0.switch_7.Z.t33 0.611304
R186 CDAC8_0.switch_7.Z.n139 CDAC8_0.switch_7.Z.t26 0.611304
R187 CDAC8_0.switch_7.Z.n137 CDAC8_0.switch_7.Z.t75 0.611304
R188 CDAC8_0.switch_7.Z.n135 CDAC8_0.switch_7.Z.t96 0.611304
R189 CDAC8_0.switch_7.Z.n133 CDAC8_0.switch_7.Z.t88 0.611304
R190 CDAC8_0.switch_7.Z.n120 CDAC8_0.switch_7.Z.t116 0.611304
R191 CDAC8_0.switch_7.Z.n117 CDAC8_0.switch_7.Z.t110 0.611304
R192 CDAC8_0.switch_7.Z.n114 CDAC8_0.switch_7.Z.t41 0.611304
R193 CDAC8_0.switch_7.Z.n112 CDAC8_0.switch_7.Z.t60 0.611304
R194 CDAC8_0.switch_7.Z.n110 CDAC8_0.switch_7.Z.t56 0.611304
R195 CDAC8_0.switch_7.Z.n108 CDAC8_0.switch_7.Z.t73 0.611304
R196 CDAC8_0.switch_7.Z.n106 CDAC8_0.switch_7.Z.t130 0.611304
R197 CDAC8_0.switch_7.Z.n131 CDAC8_0.switch_7.Z.t25 0.611304
R198 CDAC8_0.switch_7.Z.n164 CDAC8_0.switch_7.Z.t50 0.611304
R199 CDAC8_0.switch_7.Z.n127 CDAC8_0.switch_7.Z.t45 0.611304
R200 CDAC8_0.switch_7.Z.n172 CDAC8_0.switch_7.Z.t95 0.611304
R201 CDAC8_0.switch_7.Z.n123 CDAC8_0.switch_7.Z.t115 0.611304
R202 CDAC8_0.switch_7.Z.n181 CDAC8_0.switch_7.Z.t108 0.611304
R203 CDAC8_0.switch_7.Z.n116 CDAC8_0.switch_7.Z.t7 0.611304
R204 CDAC8_0.switch_7.Z.n194 CDAC8_0.switch_7.Z.t131 0.611304
R205 CDAC8_0.switch_7.Z.n93 CDAC8_0.switch_7.Z.t59 0.611304
R206 CDAC8_0.switch_7.Z.n231 CDAC8_0.switch_7.Z.t78 0.611304
R207 CDAC8_0.switch_7.Z.n94 CDAC8_0.switch_7.Z.t72 0.611304
R208 CDAC8_0.switch_7.Z.n223 CDAC8_0.switch_7.Z.t94 0.611304
R209 CDAC8_0.switch_7.Z.n154 CDAC8_0.switch_7.Z.t67 0.611304
R210 CDAC8_0.switch_7.Z.n152 CDAC8_0.switch_7.Z.t93 0.611304
R211 CDAC8_0.switch_7.Z.n150 CDAC8_0.switch_7.Z.t87 0.611304
R212 CDAC8_0.switch_7.Z.n148 CDAC8_0.switch_7.Z.t13 0.611304
R213 CDAC8_0.switch_7.Z.n146 CDAC8_0.switch_7.Z.t34 0.611304
R214 CDAC8_0.switch_7.Z.n119 CDAC8_0.switch_7.Z.t27 0.611304
R215 CDAC8_0.switch_7.Z.n186 CDAC8_0.switch_7.Z.t53 0.611304
R216 CDAC8_0.switch_7.Z.n103 CDAC8_0.switch_7.Z.t47 0.611304
R217 CDAC8_0.switch_7.Z.n199 CDAC8_0.switch_7.Z.t102 0.611304
R218 CDAC8_0.switch_7.Z.n201 CDAC8_0.switch_7.Z.t124 0.611304
R219 CDAC8_0.switch_7.Z.n203 CDAC8_0.switch_7.Z.t119 0.611304
R220 CDAC8_0.switch_7.Z.n205 CDAC8_0.switch_7.Z.t11 0.611304
R221 CDAC8_0.switch_7.Z.n207 CDAC8_0.switch_7.Z.t63 0.611304
R222 CDAC8_0.switch_7.Z.n209 CDAC8_0.switch_7.Z.t61 0.611304
R223 CDAC8_0.switch_7.Z.n98 CDAC8_0.switch_7.Z.t24 0.611304
R224 CDAC8_0.switch_7.Z.n215 CDAC8_0.switch_7.Z.t18 0.611304
R225 CDAC8_0.switch_7.Z.n104 CDAC8_0.switch_7.Z.t126 0.611304
R226 CDAC8_0.switch_7.Z.n276 CDAC8_0.switch_7.Z.n275 0.3805
R227 CDAC8_0.switch_7.Z.n279 CDAC8_0.switch_7.Z.n278 0.3805
R228 CDAC8_0.switch_7.Z.n284 CDAC8_0.switch_7.Z.n283 0.3805
R229 CDAC8_0.switch_7.Z.n287 CDAC8_0.switch_7.Z.n286 0.3805
R230 CDAC8_0.switch_7.Z.n77 CDAC8_0.switch_7.Z.n5 0.3805
R231 CDAC8_0.switch_7.Z.n69 CDAC8_0.switch_7.Z.n68 0.3805
R232 CDAC8_0.switch_7.Z.n66 CDAC8_0.switch_7.Z.n65 0.3805
R233 CDAC8_0.switch_7.Z.n60 CDAC8_0.switch_7.Z.n59 0.3805
R234 CDAC8_0.switch_7.Z.n57 CDAC8_0.switch_7.Z.n56 0.3805
R235 CDAC8_0.switch_7.Z.n52 CDAC8_0.switch_7.Z.n51 0.3805
R236 CDAC8_0.switch_7.Z.n49 CDAC8_0.switch_7.Z.n48 0.3805
R237 CDAC8_0.switch_7.Z.n271 CDAC8_0.switch_7.Z.n270 0.3805
R238 CDAC8_0.switch_7.Z.n256 CDAC8_0.switch_7.Z.n87 0.3805
R239 CDAC8_0.switch_7.Z.n254 CDAC8_0.switch_7.Z.n85 0.3805
R240 CDAC8_0.switch_7.Z.n252 CDAC8_0.switch_7.Z.n83 0.3805
R241 CDAC8_0.switch_7.Z.n250 CDAC8_0.switch_7.Z.n80 0.3805
R242 CDAC8_0.switch_7.Z.n289 CDAC8_0.switch_7.Z.n288 0.3805
R243 CDAC8_0.switch_7.Z.n292 CDAC8_0.switch_7.Z.n291 0.3805
R244 CDAC8_0.switch_7.Z.n74 CDAC8_0.switch_7.Z.n73 0.3805
R245 CDAC8_0.switch_7.Z.n71 CDAC8_0.switch_7.Z.n70 0.3805
R246 CDAC8_0.switch_7.Z.n37 CDAC8_0.switch_7.Z.n20 0.3805
R247 CDAC8_0.switch_7.Z.n39 CDAC8_0.switch_7.Z.n22 0.3805
R248 CDAC8_0.switch_7.Z.n41 CDAC8_0.switch_7.Z.n24 0.3805
R249 CDAC8_0.switch_7.Z.n43 CDAC8_0.switch_7.Z.n26 0.3805
R250 CDAC8_0.switch_7.Z.n46 CDAC8_0.switch_7.Z.n45 0.3805
R251 CDAC8_0.switch_7.Z.n258 CDAC8_0.switch_7.Z.n89 0.3805
R252 CDAC8_0.switch_7.Z.n268 CDAC8_0.switch_7.Z.n267 0.3805
R253 CDAC8_0.switch_7.Z.n263 CDAC8_0.switch_7.Z.n262 0.3805
R254 CDAC8_0.switch_7.Z.n261 CDAC8_0.switch_7.Z.n260 0.3805
R255 CDAC8_0.switch_7.Z.n204 CDAC8_0.switch_7.Z.n97 0.3805
R256 CDAC8_0.switch_7.Z.n202 CDAC8_0.switch_7.Z.n95 0.3805
R257 CDAC8_0.switch_7.Z.n200 CDAC8_0.switch_7.Z.n92 0.3805
R258 CDAC8_0.switch_7.Z.n198 CDAC8_0.switch_7.Z.n197 0.3805
R259 CDAC8_0.switch_7.Z.n188 CDAC8_0.switch_7.Z.n187 0.3805
R260 CDAC8_0.switch_7.Z.n185 CDAC8_0.switch_7.Z.n184 0.3805
R261 CDAC8_0.switch_7.Z.n145 CDAC8_0.switch_7.Z.n124 0.3805
R262 CDAC8_0.switch_7.Z.n147 CDAC8_0.switch_7.Z.n126 0.3805
R263 CDAC8_0.switch_7.Z.n149 CDAC8_0.switch_7.Z.n128 0.3805
R264 CDAC8_0.switch_7.Z.n151 CDAC8_0.switch_7.Z.n130 0.3805
R265 CDAC8_0.switch_7.Z.n153 CDAC8_0.switch_7.Z.n132 0.3805
R266 CDAC8_0.switch_7.Z.n156 CDAC8_0.switch_7.Z.n155 0.3805
R267 CDAC8_0.switch_7.Z.n206 CDAC8_0.switch_7.Z.n99 0.3805
R268 CDAC8_0.switch_7.Z.n222 CDAC8_0.switch_7.Z.n221 0.3805
R269 CDAC8_0.switch_7.Z.n225 CDAC8_0.switch_7.Z.n224 0.3805
R270 CDAC8_0.switch_7.Z.n230 CDAC8_0.switch_7.Z.n229 0.3805
R271 CDAC8_0.switch_7.Z.n233 CDAC8_0.switch_7.Z.n232 0.3805
R272 CDAC8_0.switch_7.Z.n196 CDAC8_0.switch_7.Z.n195 0.3805
R273 CDAC8_0.switch_7.Z.n193 CDAC8_0.switch_7.Z.n192 0.3805
R274 CDAC8_0.switch_7.Z.n183 CDAC8_0.switch_7.Z.n182 0.3805
R275 CDAC8_0.switch_7.Z.n180 CDAC8_0.switch_7.Z.n179 0.3805
R276 CDAC8_0.switch_7.Z.n174 CDAC8_0.switch_7.Z.n173 0.3805
R277 CDAC8_0.switch_7.Z.n171 CDAC8_0.switch_7.Z.n170 0.3805
R278 CDAC8_0.switch_7.Z.n166 CDAC8_0.switch_7.Z.n165 0.3805
R279 CDAC8_0.switch_7.Z.n163 CDAC8_0.switch_7.Z.n162 0.3805
R280 CDAC8_0.switch_7.Z.n158 CDAC8_0.switch_7.Z.n157 0.3805
R281 CDAC8_0.switch_7.Z.n217 CDAC8_0.switch_7.Z.n216 0.3805
R282 CDAC8_0.switch_7.Z.n208 CDAC8_0.switch_7.Z.n101 0.3805
R283 CDAC8_0.switch_7.Z.n211 CDAC8_0.switch_7.Z.n210 0.3805
R284 CDAC8_0.switch_7.Z.n214 CDAC8_0.switch_7.Z.n213 0.3805
R285 CDAC8_0.switch_7.Z.n1 CDAC8_0.switch_7.Z 0.259656
R286 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z 0.166261
R287 CDAC8_0.switch_7.Z.n17 CDAC8_0.switch_7.Z.n16 0.162356
R288 CDAC8_0.switch_7.Z.n50 CDAC8_0.switch_7.Z.n49 0.115412
R289 CDAC8_0.switch_7.Z.n51 CDAC8_0.switch_7.Z.n23 0.115412
R290 CDAC8_0.switch_7.Z.n58 CDAC8_0.switch_7.Z.n57 0.115412
R291 CDAC8_0.switch_7.Z.n59 CDAC8_0.switch_7.Z.n19 0.115412
R292 CDAC8_0.switch_7.Z.n67 CDAC8_0.switch_7.Z.n66 0.115412
R293 CDAC8_0.switch_7.Z.n68 CDAC8_0.switch_7.Z.n10 0.115412
R294 CDAC8_0.switch_7.Z.n76 CDAC8_0.switch_7.Z.n75 0.115412
R295 CDAC8_0.switch_7.Z.n78 CDAC8_0.switch_7.Z.n77 0.115412
R296 CDAC8_0.switch_7.Z.n286 CDAC8_0.switch_7.Z.n285 0.115412
R297 CDAC8_0.switch_7.Z.n284 CDAC8_0.switch_7.Z.n79 0.115412
R298 CDAC8_0.switch_7.Z.n278 CDAC8_0.switch_7.Z.n277 0.115412
R299 CDAC8_0.switch_7.Z.n276 CDAC8_0.switch_7.Z.n84 0.115412
R300 CDAC8_0.switch_7.Z.n270 CDAC8_0.switch_7.Z.n269 0.115412
R301 CDAC8_0.switch_7.Z.n268 CDAC8_0.switch_7.Z.n88 0.115412
R302 CDAC8_0.switch_7.Z.n45 CDAC8_0.switch_7.Z.n44 0.115412
R303 CDAC8_0.switch_7.Z.n43 CDAC8_0.switch_7.Z.n42 0.115412
R304 CDAC8_0.switch_7.Z.n41 CDAC8_0.switch_7.Z.n40 0.115412
R305 CDAC8_0.switch_7.Z.n39 CDAC8_0.switch_7.Z.n38 0.115412
R306 CDAC8_0.switch_7.Z.n37 CDAC8_0.switch_7.Z.n11 0.115412
R307 CDAC8_0.switch_7.Z.n72 CDAC8_0.switch_7.Z.n71 0.115412
R308 CDAC8_0.switch_7.Z.n73 CDAC8_0.switch_7.Z.n6 0.115412
R309 CDAC8_0.switch_7.Z.n291 CDAC8_0.switch_7.Z.n290 0.115412
R310 CDAC8_0.switch_7.Z.n289 CDAC8_0.switch_7.Z.n7 0.115412
R311 CDAC8_0.switch_7.Z.n251 CDAC8_0.switch_7.Z.n250 0.115412
R312 CDAC8_0.switch_7.Z.n253 CDAC8_0.switch_7.Z.n252 0.115412
R313 CDAC8_0.switch_7.Z.n255 CDAC8_0.switch_7.Z.n254 0.115412
R314 CDAC8_0.switch_7.Z.n257 CDAC8_0.switch_7.Z.n256 0.115412
R315 CDAC8_0.switch_7.Z.n259 CDAC8_0.switch_7.Z.n258 0.115412
R316 CDAC8_0.switch_7.Z.n47 CDAC8_0.switch_7.Z.n25 0.115412
R317 CDAC8_0.switch_7.Z.n54 CDAC8_0.switch_7.Z.n53 0.115412
R318 CDAC8_0.switch_7.Z.n55 CDAC8_0.switch_7.Z.n21 0.115412
R319 CDAC8_0.switch_7.Z.n62 CDAC8_0.switch_7.Z.n61 0.115412
R320 CDAC8_0.switch_7.Z.n64 CDAC8_0.switch_7.Z.n63 0.115412
R321 CDAC8_0.switch_7.Z.n18 CDAC8_0.switch_7.Z.n17 0.115412
R322 CDAC8_0.switch_7.Z.n15 CDAC8_0.switch_7.Z.n14 0.115412
R323 CDAC8_0.switch_7.Z.n81 CDAC8_0.switch_7.Z.n9 0.115412
R324 CDAC8_0.switch_7.Z.n282 CDAC8_0.switch_7.Z.n281 0.115412
R325 CDAC8_0.switch_7.Z.n280 CDAC8_0.switch_7.Z.n82 0.115412
R326 CDAC8_0.switch_7.Z.n274 CDAC8_0.switch_7.Z.n273 0.115412
R327 CDAC8_0.switch_7.Z.n272 CDAC8_0.switch_7.Z.n86 0.115412
R328 CDAC8_0.switch_7.Z.n266 CDAC8_0.switch_7.Z.n265 0.115412
R329 CDAC8_0.switch_7.Z.n36 CDAC8_0.switch_7.Z.n35 0.115412
R330 CDAC8_0.switch_7.Z.n34 CDAC8_0.switch_7.Z.n33 0.115412
R331 CDAC8_0.switch_7.Z.n32 CDAC8_0.switch_7.Z.n31 0.115412
R332 CDAC8_0.switch_7.Z.n30 CDAC8_0.switch_7.Z.n29 0.115412
R333 CDAC8_0.switch_7.Z.n28 CDAC8_0.switch_7.Z.n27 0.115412
R334 CDAC8_0.switch_7.Z.n13 CDAC8_0.switch_7.Z.n12 0.115412
R335 CDAC8_0.switch_7.Z.n293 CDAC8_0.switch_7.Z.n4 0.115412
R336 CDAC8_0.switch_7.Z.n240 CDAC8_0.switch_7.Z.n239 0.115412
R337 CDAC8_0.switch_7.Z.n242 CDAC8_0.switch_7.Z.n241 0.115412
R338 CDAC8_0.switch_7.Z.n244 CDAC8_0.switch_7.Z.n243 0.115412
R339 CDAC8_0.switch_7.Z.n246 CDAC8_0.switch_7.Z.n245 0.115412
R340 CDAC8_0.switch_7.Z.n248 CDAC8_0.switch_7.Z.n247 0.115412
R341 CDAC8_0.switch_7.Z.n155 CDAC8_0.switch_7.Z.n154 0.115412
R342 CDAC8_0.switch_7.Z.n153 CDAC8_0.switch_7.Z.n152 0.115412
R343 CDAC8_0.switch_7.Z.n151 CDAC8_0.switch_7.Z.n150 0.115412
R344 CDAC8_0.switch_7.Z.n149 CDAC8_0.switch_7.Z.n148 0.115412
R345 CDAC8_0.switch_7.Z.n147 CDAC8_0.switch_7.Z.n146 0.115412
R346 CDAC8_0.switch_7.Z.n145 CDAC8_0.switch_7.Z.n119 0.115412
R347 CDAC8_0.switch_7.Z.n186 CDAC8_0.switch_7.Z.n185 0.115412
R348 CDAC8_0.switch_7.Z.n187 CDAC8_0.switch_7.Z.n103 0.115412
R349 CDAC8_0.switch_7.Z.n199 CDAC8_0.switch_7.Z.n198 0.115412
R350 CDAC8_0.switch_7.Z.n201 CDAC8_0.switch_7.Z.n200 0.115412
R351 CDAC8_0.switch_7.Z.n203 CDAC8_0.switch_7.Z.n202 0.115412
R352 CDAC8_0.switch_7.Z.n205 CDAC8_0.switch_7.Z.n204 0.115412
R353 CDAC8_0.switch_7.Z.n207 CDAC8_0.switch_7.Z.n206 0.115412
R354 CDAC8_0.switch_7.Z.n209 CDAC8_0.switch_7.Z.n208 0.115412
R355 CDAC8_0.switch_7.Z.n157 CDAC8_0.switch_7.Z.n131 0.115412
R356 CDAC8_0.switch_7.Z.n164 CDAC8_0.switch_7.Z.n163 0.115412
R357 CDAC8_0.switch_7.Z.n165 CDAC8_0.switch_7.Z.n127 0.115412
R358 CDAC8_0.switch_7.Z.n172 CDAC8_0.switch_7.Z.n171 0.115412
R359 CDAC8_0.switch_7.Z.n173 CDAC8_0.switch_7.Z.n123 0.115412
R360 CDAC8_0.switch_7.Z.n181 CDAC8_0.switch_7.Z.n180 0.115412
R361 CDAC8_0.switch_7.Z.n182 CDAC8_0.switch_7.Z.n116 0.115412
R362 CDAC8_0.switch_7.Z.n194 CDAC8_0.switch_7.Z.n193 0.115412
R363 CDAC8_0.switch_7.Z.n195 CDAC8_0.switch_7.Z.n93 0.115412
R364 CDAC8_0.switch_7.Z.n232 CDAC8_0.switch_7.Z.n231 0.115412
R365 CDAC8_0.switch_7.Z.n230 CDAC8_0.switch_7.Z.n94 0.115412
R366 CDAC8_0.switch_7.Z.n224 CDAC8_0.switch_7.Z.n223 0.115412
R367 CDAC8_0.switch_7.Z.n222 CDAC8_0.switch_7.Z.n98 0.115412
R368 CDAC8_0.switch_7.Z.n216 CDAC8_0.switch_7.Z.n215 0.115412
R369 CDAC8_0.switch_7.Z.n144 CDAC8_0.switch_7.Z.n143 0.115412
R370 CDAC8_0.switch_7.Z.n142 CDAC8_0.switch_7.Z.n141 0.115412
R371 CDAC8_0.switch_7.Z.n140 CDAC8_0.switch_7.Z.n139 0.115412
R372 CDAC8_0.switch_7.Z.n138 CDAC8_0.switch_7.Z.n137 0.115412
R373 CDAC8_0.switch_7.Z.n136 CDAC8_0.switch_7.Z.n135 0.115412
R374 CDAC8_0.switch_7.Z.n134 CDAC8_0.switch_7.Z.n133 0.115412
R375 CDAC8_0.switch_7.Z.n121 CDAC8_0.switch_7.Z.n120 0.115412
R376 CDAC8_0.switch_7.Z.n118 CDAC8_0.switch_7.Z.n117 0.115412
R377 CDAC8_0.switch_7.Z.n115 CDAC8_0.switch_7.Z.n114 0.115412
R378 CDAC8_0.switch_7.Z.n113 CDAC8_0.switch_7.Z.n112 0.115412
R379 CDAC8_0.switch_7.Z.n111 CDAC8_0.switch_7.Z.n110 0.115412
R380 CDAC8_0.switch_7.Z.n109 CDAC8_0.switch_7.Z.n108 0.115412
R381 CDAC8_0.switch_7.Z.n107 CDAC8_0.switch_7.Z.n106 0.115412
R382 CDAC8_0.switch_7.Z.n105 CDAC8_0.switch_7.Z.n104 0.115412
R383 CDAC8_0.switch_7.Z.n160 CDAC8_0.switch_7.Z.n159 0.115412
R384 CDAC8_0.switch_7.Z.n161 CDAC8_0.switch_7.Z.n129 0.115412
R385 CDAC8_0.switch_7.Z.n168 CDAC8_0.switch_7.Z.n167 0.115412
R386 CDAC8_0.switch_7.Z.n169 CDAC8_0.switch_7.Z.n125 0.115412
R387 CDAC8_0.switch_7.Z.n176 CDAC8_0.switch_7.Z.n175 0.115412
R388 CDAC8_0.switch_7.Z.n178 CDAC8_0.switch_7.Z.n177 0.115412
R389 CDAC8_0.switch_7.Z.n191 CDAC8_0.switch_7.Z.n190 0.115412
R390 CDAC8_0.switch_7.Z.n234 CDAC8_0.switch_7.Z.n91 0.115412
R391 CDAC8_0.switch_7.Z.n228 CDAC8_0.switch_7.Z.n227 0.115412
R392 CDAC8_0.switch_7.Z.n226 CDAC8_0.switch_7.Z.n96 0.115412
R393 CDAC8_0.switch_7.Z.n220 CDAC8_0.switch_7.Z.n219 0.115412
R394 CDAC8_0.switch_7.Z.n218 CDAC8_0.switch_7.Z.n100 0.115412
R395 CDAC8_0.switch_7.Z.n295 CDAC8_0.switch_7.Z.n294 0.0845094
R396 CDAC8_0.switch_7.Z.n238 CDAC8_0.switch_7.Z.n237 0.0845094
R397 CDAC8_0.switch_7.Z.n189 CDAC8_0.switch_7.Z.n2 0.0845094
R398 CDAC8_0.switch_7.Z.n236 CDAC8_0.switch_7.Z.n235 0.0845094
R399 CDAC8_0.switch_7.Z.n51 CDAC8_0.switch_7.Z.n50 0.0474438
R400 CDAC8_0.switch_7.Z.n57 CDAC8_0.switch_7.Z.n23 0.0474438
R401 CDAC8_0.switch_7.Z.n59 CDAC8_0.switch_7.Z.n58 0.0474438
R402 CDAC8_0.switch_7.Z.n66 CDAC8_0.switch_7.Z.n19 0.0474438
R403 CDAC8_0.switch_7.Z.n68 CDAC8_0.switch_7.Z.n67 0.0474438
R404 CDAC8_0.switch_7.Z.n75 CDAC8_0.switch_7.Z.n10 0.0474438
R405 CDAC8_0.switch_7.Z.n77 CDAC8_0.switch_7.Z.n76 0.0474438
R406 CDAC8_0.switch_7.Z.n286 CDAC8_0.switch_7.Z.n78 0.0474438
R407 CDAC8_0.switch_7.Z.n285 CDAC8_0.switch_7.Z.n284 0.0474438
R408 CDAC8_0.switch_7.Z.n278 CDAC8_0.switch_7.Z.n79 0.0474438
R409 CDAC8_0.switch_7.Z.n277 CDAC8_0.switch_7.Z.n276 0.0474438
R410 CDAC8_0.switch_7.Z.n270 CDAC8_0.switch_7.Z.n84 0.0474438
R411 CDAC8_0.switch_7.Z.n269 CDAC8_0.switch_7.Z.n268 0.0474438
R412 CDAC8_0.switch_7.Z.n262 CDAC8_0.switch_7.Z.n88 0.0474438
R413 CDAC8_0.switch_7.Z.n44 CDAC8_0.switch_7.Z.n43 0.0474438
R414 CDAC8_0.switch_7.Z.n42 CDAC8_0.switch_7.Z.n41 0.0474438
R415 CDAC8_0.switch_7.Z.n40 CDAC8_0.switch_7.Z.n39 0.0474438
R416 CDAC8_0.switch_7.Z.n38 CDAC8_0.switch_7.Z.n37 0.0474438
R417 CDAC8_0.switch_7.Z.n71 CDAC8_0.switch_7.Z.n11 0.0474438
R418 CDAC8_0.switch_7.Z.n73 CDAC8_0.switch_7.Z.n72 0.0474438
R419 CDAC8_0.switch_7.Z.n291 CDAC8_0.switch_7.Z.n6 0.0474438
R420 CDAC8_0.switch_7.Z.n290 CDAC8_0.switch_7.Z.n289 0.0474438
R421 CDAC8_0.switch_7.Z.n250 CDAC8_0.switch_7.Z.n7 0.0474438
R422 CDAC8_0.switch_7.Z.n252 CDAC8_0.switch_7.Z.n251 0.0474438
R423 CDAC8_0.switch_7.Z.n254 CDAC8_0.switch_7.Z.n253 0.0474438
R424 CDAC8_0.switch_7.Z.n256 CDAC8_0.switch_7.Z.n255 0.0474438
R425 CDAC8_0.switch_7.Z.n258 CDAC8_0.switch_7.Z.n257 0.0474438
R426 CDAC8_0.switch_7.Z.n260 CDAC8_0.switch_7.Z.n259 0.0474438
R427 CDAC8_0.switch_7.Z.n53 CDAC8_0.switch_7.Z.n25 0.0474438
R428 CDAC8_0.switch_7.Z.n55 CDAC8_0.switch_7.Z.n54 0.0474438
R429 CDAC8_0.switch_7.Z.n61 CDAC8_0.switch_7.Z.n21 0.0474438
R430 CDAC8_0.switch_7.Z.n64 CDAC8_0.switch_7.Z.n62 0.0474438
R431 CDAC8_0.switch_7.Z.n63 CDAC8_0.switch_7.Z.n18 0.0474438
R432 CDAC8_0.switch_7.Z.n16 CDAC8_0.switch_7.Z.n15 0.0474438
R433 CDAC8_0.switch_7.Z.n14 CDAC8_0.switch_7.Z.n9 0.0474438
R434 CDAC8_0.switch_7.Z.n282 CDAC8_0.switch_7.Z.n81 0.0474438
R435 CDAC8_0.switch_7.Z.n281 CDAC8_0.switch_7.Z.n280 0.0474438
R436 CDAC8_0.switch_7.Z.n274 CDAC8_0.switch_7.Z.n82 0.0474438
R437 CDAC8_0.switch_7.Z.n273 CDAC8_0.switch_7.Z.n272 0.0474438
R438 CDAC8_0.switch_7.Z.n266 CDAC8_0.switch_7.Z.n86 0.0474438
R439 CDAC8_0.switch_7.Z.n265 CDAC8_0.switch_7.Z.n264 0.0474438
R440 CDAC8_0.switch_7.Z.n35 CDAC8_0.switch_7.Z.n34 0.0474438
R441 CDAC8_0.switch_7.Z.n33 CDAC8_0.switch_7.Z.n32 0.0474438
R442 CDAC8_0.switch_7.Z.n31 CDAC8_0.switch_7.Z.n30 0.0474438
R443 CDAC8_0.switch_7.Z.n29 CDAC8_0.switch_7.Z.n28 0.0474438
R444 CDAC8_0.switch_7.Z.n27 CDAC8_0.switch_7.Z.n13 0.0474438
R445 CDAC8_0.switch_7.Z.n12 CDAC8_0.switch_7.Z.n3 0.0474438
R446 CDAC8_0.switch_7.Z.n294 CDAC8_0.switch_7.Z.n293 0.0474438
R447 CDAC8_0.switch_7.Z.n8 CDAC8_0.switch_7.Z.n4 0.0474438
R448 CDAC8_0.switch_7.Z.n239 CDAC8_0.switch_7.Z.n238 0.0474438
R449 CDAC8_0.switch_7.Z.n241 CDAC8_0.switch_7.Z.n240 0.0474438
R450 CDAC8_0.switch_7.Z.n243 CDAC8_0.switch_7.Z.n242 0.0474438
R451 CDAC8_0.switch_7.Z.n245 CDAC8_0.switch_7.Z.n244 0.0474438
R452 CDAC8_0.switch_7.Z.n247 CDAC8_0.switch_7.Z.n246 0.0474438
R453 CDAC8_0.switch_7.Z.n249 CDAC8_0.switch_7.Z.n248 0.0474438
R454 CDAC8_0.switch_7.Z.n154 CDAC8_0.switch_7.Z.n153 0.0474438
R455 CDAC8_0.switch_7.Z.n152 CDAC8_0.switch_7.Z.n151 0.0474438
R456 CDAC8_0.switch_7.Z.n150 CDAC8_0.switch_7.Z.n149 0.0474438
R457 CDAC8_0.switch_7.Z.n148 CDAC8_0.switch_7.Z.n147 0.0474438
R458 CDAC8_0.switch_7.Z.n146 CDAC8_0.switch_7.Z.n145 0.0474438
R459 CDAC8_0.switch_7.Z.n185 CDAC8_0.switch_7.Z.n119 0.0474438
R460 CDAC8_0.switch_7.Z.n187 CDAC8_0.switch_7.Z.n186 0.0474438
R461 CDAC8_0.switch_7.Z.n198 CDAC8_0.switch_7.Z.n103 0.0474438
R462 CDAC8_0.switch_7.Z.n200 CDAC8_0.switch_7.Z.n199 0.0474438
R463 CDAC8_0.switch_7.Z.n202 CDAC8_0.switch_7.Z.n201 0.0474438
R464 CDAC8_0.switch_7.Z.n204 CDAC8_0.switch_7.Z.n203 0.0474438
R465 CDAC8_0.switch_7.Z.n206 CDAC8_0.switch_7.Z.n205 0.0474438
R466 CDAC8_0.switch_7.Z.n208 CDAC8_0.switch_7.Z.n207 0.0474438
R467 CDAC8_0.switch_7.Z.n210 CDAC8_0.switch_7.Z.n209 0.0474438
R468 CDAC8_0.switch_7.Z.n163 CDAC8_0.switch_7.Z.n131 0.0474438
R469 CDAC8_0.switch_7.Z.n165 CDAC8_0.switch_7.Z.n164 0.0474438
R470 CDAC8_0.switch_7.Z.n171 CDAC8_0.switch_7.Z.n127 0.0474438
R471 CDAC8_0.switch_7.Z.n173 CDAC8_0.switch_7.Z.n172 0.0474438
R472 CDAC8_0.switch_7.Z.n180 CDAC8_0.switch_7.Z.n123 0.0474438
R473 CDAC8_0.switch_7.Z.n182 CDAC8_0.switch_7.Z.n181 0.0474438
R474 CDAC8_0.switch_7.Z.n193 CDAC8_0.switch_7.Z.n116 0.0474438
R475 CDAC8_0.switch_7.Z.n195 CDAC8_0.switch_7.Z.n194 0.0474438
R476 CDAC8_0.switch_7.Z.n232 CDAC8_0.switch_7.Z.n93 0.0474438
R477 CDAC8_0.switch_7.Z.n231 CDAC8_0.switch_7.Z.n230 0.0474438
R478 CDAC8_0.switch_7.Z.n224 CDAC8_0.switch_7.Z.n94 0.0474438
R479 CDAC8_0.switch_7.Z.n223 CDAC8_0.switch_7.Z.n222 0.0474438
R480 CDAC8_0.switch_7.Z.n216 CDAC8_0.switch_7.Z.n98 0.0474438
R481 CDAC8_0.switch_7.Z.n215 CDAC8_0.switch_7.Z.n214 0.0474438
R482 CDAC8_0.switch_7.Z.n143 CDAC8_0.switch_7.Z.n142 0.0474438
R483 CDAC8_0.switch_7.Z.n141 CDAC8_0.switch_7.Z.n140 0.0474438
R484 CDAC8_0.switch_7.Z.n139 CDAC8_0.switch_7.Z.n138 0.0474438
R485 CDAC8_0.switch_7.Z.n137 CDAC8_0.switch_7.Z.n136 0.0474438
R486 CDAC8_0.switch_7.Z.n135 CDAC8_0.switch_7.Z.n134 0.0474438
R487 CDAC8_0.switch_7.Z.n133 CDAC8_0.switch_7.Z.n121 0.0474438
R488 CDAC8_0.switch_7.Z.n120 CDAC8_0.switch_7.Z.n118 0.0474438
R489 CDAC8_0.switch_7.Z.n117 CDAC8_0.switch_7.Z.n115 0.0474438
R490 CDAC8_0.switch_7.Z.n114 CDAC8_0.switch_7.Z.n113 0.0474438
R491 CDAC8_0.switch_7.Z.n112 CDAC8_0.switch_7.Z.n111 0.0474438
R492 CDAC8_0.switch_7.Z.n110 CDAC8_0.switch_7.Z.n109 0.0474438
R493 CDAC8_0.switch_7.Z.n108 CDAC8_0.switch_7.Z.n107 0.0474438
R494 CDAC8_0.switch_7.Z.n106 CDAC8_0.switch_7.Z.n105 0.0474438
R495 CDAC8_0.switch_7.Z.n104 CDAC8_0.switch_7.Z.n102 0.0474438
R496 CDAC8_0.switch_7.Z.n161 CDAC8_0.switch_7.Z.n160 0.0474438
R497 CDAC8_0.switch_7.Z.n167 CDAC8_0.switch_7.Z.n129 0.0474438
R498 CDAC8_0.switch_7.Z.n169 CDAC8_0.switch_7.Z.n168 0.0474438
R499 CDAC8_0.switch_7.Z.n175 CDAC8_0.switch_7.Z.n125 0.0474438
R500 CDAC8_0.switch_7.Z.n178 CDAC8_0.switch_7.Z.n176 0.0474438
R501 CDAC8_0.switch_7.Z.n177 CDAC8_0.switch_7.Z.n122 0.0474438
R502 CDAC8_0.switch_7.Z.n191 CDAC8_0.switch_7.Z.n189 0.0474438
R503 CDAC8_0.switch_7.Z.n190 CDAC8_0.switch_7.Z.n90 0.0474438
R504 CDAC8_0.switch_7.Z.n235 CDAC8_0.switch_7.Z.n234 0.0474438
R505 CDAC8_0.switch_7.Z.n228 CDAC8_0.switch_7.Z.n91 0.0474438
R506 CDAC8_0.switch_7.Z.n227 CDAC8_0.switch_7.Z.n226 0.0474438
R507 CDAC8_0.switch_7.Z.n220 CDAC8_0.switch_7.Z.n96 0.0474438
R508 CDAC8_0.switch_7.Z.n219 CDAC8_0.switch_7.Z.n218 0.0474438
R509 CDAC8_0.switch_7.Z.n212 CDAC8_0.switch_7.Z.n100 0.0474438
R510 CDAC8_0.switch_7.Z CDAC8_0.switch_7.Z.n297 0.0454219
R511 CDAC8_0.switch_7.Z.n295 CDAC8_0.switch_7.Z.n3 0.0314031
R512 CDAC8_0.switch_7.Z.n237 CDAC8_0.switch_7.Z.n8 0.0314031
R513 CDAC8_0.switch_7.Z.n122 CDAC8_0.switch_7.Z.n2 0.0314031
R514 CDAC8_0.switch_7.Z.n236 CDAC8_0.switch_7.Z.n90 0.0314031
R515 CDAC8_0.switch_7.Z.n1 CDAC8_0.switch_7.Z.n0 0.0188121
R516 EN.n61 EN.t56 158.988
R517 EN.n155 EN.t42 158.988
R518 EN EN.t13 158.581
R519 EN EN.t21 158.581
R520 EN EN.t88 158.581
R521 EN EN.t77 158.581
R522 EN EN.t9 158.581
R523 EN EN.t96 158.581
R524 EN EN.t36 158.581
R525 EN EN.t60 158.581
R526 EN EN.t35 158.581
R527 EN EN.t76 158.581
R528 EN EN.t39 158.581
R529 EN EN.t81 158.581
R530 EN EN.t79 158.581
R531 EN EN.t37 158.581
R532 EN EN.t40 158.581
R533 EN EN.t98 158.581
R534 EN.n69 EN.t6 150.293
R535 EN.n63 EN.t61 150.293
R536 EN.n145 EN.t10 150.293
R537 EN.n139 EN.t12 150.293
R538 EN.t13 EN.n181 150.293
R539 EN.t21 EN.n212 150.293
R540 EN.t88 EN.n221 150.293
R541 EN.t77 EN.n135 150.293
R542 EN.t9 EN.n244 150.293
R543 EN.t96 EN.n274 150.293
R544 EN.t36 EN.n284 150.293
R545 EN.t60 EN.n97 150.293
R546 EN.t35 EN.n106 150.293
R547 EN.t76 EN.n318 150.293
R548 EN.t39 EN.n327 150.293
R549 EN.t81 EN.n33 150.293
R550 EN.t79 EN.n350 150.293
R551 EN.t37 EN.n163 150.293
R552 EN.t40 EN.n52 150.293
R553 EN.t98 EN.n5 150.293
R554 EN.t56 EN.n60 150.273
R555 EN.t42 EN.n154 150.273
R556 EN.n186 EN.t50 150.273
R557 EN.n176 EN.t94 150.273
R558 EN.n205 EN.t71 150.273
R559 EN.n199 EN.t104 150.273
R560 EN.n226 EN.t23 150.273
R561 EN.n216 EN.t15 150.273
R562 EN.n128 EN.t89 150.273
R563 EN.n122 EN.t25 150.273
R564 EN.n249 EN.t47 150.273
R565 EN.n239 EN.t72 150.273
R566 EN.n267 EN.t46 150.273
R567 EN.n261 EN.t80 150.273
R568 EN.n289 EN.t97 150.273
R569 EN.n279 EN.t90 150.273
R570 EN.n90 EN.t66 150.273
R571 EN.n84 EN.t45 150.273
R572 EN.n111 EN.t18 150.273
R573 EN.n101 EN.t11 150.273
R574 EN.n311 EN.t17 150.273
R575 EN.n305 EN.t55 150.273
R576 EN.n332 EN.t92 150.273
R577 EN.n322 EN.t67 150.273
R578 EN.n26 EN.t29 150.273
R579 EN.n20 EN.t106 150.273
R580 EN.n355 EN.t14 150.273
R581 EN.n345 EN.t75 150.273
R582 EN.n168 EN.t101 150.273
R583 EN.n158 EN.t93 150.273
R584 EN.n45 EN.t49 150.273
R585 EN.n39 EN.t26 150.273
R586 EN.n10 EN.t38 150.273
R587 EN.n0 EN.t16 150.273
R588 EN.n194 EN.t1 115.191
R589 EN.n234 EN.t91 81.8568
R590 EN.n257 EN.t48 81.8568
R591 EN.n297 EN.t69 81.8568
R592 EN.n300 EN.t19 81.8568
R593 EN.n340 EN.t44 81.8568
R594 EN.n363 EN.t53 81.8568
R595 EN.n195 EN.t73 81.8568
R596 EN.t105 EN.n365 81.8568
R597 EN.n58 EN.t41 73.6406
R598 EN.n152 EN.t20 73.6406
R599 EN.n184 EN.t57 73.6406
R600 EN.t1 EN.n193 73.6406
R601 EN.n203 EN.t58 73.6406
R602 EN.n197 EN.t85 73.6406
R603 EN.n224 EN.t28 73.6406
R604 EN.t91 EN.n233 73.6406
R605 EN.n126 EN.t0 73.6406
R606 EN.n120 EN.t4 73.6406
R607 EN.n247 EN.t82 73.6406
R608 EN.t48 EN.n256 73.6406
R609 EN.n265 EN.t31 73.6406
R610 EN.n259 EN.t63 73.6406
R611 EN.n287 EN.t99 73.6406
R612 EN.t69 EN.n296 73.6406
R613 EN.n88 EN.t83 73.6406
R614 EN.n82 EN.t27 73.6406
R615 EN.n109 EN.t22 73.6406
R616 EN.t19 EN.n118 73.6406
R617 EN.n309 EN.t100 73.6406
R618 EN.n303 EN.t68 73.6406
R619 EN.n330 EN.t78 73.6406
R620 EN.t44 EN.n339 73.6406
R621 EN.n24 EN.t8 73.6406
R622 EN.n18 EN.t86 73.6406
R623 EN.n353 EN.t30 73.6406
R624 EN.t53 EN.n362 73.6406
R625 EN.n166 EN.t107 73.6406
R626 EN.t73 EN.n175 73.6406
R627 EN.n43 EN.t64 73.6406
R628 EN.n37 EN.t7 73.6406
R629 EN.n8 EN.t74 73.6406
R630 EN.n366 EN.t105 73.6406
R631 EN.n71 EN.t43 73.6304
R632 EN.n65 EN.t87 73.6304
R633 EN.n147 EN.t62 73.6304
R634 EN.n141 EN.t95 73.6304
R635 EN.n179 EN.t59 73.6304
R636 EN.n210 EN.t2 73.6304
R637 EN.n219 EN.t33 73.6304
R638 EN.n133 EN.t32 73.6304
R639 EN.n242 EN.t52 73.6304
R640 EN.n272 EN.t51 73.6304
R641 EN.n282 EN.t103 73.6304
R642 EN.n95 EN.t102 73.6304
R643 EN.n104 EN.t70 73.6304
R644 EN.n316 EN.t24 73.6304
R645 EN.n325 EN.t5 73.6304
R646 EN.n31 EN.t65 73.6304
R647 EN.n348 EN.t34 73.6304
R648 EN.n161 EN.t3 73.6304
R649 EN.n50 EN.t84 73.6304
R650 EN.n3 EN.t54 73.6304
R651 EN.n365 EN.n364 33.3344
R652 EN.n236 EN.n196 33.3344
R653 EN.n343 EN.n80 33.3344
R654 EN.n364 EN.n17 29.9244
R655 EN.n299 EN.n17 29.9244
R656 EN.n299 EN.n298 29.9244
R657 EN.n298 EN.n258 29.9244
R658 EN.n258 EN.n119 29.9244
R659 EN.n194 EN.n119 29.9244
R660 EN.n237 EN.n236 29.9244
R661 EN.n237 EN.n81 29.9244
R662 EN.n302 EN.n81 29.9244
R663 EN.n342 EN.n302 29.9244
R664 EN.n343 EN.n342 29.9244
R665 EN.n235 EN.n234 25.7228
R666 EN.n257 EN.n238 25.7228
R667 EN.n297 EN.n278 25.7228
R668 EN.n301 EN.n300 25.7228
R669 EN.n341 EN.n340 25.7228
R670 EN.n363 EN.n344 25.7228
R671 EN.n196 EN.n195 25.7228
R672 EN.n79 EN 23.3453
R673 EN.n77 EN.n76 20.9244
R674 EN.n75 EN.n68 15.5222
R675 EN.n151 EN.n144 15.5222
R676 EN.n191 EN.n190 15.5222
R677 EN.n209 EN.n202 15.5222
R678 EN.n231 EN.n230 15.5222
R679 EN.n132 EN.n125 15.5222
R680 EN.n254 EN.n253 15.5222
R681 EN.n271 EN.n264 15.5222
R682 EN.n294 EN.n293 15.5222
R683 EN.n94 EN.n87 15.5222
R684 EN.n116 EN.n115 15.5222
R685 EN.n315 EN.n308 15.5222
R686 EN.n337 EN.n336 15.5222
R687 EN.n30 EN.n23 15.5222
R688 EN.n360 EN.n359 15.5222
R689 EN.n173 EN.n172 15.5222
R690 EN.n49 EN.n42 15.5222
R691 EN.n15 EN.n14 15.5222
R692 EN.n78 EN 12.9568
R693 EN.n57 EN.n56 12.8934
R694 EN.n79 EN.n78 12.7234
R695 EN.n57 EN 10.1822
R696 EN.n190 EN.n183 8.26552
R697 EN.n230 EN.n223 8.26552
R698 EN.n253 EN.n246 8.26552
R699 EN.n293 EN.n286 8.26552
R700 EN.n115 EN.n108 8.26552
R701 EN.n336 EN.n329 8.26552
R702 EN.n359 EN.n352 8.26552
R703 EN.n172 EN.n165 8.26552
R704 EN.n14 EN.n7 8.26552
R705 EN.n76 EN.n75 7.83713
R706 EN.n235 EN.n215 5.58033
R707 EN.n238 EN.n138 5.58033
R708 EN.n278 EN.n277 5.58033
R709 EN.n301 EN.n100 5.58033
R710 EN.n341 EN.n321 5.58033
R711 EN.n344 EN.n36 5.58033
R712 EN.n80 EN.n55 5.58033
R713 EN.n75 EN.n74 4.5005
R714 EN.n151 EN.n150 4.5005
R715 EN.n190 EN.n189 4.5005
R716 EN.n209 EN.n208 4.5005
R717 EN.n230 EN.n229 4.5005
R718 EN.n132 EN.n131 4.5005
R719 EN.n253 EN.n252 4.5005
R720 EN.n271 EN.n270 4.5005
R721 EN.n293 EN.n292 4.5005
R722 EN.n94 EN.n93 4.5005
R723 EN.n115 EN.n114 4.5005
R724 EN.n315 EN.n314 4.5005
R725 EN.n336 EN.n335 4.5005
R726 EN.n30 EN.n29 4.5005
R727 EN.n359 EN.n358 4.5005
R728 EN.n172 EN.n171 4.5005
R729 EN.n49 EN.n48 4.5005
R730 EN.n14 EN.n13 4.5005
R731 EN.n196 EN.n157 4.31133
R732 EN.n215 EN.n214 4.20846
R733 EN.n138 EN.n137 4.20846
R734 EN.n277 EN.n276 4.20846
R735 EN.n100 EN.n99 4.20846
R736 EN.n321 EN.n320 4.20846
R737 EN.n36 EN.n35 4.20846
R738 EN.n55 EN.n54 4.20846
R739 EN.n157 EN.n151 3.98148
R740 EN.n215 EN.n209 3.98148
R741 EN.n138 EN.n132 3.98148
R742 EN.n277 EN.n271 3.98148
R743 EN.n100 EN.n94 3.98148
R744 EN.n321 EN.n315 3.98148
R745 EN.n36 EN.n30 3.98148
R746 EN.n55 EN.n49 3.98148
R747 EN.n157 EN 3.8
R748 EN.n364 EN.n363 3.4105
R749 EN.n340 EN.n17 3.4105
R750 EN.n300 EN.n299 3.4105
R751 EN.n298 EN.n297 3.4105
R752 EN.n258 EN.n257 3.4105
R753 EN.n234 EN.n119 3.4105
R754 EN.n195 EN.n194 3.4105
R755 EN.n236 EN.n235 3.4105
R756 EN.n238 EN.n237 3.4105
R757 EN.n278 EN.n81 3.4105
R758 EN.n302 EN.n301 3.4105
R759 EN.n342 EN.n341 3.4105
R760 EN.n344 EN.n343 3.4105
R761 EN.n59 EN.n58 1.19615
R762 EN.n153 EN.n152 1.19615
R763 EN.n181 EN.n180 1.19615
R764 EN.n212 EN.n211 1.19615
R765 EN.n221 EN.n220 1.19615
R766 EN.n135 EN.n134 1.19615
R767 EN.n244 EN.n243 1.19615
R768 EN.n274 EN.n273 1.19615
R769 EN.n284 EN.n283 1.19615
R770 EN.n97 EN.n96 1.19615
R771 EN.n106 EN.n105 1.19615
R772 EN.n318 EN.n317 1.19615
R773 EN.n327 EN.n326 1.19615
R774 EN.n33 EN.n32 1.19615
R775 EN.n350 EN.n349 1.19615
R776 EN.n163 EN.n162 1.19615
R777 EN.n52 EN.n51 1.19615
R778 EN.n5 EN.n4 1.19615
R779 EN.n70 EN 1.09561
R780 EN.n64 EN 1.09561
R781 EN.n146 EN 1.09561
R782 EN.n140 EN 1.09561
R783 EN.n73 EN.n72 0.796696
R784 EN.n67 EN.n66 0.796696
R785 EN.n149 EN.n148 0.796696
R786 EN.n143 EN.n142 0.796696
R787 EN.n185 EN.n184 0.796696
R788 EN.n193 EN.n192 0.796696
R789 EN.n204 EN.n203 0.796696
R790 EN.n198 EN.n197 0.796696
R791 EN.n225 EN.n224 0.796696
R792 EN.n233 EN.n232 0.796696
R793 EN.n127 EN.n126 0.796696
R794 EN.n121 EN.n120 0.796696
R795 EN.n248 EN.n247 0.796696
R796 EN.n256 EN.n255 0.796696
R797 EN.n266 EN.n265 0.796696
R798 EN.n260 EN.n259 0.796696
R799 EN.n288 EN.n287 0.796696
R800 EN.n296 EN.n295 0.796696
R801 EN.n89 EN.n88 0.796696
R802 EN.n83 EN.n82 0.796696
R803 EN.n110 EN.n109 0.796696
R804 EN.n118 EN.n117 0.796696
R805 EN.n310 EN.n309 0.796696
R806 EN.n304 EN.n303 0.796696
R807 EN.n331 EN.n330 0.796696
R808 EN.n339 EN.n338 0.796696
R809 EN.n25 EN.n24 0.796696
R810 EN.n19 EN.n18 0.796696
R811 EN.n354 EN.n353 0.796696
R812 EN.n362 EN.n361 0.796696
R813 EN.n167 EN.n166 0.796696
R814 EN.n175 EN.n174 0.796696
R815 EN.n44 EN.n43 0.796696
R816 EN.n38 EN.n37 0.796696
R817 EN.n9 EN.n8 0.796696
R818 EN.n366 EN.n16 0.796696
R819 EN.n62 EN.n61 0.783833
R820 EN.n156 EN.n155 0.783833
R821 EN.n183 EN.n182 0.783833
R822 EN.n214 EN.n213 0.783833
R823 EN.n223 EN.n222 0.783833
R824 EN.n137 EN.n136 0.783833
R825 EN.n246 EN.n245 0.783833
R826 EN.n276 EN.n275 0.783833
R827 EN.n286 EN.n285 0.783833
R828 EN.n99 EN.n98 0.783833
R829 EN.n108 EN.n107 0.783833
R830 EN.n320 EN.n319 0.783833
R831 EN.n329 EN.n328 0.783833
R832 EN.n35 EN.n34 0.783833
R833 EN.n352 EN.n351 0.783833
R834 EN.n165 EN.n164 0.783833
R835 EN.n54 EN.n53 0.783833
R836 EN.n7 EN.n6 0.783833
R837 EN.n61 EN 0.716182
R838 EN.n155 EN 0.716182
R839 EN.n183 EN 0.716182
R840 EN.n214 EN 0.716182
R841 EN.n223 EN 0.716182
R842 EN.n137 EN 0.716182
R843 EN.n246 EN 0.716182
R844 EN.n276 EN 0.716182
R845 EN.n286 EN 0.716182
R846 EN.n99 EN 0.716182
R847 EN.n108 EN 0.716182
R848 EN.n320 EN 0.716182
R849 EN.n329 EN 0.716182
R850 EN.n35 EN 0.716182
R851 EN.n352 EN 0.716182
R852 EN.n165 EN 0.716182
R853 EN.n54 EN 0.716182
R854 EN.n7 EN 0.716182
R855 EN.n73 EN 0.662609
R856 EN.n67 EN 0.662609
R857 EN.n149 EN 0.662609
R858 EN.n143 EN 0.662609
R859 EN.n185 EN 0.524957
R860 EN.n192 EN 0.524957
R861 EN.n204 EN 0.524957
R862 EN.n198 EN 0.524957
R863 EN.n225 EN 0.524957
R864 EN.n232 EN 0.524957
R865 EN.n127 EN 0.524957
R866 EN.n121 EN 0.524957
R867 EN.n248 EN 0.524957
R868 EN.n255 EN 0.524957
R869 EN.n266 EN 0.524957
R870 EN.n260 EN 0.524957
R871 EN.n288 EN 0.524957
R872 EN.n295 EN 0.524957
R873 EN.n89 EN 0.524957
R874 EN.n83 EN 0.524957
R875 EN.n110 EN 0.524957
R876 EN.n117 EN 0.524957
R877 EN.n310 EN 0.524957
R878 EN.n304 EN 0.524957
R879 EN.n331 EN 0.524957
R880 EN.n338 EN 0.524957
R881 EN.n25 EN 0.524957
R882 EN.n19 EN 0.524957
R883 EN.n354 EN 0.524957
R884 EN.n361 EN 0.524957
R885 EN.n167 EN 0.524957
R886 EN.n174 EN 0.524957
R887 EN.n44 EN 0.524957
R888 EN.n38 EN 0.524957
R889 EN.n9 EN 0.524957
R890 EN.n16 EN 0.524957
R891 EN.n69 EN 0.447191
R892 EN.n63 EN 0.447191
R893 EN.n145 EN 0.447191
R894 EN.n139 EN 0.447191
R895 EN.n181 EN 0.447191
R896 EN.n212 EN 0.447191
R897 EN.n221 EN 0.447191
R898 EN.n135 EN 0.447191
R899 EN.n244 EN 0.447191
R900 EN.n274 EN 0.447191
R901 EN.n284 EN 0.447191
R902 EN.n97 EN 0.447191
R903 EN.n106 EN 0.447191
R904 EN.n318 EN 0.447191
R905 EN.n327 EN 0.447191
R906 EN.n33 EN 0.447191
R907 EN.n350 EN 0.447191
R908 EN.n163 EN 0.447191
R909 EN.n52 EN 0.447191
R910 EN.n5 EN 0.447191
R911 EN.n188 EN 0.252453
R912 EN.n178 EN 0.252453
R913 EN.n207 EN 0.252453
R914 EN.n201 EN 0.252453
R915 EN.n228 EN 0.252453
R916 EN.n218 EN 0.252453
R917 EN.n130 EN 0.252453
R918 EN.n124 EN 0.252453
R919 EN.n251 EN 0.252453
R920 EN.n241 EN 0.252453
R921 EN.n269 EN 0.252453
R922 EN.n263 EN 0.252453
R923 EN.n291 EN 0.252453
R924 EN.n281 EN 0.252453
R925 EN.n92 EN 0.252453
R926 EN.n86 EN 0.252453
R927 EN.n113 EN 0.252453
R928 EN.n103 EN 0.252453
R929 EN.n313 EN 0.252453
R930 EN.n307 EN 0.252453
R931 EN.n334 EN 0.252453
R932 EN.n324 EN 0.252453
R933 EN.n28 EN 0.252453
R934 EN.n22 EN 0.252453
R935 EN.n357 EN 0.252453
R936 EN.n347 EN 0.252453
R937 EN.n170 EN 0.252453
R938 EN.n160 EN 0.252453
R939 EN.n47 EN 0.252453
R940 EN.n41 EN 0.252453
R941 EN.n12 EN 0.252453
R942 EN.n2 EN 0.252453
R943 EN.n70 EN.n69 0.226043
R944 EN.n64 EN.n63 0.226043
R945 EN.n146 EN.n145 0.226043
R946 EN.n140 EN.n139 0.226043
R947 EN.n188 EN.n187 0.226043
R948 EN.n178 EN.n177 0.226043
R949 EN.n207 EN.n206 0.226043
R950 EN.n201 EN.n200 0.226043
R951 EN.n228 EN.n227 0.226043
R952 EN.n218 EN.n217 0.226043
R953 EN.n130 EN.n129 0.226043
R954 EN.n124 EN.n123 0.226043
R955 EN.n251 EN.n250 0.226043
R956 EN.n241 EN.n240 0.226043
R957 EN.n269 EN.n268 0.226043
R958 EN.n263 EN.n262 0.226043
R959 EN.n291 EN.n290 0.226043
R960 EN.n281 EN.n280 0.226043
R961 EN.n92 EN.n91 0.226043
R962 EN.n86 EN.n85 0.226043
R963 EN.n113 EN.n112 0.226043
R964 EN.n103 EN.n102 0.226043
R965 EN.n313 EN.n312 0.226043
R966 EN.n307 EN.n306 0.226043
R967 EN.n334 EN.n333 0.226043
R968 EN.n324 EN.n323 0.226043
R969 EN.n28 EN.n27 0.226043
R970 EN.n22 EN.n21 0.226043
R971 EN.n357 EN.n356 0.226043
R972 EN.n347 EN.n346 0.226043
R973 EN.n170 EN.n169 0.226043
R974 EN.n160 EN.n159 0.226043
R975 EN.n47 EN.n46 0.226043
R976 EN.n41 EN.n40 0.226043
R977 EN.n12 EN.n11 0.226043
R978 EN.n2 EN.n1 0.226043
R979 EN.n58 EN 0.217464
R980 EN.n152 EN 0.217464
R981 EN.n184 EN 0.217464
R982 EN.n193 EN 0.217464
R983 EN.n203 EN 0.217464
R984 EN.n197 EN 0.217464
R985 EN.n224 EN 0.217464
R986 EN.n233 EN 0.217464
R987 EN.n126 EN 0.217464
R988 EN.n120 EN 0.217464
R989 EN.n247 EN 0.217464
R990 EN.n256 EN 0.217464
R991 EN.n265 EN 0.217464
R992 EN.n259 EN 0.217464
R993 EN.n287 EN 0.217464
R994 EN.n296 EN 0.217464
R995 EN.n88 EN 0.217464
R996 EN.n82 EN 0.217464
R997 EN.n109 EN 0.217464
R998 EN.n118 EN 0.217464
R999 EN.n309 EN 0.217464
R1000 EN.n303 EN 0.217464
R1001 EN.n330 EN 0.217464
R1002 EN.n339 EN 0.217464
R1003 EN.n24 EN 0.217464
R1004 EN.n18 EN 0.217464
R1005 EN.n353 EN 0.217464
R1006 EN.n362 EN 0.217464
R1007 EN.n166 EN 0.217464
R1008 EN.n175 EN 0.217464
R1009 EN.n43 EN 0.217464
R1010 EN.n37 EN 0.217464
R1011 EN.n8 EN 0.217464
R1012 EN EN.n366 0.217464
R1013 EN.n72 EN 0.1255
R1014 EN.n66 EN 0.1255
R1015 EN.n59 EN 0.1255
R1016 EN.n153 EN 0.1255
R1017 EN.n148 EN 0.1255
R1018 EN.n142 EN 0.1255
R1019 EN.n187 EN 0.1255
R1020 EN.n180 EN 0.1255
R1021 EN.n177 EN 0.1255
R1022 EN.n211 EN 0.1255
R1023 EN.n206 EN 0.1255
R1024 EN.n200 EN 0.1255
R1025 EN.n227 EN 0.1255
R1026 EN.n220 EN 0.1255
R1027 EN.n217 EN 0.1255
R1028 EN.n134 EN 0.1255
R1029 EN.n129 EN 0.1255
R1030 EN.n123 EN 0.1255
R1031 EN.n250 EN 0.1255
R1032 EN.n243 EN 0.1255
R1033 EN.n240 EN 0.1255
R1034 EN.n273 EN 0.1255
R1035 EN.n268 EN 0.1255
R1036 EN.n262 EN 0.1255
R1037 EN.n290 EN 0.1255
R1038 EN.n283 EN 0.1255
R1039 EN.n280 EN 0.1255
R1040 EN.n96 EN 0.1255
R1041 EN.n91 EN 0.1255
R1042 EN.n85 EN 0.1255
R1043 EN.n112 EN 0.1255
R1044 EN.n105 EN 0.1255
R1045 EN.n102 EN 0.1255
R1046 EN.n317 EN 0.1255
R1047 EN.n312 EN 0.1255
R1048 EN.n306 EN 0.1255
R1049 EN.n333 EN 0.1255
R1050 EN.n326 EN 0.1255
R1051 EN.n323 EN 0.1255
R1052 EN.n32 EN 0.1255
R1053 EN.n27 EN 0.1255
R1054 EN.n21 EN 0.1255
R1055 EN.n356 EN 0.1255
R1056 EN.n349 EN 0.1255
R1057 EN.n346 EN 0.1255
R1058 EN.n169 EN 0.1255
R1059 EN.n162 EN 0.1255
R1060 EN.n159 EN 0.1255
R1061 EN.n51 EN 0.1255
R1062 EN.n46 EN 0.1255
R1063 EN.n40 EN 0.1255
R1064 EN.n11 EN 0.1255
R1065 EN.n4 EN 0.1255
R1066 EN.n1 EN 0.1255
R1067 EN.n74 EN.n70 0.063
R1068 EN.n74 EN.n73 0.063
R1069 EN.n68 EN.n64 0.063
R1070 EN.n68 EN.n67 0.063
R1071 EN.n150 EN.n146 0.063
R1072 EN.n150 EN.n149 0.063
R1073 EN.n144 EN.n140 0.063
R1074 EN.n144 EN.n143 0.063
R1075 EN.n189 EN.n185 0.063
R1076 EN.n189 EN.n188 0.063
R1077 EN.n192 EN.n191 0.063
R1078 EN.n191 EN.n178 0.063
R1079 EN.n208 EN.n204 0.063
R1080 EN.n208 EN.n207 0.063
R1081 EN.n202 EN.n198 0.063
R1082 EN.n202 EN.n201 0.063
R1083 EN.n229 EN.n225 0.063
R1084 EN.n229 EN.n228 0.063
R1085 EN.n232 EN.n231 0.063
R1086 EN.n231 EN.n218 0.063
R1087 EN.n131 EN.n127 0.063
R1088 EN.n131 EN.n130 0.063
R1089 EN.n125 EN.n121 0.063
R1090 EN.n125 EN.n124 0.063
R1091 EN.n252 EN.n248 0.063
R1092 EN.n252 EN.n251 0.063
R1093 EN.n255 EN.n254 0.063
R1094 EN.n254 EN.n241 0.063
R1095 EN.n270 EN.n266 0.063
R1096 EN.n270 EN.n269 0.063
R1097 EN.n264 EN.n260 0.063
R1098 EN.n264 EN.n263 0.063
R1099 EN.n292 EN.n288 0.063
R1100 EN.n292 EN.n291 0.063
R1101 EN.n295 EN.n294 0.063
R1102 EN.n294 EN.n281 0.063
R1103 EN.n93 EN.n89 0.063
R1104 EN.n93 EN.n92 0.063
R1105 EN.n87 EN.n83 0.063
R1106 EN.n87 EN.n86 0.063
R1107 EN.n114 EN.n110 0.063
R1108 EN.n114 EN.n113 0.063
R1109 EN.n117 EN.n116 0.063
R1110 EN.n116 EN.n103 0.063
R1111 EN.n314 EN.n310 0.063
R1112 EN.n314 EN.n313 0.063
R1113 EN.n308 EN.n304 0.063
R1114 EN.n308 EN.n307 0.063
R1115 EN.n335 EN.n331 0.063
R1116 EN.n335 EN.n334 0.063
R1117 EN.n338 EN.n337 0.063
R1118 EN.n337 EN.n324 0.063
R1119 EN.n29 EN.n25 0.063
R1120 EN.n29 EN.n28 0.063
R1121 EN.n23 EN.n19 0.063
R1122 EN.n23 EN.n22 0.063
R1123 EN.n358 EN.n354 0.063
R1124 EN.n358 EN.n357 0.063
R1125 EN.n361 EN.n360 0.063
R1126 EN.n360 EN.n347 0.063
R1127 EN.n171 EN.n167 0.063
R1128 EN.n171 EN.n170 0.063
R1129 EN.n174 EN.n173 0.063
R1130 EN.n173 EN.n160 0.063
R1131 EN.n48 EN.n44 0.063
R1132 EN.n48 EN.n47 0.063
R1133 EN.n42 EN.n38 0.063
R1134 EN.n42 EN.n41 0.063
R1135 EN.n13 EN.n9 0.063
R1136 EN.n13 EN.n12 0.063
R1137 EN.n16 EN.n15 0.063
R1138 EN.n15 EN.n2 0.063
R1139 EN.n80 EN.n79 0.024
R1140 EN.n78 EN.n77 0.024
R1141 EN.n77 EN.n57 0.024
R1142 EN.n60 EN.n59 0.0216397
R1143 EN.n60 EN 0.0216397
R1144 EN.n154 EN.n153 0.0216397
R1145 EN.n154 EN 0.0216397
R1146 EN.n187 EN.n186 0.0216397
R1147 EN.n186 EN 0.0216397
R1148 EN.n177 EN.n176 0.0216397
R1149 EN.n176 EN 0.0216397
R1150 EN.n206 EN.n205 0.0216397
R1151 EN.n205 EN 0.0216397
R1152 EN.n200 EN.n199 0.0216397
R1153 EN.n199 EN 0.0216397
R1154 EN.n227 EN.n226 0.0216397
R1155 EN.n226 EN 0.0216397
R1156 EN.n217 EN.n216 0.0216397
R1157 EN.n216 EN 0.0216397
R1158 EN.n129 EN.n128 0.0216397
R1159 EN.n128 EN 0.0216397
R1160 EN.n123 EN.n122 0.0216397
R1161 EN.n122 EN 0.0216397
R1162 EN.n250 EN.n249 0.0216397
R1163 EN.n249 EN 0.0216397
R1164 EN.n240 EN.n239 0.0216397
R1165 EN.n239 EN 0.0216397
R1166 EN.n268 EN.n267 0.0216397
R1167 EN.n267 EN 0.0216397
R1168 EN.n262 EN.n261 0.0216397
R1169 EN.n261 EN 0.0216397
R1170 EN.n290 EN.n289 0.0216397
R1171 EN.n289 EN 0.0216397
R1172 EN.n280 EN.n279 0.0216397
R1173 EN.n279 EN 0.0216397
R1174 EN.n91 EN.n90 0.0216397
R1175 EN.n90 EN 0.0216397
R1176 EN.n85 EN.n84 0.0216397
R1177 EN.n84 EN 0.0216397
R1178 EN.n112 EN.n111 0.0216397
R1179 EN.n111 EN 0.0216397
R1180 EN.n102 EN.n101 0.0216397
R1181 EN.n101 EN 0.0216397
R1182 EN.n312 EN.n311 0.0216397
R1183 EN.n311 EN 0.0216397
R1184 EN.n306 EN.n305 0.0216397
R1185 EN.n305 EN 0.0216397
R1186 EN.n333 EN.n332 0.0216397
R1187 EN.n332 EN 0.0216397
R1188 EN.n323 EN.n322 0.0216397
R1189 EN.n322 EN 0.0216397
R1190 EN.n27 EN.n26 0.0216397
R1191 EN.n26 EN 0.0216397
R1192 EN.n21 EN.n20 0.0216397
R1193 EN.n20 EN 0.0216397
R1194 EN.n356 EN.n355 0.0216397
R1195 EN.n355 EN 0.0216397
R1196 EN.n346 EN.n345 0.0216397
R1197 EN.n345 EN 0.0216397
R1198 EN.n169 EN.n168 0.0216397
R1199 EN.n168 EN 0.0216397
R1200 EN.n159 EN.n158 0.0216397
R1201 EN.n158 EN 0.0216397
R1202 EN.n46 EN.n45 0.0216397
R1203 EN.n45 EN 0.0216397
R1204 EN.n40 EN.n39 0.0216397
R1205 EN.n39 EN 0.0216397
R1206 EN.n11 EN.n10 0.0216397
R1207 EN.n10 EN 0.0216397
R1208 EN.n1 EN.n0 0.0216397
R1209 EN.n0 EN 0.0216397
R1210 EN.n76 EN 0.0204394
R1211 EN.n365 EN 0.0204394
R1212 EN.n72 EN.n71 0.0107679
R1213 EN.n71 EN 0.0107679
R1214 EN.n66 EN.n65 0.0107679
R1215 EN.n65 EN 0.0107679
R1216 EN.n148 EN.n147 0.0107679
R1217 EN.n147 EN 0.0107679
R1218 EN.n142 EN.n141 0.0107679
R1219 EN.n141 EN 0.0107679
R1220 EN.n180 EN.n179 0.0107679
R1221 EN.n179 EN 0.0107679
R1222 EN.n211 EN.n210 0.0107679
R1223 EN.n210 EN 0.0107679
R1224 EN.n220 EN.n219 0.0107679
R1225 EN.n219 EN 0.0107679
R1226 EN.n134 EN.n133 0.0107679
R1227 EN.n133 EN 0.0107679
R1228 EN.n243 EN.n242 0.0107679
R1229 EN.n242 EN 0.0107679
R1230 EN.n273 EN.n272 0.0107679
R1231 EN.n272 EN 0.0107679
R1232 EN.n283 EN.n282 0.0107679
R1233 EN.n282 EN 0.0107679
R1234 EN.n96 EN.n95 0.0107679
R1235 EN.n95 EN 0.0107679
R1236 EN.n105 EN.n104 0.0107679
R1237 EN.n104 EN 0.0107679
R1238 EN.n317 EN.n316 0.0107679
R1239 EN.n316 EN 0.0107679
R1240 EN.n326 EN.n325 0.0107679
R1241 EN.n325 EN 0.0107679
R1242 EN.n32 EN.n31 0.0107679
R1243 EN.n31 EN 0.0107679
R1244 EN.n349 EN.n348 0.0107679
R1245 EN.n348 EN 0.0107679
R1246 EN.n162 EN.n161 0.0107679
R1247 EN.n161 EN 0.0107679
R1248 EN.n51 EN.n50 0.0107679
R1249 EN.n50 EN 0.0107679
R1250 EN.n4 EN.n3 0.0107679
R1251 EN.n3 EN 0.0107679
R1252 EN.n62 EN 0.00441667
R1253 EN.n156 EN 0.00441667
R1254 EN.n182 EN 0.00441667
R1255 EN.n213 EN 0.00441667
R1256 EN.n222 EN 0.00441667
R1257 EN.n136 EN 0.00441667
R1258 EN.n245 EN 0.00441667
R1259 EN.n275 EN 0.00441667
R1260 EN.n285 EN 0.00441667
R1261 EN.n98 EN 0.00441667
R1262 EN.n107 EN 0.00441667
R1263 EN.n319 EN 0.00441667
R1264 EN.n328 EN 0.00441667
R1265 EN.n34 EN 0.00441667
R1266 EN.n351 EN 0.00441667
R1267 EN.n164 EN 0.00441667
R1268 EN.n53 EN 0.00441667
R1269 EN.n56 EN 0.00441667
R1270 EN.n6 EN 0.00441667
R1271 EN EN.n62 0.00406061
R1272 EN EN.n156 0.00406061
R1273 EN.n182 EN 0.00406061
R1274 EN.n213 EN 0.00406061
R1275 EN.n222 EN 0.00406061
R1276 EN.n136 EN 0.00406061
R1277 EN.n245 EN 0.00406061
R1278 EN.n275 EN 0.00406061
R1279 EN.n285 EN 0.00406061
R1280 EN.n98 EN 0.00406061
R1281 EN.n107 EN 0.00406061
R1282 EN.n319 EN 0.00406061
R1283 EN.n328 EN 0.00406061
R1284 EN.n34 EN 0.00406061
R1285 EN.n351 EN 0.00406061
R1286 EN.n164 EN 0.00406061
R1287 EN.n53 EN 0.00406061
R1288 EN.n6 EN 0.00406061
R1289 EN.n56 EN 0.00406061
R1290 GND.n3527 GND.n3526 49144.5
R1291 GND.n3269 GND.n3268 49144.5
R1292 GND.n2063 GND.n697 45562.9
R1293 GND.n1143 GND.n1068 45562.9
R1294 GND.n1568 GND.n1567 45562.9
R1295 GND.n1980 GND.n828 45562.9
R1296 GND.n3445 GND.n3444 45562.9
R1297 GND.n4259 GND.n4258 45562.9
R1298 GND.n2144 GND.n640 45562.9
R1299 GND.n2065 GND.n2064 45562.9
R1300 GND.n1982 GND.n1981 45562.9
R1301 GND.n2991 GND.n2990 21012.4
R1302 GND.n2772 GND.n2771 19588.1
R1303 GND.n2988 GND.n2987 18646.4
R1304 GND.n1622 GND.n1621 18472.2
R1305 GND.n2989 GND.n2170 15564.8
R1306 GND.n2987 GND.n2171 14136.5
R1307 GND.n2991 GND.n2170 14058
R1308 GND.n2990 GND.n2171 13948.5
R1309 GND.n3398 GND.n3397 12551.1
R1310 GND.n3598 GND.n3597 12551.1
R1311 GND.n3121 GND.n3120 10572.6
R1312 GND.n2772 GND.n2171 10045.2
R1313 GND.n3120 GND.n576 9469.68
R1314 GND.n2771 GND.n576 9469.68
R1315 GND.n3050 GND.n2144 8982.04
R1316 GND.n2017 GND.n805 8969.43
R1317 GND.n1669 GND.n907 8969.43
R1318 GND.n1670 GND.n1669 8969.43
R1319 GND.n1532 GND.n858 8969.43
R1320 GND.n1503 GND.n858 8969.43
R1321 GND.n3573 GND.n3572 8969.43
R1322 GND.n3344 GND.n412 8969.43
R1323 GND.n2100 GND.n674 8969.43
R1324 GND.n2100 GND.n2099 8969.43
R1325 GND.n2017 GND.n2016 8969.43
R1326 GND.n2990 GND.n2989 8048.91
R1327 GND.n3968 GND.n222 6971.5
R1328 GND.n3964 GND.n222 6971.5
R1329 GND.n3968 GND.n223 6971.5
R1330 GND.n3964 GND.n223 6971.5
R1331 GND.n3982 GND.n212 6971.5
R1332 GND.n3978 GND.n212 6971.5
R1333 GND.n3982 GND.n213 6971.5
R1334 GND.n3978 GND.n213 6971.5
R1335 GND.n3989 GND.n208 6971.5
R1336 GND.n3985 GND.n208 6971.5
R1337 GND.n3989 GND.n209 6971.5
R1338 GND.n3985 GND.n209 6971.5
R1339 GND.n4013 GND.n195 6971.5
R1340 GND.n4009 GND.n195 6971.5
R1341 GND.n4013 GND.n196 6971.5
R1342 GND.n4009 GND.n196 6971.5
R1343 GND.n4027 GND.n184 6971.5
R1344 GND.n4023 GND.n184 6971.5
R1345 GND.n4027 GND.n185 6971.5
R1346 GND.n4023 GND.n185 6971.5
R1347 GND.n4034 GND.n180 6971.5
R1348 GND.n4030 GND.n180 6971.5
R1349 GND.n4034 GND.n181 6971.5
R1350 GND.n4030 GND.n181 6971.5
R1351 GND.n4063 GND.n164 6971.5
R1352 GND.n4059 GND.n164 6971.5
R1353 GND.n4063 GND.n165 6971.5
R1354 GND.n4059 GND.n165 6971.5
R1355 GND.n4077 GND.n154 6971.5
R1356 GND.n4073 GND.n154 6971.5
R1357 GND.n4077 GND.n155 6971.5
R1358 GND.n4073 GND.n155 6971.5
R1359 GND.n4084 GND.n150 6971.5
R1360 GND.n4080 GND.n150 6971.5
R1361 GND.n4084 GND.n151 6971.5
R1362 GND.n4080 GND.n151 6971.5
R1363 GND.n4108 GND.n137 6971.5
R1364 GND.n4104 GND.n137 6971.5
R1365 GND.n4108 GND.n138 6971.5
R1366 GND.n4104 GND.n138 6971.5
R1367 GND.n4122 GND.n126 6971.5
R1368 GND.n4118 GND.n126 6971.5
R1369 GND.n4122 GND.n127 6971.5
R1370 GND.n4118 GND.n127 6971.5
R1371 GND.n4129 GND.n122 6971.5
R1372 GND.n4125 GND.n122 6971.5
R1373 GND.n4129 GND.n123 6971.5
R1374 GND.n4125 GND.n123 6971.5
R1375 GND.n4158 GND.n105 6971.5
R1376 GND.n4154 GND.n105 6971.5
R1377 GND.n4158 GND.n106 6971.5
R1378 GND.n4154 GND.n106 6971.5
R1379 GND.n3635 GND.n317 6971.5
R1380 GND.n3675 GND.n317 6971.5
R1381 GND.n3635 GND.n318 6971.5
R1382 GND.n3675 GND.n318 6971.5
R1383 GND.n3608 GND.n334 6971.5
R1384 GND.n3613 GND.n334 6971.5
R1385 GND.n3608 GND.n335 6971.5
R1386 GND.n3613 GND.n335 6971.5
R1387 GND.n341 GND.n340 6971.5
R1388 GND.n3600 GND.n340 6971.5
R1389 GND.n3599 GND.n341 6971.5
R1390 GND.n3600 GND.n3599 6971.5
R1391 GND.n4176 GND.n84 6971.5
R1392 GND.n4176 GND.n85 6971.5
R1393 GND.n84 GND.n83 6971.5
R1394 GND.n85 GND.n83 6971.5
R1395 GND.n4252 GND.n25 6971.5
R1396 GND.n4256 GND.n25 6971.5
R1397 GND.n4252 GND.n26 6971.5
R1398 GND.n4256 GND.n26 6971.5
R1399 GND.n4237 GND.n34 6971.5
R1400 GND.n4241 GND.n34 6971.5
R1401 GND.n4237 GND.n35 6971.5
R1402 GND.n4241 GND.n35 6971.5
R1403 GND.n540 GND.n539 6971.5
R1404 GND.n3192 GND.n539 6971.5
R1405 GND.n3191 GND.n540 6971.5
R1406 GND.n3192 GND.n3191 6971.5
R1407 GND.n3158 GND.n551 6971.5
R1408 GND.n3166 GND.n551 6971.5
R1409 GND.n3158 GND.n552 6971.5
R1410 GND.n3166 GND.n552 6971.5
R1411 GND.n3131 GND.n568 6971.5
R1412 GND.n3136 GND.n568 6971.5
R1413 GND.n3131 GND.n569 6971.5
R1414 GND.n3136 GND.n569 6971.5
R1415 GND.n575 GND.n574 6971.5
R1416 GND.n3123 GND.n574 6971.5
R1417 GND.n3122 GND.n575 6971.5
R1418 GND.n3123 GND.n3122 6971.5
R1419 GND.n3062 GND.n622 6971.5
R1420 GND.n3052 GND.n622 6971.5
R1421 GND.n3062 GND.n623 6971.5
R1422 GND.n3052 GND.n623 6971.5
R1423 GND.n3098 GND.n593 6971.5
R1424 GND.n3088 GND.n593 6971.5
R1425 GND.n3098 GND.n594 6971.5
R1426 GND.n3088 GND.n594 6971.5
R1427 GND.n3111 GND.n581 6971.5
R1428 GND.n3101 GND.n581 6971.5
R1429 GND.n3111 GND.n582 6971.5
R1430 GND.n3101 GND.n582 6971.5
R1431 GND.n629 GND.n621 6971.5
R1432 GND.n632 GND.n629 6971.5
R1433 GND.n631 GND.n621 6971.5
R1434 GND.n632 GND.n631 6971.5
R1435 GND.n600 GND.n592 6971.5
R1436 GND.n603 GND.n600 6971.5
R1437 GND.n602 GND.n592 6971.5
R1438 GND.n603 GND.n602 6971.5
R1439 GND.n588 GND.n580 6971.5
R1440 GND.n591 GND.n588 6971.5
R1441 GND.n590 GND.n580 6971.5
R1442 GND.n591 GND.n590 6971.5
R1443 GND.n1915 GND.n1902 6971.5
R1444 GND.n1915 GND.n1903 6971.5
R1445 GND.n1916 GND.n1902 6971.5
R1446 GND.n1916 GND.n1903 6971.5
R1447 GND.n1793 GND.n1784 6971.5
R1448 GND.n1790 GND.n1784 6971.5
R1449 GND.n1793 GND.n1785 6971.5
R1450 GND.n1790 GND.n1785 6971.5
R1451 GND.n1823 GND.n1814 6971.5
R1452 GND.n1820 GND.n1814 6971.5
R1453 GND.n1823 GND.n1815 6971.5
R1454 GND.n1820 GND.n1815 6971.5
R1455 GND.n1853 GND.n1844 6971.5
R1456 GND.n1850 GND.n1844 6971.5
R1457 GND.n1853 GND.n1845 6971.5
R1458 GND.n1850 GND.n1845 6971.5
R1459 GND.n1838 GND.n1829 6971.5
R1460 GND.n1835 GND.n1829 6971.5
R1461 GND.n1838 GND.n1830 6971.5
R1462 GND.n1835 GND.n1830 6971.5
R1463 GND.n1808 GND.n1799 6971.5
R1464 GND.n1805 GND.n1799 6971.5
R1465 GND.n1808 GND.n1800 6971.5
R1466 GND.n1805 GND.n1800 6971.5
R1467 GND.n1778 GND.n1769 6971.5
R1468 GND.n1775 GND.n1769 6971.5
R1469 GND.n1778 GND.n1770 6971.5
R1470 GND.n1775 GND.n1770 6971.5
R1471 GND.n1978 GND.n829 6971.5
R1472 GND.n1970 GND.n829 6971.5
R1473 GND.n1978 GND.n830 6971.5
R1474 GND.n1970 GND.n830 6971.5
R1475 GND.n1397 GND.n1382 6971.5
R1476 GND.n1389 GND.n1382 6971.5
R1477 GND.n1397 GND.n1383 6971.5
R1478 GND.n1389 GND.n1383 6971.5
R1479 GND.n1402 GND.n1380 6971.5
R1480 GND.n1402 GND.n1381 6971.5
R1481 GND.n1403 GND.n1380 6971.5
R1482 GND.n1403 GND.n1381 6971.5
R1483 GND.n1426 GND.n1361 6971.5
R1484 GND.n1426 GND.n1362 6971.5
R1485 GND.n1427 GND.n1361 6971.5
R1486 GND.n1427 GND.n1362 6971.5
R1487 GND.n1994 GND.n820 6971.5
R1488 GND.n1990 GND.n820 6971.5
R1489 GND.n1994 GND.n821 6971.5
R1490 GND.n1990 GND.n821 6971.5
R1491 GND.n2001 GND.n816 6971.5
R1492 GND.n1997 GND.n816 6971.5
R1493 GND.n2001 GND.n817 6971.5
R1494 GND.n1997 GND.n817 6971.5
R1495 GND.n2015 GND.n806 6971.5
R1496 GND.n2011 GND.n806 6971.5
R1497 GND.n2015 GND.n807 6971.5
R1498 GND.n2011 GND.n807 6971.5
R1499 GND.n2028 GND.n797 6971.5
R1500 GND.n2020 GND.n797 6971.5
R1501 GND.n2028 GND.n798 6971.5
R1502 GND.n2020 GND.n798 6971.5
R1503 GND.n794 GND.n793 6971.5
R1504 GND.n2031 GND.n794 6971.5
R1505 GND.n2032 GND.n793 6971.5
R1506 GND.n2032 GND.n2031 6971.5
R1507 GND.n2061 GND.n698 6971.5
R1508 GND.n2053 GND.n698 6971.5
R1509 GND.n2061 GND.n699 6971.5
R1510 GND.n2053 GND.n699 6971.5
R1511 GND.n706 GND.n705 6971.5
R1512 GND.n770 GND.n705 6971.5
R1513 GND.n769 GND.n706 6971.5
R1514 GND.n770 GND.n769 6971.5
R1515 GND.n754 GND.n707 6971.5
R1516 GND.n766 GND.n707 6971.5
R1517 GND.n754 GND.n708 6971.5
R1518 GND.n766 GND.n708 6971.5
R1519 GND.n723 GND.n719 6971.5
R1520 GND.n732 GND.n719 6971.5
R1521 GND.n723 GND.n720 6971.5
R1522 GND.n732 GND.n720 6971.5
R1523 GND.n2077 GND.n689 6971.5
R1524 GND.n2073 GND.n689 6971.5
R1525 GND.n2077 GND.n690 6971.5
R1526 GND.n2073 GND.n690 6971.5
R1527 GND.n2084 GND.n685 6971.5
R1528 GND.n2080 GND.n685 6971.5
R1529 GND.n2084 GND.n686 6971.5
R1530 GND.n2080 GND.n686 6971.5
R1531 GND.n2098 GND.n675 6971.5
R1532 GND.n2094 GND.n675 6971.5
R1533 GND.n2098 GND.n676 6971.5
R1534 GND.n2094 GND.n676 6971.5
R1535 GND.n2111 GND.n666 6971.5
R1536 GND.n2103 GND.n666 6971.5
R1537 GND.n2111 GND.n667 6971.5
R1538 GND.n2103 GND.n667 6971.5
R1539 GND.n663 GND.n662 6971.5
R1540 GND.n2114 GND.n663 6971.5
R1541 GND.n2115 GND.n662 6971.5
R1542 GND.n2115 GND.n2114 6971.5
R1543 GND.n2142 GND.n641 6971.5
R1544 GND.n2136 GND.n641 6971.5
R1545 GND.n2142 GND.n642 6971.5
R1546 GND.n2136 GND.n642 6971.5
R1547 GND.n1265 GND.n1210 6971.5
R1548 GND.n1269 GND.n1210 6971.5
R1549 GND.n1265 GND.n1211 6971.5
R1550 GND.n1269 GND.n1211 6971.5
R1551 GND.n1258 GND.n1214 6971.5
R1552 GND.n1262 GND.n1214 6971.5
R1553 GND.n1258 GND.n1215 6971.5
R1554 GND.n1262 GND.n1215 6971.5
R1555 GND.n1243 GND.n1223 6971.5
R1556 GND.n1247 GND.n1223 6971.5
R1557 GND.n1243 GND.n1224 6971.5
R1558 GND.n1247 GND.n1224 6971.5
R1559 GND.n1344 GND.n1189 6971.5
R1560 GND.n1348 GND.n1189 6971.5
R1561 GND.n1344 GND.n1190 6971.5
R1562 GND.n1348 GND.n1190 6971.5
R1563 GND.n1337 GND.n1193 6971.5
R1564 GND.n1341 GND.n1193 6971.5
R1565 GND.n1337 GND.n1194 6971.5
R1566 GND.n1341 GND.n1194 6971.5
R1567 GND.n1326 GND.n1202 6971.5
R1568 GND.n1326 GND.n1203 6971.5
R1569 GND.n1322 GND.n1203 6971.5
R1570 GND.n1322 GND.n1202 6971.5
R1571 GND.n1754 GND.n851 6971.5
R1572 GND.n1746 GND.n851 6971.5
R1573 GND.n1754 GND.n852 6971.5
R1574 GND.n1746 GND.n852 6971.5
R1575 GND.n1571 GND.n1570 6971.5
R1576 GND.n1570 GND.n1060 6971.5
R1577 GND.n1571 GND.n881 6971.5
R1578 GND.n1060 GND.n881 6971.5
R1579 GND.n1576 GND.n1059 6971.5
R1580 GND.n1576 GND.n1574 6971.5
R1581 GND.n1059 GND.n877 6971.5
R1582 GND.n1574 GND.n877 6971.5
R1583 GND.n1742 GND.n859 6971.5
R1584 GND.n1734 GND.n859 6971.5
R1585 GND.n1742 GND.n860 6971.5
R1586 GND.n1734 GND.n860 6971.5
R1587 GND.n1105 GND.n1095 6971.5
R1588 GND.n1106 GND.n1105 6971.5
R1589 GND.n1095 GND.n1093 6971.5
R1590 GND.n1106 GND.n1093 6971.5
R1591 GND.n1101 GND.n1099 6971.5
R1592 GND.n1102 GND.n1101 6971.5
R1593 GND.n1099 GND.n1089 6971.5
R1594 GND.n1102 GND.n1089 6971.5
R1595 GND.n1141 GND.n1069 6971.5
R1596 GND.n1079 GND.n1069 6971.5
R1597 GND.n1141 GND.n1070 6971.5
R1598 GND.n1079 GND.n1070 6971.5
R1599 GND.n1028 GND.n1017 6971.5
R1600 GND.n1029 GND.n1028 6971.5
R1601 GND.n1017 GND.n931 6971.5
R1602 GND.n1029 GND.n931 6971.5
R1603 GND.n1024 GND.n1019 6971.5
R1604 GND.n1025 GND.n1024 6971.5
R1605 GND.n1019 GND.n927 6971.5
R1606 GND.n1025 GND.n927 6971.5
R1607 GND.n1666 GND.n909 6971.5
R1608 GND.n1658 GND.n909 6971.5
R1609 GND.n1666 GND.n910 6971.5
R1610 GND.n1658 GND.n910 6971.5
R1611 GND.n1009 GND.n937 6971.5
R1612 GND.n1013 GND.n937 6971.5
R1613 GND.n1009 GND.n938 6971.5
R1614 GND.n1013 GND.n938 6971.5
R1615 GND.n1002 GND.n941 6971.5
R1616 GND.n1006 GND.n941 6971.5
R1617 GND.n1002 GND.n942 6971.5
R1618 GND.n1006 GND.n942 6971.5
R1619 GND.n987 GND.n950 6971.5
R1620 GND.n991 GND.n950 6971.5
R1621 GND.n987 GND.n951 6971.5
R1622 GND.n991 GND.n951 6971.5
R1623 GND.n1682 GND.n900 6971.5
R1624 GND.n1678 GND.n900 6971.5
R1625 GND.n1682 GND.n901 6971.5
R1626 GND.n1678 GND.n901 6971.5
R1627 GND.n1689 GND.n896 6971.5
R1628 GND.n1685 GND.n896 6971.5
R1629 GND.n1689 GND.n897 6971.5
R1630 GND.n1685 GND.n897 6971.5
R1631 GND.n1067 GND.n886 6971.5
R1632 GND.n1062 GND.n886 6971.5
R1633 GND.n1067 GND.n1066 6971.5
R1634 GND.n1066 GND.n1062 6971.5
R1635 GND.n1555 GND.n1147 6971.5
R1636 GND.n1559 GND.n1147 6971.5
R1637 GND.n1555 GND.n1148 6971.5
R1638 GND.n1559 GND.n1148 6971.5
R1639 GND.n1548 GND.n1151 6971.5
R1640 GND.n1552 GND.n1151 6971.5
R1641 GND.n1548 GND.n1152 6971.5
R1642 GND.n1552 GND.n1152 6971.5
R1643 GND.n1533 GND.n1160 6971.5
R1644 GND.n1537 GND.n1160 6971.5
R1645 GND.n1533 GND.n1161 6971.5
R1646 GND.n1537 GND.n1161 6971.5
R1647 GND.n1495 GND.n1168 6971.5
R1648 GND.n1499 GND.n1168 6971.5
R1649 GND.n1495 GND.n1169 6971.5
R1650 GND.n1499 GND.n1169 6971.5
R1651 GND.n1488 GND.n1172 6971.5
R1652 GND.n1492 GND.n1172 6971.5
R1653 GND.n1488 GND.n1173 6971.5
R1654 GND.n1492 GND.n1173 6971.5
R1655 GND.n1473 GND.n1181 6971.5
R1656 GND.n1477 GND.n1181 6971.5
R1657 GND.n1473 GND.n1182 6971.5
R1658 GND.n1477 GND.n1182 6971.5
R1659 GND.n1948 GND.n849 6971.5
R1660 GND.n1948 GND.n850 6971.5
R1661 GND.n1949 GND.n849 6971.5
R1662 GND.n1949 GND.n850 6971.5
R1663 GND.n3338 GND.n413 6971.5
R1664 GND.n3342 GND.n413 6971.5
R1665 GND.n3338 GND.n414 6971.5
R1666 GND.n3342 GND.n414 6971.5
R1667 GND.n3236 GND.n3218 6971.5
R1668 GND.n3232 GND.n3218 6971.5
R1669 GND.n3236 GND.n3219 6971.5
R1670 GND.n3232 GND.n3219 6971.5
R1671 GND.n3243 GND.n3214 6971.5
R1672 GND.n3239 GND.n3214 6971.5
R1673 GND.n3243 GND.n3215 6971.5
R1674 GND.n3239 GND.n3215 6971.5
R1675 GND.n492 GND.n491 6971.5
R1676 GND.n3311 GND.n491 6971.5
R1677 GND.n3310 GND.n492 6971.5
R1678 GND.n3311 GND.n3310 6971.5
R1679 GND.n3279 GND.n505 6971.5
R1680 GND.n3284 GND.n505 6971.5
R1681 GND.n3279 GND.n506 6971.5
R1682 GND.n3284 GND.n506 6971.5
R1683 GND.n512 GND.n511 6971.5
R1684 GND.n3271 GND.n511 6971.5
R1685 GND.n3270 GND.n512 6971.5
R1686 GND.n3271 GND.n3270 6971.5
R1687 GND.n3488 GND.n348 6971.5
R1688 GND.n3574 GND.n348 6971.5
R1689 GND.n3488 GND.n349 6971.5
R1690 GND.n3574 GND.n349 6971.5
R1691 GND.n3514 GND.n3466 6971.5
R1692 GND.n3506 GND.n3466 6971.5
R1693 GND.n3514 GND.n3467 6971.5
R1694 GND.n3506 GND.n3467 6971.5
R1695 GND.n3566 GND.n351 6971.5
R1696 GND.n3570 GND.n351 6971.5
R1697 GND.n3566 GND.n352 6971.5
R1698 GND.n3570 GND.n352 6971.5
R1699 GND.n363 GND.n362 6971.5
R1700 GND.n3544 GND.n362 6971.5
R1701 GND.n3543 GND.n363 6971.5
R1702 GND.n3544 GND.n3543 6971.5
R1703 GND.n3536 GND.n364 6971.5
R1704 GND.n3540 GND.n364 6971.5
R1705 GND.n3536 GND.n365 6971.5
R1706 GND.n3540 GND.n365 6971.5
R1707 GND.n458 GND.n379 6971.5
R1708 GND.n3447 GND.n379 6971.5
R1709 GND.n458 GND.n380 6971.5
R1710 GND.n3447 GND.n380 6971.5
R1711 GND.n472 GND.n431 6971.5
R1712 GND.n468 GND.n431 6971.5
R1713 GND.n472 GND.n432 6971.5
R1714 GND.n468 GND.n432 6971.5
R1715 GND.n479 GND.n427 6971.5
R1716 GND.n475 GND.n427 6971.5
R1717 GND.n479 GND.n428 6971.5
R1718 GND.n475 GND.n428 6971.5
R1719 GND.n3435 GND.n382 6971.5
R1720 GND.n3443 GND.n382 6971.5
R1721 GND.n3435 GND.n383 6971.5
R1722 GND.n3443 GND.n383 6971.5
R1723 GND.n3408 GND.n399 6971.5
R1724 GND.n3413 GND.n399 6971.5
R1725 GND.n3408 GND.n400 6971.5
R1726 GND.n3413 GND.n400 6971.5
R1727 GND.n406 GND.n405 6971.5
R1728 GND.n3400 GND.n405 6971.5
R1729 GND.n3399 GND.n406 6971.5
R1730 GND.n3400 GND.n3399 6971.5
R1731 GND.n3525 GND.n372 6971.5
R1732 GND.n3525 GND.n373 6971.5
R1733 GND.n3517 GND.n372 6971.5
R1734 GND.n3517 GND.n373 6971.5
R1735 GND.n3911 GND.n3898 6971.5
R1736 GND.n3903 GND.n3898 6971.5
R1737 GND.n3911 GND.n3899 6971.5
R1738 GND.n3903 GND.n3899 6971.5
R1739 GND.n3887 GND.n238 6971.5
R1740 GND.n3888 GND.n3887 6971.5
R1741 GND.n238 GND.n232 6971.5
R1742 GND.n3888 GND.n232 6971.5
R1743 GND.n3871 GND.n242 6971.5
R1744 GND.n3879 GND.n242 6971.5
R1745 GND.n3871 GND.n243 6971.5
R1746 GND.n3879 GND.n243 6971.5
R1747 GND.n3844 GND.n259 6971.5
R1748 GND.n3849 GND.n259 6971.5
R1749 GND.n3844 GND.n260 6971.5
R1750 GND.n3849 GND.n260 6971.5
R1751 GND.n266 GND.n265 6971.5
R1752 GND.n3836 GND.n265 6971.5
R1753 GND.n3835 GND.n266 6971.5
R1754 GND.n3836 GND.n3835 6971.5
R1755 GND.n3749 GND.n267 6971.5
R1756 GND.n3828 GND.n267 6971.5
R1757 GND.n3749 GND.n268 6971.5
R1758 GND.n3828 GND.n268 6971.5
R1759 GND.n3734 GND.n288 6971.5
R1760 GND.n3735 GND.n3734 6971.5
R1761 GND.n288 GND.n282 6971.5
R1762 GND.n3735 GND.n282 6971.5
R1763 GND.n3730 GND.n290 6971.5
R1764 GND.n3731 GND.n3730 6971.5
R1765 GND.n290 GND.n278 6971.5
R1766 GND.n3731 GND.n278 6971.5
R1767 GND.n3718 GND.n292 6971.5
R1768 GND.n3726 GND.n292 6971.5
R1769 GND.n3718 GND.n293 6971.5
R1770 GND.n3726 GND.n293 6971.5
R1771 GND.n3691 GND.n309 6971.5
R1772 GND.n3696 GND.n309 6971.5
R1773 GND.n3691 GND.n310 6971.5
R1774 GND.n3696 GND.n310 6971.5
R1775 GND.n316 GND.n315 6971.5
R1776 GND.n3683 GND.n315 6971.5
R1777 GND.n3682 GND.n316 6971.5
R1778 GND.n3683 GND.n3682 6971.5
R1779 GND.n3883 GND.n240 6971.5
R1780 GND.n240 GND.n228 6971.5
R1781 GND.n3884 GND.n3883 6971.5
R1782 GND.n3884 GND.n228 6971.5
R1783 GND.n4268 GND.n19 6971.5
R1784 GND.n4260 GND.n19 6971.5
R1785 GND.n4268 GND.n20 6971.5
R1786 GND.n4260 GND.n20 6971.5
R1787 GND.n3176 GND.n3175 6971.5
R1788 GND.n3175 GND.n3170 6971.5
R1789 GND.n3176 GND.n7 6971.5
R1790 GND.n3170 GND.n7 6971.5
R1791 GND.n3180 GND.n3179 6971.5
R1792 GND.n3180 GND.n3 6971.5
R1793 GND.n3179 GND.n3168 6971.5
R1794 GND.n3168 GND.n3 6971.5
R1795 GND.n2153 GND.n2152 6971.5
R1796 GND.n3023 GND.n2152 6971.5
R1797 GND.n3022 GND.n2153 6971.5
R1798 GND.n3023 GND.n3022 6971.5
R1799 GND.n3007 GND.n2159 6971.5
R1800 GND.n3011 GND.n2159 6971.5
R1801 GND.n3007 GND.n2160 6971.5
R1802 GND.n3011 GND.n2160 6971.5
R1803 GND.n3000 GND.n2163 6971.5
R1804 GND.n3004 GND.n2163 6971.5
R1805 GND.n3000 GND.n2164 6971.5
R1806 GND.n3004 GND.n2164 6971.5
R1807 GND.n2823 GND.n2811 6971.5
R1808 GND.n2823 GND.n2812 6971.5
R1809 GND.n2811 GND.n2808 6971.5
R1810 GND.n2812 GND.n2808 6971.5
R1811 GND.n2856 GND.n2467 6971.5
R1812 GND.n2848 GND.n2467 6971.5
R1813 GND.n2856 GND.n2468 6971.5
R1814 GND.n2848 GND.n2468 6971.5
R1815 GND.n2861 GND.n2461 6971.5
R1816 GND.n2861 GND.n2462 6971.5
R1817 GND.n2862 GND.n2461 6971.5
R1818 GND.n2862 GND.n2462 6971.5
R1819 GND.n2824 GND.n2803 6971.5
R1820 GND.n2824 GND.n2804 6971.5
R1821 GND.n2807 GND.n2803 6971.5
R1822 GND.n2807 GND.n2804 6971.5
R1823 GND.n2791 GND.n2466 6971.5
R1824 GND.n2791 GND.n2473 6971.5
R1825 GND.n2792 GND.n2466 6971.5
R1826 GND.n2792 GND.n2473 6971.5
R1827 GND.n2781 GND.n2463 6971.5
R1828 GND.n2465 GND.n2463 6971.5
R1829 GND.n2781 GND.n2464 6971.5
R1830 GND.n2465 GND.n2464 6971.5
R1831 GND.n2929 GND.n2908 6971.5
R1832 GND.n2919 GND.n2908 6971.5
R1833 GND.n2929 GND.n2909 6971.5
R1834 GND.n2919 GND.n2909 6971.5
R1835 GND.n2965 GND.n2879 6971.5
R1836 GND.n2955 GND.n2879 6971.5
R1837 GND.n2965 GND.n2880 6971.5
R1838 GND.n2955 GND.n2880 6971.5
R1839 GND.n2978 GND.n2177 6971.5
R1840 GND.n2968 GND.n2177 6971.5
R1841 GND.n2978 GND.n2178 6971.5
R1842 GND.n2968 GND.n2178 6971.5
R1843 GND.n2915 GND.n2907 6971.5
R1844 GND.n2917 GND.n2915 6971.5
R1845 GND.n2916 GND.n2907 6971.5
R1846 GND.n2917 GND.n2916 6971.5
R1847 GND.n2886 GND.n2878 6971.5
R1848 GND.n2889 GND.n2886 6971.5
R1849 GND.n2888 GND.n2878 6971.5
R1850 GND.n2889 GND.n2888 6971.5
R1851 GND.n2874 GND.n2176 6971.5
R1852 GND.n2877 GND.n2874 6971.5
R1853 GND.n2876 GND.n2176 6971.5
R1854 GND.n2877 GND.n2876 6971.5
R1855 GND.n2397 GND.n2376 6971.5
R1856 GND.n2387 GND.n2376 6971.5
R1857 GND.n2397 GND.n2377 6971.5
R1858 GND.n2387 GND.n2377 6971.5
R1859 GND.n2433 GND.n2347 6971.5
R1860 GND.n2423 GND.n2347 6971.5
R1861 GND.n2433 GND.n2348 6971.5
R1862 GND.n2423 GND.n2348 6971.5
R1863 GND.n2446 GND.n2335 6971.5
R1864 GND.n2436 GND.n2335 6971.5
R1865 GND.n2446 GND.n2336 6971.5
R1866 GND.n2436 GND.n2336 6971.5
R1867 GND.n2383 GND.n2375 6971.5
R1868 GND.n2385 GND.n2383 6971.5
R1869 GND.n2384 GND.n2375 6971.5
R1870 GND.n2385 GND.n2384 6971.5
R1871 GND.n2354 GND.n2346 6971.5
R1872 GND.n2357 GND.n2354 6971.5
R1873 GND.n2356 GND.n2346 6971.5
R1874 GND.n2357 GND.n2356 6971.5
R1875 GND.n2342 GND.n2334 6971.5
R1876 GND.n2345 GND.n2342 6971.5
R1877 GND.n2344 GND.n2334 6971.5
R1878 GND.n2345 GND.n2344 6971.5
R1879 GND.n2270 GND.n2249 6971.5
R1880 GND.n2260 GND.n2249 6971.5
R1881 GND.n2270 GND.n2250 6971.5
R1882 GND.n2260 GND.n2250 6971.5
R1883 GND.n2306 GND.n2220 6971.5
R1884 GND.n2296 GND.n2220 6971.5
R1885 GND.n2306 GND.n2221 6971.5
R1886 GND.n2296 GND.n2221 6971.5
R1887 GND.n2319 GND.n2208 6971.5
R1888 GND.n2309 GND.n2208 6971.5
R1889 GND.n2319 GND.n2209 6971.5
R1890 GND.n2309 GND.n2209 6971.5
R1891 GND.n2256 GND.n2248 6971.5
R1892 GND.n2258 GND.n2256 6971.5
R1893 GND.n2257 GND.n2248 6971.5
R1894 GND.n2258 GND.n2257 6971.5
R1895 GND.n2227 GND.n2219 6971.5
R1896 GND.n2230 GND.n2227 6971.5
R1897 GND.n2229 GND.n2219 6971.5
R1898 GND.n2230 GND.n2229 6971.5
R1899 GND.n2215 GND.n2207 6971.5
R1900 GND.n2218 GND.n2215 6971.5
R1901 GND.n2217 GND.n2207 6971.5
R1902 GND.n2218 GND.n2217 6971.5
R1903 GND.n2592 GND.n2571 6971.5
R1904 GND.n2582 GND.n2571 6971.5
R1905 GND.n2592 GND.n2572 6971.5
R1906 GND.n2582 GND.n2572 6971.5
R1907 GND.n2628 GND.n2542 6971.5
R1908 GND.n2618 GND.n2542 6971.5
R1909 GND.n2628 GND.n2543 6971.5
R1910 GND.n2618 GND.n2543 6971.5
R1911 GND.n2641 GND.n2530 6971.5
R1912 GND.n2631 GND.n2530 6971.5
R1913 GND.n2641 GND.n2531 6971.5
R1914 GND.n2631 GND.n2531 6971.5
R1915 GND.n2578 GND.n2570 6971.5
R1916 GND.n2580 GND.n2578 6971.5
R1917 GND.n2579 GND.n2570 6971.5
R1918 GND.n2580 GND.n2579 6971.5
R1919 GND.n2549 GND.n2541 6971.5
R1920 GND.n2552 GND.n2549 6971.5
R1921 GND.n2551 GND.n2541 6971.5
R1922 GND.n2552 GND.n2551 6971.5
R1923 GND.n2537 GND.n2529 6971.5
R1924 GND.n2540 GND.n2537 6971.5
R1925 GND.n2539 GND.n2529 6971.5
R1926 GND.n2540 GND.n2539 6971.5
R1927 GND.n2713 GND.n2692 6971.5
R1928 GND.n2703 GND.n2692 6971.5
R1929 GND.n2713 GND.n2693 6971.5
R1930 GND.n2703 GND.n2693 6971.5
R1931 GND.n2749 GND.n2663 6971.5
R1932 GND.n2739 GND.n2663 6971.5
R1933 GND.n2749 GND.n2664 6971.5
R1934 GND.n2739 GND.n2664 6971.5
R1935 GND.n2762 GND.n2511 6971.5
R1936 GND.n2752 GND.n2511 6971.5
R1937 GND.n2762 GND.n2512 6971.5
R1938 GND.n2752 GND.n2512 6971.5
R1939 GND.n2699 GND.n2691 6971.5
R1940 GND.n2701 GND.n2699 6971.5
R1941 GND.n2700 GND.n2691 6971.5
R1942 GND.n2701 GND.n2700 6971.5
R1943 GND.n2670 GND.n2662 6971.5
R1944 GND.n2673 GND.n2670 6971.5
R1945 GND.n2672 GND.n2662 6971.5
R1946 GND.n2673 GND.n2672 6971.5
R1947 GND.n2658 GND.n2510 6971.5
R1948 GND.n2661 GND.n2658 6971.5
R1949 GND.n2660 GND.n2510 6971.5
R1950 GND.n2661 GND.n2660 6971.5
R1951 GND.n1944 GND.n1759 6971.5
R1952 GND.n1944 GND.n1760 6971.5
R1953 GND.n1940 GND.n1760 6971.5
R1954 GND.n1940 GND.n1759 6971.5
R1955 GND.n1907 GND.n94 6971.5
R1956 GND.n1911 GND.n94 6971.5
R1957 GND.n1910 GND.n1907 6971.5
R1958 GND.n1911 GND.n1910 6971.5
R1959 GND.n3182 GND.n3181 5897.47
R1960 GND.n3681 GND.n3680 5734.32
R1961 GND.n3729 GND.n3728 5734.32
R1962 GND.n3834 GND.n3833 5734.32
R1963 GND.n3882 GND.n3881 5734.32
R1964 GND.n4006 GND.n199 5246.88
R1965 GND.n3999 GND.n199 5246.88
R1966 GND.n4006 GND.n200 5246.88
R1967 GND.n3999 GND.n200 5246.88
R1968 GND.n4046 GND.n175 5246.88
R1969 GND.n4046 GND.n176 5246.88
R1970 GND.n4048 GND.n175 5246.88
R1971 GND.n4048 GND.n176 5246.88
R1972 GND.n4101 GND.n141 5246.88
R1973 GND.n4094 GND.n141 5246.88
R1974 GND.n4101 GND.n142 5246.88
R1975 GND.n4094 GND.n142 5246.88
R1976 GND.n4141 GND.n117 5246.88
R1977 GND.n4141 GND.n118 5246.88
R1978 GND.n4143 GND.n117 5246.88
R1979 GND.n4143 GND.n118 5246.88
R1980 GND.n3975 GND.n216 5246.88
R1981 GND.n3971 GND.n216 5246.88
R1982 GND.n3975 GND.n217 5246.88
R1983 GND.n3971 GND.n217 5246.88
R1984 GND.n4020 GND.n189 5246.88
R1985 GND.n4016 GND.n189 5246.88
R1986 GND.n4020 GND.n190 5246.88
R1987 GND.n4016 GND.n190 5246.88
R1988 GND.n4070 GND.n158 5246.88
R1989 GND.n4066 GND.n158 5246.88
R1990 GND.n4070 GND.n159 5246.88
R1991 GND.n4066 GND.n159 5246.88
R1992 GND.n4115 GND.n131 5246.88
R1993 GND.n4111 GND.n131 5246.88
R1994 GND.n4115 GND.n132 5246.88
R1995 GND.n4111 GND.n132 5246.88
R1996 GND.n4162 GND.n99 5246.88
R1997 GND.n4162 GND.n100 5246.88
R1998 GND.n103 GND.n99 5246.88
R1999 GND.n103 GND.n100 5246.88
R2000 GND.n3625 GND.n322 5246.88
R2001 GND.n3632 GND.n322 5246.88
R2002 GND.n3625 GND.n323 5246.88
R2003 GND.n3632 GND.n323 5246.88
R2004 GND.n4181 GND.n77 5246.88
R2005 GND.n4181 GND.n78 5246.88
R2006 GND.n4183 GND.n77 5246.88
R2007 GND.n4183 GND.n78 5246.88
R2008 GND.n4203 GND.n61 5246.88
R2009 GND.n4196 GND.n61 5246.88
R2010 GND.n4203 GND.n62 5246.88
R2011 GND.n4196 GND.n62 5246.88
R2012 GND.n4210 GND.n56 5246.88
R2013 GND.n4210 GND.n57 5246.88
R2014 GND.n4212 GND.n56 5246.88
R2015 GND.n4212 GND.n57 5246.88
R2016 GND.n4232 GND.n40 5246.88
R2017 GND.n4225 GND.n40 5246.88
R2018 GND.n4232 GND.n41 5246.88
R2019 GND.n4225 GND.n41 5246.88
R2020 GND.n3038 GND.n3031 5246.88
R2021 GND.n3038 GND.n3032 5246.88
R2022 GND.n3040 GND.n3031 5246.88
R2023 GND.n3040 GND.n3032 5246.88
R2024 GND.n4245 GND.n29 5246.88
R2025 GND.n4249 GND.n29 5246.88
R2026 GND.n4245 GND.n30 5246.88
R2027 GND.n4249 GND.n30 5246.88
R2028 GND.n3148 GND.n556 5246.88
R2029 GND.n3155 GND.n556 5246.88
R2030 GND.n3148 GND.n557 5246.88
R2031 GND.n3155 GND.n557 5246.88
R2032 GND.n3074 GND.n620 5246.88
R2033 GND.n3074 GND.n3065 5246.88
R2034 GND.n620 GND.n615 5246.88
R2035 GND.n3065 GND.n615 5246.88
R2036 GND.n3076 GND.n613 5246.88
R2037 GND.n3076 GND.n614 5246.88
R2038 GND.n616 GND.n613 5246.88
R2039 GND.n616 GND.n614 5246.88
R2040 GND.n1609 GND.n1031 5246.88
R2041 GND.n1617 GND.n1031 5246.88
R2042 GND.n1609 GND.n1032 5246.88
R2043 GND.n1617 GND.n1032 5246.88
R2044 GND.n1595 GND.n1036 5246.88
R2045 GND.n1603 GND.n1036 5246.88
R2046 GND.n1595 GND.n1037 5246.88
R2047 GND.n1603 GND.n1037 5246.88
R2048 GND.n1967 GND.n835 5246.88
R2049 GND.n1960 GND.n835 5246.88
R2050 GND.n1967 GND.n836 5246.88
R2051 GND.n1960 GND.n836 5246.88
R2052 GND.n1421 GND.n1363 5246.88
R2053 GND.n1414 GND.n1363 5246.88
R2054 GND.n1421 GND.n1364 5246.88
R2055 GND.n1414 GND.n1364 5246.88
R2056 GND.n2008 GND.n810 5246.88
R2057 GND.n2004 GND.n810 5246.88
R2058 GND.n2008 GND.n811 5246.88
R2059 GND.n2004 GND.n811 5246.88
R2060 GND.n2050 GND.n777 5246.88
R2061 GND.n2043 GND.n777 5246.88
R2062 GND.n2050 GND.n778 5246.88
R2063 GND.n2043 GND.n778 5246.88
R2064 GND.n736 GND.n715 5246.88
R2065 GND.n744 GND.n715 5246.88
R2066 GND.n736 GND.n716 5246.88
R2067 GND.n744 GND.n716 5246.88
R2068 GND.n2091 GND.n679 5246.88
R2069 GND.n2087 GND.n679 5246.88
R2070 GND.n2091 GND.n680 5246.88
R2071 GND.n2087 GND.n680 5246.88
R2072 GND.n2133 GND.n646 5246.88
R2073 GND.n2126 GND.n646 5246.88
R2074 GND.n2133 GND.n647 5246.88
R2075 GND.n2126 GND.n647 5246.88
R2076 GND.n1251 GND.n1218 5246.88
R2077 GND.n1255 GND.n1218 5246.88
R2078 GND.n1251 GND.n1219 5246.88
R2079 GND.n1255 GND.n1219 5246.88
R2080 GND.n1330 GND.n1197 5246.88
R2081 GND.n1334 GND.n1197 5246.88
R2082 GND.n1330 GND.n1198 5246.88
R2083 GND.n1334 GND.n1198 5246.88
R2084 GND.n1731 GND.n865 5246.88
R2085 GND.n1724 GND.n865 5246.88
R2086 GND.n1731 GND.n866 5246.88
R2087 GND.n1724 GND.n866 5246.88
R2088 GND.n1129 GND.n1076 5246.88
R2089 GND.n1129 GND.n1077 5246.88
R2090 GND.n1131 GND.n1076 5246.88
R2091 GND.n1131 GND.n1077 5246.88
R2092 GND.n1655 GND.n915 5246.88
R2093 GND.n1648 GND.n915 5246.88
R2094 GND.n1655 GND.n916 5246.88
R2095 GND.n1648 GND.n916 5246.88
R2096 GND.n995 GND.n945 5246.88
R2097 GND.n999 GND.n945 5246.88
R2098 GND.n995 GND.n946 5246.88
R2099 GND.n999 GND.n946 5246.88
R2100 GND.n1693 GND.n891 5246.88
R2101 GND.n1693 GND.n892 5246.88
R2102 GND.n895 GND.n891 5246.88
R2103 GND.n895 GND.n892 5246.88
R2104 GND.n1541 GND.n1155 5246.88
R2105 GND.n1545 GND.n1155 5246.88
R2106 GND.n1541 GND.n1156 5246.88
R2107 GND.n1545 GND.n1156 5246.88
R2108 GND.n1481 GND.n1176 5246.88
R2109 GND.n1485 GND.n1176 5246.88
R2110 GND.n1481 GND.n1177 5246.88
R2111 GND.n1485 GND.n1177 5246.88
R2112 GND.n530 GND.n514 5246.88
R2113 GND.n3266 GND.n514 5246.88
R2114 GND.n530 GND.n515 5246.88
R2115 GND.n3266 GND.n515 5246.88
R2116 GND.n3331 GND.n417 5246.88
R2117 GND.n3335 GND.n417 5246.88
R2118 GND.n3331 GND.n418 5246.88
R2119 GND.n3335 GND.n418 5246.88
R2120 GND.n3296 GND.n493 5246.88
R2121 GND.n3307 GND.n493 5246.88
R2122 GND.n3296 GND.n494 5246.88
R2123 GND.n3307 GND.n494 5246.88
R2124 GND.n3493 GND.n3479 5246.88
R2125 GND.n3493 GND.n3480 5246.88
R2126 GND.n3495 GND.n3479 5246.88
R2127 GND.n3495 GND.n3480 5246.88
R2128 GND.n3559 GND.n355 5246.88
R2129 GND.n3563 GND.n355 5246.88
R2130 GND.n3559 GND.n356 5246.88
R2131 GND.n3563 GND.n356 5246.88
R2132 GND.n3370 GND.n3366 5246.88
R2133 GND.n3370 GND.n3367 5246.88
R2134 GND.n3372 GND.n3366 5246.88
R2135 GND.n3372 GND.n3367 5246.88
R2136 GND.n465 GND.n435 5246.88
R2137 GND.n461 GND.n435 5246.88
R2138 GND.n465 GND.n436 5246.88
R2139 GND.n461 GND.n436 5246.88
R2140 GND.n3384 GND.n3357 5246.88
R2141 GND.n3377 GND.n3357 5246.88
R2142 GND.n3384 GND.n3359 5246.88
R2143 GND.n3377 GND.n3359 5246.88
R2144 GND.n3425 GND.n387 5246.88
R2145 GND.n3432 GND.n387 5246.88
R2146 GND.n3425 GND.n388 5246.88
R2147 GND.n3432 GND.n388 5246.88
R2148 GND.n3347 GND.n408 5246.88
R2149 GND.n3347 GND.n409 5246.88
R2150 GND.n3395 GND.n408 5246.88
R2151 GND.n3395 GND.n409 5246.88
R2152 GND.n3921 GND.n3892 5246.88
R2153 GND.n3914 GND.n3892 5246.88
R2154 GND.n3921 GND.n3893 5246.88
R2155 GND.n3914 GND.n3893 5246.88
R2156 GND.n3861 GND.n247 5246.88
R2157 GND.n3868 GND.n247 5246.88
R2158 GND.n3861 GND.n248 5246.88
R2159 GND.n3868 GND.n248 5246.88
R2160 GND.n3759 GND.n3739 5246.88
R2161 GND.n3752 GND.n3739 5246.88
R2162 GND.n3759 GND.n3740 5246.88
R2163 GND.n3752 GND.n3740 5246.88
R2164 GND.n3708 GND.n297 5246.88
R2165 GND.n3715 GND.n297 5246.88
R2166 GND.n3708 GND.n298 5246.88
R2167 GND.n3715 GND.n298 5246.88
R2168 GND.n4278 GND.n13 5246.88
R2169 GND.n4271 GND.n13 5246.88
R2170 GND.n4278 GND.n14 5246.88
R2171 GND.n4271 GND.n14 5246.88
R2172 GND.n3015 GND.n2154 5246.88
R2173 GND.n3019 GND.n2154 5246.88
R2174 GND.n3015 GND.n2155 5246.88
R2175 GND.n3019 GND.n2155 5246.88
R2176 GND.n2835 GND.n2482 5246.88
R2177 GND.n2835 GND.n2483 5246.88
R2178 GND.n2837 GND.n2482 5246.88
R2179 GND.n2837 GND.n2483 5246.88
R2180 GND.n2832 GND.n2488 5246.88
R2181 GND.n2832 GND.n2489 5246.88
R2182 GND.n2488 GND.n2484 5246.88
R2183 GND.n2489 GND.n2484 5246.88
R2184 GND.n2941 GND.n2906 5246.88
R2185 GND.n2941 GND.n2932 5246.88
R2186 GND.n2906 GND.n2901 5246.88
R2187 GND.n2932 GND.n2901 5246.88
R2188 GND.n2943 GND.n2899 5246.88
R2189 GND.n2943 GND.n2900 5246.88
R2190 GND.n2902 GND.n2899 5246.88
R2191 GND.n2902 GND.n2900 5246.88
R2192 GND.n2409 GND.n2374 5246.88
R2193 GND.n2409 GND.n2400 5246.88
R2194 GND.n2374 GND.n2369 5246.88
R2195 GND.n2400 GND.n2369 5246.88
R2196 GND.n2411 GND.n2367 5246.88
R2197 GND.n2411 GND.n2368 5246.88
R2198 GND.n2370 GND.n2367 5246.88
R2199 GND.n2370 GND.n2368 5246.88
R2200 GND.n2282 GND.n2247 5246.88
R2201 GND.n2282 GND.n2273 5246.88
R2202 GND.n2247 GND.n2242 5246.88
R2203 GND.n2273 GND.n2242 5246.88
R2204 GND.n2284 GND.n2240 5246.88
R2205 GND.n2284 GND.n2241 5246.88
R2206 GND.n2243 GND.n2240 5246.88
R2207 GND.n2243 GND.n2241 5246.88
R2208 GND.n2604 GND.n2569 5246.88
R2209 GND.n2604 GND.n2595 5246.88
R2210 GND.n2569 GND.n2564 5246.88
R2211 GND.n2595 GND.n2564 5246.88
R2212 GND.n2606 GND.n2562 5246.88
R2213 GND.n2606 GND.n2563 5246.88
R2214 GND.n2565 GND.n2562 5246.88
R2215 GND.n2565 GND.n2563 5246.88
R2216 GND.n2725 GND.n2690 5246.88
R2217 GND.n2725 GND.n2716 5246.88
R2218 GND.n2690 GND.n2685 5246.88
R2219 GND.n2716 GND.n2685 5246.88
R2220 GND.n2727 GND.n2683 5246.88
R2221 GND.n2727 GND.n2684 5246.88
R2222 GND.n2686 GND.n2683 5246.88
R2223 GND.n2686 GND.n2684 5246.88
R2224 GND.n1053 GND.n1048 5246.88
R2225 GND.n1053 GND.n1049 5246.88
R2226 GND.n1582 GND.n1048 5246.88
R2227 GND.n1582 GND.n1049 5246.88
R2228 GND.n1336 GND.n1335 4207.44
R2229 GND.n1001 GND.n1000 4207.44
R2230 GND.n1691 GND.n1690 4207.44
R2231 GND.n1547 GND.n1546 4207.44
R2232 GND.n1487 GND.n1486 4207.44
R2233 GND.n1257 GND.n1256 4207.44
R2234 GND.n2086 GND.n2085 4207.44
R2235 GND.n2003 GND.n2002 4207.44
R2236 GND.n4056 GND.n168 3522.26
R2237 GND.n3830 GND.n168 3522.26
R2238 GND.n4056 GND.n169 3522.26
R2239 GND.n3830 GND.n169 3522.26
R2240 GND.n4151 GND.n109 3522.26
R2241 GND.n3677 GND.n109 3522.26
R2242 GND.n4151 GND.n110 3522.26
R2243 GND.n3677 GND.n110 3522.26
R2244 GND.n4041 GND.n177 3522.26
R2245 GND.n4037 GND.n177 3522.26
R2246 GND.n4041 GND.n178 3522.26
R2247 GND.n4037 GND.n178 3522.26
R2248 GND.n4091 GND.n147 3522.26
R2249 GND.n4087 GND.n147 3522.26
R2250 GND.n4091 GND.n148 3522.26
R2251 GND.n4087 GND.n148 3522.26
R2252 GND.n4136 GND.n119 3522.26
R2253 GND.n4132 GND.n119 3522.26
R2254 GND.n4136 GND.n120 3522.26
R2255 GND.n4132 GND.n120 3522.26
R2256 GND.n3610 GND.n327 3522.26
R2257 GND.n3621 GND.n327 3522.26
R2258 GND.n3610 GND.n328 3522.26
R2259 GND.n3621 GND.n328 3522.26
R2260 GND.n3595 GND.n343 3522.26
R2261 GND.n3591 GND.n343 3522.26
R2262 GND.n3595 GND.n344 3522.26
R2263 GND.n3591 GND.n344 3522.26
R2264 GND.n4191 GND.n70 3522.26
R2265 GND.n79 GND.n70 3522.26
R2266 GND.n4191 GND.n71 3522.26
R2267 GND.n79 GND.n71 3522.26
R2268 GND.n4220 GND.n49 3522.26
R2269 GND.n58 GND.n49 3522.26
R2270 GND.n4220 GND.n50 3522.26
R2271 GND.n58 GND.n50 3522.26
R2272 GND.n3048 GND.n2145 3522.26
R2273 GND.n3033 GND.n2145 3522.26
R2274 GND.n3048 GND.n2146 3522.26
R2275 GND.n3033 GND.n2146 3522.26
R2276 GND.n3184 GND.n541 3522.26
R2277 GND.n3188 GND.n541 3522.26
R2278 GND.n3184 GND.n542 3522.26
R2279 GND.n3188 GND.n542 3522.26
R2280 GND.n3133 GND.n561 3522.26
R2281 GND.n3144 GND.n561 3522.26
R2282 GND.n3133 GND.n562 3522.26
R2283 GND.n3144 GND.n562 3522.26
R2284 GND.n3085 GND.n604 3522.26
R2285 GND.n617 GND.n604 3522.26
R2286 GND.n3085 GND.n605 3522.26
R2287 GND.n617 GND.n605 3522.26
R2288 GND.n3118 GND.n577 3522.26
R2289 GND.n3114 GND.n577 3522.26
R2290 GND.n3118 GND.n578 3522.26
R2291 GND.n3114 GND.n578 3522.26
R2292 GND.n1577 GND.n1040 3522.26
R2293 GND.n1591 GND.n1040 3522.26
R2294 GND.n1577 GND.n1041 3522.26
R2295 GND.n1591 GND.n1041 3522.26
R2296 GND.n1957 GND.n842 3522.26
R2297 GND.n1937 GND.n842 3522.26
R2298 GND.n1937 GND.n843 3522.26
R2299 GND.n1957 GND.n843 3522.26
R2300 GND.n1411 GND.n1371 3522.26
R2301 GND.n1375 GND.n1371 3522.26
R2302 GND.n1411 GND.n1372 3522.26
R2303 GND.n1375 GND.n1372 3522.26
R2304 GND.n1987 GND.n824 3522.26
R2305 GND.n1983 GND.n824 3522.26
R2306 GND.n1987 GND.n825 3522.26
R2307 GND.n1983 GND.n825 3522.26
R2308 GND.n2040 GND.n783 3522.26
R2309 GND.n790 GND.n783 3522.26
R2310 GND.n2040 GND.n784 3522.26
R2311 GND.n790 GND.n784 3522.26
R2312 GND.n746 GND.n714 3522.26
R2313 GND.n749 GND.n714 3522.26
R2314 GND.n746 GND.n712 3522.26
R2315 GND.n749 GND.n712 3522.26
R2316 GND.n2070 GND.n693 3522.26
R2317 GND.n2066 GND.n693 3522.26
R2318 GND.n2070 GND.n694 3522.26
R2319 GND.n2066 GND.n694 3522.26
R2320 GND.n2123 GND.n652 3522.26
R2321 GND.n659 GND.n652 3522.26
R2322 GND.n2123 GND.n653 3522.26
R2323 GND.n659 GND.n653 3522.26
R2324 GND.n1209 GND.n1207 3522.26
R2325 GND.n1273 GND.n1207 3522.26
R2326 GND.n1272 GND.n1209 3522.26
R2327 GND.n1273 GND.n1272 3522.26
R2328 GND.n1188 GND.n1186 3522.26
R2329 GND.n1352 GND.n1186 3522.26
R2330 GND.n1351 GND.n1188 3522.26
R2331 GND.n1352 GND.n1351 3522.26
R2332 GND.n1721 GND.n871 3522.26
R2333 GND.n1056 GND.n871 3522.26
R2334 GND.n1721 GND.n872 3522.26
R2335 GND.n1056 GND.n872 3522.26
R2336 GND.n1124 GND.n1082 3522.26
R2337 GND.n1096 GND.n1082 3522.26
R2338 GND.n1124 GND.n1083 3522.26
R2339 GND.n1096 GND.n1083 3522.26
R2340 GND.n1645 GND.n921 3522.26
R2341 GND.n1021 GND.n921 3522.26
R2342 GND.n1645 GND.n922 3522.26
R2343 GND.n1021 GND.n922 3522.26
R2344 GND.n1015 GND.n934 3522.26
R2345 GND.n1623 GND.n934 3522.26
R2346 GND.n1015 GND.n936 3522.26
R2347 GND.n1623 GND.n936 3522.26
R2348 GND.n1675 GND.n904 3522.26
R2349 GND.n1671 GND.n904 3522.26
R2350 GND.n1675 GND.n905 3522.26
R2351 GND.n1671 GND.n905 3522.26
R2352 GND.n1562 GND.n1144 3522.26
R2353 GND.n1566 GND.n1144 3522.26
R2354 GND.n1562 GND.n1145 3522.26
R2355 GND.n1566 GND.n1145 3522.26
R2356 GND.n1501 GND.n1165 3522.26
R2357 GND.n1504 GND.n1165 3522.26
R2358 GND.n1501 GND.n1167 3522.26
R2359 GND.n1504 GND.n1167 3522.26
R2360 GND.n3212 GND.n3210 3522.26
R2361 GND.n3246 GND.n3210 3522.26
R2362 GND.n3213 GND.n3212 3522.26
R2363 GND.n3246 GND.n3213 3522.26
R2364 GND.n3281 GND.n498 3522.26
R2365 GND.n3292 GND.n498 3522.26
R2366 GND.n3281 GND.n499 3522.26
R2367 GND.n3292 GND.n499 3522.26
R2368 GND.n3503 GND.n3471 3522.26
R2369 GND.n3481 GND.n3471 3522.26
R2370 GND.n3503 GND.n3472 3522.26
R2371 GND.n3481 GND.n3472 3522.26
R2372 GND.n3529 GND.n368 3522.26
R2373 GND.n3533 GND.n368 3522.26
R2374 GND.n3529 GND.n369 3522.26
R2375 GND.n3533 GND.n369 3522.26
R2376 GND.n425 GND.n423 3522.26
R2377 GND.n482 GND.n423 3522.26
R2378 GND.n426 GND.n425 3522.26
R2379 GND.n482 GND.n426 3522.26
R2380 GND.n3356 GND.n3355 3522.26
R2381 GND.n3387 GND.n3356 3522.26
R2382 GND.n3355 GND.n3353 3522.26
R2383 GND.n3387 GND.n3353 3522.26
R2384 GND.n3410 GND.n392 3522.26
R2385 GND.n3421 GND.n392 3522.26
R2386 GND.n3410 GND.n393 3522.26
R2387 GND.n3421 GND.n393 3522.26
R2388 GND.n3890 GND.n237 3522.26
R2389 GND.n3924 GND.n237 3522.26
R2390 GND.n3890 GND.n235 3522.26
R2391 GND.n3924 GND.n235 3522.26
R2392 GND.n3846 GND.n252 3522.26
R2393 GND.n3857 GND.n252 3522.26
R2394 GND.n3846 GND.n253 3522.26
R2395 GND.n3857 GND.n253 3522.26
R2396 GND.n3737 GND.n287 3522.26
R2397 GND.n3762 GND.n287 3522.26
R2398 GND.n3737 GND.n285 3522.26
R2399 GND.n3762 GND.n285 3522.26
R2400 GND.n3693 GND.n302 3522.26
R2401 GND.n3704 GND.n302 3522.26
R2402 GND.n3693 GND.n303 3522.26
R2403 GND.n3704 GND.n303 3522.26
R2404 GND.n3172 GND.n12 3522.26
R2405 GND.n4281 GND.n12 3522.26
R2406 GND.n3172 GND.n10 3522.26
R2407 GND.n4281 GND.n10 3522.26
R2408 GND.n521 GND.n518 3522.26
R2409 GND.n526 GND.n518 3522.26
R2410 GND.n521 GND.n519 3522.26
R2411 GND.n526 GND.n519 3522.26
R2412 GND.n2993 GND.n2167 3522.26
R2413 GND.n2997 GND.n2167 3522.26
R2414 GND.n2993 GND.n2168 3522.26
R2415 GND.n2997 GND.n2168 3522.26
R2416 GND.n2845 GND.n2474 3522.26
R2417 GND.n2485 GND.n2474 3522.26
R2418 GND.n2845 GND.n2475 3522.26
R2419 GND.n2485 GND.n2475 3522.26
R2420 GND.n2774 GND.n2499 3522.26
R2421 GND.n2778 GND.n2499 3522.26
R2422 GND.n2774 GND.n2500 3522.26
R2423 GND.n2778 GND.n2500 3522.26
R2424 GND.n2952 GND.n2890 3522.26
R2425 GND.n2903 GND.n2890 3522.26
R2426 GND.n2952 GND.n2891 3522.26
R2427 GND.n2903 GND.n2891 3522.26
R2428 GND.n2985 GND.n2173 3522.26
R2429 GND.n2981 GND.n2173 3522.26
R2430 GND.n2985 GND.n2174 3522.26
R2431 GND.n2981 GND.n2174 3522.26
R2432 GND.n2420 GND.n2358 3522.26
R2433 GND.n2371 GND.n2358 3522.26
R2434 GND.n2420 GND.n2359 3522.26
R2435 GND.n2371 GND.n2359 3522.26
R2436 GND.n2451 GND.n2332 3522.26
R2437 GND.n2451 GND.n2333 3522.26
R2438 GND.n2450 GND.n2332 3522.26
R2439 GND.n2450 GND.n2333 3522.26
R2440 GND.n2293 GND.n2231 3522.26
R2441 GND.n2244 GND.n2231 3522.26
R2442 GND.n2293 GND.n2232 3522.26
R2443 GND.n2244 GND.n2232 3522.26
R2444 GND.n2324 GND.n2204 3522.26
R2445 GND.n2324 GND.n2205 3522.26
R2446 GND.n2323 GND.n2204 3522.26
R2447 GND.n2323 GND.n2205 3522.26
R2448 GND.n2615 GND.n2553 3522.26
R2449 GND.n2566 GND.n2553 3522.26
R2450 GND.n2615 GND.n2554 3522.26
R2451 GND.n2566 GND.n2554 3522.26
R2452 GND.n2646 GND.n2526 3522.26
R2453 GND.n2646 GND.n2527 3522.26
R2454 GND.n2645 GND.n2526 3522.26
R2455 GND.n2645 GND.n2527 3522.26
R2456 GND.n2736 GND.n2674 3522.26
R2457 GND.n2687 GND.n2674 3522.26
R2458 GND.n2736 GND.n2675 3522.26
R2459 GND.n2687 GND.n2675 3522.26
R2460 GND.n2769 GND.n2507 3522.26
R2461 GND.n2765 GND.n2507 3522.26
R2462 GND.n2769 GND.n2508 3522.26
R2463 GND.n2765 GND.n2508 3522.26
R2464 GND.n3996 GND.n205 3522.26
R2465 GND.n3992 GND.n205 3522.26
R2466 GND.n3996 GND.n206 3522.26
R2467 GND.n3992 GND.n206 3522.26
R2468 GND.n1621 GND.n1030 3443.83
R2469 GND.n1669 GND.n1668 3097.63
R2470 GND.n1744 GND.n858 3097.63
R2471 GND.n2101 GND.n2100 3097.63
R2472 GND.n2018 GND.n2017 3097.63
R2473 GND.n2989 GND.n2988 3081.57
R2474 GND.t626 GND.t360 2955.8
R2475 GND.t626 GND.t511 2955.8
R2476 GND.t32 GND.t659 2955.8
R2477 GND.t659 GND.t489 2955.8
R2478 GND.t301 GND.t720 2955.8
R2479 GND.t720 GND.t825 2955.8
R2480 GND.t41 GND.t708 2955.8
R2481 GND.t41 GND.t166 2955.8
R2482 GND.t372 GND.t760 2955.8
R2483 GND.t760 GND.t126 2955.8
R2484 GND.t17 GND.t676 2955.8
R2485 GND.t676 GND.t562 2955.8
R2486 GND.t471 GND.t188 2955.8
R2487 GND.t471 GND.t499 2955.8
R2488 GND.t214 GND.t369 2955.8
R2489 GND.t525 GND.t214 2955.8
R2490 GND.t762 GND.t843 2955.8
R2491 GND.t174 GND.t762 2955.8
R2492 GND.t403 GND.t276 2955.8
R2493 GND.t276 GND.t574 2955.8
R2494 GND.t310 GND.t93 2955.8
R2495 GND.t93 GND.t580 2955.8
R2496 GND.t450 GND.t797 2955.8
R2497 GND.t797 GND.t831 2955.8
R2498 GND.t280 GND.t42 2955.8
R2499 GND.t280 GND.t519 2955.8
R2500 GND.t285 GND.t866 2955.8
R2501 GND.t866 GND.t550 2955.8
R2502 GND.t415 GND.t638 2955.8
R2503 GND.t638 GND.t114 2955.8
R2504 GND.t441 GND.t570 2955.8
R2505 GND.t441 GND.t77 2955.8
R2506 GND.t182 GND.t827 2955.8
R2507 GND.t315 GND.t182 2955.8
R2508 GND.t162 GND.t745 2955.8
R2509 GND.t745 GND.t810 2955.8
R2510 GND.t731 GND.t509 2955.8
R2511 GND.t381 GND.t731 2955.8
R2512 GND.t710 GND.t146 2955.8
R2513 GND.t243 GND.t710 2955.8
R2514 GND.t144 GND.t775 2955.8
R2515 GND.t775 GND.t686 2955.8
R2516 GND.t623 GND.t533 2955.8
R2517 GND.t623 GND.t297 2955.8
R2518 GND.t770 GND.t833 2955.8
R2519 GND.t54 GND.t770 2955.8
R2520 GND.t164 GND.t769 2955.8
R2521 GND.t769 GND.t99 2955.8
R2522 GND.t258 GND.t546 2955.8
R2523 GND.t258 GND.t382 2955.8
R2524 GND.t634 GND.t148 2955.8
R2525 GND.t634 GND.t61 2955.8
R2526 GND.t102 GND.t217 2955.8
R2527 GND.t217 GND.t194 2955.8
R2528 GND.t809 GND.t578 2955.8
R2529 GND.t809 GND.t76 2955.8
R2530 GND.t591 GND.t120 2955.8
R2531 GND.t881 GND.t591 2955.8
R2532 GND.t813 GND.t220 2955.8
R2533 GND.t220 GND.t592 2955.8
R2534 GND.t191 GND.t523 2955.8
R2535 GND.t191 GND.t300 2955.8
R2536 GND.t759 GND.t170 2955.8
R2537 GND.t759 GND.t609 2955.8
R2538 GND.t71 GND.t122 2955.8
R2539 GND.t677 GND.t71 2955.8
R2540 GND.t611 GND.t529 2955.8
R2541 GND.t611 GND.t298 2955.8
R2542 GND.t190 GND.t815 2955.8
R2543 GND.t190 GND.t85 2955.8
R2544 GND.t218 GND.t118 2955.8
R2545 GND.t359 GND.t218 2955.8
R2546 GND.t867 GND.t544 2955.8
R2547 GND.t867 GND.t322 2955.8
R2548 GND.t287 GND.t150 2955.8
R2549 GND.t600 GND.t287 2955.8
R2550 GND.t647 GND.t168 2955.8
R2551 GND.t647 GND.t706 2955.8
R2552 GND.t211 GND.t212 2955.8
R2553 GND.t211 GND.t568 2955.8
R2554 GND.t348 GND.t286 2955.8
R2555 GND.t286 GND.t517 2955.8
R2556 GND.t417 GND.t395 2955.8
R2557 GND.t395 GND.t158 2955.8
R2558 GND.t474 GND.t805 2955.8
R2559 GND.t497 GND.t474 2955.8
R2560 GND.t198 GND.t342 2955.8
R2561 GND.t566 GND.t198 2955.8
R2562 GND.t800 GND.t68 2955.8
R2563 GND.t134 GND.t800 2955.8
R2564 GND.t38 GND.t364 2955.8
R2565 GND.t556 GND.t38 2955.8
R2566 GND.t321 GND.t234 2955.8
R2567 GND.t479 GND.t321 2955.8
R2568 GND.t692 GND.t327 2955.8
R2569 GND.t172 GND.t692 2955.8
R2570 GND.t755 GND.t485 2955.8
R2571 GND.t755 GND.t307 2955.8
R2572 GND.t733 GND.t116 2955.8
R2573 GND.t628 GND.t733 2955.8
R2574 GND.t178 GND.t94 2955.8
R2575 GND.t94 GND.t272 2955.8
R2576 GND.n1668 GND.n908 2528.02
R2577 GND.n1745 GND.n1744 2528.02
R2578 GND.n2102 GND.n2101 2528.02
R2579 GND.n2019 GND.n2018 2528.02
R2580 GND.n1568 GND.n1143 2291.01
R2581 GND.n2064 GND.n2063 2291.01
R2582 GND.n1981 GND.n1980 2291.01
R2583 GND.n3728 GND.n3727 2152.7
R2584 GND.n3833 GND.n3829 2152.7
R2585 GND.n3881 GND.n3880 2152.7
R2586 GND.n3680 GND.n3676 2152.7
R2587 GND.n3183 GND.n3182 1937.25
R2588 GND.n4117 GND.n4116 1847.07
R2589 GND.n4072 GND.n4071 1847.07
R2590 GND.n4022 GND.n4021 1847.07
R2591 GND.n3977 GND.n3976 1847.07
R2592 GND.n1569 GND.n1568 1797.97
R2593 GND.n2064 GND.n696 1797.97
R2594 GND.n1981 GND.n827 1797.97
R2595 GND.n3903 GND.t677 1542.9
R2596 GND.t438 GND.t542 1540.25
R2597 GND.t438 GND.t330 1540.25
R2598 GND.t465 GND.t237 1540.25
R2599 GND.t465 GND.t368 1540.25
R2600 GND.t365 GND.t384 1540.25
R2601 GND.t365 GND.t90 1540.25
R2602 GND.t95 GND.t239 1540.25
R2603 GND.t95 GND.t622 1540.25
R2604 GND.t713 GND.t749 1540.25
R2605 GND.t713 GND.t199 1540.25
R2606 GND.t350 GND.t235 1540.25
R2607 GND.t350 GND.t207 1540.25
R2608 GND.t383 GND.t389 1540.25
R2609 GND.t383 GND.t596 1540.25
R2610 GND.t87 GND.t427 1540.25
R2611 GND.t87 GND.t267 1540.25
R2612 GND.t55 GND.t651 1540.25
R2613 GND.t55 GND.t375 1540.25
R2614 GND.t437 GND.t241 1540.25
R2615 GND.t437 GND.t251 1540.25
R2616 GND.t711 GND.t273 1540.25
R2617 GND.t711 GND.t37 1540.25
R2618 GND.t725 GND.t5 1540.25
R2619 GND.t725 GND.t50 1540.25
R2620 GND.t633 GND.t649 1540.25
R2621 GND.t633 GND.t46 1540.25
R2622 GND.t75 GND.t27 1540.25
R2623 GND.t75 GND.t803 1540.25
R2624 GND.t470 GND.t422 1540.25
R2625 GND.t470 GND.t288 1540.25
R2626 GND.t699 GND.t270 1540.25
R2627 GND.t699 GND.t792 1540.25
R2628 GND.t255 GND.t338 1540.25
R2629 GND.t255 GND.t254 1540.25
R2630 GND.t462 GND.t9 1540.25
R2631 GND.t462 GND.t754 1540.25
R2632 GND.t360 GND.n697 1477.9
R2633 GND.n1327 GND.t511 1477.9
R2634 GND.n1329 GND.t413 1477.9
R2635 GND.t413 GND.n1328 1477.9
R2636 GND.n1328 GND.t410 1477.9
R2637 GND.n1335 GND.t410 1477.9
R2638 GND.n1336 GND.t32 1477.9
R2639 GND.n1342 GND.t489 1477.9
R2640 GND.n1343 GND.t301 1477.9
R2641 GND.n1349 GND.t825 1477.9
R2642 GND.t721 GND.n1350 1477.9
R2643 GND.t721 GND.n805 1477.9
R2644 GND.t708 GND.n907 1477.9
R2645 GND.n992 GND.t166 1477.9
R2646 GND.n994 GND.t351 1477.9
R2647 GND.t351 GND.n993 1477.9
R2648 GND.n993 GND.t859 1477.9
R2649 GND.n1000 GND.t859 1477.9
R2650 GND.n1001 GND.t372 1477.9
R2651 GND.n1007 GND.t126 1477.9
R2652 GND.n1008 GND.t17 1477.9
R2653 GND.n1014 GND.t562 1477.9
R2654 GND.t641 GND.n1016 1477.9
R2655 GND.n1622 GND.t641 1477.9
R2656 GND.n1068 GND.t188 1477.9
R2657 GND.t499 GND.n1065 1477.9
R2658 GND.n1064 GND.t715 1477.9
R2659 GND.n1692 GND.t715 1477.9
R2660 GND.n1692 GND.t870 1477.9
R2661 GND.t870 GND.n1691 1477.9
R2662 GND.n1690 GND.t369 1477.9
R2663 GND.n1684 GND.t525 1477.9
R2664 GND.n1683 GND.t843 1477.9
R2665 GND.n1677 GND.t174 1477.9
R2666 GND.n1676 GND.t386 1477.9
R2667 GND.n1670 GND.t386 1477.9
R2668 GND.n1532 GND.t403 1477.9
R2669 GND.n1538 GND.t574 1477.9
R2670 GND.n1540 GND.t588 1477.9
R2671 GND.t588 GND.n1539 1477.9
R2672 GND.n1539 GND.t311 1477.9
R2673 GND.n1546 GND.t311 1477.9
R2674 GND.n1547 GND.t310 1477.9
R2675 GND.n1553 GND.t580 1477.9
R2676 GND.n1554 GND.t450 1477.9
R2677 GND.n1560 GND.t831 1477.9
R2678 GND.n1561 GND.t406 1477.9
R2679 GND.n1567 GND.t406 1477.9
R2680 GND.t42 GND.n828 1477.9
R2681 GND.n1478 GND.t519 1477.9
R2682 GND.n1480 GND.t269 1477.9
R2683 GND.t269 GND.n1479 1477.9
R2684 GND.n1479 GND.t787 1477.9
R2685 GND.n1486 GND.t787 1477.9
R2686 GND.n1487 GND.t285 1477.9
R2687 GND.n1493 GND.t550 1477.9
R2688 GND.n1494 GND.t415 1477.9
R2689 GND.n1500 GND.t114 1477.9
R2690 GND.t751 GND.n1502 1477.9
R2691 GND.n1503 GND.t751 1477.9
R2692 GND.t570 GND.n3398 1477.9
R2693 GND.t77 GND.n401 1477.9
R2694 GND.t827 GND.n3409 1477.9
R2695 GND.n3412 GND.t315 1477.9
R2696 GND.n3411 GND.t446 1477.9
R2697 GND.n3422 GND.t446 1477.9
R2698 GND.n3424 GND.t281 1477.9
R2699 GND.t281 GND.n3423 1477.9
R2700 GND.n3423 GND.t808 1477.9
R2701 GND.n3433 GND.t808 1477.9
R2702 GND.n3434 GND.t162 1477.9
R2703 GND.n3444 GND.t810 1477.9
R2704 GND.n3526 GND.t509 1477.9
R2705 GND.n3516 GND.t381 1477.9
R2706 GND.n3515 GND.t146 1477.9
R2707 GND.n3505 GND.t243 1477.9
R2708 GND.n3504 GND.t840 1477.9
R2709 GND.n3482 GND.t840 1477.9
R2710 GND.t246 GND.n3483 1477.9
R2711 GND.n3494 GND.t246 1477.9
R2712 GND.n3494 GND.t637 1477.9
R2713 GND.t637 GND.n3490 1477.9
R2714 GND.n3489 GND.t144 1477.9
R2715 GND.n3573 GND.t686 1477.9
R2716 GND.t533 GND.n3681 1477.9
R2717 GND.t297 GND.n311 1477.9
R2718 GND.t833 GND.n3692 1477.9
R2719 GND.n3695 GND.t54 1477.9
R2720 GND.n3694 GND.t453 1477.9
R2721 GND.n3705 GND.t453 1477.9
R2722 GND.n3707 GND.t682 1477.9
R2723 GND.t682 GND.n3706 1477.9
R2724 GND.n3706 GND.t392 1477.9
R2725 GND.n3716 GND.t392 1477.9
R2726 GND.n3717 GND.t164 1477.9
R2727 GND.n3727 GND.t99 1477.9
R2728 GND.t546 GND.n3729 1477.9
R2729 GND.n3732 GND.t382 1477.9
R2730 GND.t148 GND.n3733 1477.9
R2731 GND.n3736 GND.t61 1477.9
R2732 GND.t224 GND.n3738 1477.9
R2733 GND.n3761 GND.t224 1477.9
R2734 GND.n3760 GND.t227 1477.9
R2735 GND.n3744 GND.t227 1477.9
R2736 GND.t376 GND.n3744 1477.9
R2737 GND.n3751 GND.t376 1477.9
R2738 GND.n3750 GND.t102 1477.9
R2739 GND.n3829 GND.t194 1477.9
R2740 GND.t578 GND.n3834 1477.9
R2741 GND.t76 GND.n261 1477.9
R2742 GND.t120 GND.n3845 1477.9
R2743 GND.n3848 GND.t881 1477.9
R2744 GND.n3847 GND.t18 1477.9
R2745 GND.n3858 GND.t18 1477.9
R2746 GND.n3860 GND.t362 1477.9
R2747 GND.t362 GND.n3859 1477.9
R2748 GND.n3859 GND.t63 1477.9
R2749 GND.n3869 GND.t63 1477.9
R2750 GND.n3870 GND.t813 1477.9
R2751 GND.n3880 GND.t592 1477.9
R2752 GND.t523 GND.n3882 1477.9
R2753 GND.n3885 GND.t300 1477.9
R2754 GND.t170 GND.n3886 1477.9
R2755 GND.n3889 GND.t609 1477.9
R2756 GND.t457 GND.n3891 1477.9
R2757 GND.n3923 GND.t457 1477.9
R2758 GND.n3922 GND.t277 1477.9
R2759 GND.n3897 GND.t277 1477.9
R2760 GND.t599 GND.n3897 1477.9
R2761 GND.n3913 GND.t599 1477.9
R2762 GND.n3912 GND.t122 1477.9
R2763 GND.n3181 GND.t529 1477.9
R2764 GND.t298 GND.n3178 1477.9
R2765 GND.n3177 GND.t815 1477.9
R2766 GND.t85 GND.n3174 1477.9
R2767 GND.n3173 GND.t295 1477.9
R2768 GND.n4280 GND.t295 1477.9
R2769 GND.n4279 GND.t39 1477.9
R2770 GND.n18 GND.t39 1477.9
R2771 GND.t879 GND.n18 1477.9
R2772 GND.n4270 GND.t879 1477.9
R2773 GND.n4269 GND.t118 1477.9
R2774 GND.n4259 GND.t359 1477.9
R2775 GND.t544 GND.n3269 1477.9
R2776 GND.t322 GND.n507 1477.9
R2777 GND.t150 GND.n3280 1477.9
R2778 GND.n3283 GND.t600 1477.9
R2779 GND.n3282 GND.t459 1477.9
R2780 GND.n3293 GND.t459 1477.9
R2781 GND.n3295 GND.t601 1477.9
R2782 GND.t601 GND.n3294 1477.9
R2783 GND.n3294 GND.t882 1477.9
R2784 GND.n3308 GND.t882 1477.9
R2785 GND.t168 GND.n3309 1477.9
R2786 GND.t706 GND.n412 1477.9
R2787 GND.t212 GND.n640 1477.9
R2788 GND.n1248 GND.t568 1477.9
R2789 GND.n1250 GND.t337 1477.9
R2790 GND.t337 GND.n1249 1477.9
R2791 GND.n1249 GND.t64 1477.9
R2792 GND.n1256 GND.t64 1477.9
R2793 GND.n1257 GND.t348 1477.9
R2794 GND.n1263 GND.t517 1477.9
R2795 GND.n1264 GND.t417 1477.9
R2796 GND.n1270 GND.t158 1477.9
R2797 GND.t612 GND.n1271 1477.9
R2798 GND.t612 GND.n674 1477.9
R2799 GND.n2099 GND.t805 1477.9
R2800 GND.n2093 GND.t497 1477.9
R2801 GND.n2092 GND.t378 1477.9
R2802 GND.n684 GND.t378 1477.9
R2803 GND.t256 GND.n684 1477.9
R2804 GND.n2086 GND.t256 1477.9
R2805 GND.n2085 GND.t342 1477.9
R2806 GND.n2079 GND.t566 1477.9
R2807 GND.n2078 GND.t68 1477.9
R2808 GND.n2072 GND.t134 1477.9
R2809 GND.n2071 GND.t798 1477.9
R2810 GND.n2065 GND.t798 1477.9
R2811 GND.n2016 GND.t364 1477.9
R2812 GND.n2010 GND.t556 1477.9
R2813 GND.n2009 GND.t586 1477.9
R2814 GND.n815 GND.t586 1477.9
R2815 GND.t689 GND.n815 1477.9
R2816 GND.n2003 GND.t689 1477.9
R2817 GND.n2002 GND.t234 1477.9
R2818 GND.n1996 GND.t479 1477.9
R2819 GND.n1995 GND.t327 1477.9
R2820 GND.n1989 GND.t172 1477.9
R2821 GND.n1988 GND.t23 1477.9
R2822 GND.n1982 GND.t23 1477.9
R2823 GND.t485 GND.n3598 1477.9
R2824 GND.t307 GND.n336 1477.9
R2825 GND.t116 GND.n3609 1477.9
R2826 GND.n3612 GND.t628 1477.9
R2827 GND.n3611 GND.t13 1477.9
R2828 GND.n3622 GND.t13 1477.9
R2829 GND.n3624 GND.t782 1477.9
R2830 GND.t782 GND.n3623 1477.9
R2831 GND.n3623 GND.t223 1477.9
R2832 GND.n3633 GND.t223 1477.9
R2833 GND.n3634 GND.t178 1477.9
R2834 GND.n3676 GND.t272 1477.9
R2835 GND.t643 GND.t513 1297.6
R2836 GND.t409 GND.t643 1297.6
R2837 GND.t662 GND.t124 1297.6
R2838 GND.t323 GND.t662 1297.6
R2839 GND.t36 GND.t477 1297.6
R2840 GND.t684 GND.t36 1297.6
R2841 GND.t880 GND.t537 1297.6
R2842 GND.t776 GND.t880 1297.6
R2843 GND.t98 GND.t104 1297.6
R2844 GND.t261 GND.t98 1297.6
R2845 GND.t408 GND.t554 1297.6
R2846 GND.t734 GND.t493 1297.6
R2847 GND.t349 GND.t734 1297.6
R2848 GND.t855 GND.t817 1297.6
R2849 GND.t448 GND.t855 1297.6
R2850 GND.t839 GND.t475 1297.6
R2851 GND.t208 GND.t839 1297.6
R2852 GND.t352 GND.t507 1297.6
R2853 GND.t640 GND.t352 1297.6
R2854 GND.t291 GND.t132 1297.6
R2855 GND.t842 GND.t291 1297.6
R2856 GND.t45 GND.t527 1297.6
R2857 GND.t473 GND.t576 1297.6
R2858 GND.t268 GND.t473 1297.6
R2859 GND.n467 GND.n466 1297.44
R2860 GND.n3558 GND.n69 1297.44
R2861 GND.n3330 GND.n48 1297.44
R2862 GND.n4244 GND.n4242 1297.44
R2863 GND.n4103 GND.n4102 1246.88
R2864 GND.n4093 GND.n4092 1246.88
R2865 GND.n4008 GND.n4007 1246.88
R2866 GND.n3998 GND.n3997 1246.88
R2867 GND.n1621 GND.n1620 1235.69
R2868 GND.t464 GND.t388 1230.8
R2869 GND.t491 GND.t464 1230.8
R2870 GND.t732 GND.t878 1230.8
R2871 GND.t732 GND.t521 1230.8
R2872 GND.t213 GND.t262 1230.8
R2873 GND.t213 GND.t154 1230.8
R2874 GND.t691 GND.t796 1230.8
R2875 GND.t110 GND.t691 1230.8
R2876 GND.t176 GND.t712 1230.8
R2877 GND.t466 GND.t304 1230.8
R2878 GND.t466 GND.t572 1230.8
R2879 GND.t88 GND.t753 1230.8
R2880 GND.t138 GND.t88 1230.8
R2881 GND.t709 GND.t219 1230.8
R2882 GND.t219 GND.t136 1230.8
R2883 GND.t864 GND.t67 1230.8
R2884 GND.t864 GND.t548 1230.8
R2885 GND.t767 GND.t292 1230.8
R2886 GND.t660 GND.t875 1230.8
R2887 GND.t140 GND.t660 1230.8
R2888 GND.t823 GND.t774 1230.8
R2889 GND.t345 GND.t293 1230.8
R2890 GND.t501 GND.t345 1230.8
R2891 GND.t730 GND.t60 1230.8
R2892 GND.t730 GND.t112 1230.8
R2893 GND.t635 GND.t405 1230.8
R2894 GND.t635 GND.t142 1230.8
R2895 GND.t433 GND.t380 1230.8
R2896 GND.t433 GND.t515 1230.8
R2897 GND.t440 GND.t802 1230.8
R2898 GND.t829 GND.t440 1230.8
R2899 GND.t130 GND.t404 1230.8
R2900 GND.t780 GND.t20 1230.8
R2901 GND.t558 GND.t780 1230.8
R2902 GND.t221 GND.t724 1230.8
R2903 GND.t221 GND.t156 1230.8
R2904 GND.t56 GND.t688 1230.8
R2905 GND.t56 GND.t108 1230.8
R2906 GND.t472 GND.t461 1230.8
R2907 GND.t472 GND.t487 1230.8
R2908 GND.t604 GND.t693 1230.8
R2909 GND.t604 GND.t821 1230.8
R2910 GND.n2528 GND.n576 1216.65
R2911 GND.n2771 GND.n2770 1216.65
R2912 GND.n3120 GND.n3119 1216.65
R2913 GND.t204 GND.t206 1201.24
R2914 GND.t206 GND.t868 1201.24
R2915 GND.n1035 GND.t408 1041.88
R2916 GND.n2101 GND.n673 1036.63
R2917 GND.n2018 GND.n804 1036.63
R2918 GND.n1668 GND.n1667 1036.63
R2919 GND.n1744 GND.n1743 1036.63
R2920 GND.n3182 GND.n3167 1017.54
R2921 GND.t316 GND.t318 1004.31
R2922 GND.t318 GND.t765 1004.31
R2923 GND.t47 GND.t49 1004.31
R2924 GND.t49 GND.t185 1004.31
R2925 GND.t701 GND.t703 1004.31
R2926 GND.t703 GND.t100 1004.31
R2927 GND.t777 GND.t779 1002.82
R2928 GND.t779 GND.t605 1002.82
R2929 GND.n1606 GND.t712 988.246
R2930 GND.n4234 GND.t774 988.246
R2931 GND.n4205 GND.t404 988.246
R2932 GND.n1620 GND.t45 948.895
R2933 GND.t670 GND.t819 911.471
R2934 GND.t449 GND.t670 911.471
R2935 GND.t503 GND.t354 911.471
R2936 GND.t539 GND.t582 911.471
R2937 GND.t582 GND.t773 911.471
R2938 GND.t152 GND.t26 911.471
R2939 GND.t26 GND.t226 911.471
R2940 GND.t617 GND.t560 911.471
R2941 GND.t617 GND.t248 911.471
R2942 GND.t564 GND.t197 911.471
R2943 GND.t197 GND.t627 911.471
R2944 GND.t357 GND.t106 911.471
R2945 GND.t414 GND.t357 911.471
R2946 GND.t756 GND.t552 911.471
R2947 GND.t756 GND.t603 911.471
R2948 GND.t531 GND.t707 911.471
R2949 GND.t707 GND.t585 911.471
R2950 GND.t654 GND.t128 911.471
R2951 GND.t654 GND.t326 911.471
R2952 GND.t610 GND.t86 911.471
R2953 GND.t483 GND.t361 911.471
R2954 GND.t361 GND.t584 911.471
R2955 GND.t80 GND.t299 911.471
R2956 GND.n3397 GND.n407 770.634
R2957 GND.n3572 GND.n3571 770.634
R2958 GND.n3344 GND.n3343 770.634
R2959 GND.n3597 GND.n3596 770.634
R2960 GND.n2986 GND.t739 770.125
R2961 GND.n2980 GND.t739 770.125
R2962 GND.n2979 GND.t542 770.125
R2963 GND.n2967 GND.t330 770.125
R2964 GND.n2966 GND.t237 770.125
R2965 GND.n2954 GND.t368 770.125
R2966 GND.n2953 GND.t657 770.125
R2967 GND.n2904 GND.t657 770.125
R2968 GND.n2905 GND.t789 770.125
R2969 GND.n2942 GND.t789 770.125
R2970 GND.n2942 GND.t209 770.125
R2971 GND.n2931 GND.t209 770.125
R2972 GND.n2930 GND.t384 770.125
R2973 GND.t90 GND.n634 770.125
R2974 GND.t735 GND.n2172 770.125
R2975 GND.t735 GND.n2448 770.125
R2976 GND.n2447 GND.t239 770.125
R2977 GND.n2435 GND.t622 770.125
R2978 GND.n2434 GND.t749 770.125
R2979 GND.n2422 GND.t199 770.125
R2980 GND.n2421 GND.t620 770.125
R2981 GND.n2372 GND.t620 770.125
R2982 GND.n2373 GND.t366 770.125
R2983 GND.n2410 GND.t366 770.125
R2984 GND.n2410 GND.t52 770.125
R2985 GND.n2399 GND.t52 770.125
R2986 GND.n2398 GND.t235 770.125
R2987 GND.t207 GND.n635 770.125
R2988 GND.t849 GND.n2206 770.125
R2989 GND.t849 GND.n2321 770.125
R2990 GND.n2320 GND.t389 770.125
R2991 GND.n2308 GND.t596 770.125
R2992 GND.n2307 GND.t427 770.125
R2993 GND.n2295 GND.t267 770.125
R2994 GND.n2294 GND.t594 770.125
R2995 GND.n2245 GND.t594 770.125
R2996 GND.n2246 GND.t319 770.125
R2997 GND.n2283 GND.t319 770.125
R2998 GND.n2283 GND.t53 770.125
R2999 GND.n2272 GND.t53 770.125
R3000 GND.n2271 GND.t651 770.125
R3001 GND.t375 GND.n636 770.125
R3002 GND.t737 GND.n2528 770.125
R3003 GND.t737 GND.n2643 770.125
R3004 GND.n2642 GND.t241 770.125
R3005 GND.n2630 GND.t251 770.125
R3006 GND.n2629 GND.t273 770.125
R3007 GND.n2617 GND.t37 770.125
R3008 GND.n2616 GND.t249 770.125
R3009 GND.n2567 GND.t249 770.125
R3010 GND.n2568 GND.t607 770.125
R3011 GND.n2605 GND.t607 770.125
R3012 GND.n2605 GND.t195 770.125
R3013 GND.n2594 GND.t195 770.125
R3014 GND.n2593 GND.t5 770.125
R3015 GND.t50 GND.n637 770.125
R3016 GND.n2770 GND.t697 770.125
R3017 GND.n2764 GND.t697 770.125
R3018 GND.n2763 GND.t649 770.125
R3019 GND.n2751 GND.t46 770.125
R3020 GND.n2750 GND.t27 770.125
R3021 GND.n2738 GND.t803 770.125
R3022 GND.n2737 GND.t3 770.125
R3023 GND.n2688 GND.t3 770.125
R3024 GND.n2689 GND.t631 770.125
R3025 GND.n2726 GND.t631 770.125
R3026 GND.n2726 GND.t196 770.125
R3027 GND.n2715 GND.t196 770.125
R3028 GND.n2714 GND.t422 770.125
R3029 GND.t288 GND.n638 770.125
R3030 GND.n3119 GND.t851 770.125
R3031 GND.n3113 GND.t851 770.125
R3032 GND.n3112 GND.t270 770.125
R3033 GND.n3100 GND.t792 770.125
R3034 GND.n3099 GND.t338 770.125
R3035 GND.n3087 GND.t254 770.125
R3036 GND.n3086 GND.t883 770.125
R3037 GND.n618 GND.t883 770.125
R3038 GND.n619 GND.t340 770.125
R3039 GND.n3075 GND.t340 770.125
R3040 GND.n3075 GND.t44 770.125
R3041 GND.n3064 GND.t44 770.125
R3042 GND.n3063 GND.t9 770.125
R3043 GND.n3051 GND.t754 770.125
R3044 GND.n4235 GND.t610 767.476
R3045 GND.n1621 GND.n1619 753.46
R3046 GND.n1619 GND.n1618 751.688
R3047 GND.n4206 GND.t354 731.85
R3048 GND.n3964 GND.t268 713.799
R3049 GND.t648 GND.t7 698.269
R3050 GND.t648 GND.t2 698.269
R3051 GND.t434 GND.t467 698.269
R3052 GND.t434 GND.t668 698.269
R3053 GND.t353 GND.t495 698.269
R3054 GND.t353 GND.t284 698.269
R3055 GND.n1581 GND.n1580 696.773
R3056 GND.n1608 GND.n1606 696.773
R3057 GND.n4234 GND.n4233 696.773
R3058 GND.n4224 GND.n4223 696.773
R3059 GND.n4205 GND.n4204 696.773
R3060 GND.n4195 GND.n4194 696.773
R3061 GND.n1050 GND.t535 659.5
R3062 GND.n1757 GND.t629 648.799
R3063 GND.n4161 GND.t629 648.799
R3064 GND.n4161 GND.t222 648.799
R3065 GND.t222 GND.n4160 648.799
R3066 GND.n4153 GND.t409 648.799
R3067 GND.n4152 GND.t215 648.799
R3068 GND.n3678 GND.t215 648.799
R3069 GND.n4142 GND.t469 648.799
R3070 GND.n4142 GND.t69 648.799
R3071 GND.t69 GND.n4138 648.799
R3072 GND.n4137 GND.t664 648.799
R3073 GND.n4131 GND.t664 648.799
R3074 GND.n4130 GND.t124 648.799
R3075 GND.n4124 GND.t323 648.799
R3076 GND.n4123 GND.t477 648.799
R3077 GND.n4116 GND.t429 648.799
R3078 GND.n136 GND.t429 648.799
R3079 GND.t391 GND.n136 648.799
R3080 GND.n4110 GND.t391 648.799
R3081 GND.n4109 GND.t537 648.799
R3082 GND.n4103 GND.t776 648.799
R3083 GND.n4102 GND.t661 648.799
R3084 GND.n3728 GND.t661 648.799
R3085 GND.n3728 GND.t431 648.799
R3086 GND.n4093 GND.t431 648.799
R3087 GND.n4092 GND.t0 648.799
R3088 GND.n4086 GND.t0 648.799
R3089 GND.n4085 GND.t104 648.799
R3090 GND.n4079 GND.t261 648.799
R3091 GND.n4078 GND.t554 648.799
R3092 GND.n4072 GND.t229 648.799
R3093 GND.n4071 GND.t624 648.799
R3094 GND.n163 GND.t624 648.799
R3095 GND.t200 GND.n163 648.799
R3096 GND.n4065 GND.t200 648.799
R3097 GND.n4064 GND.t493 648.799
R3098 GND.n4058 GND.t349 648.799
R3099 GND.n4057 GND.t806 648.799
R3100 GND.n3831 GND.t806 648.799
R3101 GND.n4047 GND.t838 648.799
R3102 GND.n4047 GND.t78 648.799
R3103 GND.t78 GND.n4043 648.799
R3104 GND.n4042 GND.t856 648.799
R3105 GND.n4036 GND.t856 648.799
R3106 GND.n4035 GND.t817 648.799
R3107 GND.n4029 GND.t448 648.799
R3108 GND.n4028 GND.t475 648.799
R3109 GND.n4021 GND.t444 648.799
R3110 GND.n194 GND.t444 648.799
R3111 GND.t62 GND.n194 648.799
R3112 GND.n4015 GND.t62 648.799
R3113 GND.n4014 GND.t507 648.799
R3114 GND.n4008 GND.t640 648.799
R3115 GND.n4007 GND.t193 648.799
R3116 GND.n3881 GND.t193 648.799
R3117 GND.n3881 GND.t289 648.799
R3118 GND.n3998 GND.t289 648.799
R3119 GND.n3997 GND.t91 648.799
R3120 GND.n3991 GND.t91 648.799
R3121 GND.n3990 GND.t132 648.799
R3122 GND.n3984 GND.t842 648.799
R3123 GND.n3983 GND.t527 648.799
R3124 GND.n3977 GND.t279 648.799
R3125 GND.n3976 GND.t263 648.799
R3126 GND.n221 GND.t263 648.799
R3127 GND.t598 GND.n221 648.799
R3128 GND.n3970 GND.t598 648.799
R3129 GND.n3969 GND.t576 648.799
R3130 GND.n1579 GND.n1578 641.857
R3131 GND.n1605 GND.n1604 641.857
R3132 GND.n4222 GND.n4221 641.857
R3133 GND.n4207 GND.n4206 641.857
R3134 GND.n4193 GND.n4192 641.857
R3135 GND.n1329 GND.n1327 625.822
R3136 GND.n1343 GND.n1342 625.822
R3137 GND.n1350 GND.n1349 625.822
R3138 GND.n994 GND.n992 625.822
R3139 GND.n1008 GND.n1007 625.822
R3140 GND.n1016 GND.n1014 625.822
R3141 GND.n1065 GND.n1064 625.822
R3142 GND.n1684 GND.n1683 625.822
R3143 GND.n1677 GND.n1676 625.822
R3144 GND.n1540 GND.n1538 625.822
R3145 GND.n1554 GND.n1553 625.822
R3146 GND.n1561 GND.n1560 625.822
R3147 GND.n1480 GND.n1478 625.822
R3148 GND.n1494 GND.n1493 625.822
R3149 GND.n1502 GND.n1500 625.822
R3150 GND.n3409 GND.n401 625.822
R3151 GND.n3412 GND.n3411 625.822
R3152 GND.n3424 GND.n3422 625.822
R3153 GND.n3434 GND.n3433 625.822
R3154 GND.n3516 GND.n3515 625.822
R3155 GND.n3505 GND.n3504 625.822
R3156 GND.n3483 GND.n3482 625.822
R3157 GND.n3490 GND.n3489 625.822
R3158 GND.n3692 GND.n311 625.822
R3159 GND.n3695 GND.n3694 625.822
R3160 GND.n3707 GND.n3705 625.822
R3161 GND.n3717 GND.n3716 625.822
R3162 GND.n3733 GND.n3732 625.822
R3163 GND.n3738 GND.n3736 625.822
R3164 GND.n3761 GND.n3760 625.822
R3165 GND.n3751 GND.n3750 625.822
R3166 GND.n3845 GND.n261 625.822
R3167 GND.n3848 GND.n3847 625.822
R3168 GND.n3860 GND.n3858 625.822
R3169 GND.n3870 GND.n3869 625.822
R3170 GND.n3886 GND.n3885 625.822
R3171 GND.n3891 GND.n3889 625.822
R3172 GND.n3923 GND.n3922 625.822
R3173 GND.n3913 GND.n3912 625.822
R3174 GND.n3178 GND.n3177 625.822
R3175 GND.n3174 GND.n3173 625.822
R3176 GND.n4280 GND.n4279 625.822
R3177 GND.n4270 GND.n4269 625.822
R3178 GND.n3280 GND.n507 625.822
R3179 GND.n3283 GND.n3282 625.822
R3180 GND.n3295 GND.n3293 625.822
R3181 GND.n3309 GND.n3308 625.822
R3182 GND.n1250 GND.n1248 625.822
R3183 GND.n1264 GND.n1263 625.822
R3184 GND.n1271 GND.n1270 625.822
R3185 GND.n2093 GND.n2092 625.822
R3186 GND.n2079 GND.n2078 625.822
R3187 GND.n2072 GND.n2071 625.822
R3188 GND.n2010 GND.n2009 625.822
R3189 GND.n1996 GND.n1995 625.822
R3190 GND.n1989 GND.n1988 625.822
R3191 GND.n3609 GND.n336 625.822
R3192 GND.n3612 GND.n3611 625.822
R3193 GND.n3624 GND.n3622 625.822
R3194 GND.n3634 GND.n3633 625.822
R3195 GND.n1667 GND.t388 615.399
R3196 GND.n1657 GND.t491 615.399
R3197 GND.n1656 GND.t51 615.399
R3198 GND.n920 GND.t51 615.399
R3199 GND.t370 GND.n920 615.399
R3200 GND.n1647 GND.t370 615.399
R3201 GND.n1646 GND.t844 615.399
R3202 GND.n1022 GND.t844 615.399
R3203 GND.t878 GND.n1023 615.399
R3204 GND.n1026 GND.t521 615.399
R3205 GND.t262 GND.n1027 615.399
R3206 GND.n1030 GND.t154 615.399
R3207 GND.n1142 GND.t796 615.399
R3208 GND.n1080 GND.t110 615.399
R3209 GND.t714 GND.n1081 615.399
R3210 GND.n1130 GND.t714 615.399
R3211 GND.n1130 GND.t811 615.399
R3212 GND.t811 GND.n1126 615.399
R3213 GND.n1125 GND.t451 615.399
R3214 GND.n1097 GND.t451 615.399
R3215 GND.n1098 GND.t646 615.399
R3216 GND.n1103 GND.t176 615.399
R3217 GND.t304 GND.n1104 615.399
R3218 GND.t572 GND.n908 615.399
R3219 GND.n1743 GND.t753 615.399
R3220 GND.n1733 GND.t138 615.399
R3221 GND.n1732 GND.t587 615.399
R3222 GND.n870 GND.t587 615.399
R3223 GND.t308 GND.n870 615.399
R3224 GND.n1723 GND.t308 615.399
R3225 GND.n1722 GND.t11 615.399
R3226 GND.n1057 GND.t11 615.399
R3227 GND.n1573 GND.t136 615.399
R3228 GND.n1572 GND.t67 615.399
R3229 GND.t548 GND.n1569 615.399
R3230 GND.t160 GND.n1756 615.399
R3231 GND.n1755 GND.t292 615.399
R3232 GND.n1745 GND.t535 615.399
R3233 GND.n2143 GND.t875 615.399
R3234 GND.n2135 GND.t140 615.399
R3235 GND.n2134 GND.t419 615.399
R3236 GND.n651 GND.t419 615.399
R3237 GND.t346 GND.n651 615.399
R3238 GND.n2125 GND.t346 615.399
R3239 GND.n2124 GND.t15 615.399
R3240 GND.n660 GND.t15 615.399
R3241 GND.n661 GND.t66 615.399
R3242 GND.n2113 GND.t823 615.399
R3243 GND.n2112 GND.t293 615.399
R3244 GND.n2102 GND.t501 615.399
R3245 GND.t60 GND.n673 615.399
R3246 GND.n733 GND.t112 615.399
R3247 GND.n735 GND.t729 615.399
R3248 GND.t729 GND.n734 615.399
R3249 GND.n734 GND.t343 615.399
R3250 GND.n745 GND.t343 615.399
R3251 GND.t455 GND.n747 615.399
R3252 GND.n748 GND.t455 615.399
R3253 GND.n767 GND.t142 615.399
R3254 GND.t380 GND.n768 615.399
R3255 GND.t515 GND.n696 615.399
R3256 GND.n2062 GND.t802 615.399
R3257 GND.n2052 GND.t829 615.399
R3258 GND.n2051 GND.t583 615.399
R3259 GND.n782 GND.t583 615.399
R3260 GND.t33 GND.n782 615.399
R3261 GND.n2042 GND.t33 615.399
R3262 GND.n2041 GND.t259 615.399
R3263 GND.n791 GND.t259 615.399
R3264 GND.n792 GND.t412 615.399
R3265 GND.n2030 GND.t130 615.399
R3266 GND.n2029 GND.t20 615.399
R3267 GND.n2019 GND.t558 615.399
R3268 GND.t724 GND.n804 615.399
R3269 GND.t156 GND.n1423 615.399
R3270 GND.n1422 GND.t187 615.399
R3271 GND.n1370 GND.t187 615.399
R3272 GND.t232 GND.n1370 615.399
R3273 GND.n1413 GND.t232 615.399
R3274 GND.n1412 GND.t302 615.399
R3275 GND.n1374 GND.t302 615.399
R3276 GND.t108 GND.n1399 615.399
R3277 GND.n1398 GND.t461 615.399
R3278 GND.t487 GND.n827 615.399
R3279 GND.n1979 GND.t693 615.399
R3280 GND.n1968 GND.t848 615.399
R3281 GND.n840 GND.t848 615.399
R3282 GND.t183 GND.n840 615.399
R3283 GND.n1959 GND.t183 615.399
R3284 GND.n1777 GND.t204 600.622
R3285 GND.t868 GND.n1776 600.622
R3286 GND.n4159 GND.n104 583.285
R3287 GND.n3014 GND.n3012 579.418
R3288 GND.n1050 GND.t767 571.298
R3289 GND.t768 GND.t230 569.819
R3290 GND.n4177 GND.t180 555.197
R3291 GND.t694 GND.t781 554.254
R3292 GND.t865 GND.t836 551.01
R3293 GND.t865 GND.t791 551.01
R3294 GND.t89 GND.t397 551.01
R3295 GND.t858 GND.t89 551.01
R3296 GND.t420 GND.t687 551.01
R3297 GND.t687 GND.t72 551.01
R3298 GND.n130 GND.t684 530.452
R3299 GND.n188 GND.t208 530.452
R3300 GND.n1758 GND.t160 527.198
R3301 GND.t481 GND.n841 521.053
R3302 GND.n3680 GND.n3679 511.432
R3303 GND.n3833 GND.n3832 511.432
R3304 GND.n1580 GND.t709 503.144
R3305 GND.n4223 GND.t405 503.144
R3306 GND.n4194 GND.t688 503.144
R3307 GND.n1807 GND.t316 502.156
R3308 GND.t765 GND.n1806 502.156
R3309 GND.n1837 GND.t47 502.156
R3310 GND.t185 GND.n1836 502.156
R3311 GND.n1792 GND.t701 502.156
R3312 GND.t100 GND.n1791 502.156
R3313 GND.n1852 GND.t777 501.411
R3314 GND.t605 GND.n1851 501.411
R3315 GND.n4235 GND.n39 492.76
R3316 GND.n3967 GND.n3966 467.2
R3317 GND.n3966 GND.n3965 467.2
R3318 GND.n3981 GND.n3980 467.2
R3319 GND.n3980 GND.n3979 467.2
R3320 GND.n3988 GND.n3987 467.2
R3321 GND.n3987 GND.n3986 467.2
R3322 GND.n4012 GND.n4011 467.2
R3323 GND.n4011 GND.n4010 467.2
R3324 GND.n4026 GND.n4025 467.2
R3325 GND.n4025 GND.n4024 467.2
R3326 GND.n4033 GND.n4032 467.2
R3327 GND.n4032 GND.n4031 467.2
R3328 GND.n4062 GND.n4061 467.2
R3329 GND.n4061 GND.n4060 467.2
R3330 GND.n4076 GND.n4075 467.2
R3331 GND.n4075 GND.n4074 467.2
R3332 GND.n4083 GND.n4082 467.2
R3333 GND.n4082 GND.n4081 467.2
R3334 GND.n4107 GND.n4106 467.2
R3335 GND.n4106 GND.n4105 467.2
R3336 GND.n4121 GND.n4120 467.2
R3337 GND.n4120 GND.n4119 467.2
R3338 GND.n4128 GND.n4127 467.2
R3339 GND.n4127 GND.n4126 467.2
R3340 GND.n4157 GND.n4156 467.2
R3341 GND.n4156 GND.n4155 467.2
R3342 GND.n88 GND.n87 467.2
R3343 GND.n89 GND.n88 467.2
R3344 GND.n4254 GND.n4253 467.2
R3345 GND.n4255 GND.n4254 467.2
R3346 GND.n4239 GND.n4238 467.2
R3347 GND.n4240 GND.n4239 467.2
R3348 GND.n545 GND.n538 467.2
R3349 GND.n3193 GND.n538 467.2
R3350 GND.n630 GND.n625 467.2
R3351 GND.n630 GND.n628 467.2
R3352 GND.n3053 GND.n624 467.2
R3353 GND.n3061 GND.n624 467.2
R3354 GND.n601 GND.n596 467.2
R3355 GND.n601 GND.n599 467.2
R3356 GND.n3089 GND.n595 467.2
R3357 GND.n3097 GND.n595 467.2
R3358 GND.n589 GND.n584 467.2
R3359 GND.n589 GND.n587 467.2
R3360 GND.n3102 GND.n583 467.2
R3361 GND.n3110 GND.n583 467.2
R3362 GND.n1789 GND.n1783 467.2
R3363 GND.n1794 GND.n1783 467.2
R3364 GND.n1804 GND.n1798 467.2
R3365 GND.n1809 GND.n1798 467.2
R3366 GND.n1819 GND.n1813 467.2
R3367 GND.n1824 GND.n1813 467.2
R3368 GND.n1834 GND.n1828 467.2
R3369 GND.n1839 GND.n1828 467.2
R3370 GND.n1849 GND.n1843 467.2
R3371 GND.n1854 GND.n1843 467.2
R3372 GND.n1779 GND.n1768 467.2
R3373 GND.n1774 GND.n1768 467.2
R3374 GND.n1268 GND.n1267 467.2
R3375 GND.n1267 GND.n1266 467.2
R3376 GND.n1261 GND.n1260 467.2
R3377 GND.n1260 GND.n1259 467.2
R3378 GND.n2075 GND.n2074 467.2
R3379 GND.n2076 GND.n2075 467.2
R3380 GND.n2082 GND.n2081 467.2
R3381 GND.n2083 GND.n2082 467.2
R3382 GND.n2096 GND.n2095 467.2
R3383 GND.n2097 GND.n2096 467.2
R3384 GND.n1346 GND.n1345 467.2
R3385 GND.n1347 GND.n1346 467.2
R3386 GND.n1339 GND.n1338 467.2
R3387 GND.n1340 GND.n1339 467.2
R3388 GND.n1325 GND.n1324 467.2
R3389 GND.n1324 GND.n1323 467.2
R3390 GND.n1992 GND.n1991 467.2
R3391 GND.n1993 GND.n1992 467.2
R3392 GND.n1999 GND.n1998 467.2
R3393 GND.n2000 GND.n1999 467.2
R3394 GND.n2013 GND.n2012 467.2
R3395 GND.n2014 GND.n2013 467.2
R3396 GND.n1753 GND.n853 467.2
R3397 GND.n1747 GND.n853 467.2
R3398 GND.n1061 GND.n880 467.2
R3399 GND.n1061 GND.n882 467.2
R3400 GND.n1575 GND.n876 467.2
R3401 GND.n1575 GND.n878 467.2
R3402 GND.n1741 GND.n861 467.2
R3403 GND.n1735 GND.n861 467.2
R3404 GND.n1094 GND.n1092 467.2
R3405 GND.n1107 GND.n1094 467.2
R3406 GND.n1100 GND.n1088 467.2
R3407 GND.n1100 GND.n1090 467.2
R3408 GND.n1140 GND.n1071 467.2
R3409 GND.n1078 GND.n1071 467.2
R3410 GND.n1018 GND.n930 467.2
R3411 GND.n1018 GND.n932 467.2
R3412 GND.n1020 GND.n926 467.2
R3413 GND.n1020 GND.n928 467.2
R3414 GND.n1665 GND.n911 467.2
R3415 GND.n1659 GND.n911 467.2
R3416 GND.n1011 GND.n1010 467.2
R3417 GND.n1012 GND.n1011 467.2
R3418 GND.n1004 GND.n1003 467.2
R3419 GND.n1005 GND.n1004 467.2
R3420 GND.n989 GND.n988 467.2
R3421 GND.n990 GND.n989 467.2
R3422 GND.n1681 GND.n1680 467.2
R3423 GND.n1680 GND.n1679 467.2
R3424 GND.n1688 GND.n1687 467.2
R3425 GND.n1687 GND.n1686 467.2
R3426 GND.n1063 GND.n885 467.2
R3427 GND.n1063 GND.n887 467.2
R3428 GND.n1557 GND.n1556 467.2
R3429 GND.n1558 GND.n1557 467.2
R3430 GND.n1550 GND.n1549 467.2
R3431 GND.n1551 GND.n1550 467.2
R3432 GND.n1535 GND.n1534 467.2
R3433 GND.n1536 GND.n1535 467.2
R3434 GND.n1497 GND.n1496 467.2
R3435 GND.n1498 GND.n1497 467.2
R3436 GND.n1490 GND.n1489 467.2
R3437 GND.n1491 GND.n1490 467.2
R3438 GND.n1475 GND.n1474 467.2
R3439 GND.n1476 GND.n1475 467.2
R3440 GND.n1947 GND.n1946 467.2
R3441 GND.n1947 GND.n847 467.2
R3442 GND.n1971 GND.n831 467.2
R3443 GND.n1977 GND.n831 467.2
R3444 GND.n1390 GND.n1384 467.2
R3445 GND.n1396 GND.n1384 467.2
R3446 GND.n1401 GND.n1400 467.2
R3447 GND.n1401 GND.n1378 467.2
R3448 GND.n1425 GND.n1424 467.2
R3449 GND.n1425 GND.n1359 467.2
R3450 GND.n2021 GND.n799 467.2
R3451 GND.n2027 GND.n799 467.2
R3452 GND.n796 GND.n795 467.2
R3453 GND.n795 GND.n788 467.2
R3454 GND.n2054 GND.n700 467.2
R3455 GND.n2060 GND.n700 467.2
R3456 GND.n771 GND.n704 467.2
R3457 GND.n759 GND.n704 467.2
R3458 GND.n765 GND.n709 467.2
R3459 GND.n755 GND.n709 467.2
R3460 GND.n731 GND.n721 467.2
R3461 GND.n724 GND.n721 467.2
R3462 GND.n3340 GND.n3339 467.2
R3463 GND.n3341 GND.n3340 467.2
R3464 GND.n3235 GND.n3234 467.2
R3465 GND.n3234 GND.n3233 467.2
R3466 GND.n3242 GND.n3241 467.2
R3467 GND.n3241 GND.n3240 467.2
R3468 GND.n3312 GND.n490 467.2
R3469 GND.n3300 GND.n490 467.2
R3470 GND.n3285 GND.n504 467.2
R3471 GND.n3278 GND.n504 467.2
R3472 GND.n3487 GND.n347 467.2
R3473 GND.n3575 GND.n347 467.2
R3474 GND.n3513 GND.n3468 467.2
R3475 GND.n3507 GND.n3468 467.2
R3476 GND.n3568 GND.n3567 467.2
R3477 GND.n3569 GND.n3568 467.2
R3478 GND.n3451 GND.n361 467.2
R3479 GND.n3545 GND.n361 467.2
R3480 GND.n3538 GND.n3537 467.2
R3481 GND.n3539 GND.n3538 467.2
R3482 GND.n457 GND.n378 467.2
R3483 GND.n3448 GND.n378 467.2
R3484 GND.n471 GND.n470 467.2
R3485 GND.n470 GND.n469 467.2
R3486 GND.n478 GND.n477 467.2
R3487 GND.n477 GND.n476 467.2
R3488 GND.n3436 GND.n384 467.2
R3489 GND.n3442 GND.n384 467.2
R3490 GND.n3407 GND.n398 467.2
R3491 GND.n3414 GND.n398 467.2
R3492 GND.n3315 GND.n404 467.2
R3493 GND.n3401 GND.n404 467.2
R3494 GND.n3518 GND.n374 467.2
R3495 GND.n3524 GND.n374 467.2
R3496 GND.n3674 GND.n319 467.2
R3497 GND.n3636 GND.n319 467.2
R3498 GND.n3614 GND.n333 467.2
R3499 GND.n3607 GND.n333 467.2
R3500 GND.n3601 GND.n339 467.2
R3501 GND.n3578 GND.n339 467.2
R3502 GND.n3910 GND.n3900 467.2
R3503 GND.n3904 GND.n3900 467.2
R3504 GND.n239 GND.n231 467.2
R3505 GND.n239 GND.n233 467.2
R3506 GND.n3872 GND.n244 467.2
R3507 GND.n3878 GND.n244 467.2
R3508 GND.n3843 GND.n258 467.2
R3509 GND.n3850 GND.n258 467.2
R3510 GND.n272 GND.n264 467.2
R3511 GND.n3837 GND.n264 467.2
R3512 GND.n3748 GND.n269 467.2
R3513 GND.n3827 GND.n269 467.2
R3514 GND.n289 GND.n281 467.2
R3515 GND.n289 GND.n283 467.2
R3516 GND.n291 GND.n277 467.2
R3517 GND.n291 GND.n279 467.2
R3518 GND.n3719 GND.n294 467.2
R3519 GND.n3725 GND.n294 467.2
R3520 GND.n3690 GND.n308 467.2
R3521 GND.n3697 GND.n308 467.2
R3522 GND.n3640 GND.n314 467.2
R3523 GND.n3684 GND.n314 467.2
R3524 GND.n241 GND.n229 467.2
R3525 GND.n241 GND.n227 467.2
R3526 GND.n4267 GND.n21 467.2
R3527 GND.n4261 GND.n21 467.2
R3528 GND.n3171 GND.n6 467.2
R3529 GND.n3171 GND.n8 467.2
R3530 GND.n3169 GND.n4 467.2
R3531 GND.n3169 GND.n2 467.2
R3532 GND.n3252 GND.n510 467.2
R3533 GND.n3272 GND.n510 467.2
R3534 GND.n2104 GND.n668 467.2
R3535 GND.n2110 GND.n668 467.2
R3536 GND.n665 GND.n664 467.2
R3537 GND.n664 GND.n657 467.2
R3538 GND.n2137 GND.n643 467.2
R3539 GND.n2141 GND.n643 467.2
R3540 GND.n1245 GND.n1244 467.2
R3541 GND.n1246 GND.n1245 467.2
R3542 GND.n2182 GND.n2151 467.2
R3543 GND.n3024 GND.n2151 467.2
R3544 GND.n3009 GND.n3008 467.2
R3545 GND.n3010 GND.n3009 467.2
R3546 GND.n3002 GND.n3001 467.2
R3547 GND.n3003 GND.n3002 467.2
R3548 GND.n2822 GND.n2821 467.2
R3549 GND.n2822 GND.n2813 467.2
R3550 GND.n2849 GND.n2469 467.2
R3551 GND.n2855 GND.n2469 467.2
R3552 GND.n2860 GND.n2459 467.2
R3553 GND.n2860 GND.n2859 467.2
R3554 GND.n2806 GND.n2805 467.2
R3555 GND.n2806 GND.n2800 467.2
R3556 GND.n2794 GND.n2793 467.2
R3557 GND.n2793 GND.n2790 467.2
R3558 GND.n2784 GND.n2783 467.2
R3559 GND.n2783 GND.n2782 467.2
R3560 GND.n2914 GND.n2911 467.2
R3561 GND.n2918 GND.n2914 467.2
R3562 GND.n2920 GND.n2910 467.2
R3563 GND.n2928 GND.n2910 467.2
R3564 GND.n2887 GND.n2882 467.2
R3565 GND.n2887 GND.n2885 467.2
R3566 GND.n2956 GND.n2881 467.2
R3567 GND.n2964 GND.n2881 467.2
R3568 GND.n2875 GND.n2180 467.2
R3569 GND.n2875 GND.n2873 467.2
R3570 GND.n2969 GND.n2179 467.2
R3571 GND.n2977 GND.n2179 467.2
R3572 GND.n2382 GND.n2379 467.2
R3573 GND.n2386 GND.n2382 467.2
R3574 GND.n2388 GND.n2378 467.2
R3575 GND.n2396 GND.n2378 467.2
R3576 GND.n2355 GND.n2350 467.2
R3577 GND.n2355 GND.n2353 467.2
R3578 GND.n2424 GND.n2349 467.2
R3579 GND.n2432 GND.n2349 467.2
R3580 GND.n2343 GND.n2338 467.2
R3581 GND.n2343 GND.n2341 467.2
R3582 GND.n2437 GND.n2337 467.2
R3583 GND.n2445 GND.n2337 467.2
R3584 GND.n2255 GND.n2252 467.2
R3585 GND.n2259 GND.n2255 467.2
R3586 GND.n2261 GND.n2251 467.2
R3587 GND.n2269 GND.n2251 467.2
R3588 GND.n2228 GND.n2223 467.2
R3589 GND.n2228 GND.n2226 467.2
R3590 GND.n2297 GND.n2222 467.2
R3591 GND.n2305 GND.n2222 467.2
R3592 GND.n2216 GND.n2211 467.2
R3593 GND.n2216 GND.n2214 467.2
R3594 GND.n2310 GND.n2210 467.2
R3595 GND.n2318 GND.n2210 467.2
R3596 GND.n2577 GND.n2574 467.2
R3597 GND.n2581 GND.n2577 467.2
R3598 GND.n2583 GND.n2573 467.2
R3599 GND.n2591 GND.n2573 467.2
R3600 GND.n2550 GND.n2545 467.2
R3601 GND.n2550 GND.n2548 467.2
R3602 GND.n2619 GND.n2544 467.2
R3603 GND.n2627 GND.n2544 467.2
R3604 GND.n2538 GND.n2533 467.2
R3605 GND.n2538 GND.n2536 467.2
R3606 GND.n2632 GND.n2532 467.2
R3607 GND.n2640 GND.n2532 467.2
R3608 GND.n2698 GND.n2695 467.2
R3609 GND.n2702 GND.n2698 467.2
R3610 GND.n2704 GND.n2694 467.2
R3611 GND.n2712 GND.n2694 467.2
R3612 GND.n2671 GND.n2666 467.2
R3613 GND.n2671 GND.n2669 467.2
R3614 GND.n2740 GND.n2665 467.2
R3615 GND.n2748 GND.n2665 467.2
R3616 GND.n2659 GND.n2514 467.2
R3617 GND.n2659 GND.n2657 467.2
R3618 GND.n2753 GND.n2513 467.2
R3619 GND.n2761 GND.n2513 467.2
R3620 GND.n1943 GND.n1942 467.2
R3621 GND.n1942 GND.n1941 467.2
R3622 GND.n1914 GND.n1857 467.2
R3623 GND.n1914 GND.n1913 467.2
R3624 GND.n1908 GND.n93 467.2
R3625 GND.n1908 GND.n95 467.2
R3626 GND.n3165 GND.n553 467.2
R3627 GND.n3159 GND.n553 467.2
R3628 GND.n3137 GND.n567 467.2
R3629 GND.n3130 GND.n567 467.2
R3630 GND.n3124 GND.n573 467.2
R3631 GND.n2516 GND.n573 467.2
R3632 GND.n1969 GND.n82 463.053
R3633 GND.n4153 GND.n4152 460.712
R3634 GND.n4138 GND.n4137 460.712
R3635 GND.n4058 GND.n4057 460.712
R3636 GND.n4043 GND.n4042 460.712
R3637 GND.n1912 GND.t21 456.574
R3638 GND.t704 GND.n407 455.736
R3639 GND.n481 GND.t704 455.736
R3640 GND.n480 GND.t819 455.736
R3641 GND.n474 GND.t449 455.736
R3642 GND.n473 GND.t503 455.736
R3643 GND.n467 GND.t673 455.736
R3644 GND.n466 GND.t313 455.736
R3645 GND.n440 GND.t313 455.736
R3646 GND.t189 GND.n440 455.736
R3647 GND.n460 GND.t189 455.736
R3648 GND.n459 GND.t539 455.736
R3649 GND.n3446 GND.t773 455.736
R3650 GND.n3528 GND.t30 455.736
R3651 GND.n3534 GND.t30 455.736
R3652 GND.n3535 GND.t152 455.736
R3653 GND.n3541 GND.t226 455.736
R3654 GND.t560 GND.n3542 455.736
R3655 GND.n3558 GND.t244 455.736
R3656 GND.t244 GND.n3557 455.736
R3657 GND.n3557 GND.t74 455.736
R3658 GND.n3564 GND.t74 455.736
R3659 GND.n3565 GND.t564 455.736
R3660 GND.n3571 GND.t627 455.736
R3661 GND.t335 GND.n513 455.736
R3662 GND.n3245 GND.t335 455.736
R3663 GND.n3244 GND.t106 455.736
R3664 GND.n3238 GND.t414 455.736
R3665 GND.n3237 GND.t552 455.736
R3666 GND.n3330 GND.t784 455.736
R3667 GND.t784 GND.n3329 455.736
R3668 GND.n3329 GND.t728 455.736
R3669 GND.n3336 GND.t728 455.736
R3670 GND.n3337 GND.t531 455.736
R3671 GND.n3343 GND.t585 455.736
R3672 GND.n3183 GND.t655 455.736
R3673 GND.n3189 GND.t655 455.736
R3674 GND.t128 GND.n3190 455.736
R3675 GND.t326 GND.n38 455.736
R3676 GND.n4236 GND.t505 455.736
R3677 GND.n4242 GND.t86 455.736
R3678 GND.n4244 GND.t666 455.736
R3679 GND.t666 GND.n4243 455.736
R3680 GND.n4243 GND.t35 455.736
R3681 GND.n4250 GND.t35 455.736
R3682 GND.n4251 GND.t483 455.736
R3683 GND.n4257 GND.t584 455.736
R3684 GND.n3596 GND.t83 455.736
R3685 GND.n3590 GND.t83 455.736
R3686 GND.n3589 GND.t180 455.736
R3687 GND.n1905 GND.t299 455.736
R3688 GND.n1906 GND.t481 455.736
R3689 GND.t589 GND.t876 431.428
R3690 GND.t876 GND.t96 431.428
R3691 GND.n1619 GND.n188 416.842
R3692 GND.n1605 GND.n1035 416.842
R3693 GND.n1579 GND.n130 416.842
R3694 GND.t424 GND.t439 407.051
R3695 GND.t439 GND.t593 407.051
R3696 GND.t393 GND.t57 407.051
R3697 GND.t57 GND.t861 407.051
R3698 GND.t442 GND.t614 407.051
R3699 GND.t442 GND.t402 407.051
R3700 GND.n4193 GND.t248 372.606
R3701 GND.n4222 GND.t603 372.606
R3702 GND.n4177 GND.t80 356.276
R3703 GND.n3974 GND.n3973 351.625
R3704 GND.n3973 GND.n3972 351.625
R3705 GND.n4019 GND.n4018 351.625
R3706 GND.n4018 GND.n4017 351.625
R3707 GND.n4069 GND.n4068 351.625
R3708 GND.n4068 GND.n4067 351.625
R3709 GND.n4114 GND.n4113 351.625
R3710 GND.n4113 GND.n4112 351.625
R3711 GND.n102 GND.n97 351.625
R3712 GND.n102 GND.n101 351.625
R3713 GND.n4247 GND.n4246 351.625
R3714 GND.n4248 GND.n4247 351.625
R3715 GND.n3068 GND.n3067 351.625
R3716 GND.n3069 GND.n3068 351.625
R3717 GND.n3073 GND.n3072 351.625
R3718 GND.n3073 GND.n3066 351.625
R3719 GND.n3037 GND.n3036 351.625
R3720 GND.n3037 GND.n3029 351.625
R3721 GND.n1610 GND.n1033 351.625
R3722 GND.n1616 GND.n1033 351.625
R3723 GND.n1596 GND.n1038 351.625
R3724 GND.n1602 GND.n1038 351.625
R3725 GND.n1254 GND.n1253 351.625
R3726 GND.n1253 GND.n1252 351.625
R3727 GND.n2089 GND.n2088 351.625
R3728 GND.n2090 GND.n2089 351.625
R3729 GND.n1332 GND.n1331 351.625
R3730 GND.n1333 GND.n1332 351.625
R3731 GND.n2006 GND.n2005 351.625
R3732 GND.n2007 GND.n2006 351.625
R3733 GND.n1730 GND.n867 351.625
R3734 GND.n1725 GND.n867 351.625
R3735 GND.n1128 GND.n1074 351.625
R3736 GND.n1128 GND.n1127 351.625
R3737 GND.n1654 GND.n917 351.625
R3738 GND.n1649 GND.n917 351.625
R3739 GND.n997 GND.n996 351.625
R3740 GND.n998 GND.n997 351.625
R3741 GND.n894 GND.n889 351.625
R3742 GND.n894 GND.n893 351.625
R3743 GND.n1543 GND.n1542 351.625
R3744 GND.n1544 GND.n1543 351.625
R3745 GND.n1483 GND.n1482 351.625
R3746 GND.n1484 GND.n1483 351.625
R3747 GND.n1961 GND.n837 351.625
R3748 GND.n1966 GND.n837 351.625
R3749 GND.n1415 GND.n1365 351.625
R3750 GND.n1420 GND.n1365 351.625
R3751 GND.n2044 GND.n779 351.625
R3752 GND.n2049 GND.n779 351.625
R3753 GND.n743 GND.n717 351.625
R3754 GND.n737 GND.n717 351.625
R3755 GND.n3333 GND.n3332 351.625
R3756 GND.n3334 GND.n3333 351.625
R3757 GND.n3306 GND.n495 351.625
R3758 GND.n3297 GND.n495 351.625
R3759 GND.n3492 GND.n3477 351.625
R3760 GND.n3492 GND.n3491 351.625
R3761 GND.n3561 GND.n3560 351.625
R3762 GND.n3562 GND.n3561 351.625
R3763 GND.n464 GND.n463 351.625
R3764 GND.n463 GND.n462 351.625
R3765 GND.n3383 GND.n3360 351.625
R3766 GND.n3378 GND.n3360 351.625
R3767 GND.n3426 GND.n389 351.625
R3768 GND.n3431 GND.n389 351.625
R3769 GND.n3394 GND.n410 351.625
R3770 GND.n3348 GND.n410 351.625
R3771 GND.n3265 GND.n516 351.625
R3772 GND.n531 GND.n516 351.625
R3773 GND.n4000 GND.n201 351.625
R3774 GND.n4005 GND.n201 351.625
R3775 GND.n4045 GND.n4044 351.625
R3776 GND.n4045 GND.n173 351.625
R3777 GND.n4095 GND.n143 351.625
R3778 GND.n4100 GND.n143 351.625
R3779 GND.n4140 GND.n4139 351.625
R3780 GND.n4140 GND.n115 351.625
R3781 GND.n3369 GND.n3364 351.625
R3782 GND.n3369 GND.n3368 351.625
R3783 GND.n3631 GND.n324 351.625
R3784 GND.n3626 GND.n324 351.625
R3785 GND.n3920 GND.n3894 351.625
R3786 GND.n3915 GND.n3894 351.625
R3787 GND.n3862 GND.n249 351.625
R3788 GND.n3867 GND.n249 351.625
R3789 GND.n3758 GND.n3741 351.625
R3790 GND.n3753 GND.n3741 351.625
R3791 GND.n3709 GND.n299 351.625
R3792 GND.n3714 GND.n299 351.625
R3793 GND.n4277 GND.n15 351.625
R3794 GND.n4272 GND.n15 351.625
R3795 GND.n2127 GND.n648 351.625
R3796 GND.n2132 GND.n648 351.625
R3797 GND.n3017 GND.n3016 351.625
R3798 GND.n3018 GND.n3017 351.625
R3799 GND.n2834 GND.n2833 351.625
R3800 GND.n2834 GND.n2480 351.625
R3801 GND.n2493 GND.n2492 351.625
R3802 GND.n2492 GND.n2491 351.625
R3803 GND.n2935 GND.n2934 351.625
R3804 GND.n2936 GND.n2935 351.625
R3805 GND.n2940 GND.n2939 351.625
R3806 GND.n2940 GND.n2933 351.625
R3807 GND.n2403 GND.n2402 351.625
R3808 GND.n2404 GND.n2403 351.625
R3809 GND.n2408 GND.n2407 351.625
R3810 GND.n2408 GND.n2401 351.625
R3811 GND.n2276 GND.n2275 351.625
R3812 GND.n2277 GND.n2276 351.625
R3813 GND.n2281 GND.n2280 351.625
R3814 GND.n2281 GND.n2274 351.625
R3815 GND.n2598 GND.n2597 351.625
R3816 GND.n2599 GND.n2598 351.625
R3817 GND.n2603 GND.n2602 351.625
R3818 GND.n2603 GND.n2596 351.625
R3819 GND.n2719 GND.n2718 351.625
R3820 GND.n2720 GND.n2719 351.625
R3821 GND.n2724 GND.n2723 351.625
R3822 GND.n2724 GND.n2717 351.625
R3823 GND.n1583 GND.n1047 351.625
R3824 GND.n1052 GND.n1047 351.625
R3825 GND.n4180 GND.n4179 351.625
R3826 GND.n4180 GND.n75 351.625
R3827 GND.n4197 GND.n63 351.625
R3828 GND.n4202 GND.n63 351.625
R3829 GND.n4209 GND.n4208 351.625
R3830 GND.n4209 GND.n54 351.625
R3831 GND.n4226 GND.n42 351.625
R3832 GND.n4231 GND.n42 351.625
R3833 GND.n3154 GND.n558 351.625
R3834 GND.n3149 GND.n558 351.625
R3835 GND.n2773 GND.t435 349.135
R3836 GND.n2779 GND.t435 349.135
R3837 GND.n2780 GND.t7 349.135
R3838 GND.t2 GND.n2858 349.135
R3839 GND.n2857 GND.t467 349.135
R3840 GND.n2847 GND.t668 349.135
R3841 GND.n2846 GND.t331 349.135
R3842 GND.n2486 GND.t331 349.135
R3843 GND.n2487 GND.t674 349.135
R3844 GND.n2836 GND.t674 349.135
R3845 GND.n2836 GND.t210 349.135
R3846 GND.n2809 GND.t210 349.135
R3847 GND.n2810 GND.t495 349.135
R3848 GND.t284 GND.n633 349.135
R3849 GND.n1620 GND.t279 348.704
R3850 GND.t21 GND.n1904 336.942
R3851 GND.n2980 GND.n2979 326.113
R3852 GND.n2967 GND.n2966 326.113
R3853 GND.n2954 GND.n2953 326.113
R3854 GND.n2905 GND.n2904 326.113
R3855 GND.n2931 GND.n2930 326.113
R3856 GND.n2448 GND.n2447 326.113
R3857 GND.n2435 GND.n2434 326.113
R3858 GND.n2422 GND.n2421 326.113
R3859 GND.n2373 GND.n2372 326.113
R3860 GND.n2399 GND.n2398 326.113
R3861 GND.n2321 GND.n2320 326.113
R3862 GND.n2308 GND.n2307 326.113
R3863 GND.n2295 GND.n2294 326.113
R3864 GND.n2246 GND.n2245 326.113
R3865 GND.n2272 GND.n2271 326.113
R3866 GND.n2643 GND.n2642 326.113
R3867 GND.n2630 GND.n2629 326.113
R3868 GND.n2617 GND.n2616 326.113
R3869 GND.n2568 GND.n2567 326.113
R3870 GND.n2594 GND.n2593 326.113
R3871 GND.n2764 GND.n2763 326.113
R3872 GND.n2751 GND.n2750 326.113
R3873 GND.n2738 GND.n2737 326.113
R3874 GND.n2689 GND.n2688 326.113
R3875 GND.n2715 GND.n2714 326.113
R3876 GND.n3113 GND.n3112 326.113
R3877 GND.n3100 GND.n3099 326.113
R3878 GND.n3087 GND.n3086 326.113
R3879 GND.n619 GND.n618 326.113
R3880 GND.n3064 GND.n3063 326.113
R3881 GND.n2992 GND.n2991 321.531
R3882 GND.n1143 GND.n1142 306.584
R3883 GND.n2144 GND.n2143 306.584
R3884 GND.n2063 GND.n2062 306.584
R3885 GND.n1980 GND.n1979 306.584
R3886 GND.n1054 GND.n1050 290.815
R3887 GND.t618 GND.n381 281.065
R3888 GND.n3386 GND.t618 281.065
R3889 GND.n3385 GND.t443 281.065
R3890 GND.n3358 GND.t443 281.065
R3891 GND.n3358 GND.t305 281.065
R3892 GND.t305 GND.n371 281.065
R3893 GND.n3346 GND.t358 281.065
R3894 GND.t358 GND.n3345 281.065
R3895 GND.n3345 GND.t671 281.065
R3896 GND.n3396 GND.t671 281.065
R3897 GND.t29 GND.n350 281.065
R3898 GND.n3371 GND.t29 281.065
R3899 GND.n3371 GND.t81 281.065
R3900 GND.t81 GND.n342 281.065
R3901 GND.t355 GND.n24 281.065
R3902 GND.n527 GND.t355 281.065
R3903 GND.n529 GND.t835 281.065
R3904 GND.t835 GND.n528 281.065
R3905 GND.n528 GND.t324 281.065
R3906 GND.n3267 GND.t324 281.065
R3907 GND.t836 GND.n3121 275.505
R3908 GND.t791 GND.n570 275.505
R3909 GND.t397 GND.n3132 275.505
R3910 GND.n3135 GND.t858 275.505
R3911 GND.n3134 GND.t793 275.505
R3912 GND.n3145 GND.t793 275.505
R3913 GND.n3147 GND.t252 275.505
R3914 GND.t252 GND.n3146 275.505
R3915 GND.n3146 GND.t43 275.505
R3916 GND.n3156 GND.t43 275.505
R3917 GND.n3157 GND.t420 275.505
R3918 GND.n3167 GND.t72 275.505
R3919 GND.n1936 GND.t678 274.82
R3920 GND.t685 GND.n1945 274.82
R3921 GND.n4160 GND.n4159 274.736
R3922 GND.n3679 GND.n3678 274.736
R3923 GND.n4131 GND.n4130 274.736
R3924 GND.n4124 GND.n4123 274.736
R3925 GND.n4110 GND.n4109 274.736
R3926 GND.n4086 GND.n4085 274.736
R3927 GND.n4079 GND.n4078 274.736
R3928 GND.n4065 GND.n4064 274.736
R3929 GND.n3832 GND.n3831 274.736
R3930 GND.n4036 GND.n4035 274.736
R3931 GND.n4029 GND.n4028 274.736
R3932 GND.n4015 GND.n4014 274.736
R3933 GND.n3991 GND.n3990 274.736
R3934 GND.n3984 GND.n3983 274.736
R3935 GND.n3970 GND.n3969 274.736
R3936 GND.n1657 GND.n1656 260.592
R3937 GND.n1647 GND.n1646 260.592
R3938 GND.n1023 GND.n1022 260.592
R3939 GND.n1027 GND.n1026 260.592
R3940 GND.n1081 GND.n1080 260.592
R3941 GND.n1126 GND.n1125 260.592
R3942 GND.n1098 GND.n1097 260.592
R3943 GND.n1104 GND.n1103 260.592
R3944 GND.n1733 GND.n1732 260.592
R3945 GND.n1723 GND.n1722 260.592
R3946 GND.n1058 GND.n1057 260.592
R3947 GND.n1573 GND.n1572 260.592
R3948 GND.n1756 GND.n1755 260.592
R3949 GND.n2135 GND.n2134 260.592
R3950 GND.n2125 GND.n2124 260.592
R3951 GND.n661 GND.n660 260.592
R3952 GND.n2113 GND.n2112 260.592
R3953 GND.n735 GND.n733 260.592
R3954 GND.n747 GND.n745 260.592
R3955 GND.n748 GND.n47 260.592
R3956 GND.n768 GND.n767 260.592
R3957 GND.n2052 GND.n2051 260.592
R3958 GND.n2042 GND.n2041 260.592
R3959 GND.n792 GND.n791 260.592
R3960 GND.n2030 GND.n2029 260.592
R3961 GND.n1423 GND.n1422 260.592
R3962 GND.n1413 GND.n1412 260.592
R3963 GND.n1374 GND.n68 260.592
R3964 GND.n1399 GND.n1398 260.592
R3965 GND.n1969 GND.n1968 260.592
R3966 GND.n1959 GND.n1958 260.592
R3967 GND.n841 GND.n82 260.257
R3968 GND.n1035 GND.t229 255.716
R3969 GND.n1758 GND.n104 246.612
R3970 GND.n1606 GND.t646 242.552
R3971 GND.n4234 GND.t66 242.552
R3972 GND.n4205 GND.t412 242.552
R3973 GND.n4178 GND.n4177 242.542
R3974 GND.n4040 GND.n4039 236.048
R3975 GND.n4039 GND.n4038 236.048
R3976 GND.n4090 GND.n4089 236.048
R3977 GND.n4089 GND.n4088 236.048
R3978 GND.n4135 GND.n4134 236.048
R3979 GND.n4134 GND.n4133 236.048
R3980 GND.n3594 GND.n3593 236.048
R3981 GND.n3593 GND.n3592 236.048
R3982 GND.n3186 GND.n3185 236.048
R3983 GND.n3187 GND.n3186 236.048
R3984 GND.n607 GND.n606 236.048
R3985 GND.n3084 GND.n606 236.048
R3986 GND.n2148 GND.n2147 236.048
R3987 GND.n3047 GND.n2147 236.048
R3988 GND.n1043 GND.n1042 236.048
R3989 GND.n1590 GND.n1042 236.048
R3990 GND.n1274 GND.n1208 236.048
R3991 GND.n1208 GND.n1206 236.048
R3992 GND.n2068 GND.n2067 236.048
R3993 GND.n2069 GND.n2068 236.048
R3994 GND.n1187 GND.n1185 236.048
R3995 GND.n1353 GND.n1187 236.048
R3996 GND.n1985 GND.n1984 236.048
R3997 GND.n1986 GND.n1985 236.048
R3998 GND.n1720 GND.n873 236.048
R3999 GND.n874 GND.n873 236.048
R4000 GND.n1123 GND.n1084 236.048
R4001 GND.n1085 GND.n1084 236.048
R4002 GND.n1644 GND.n923 236.048
R4003 GND.n924 GND.n923 236.048
R4004 GND.n935 GND.n933 236.048
R4005 GND.n1624 GND.n935 236.048
R4006 GND.n1674 GND.n1673 236.048
R4007 GND.n1673 GND.n1672 236.048
R4008 GND.n1564 GND.n1563 236.048
R4009 GND.n1565 GND.n1564 236.048
R4010 GND.n1166 GND.n1164 236.048
R4011 GND.n1505 GND.n1166 236.048
R4012 GND.n845 GND.n844 236.048
R4013 GND.n1956 GND.n844 236.048
R4014 GND.n1376 GND.n1373 236.048
R4015 GND.n1410 GND.n1373 236.048
R4016 GND.n786 GND.n785 236.048
R4017 GND.n2039 GND.n785 236.048
R4018 GND.n750 GND.n713 236.048
R4019 GND.n713 GND.n711 236.048
R4020 GND.n3211 GND.n3209 236.048
R4021 GND.n3247 GND.n3211 236.048
R4022 GND.n3291 GND.n500 236.048
R4023 GND.n501 GND.n500 236.048
R4024 GND.n3502 GND.n3473 236.048
R4025 GND.n3474 GND.n3473 236.048
R4026 GND.n3531 GND.n3530 236.048
R4027 GND.n3532 GND.n3531 236.048
R4028 GND.n424 GND.n422 236.048
R4029 GND.n483 GND.n424 236.048
R4030 GND.n3354 GND.n3352 236.048
R4031 GND.n3388 GND.n3354 236.048
R4032 GND.n395 GND.n394 236.048
R4033 GND.n3420 GND.n394 236.048
R4034 GND.n171 GND.n170 236.048
R4035 GND.n4055 GND.n170 236.048
R4036 GND.n112 GND.n111 236.048
R4037 GND.n4150 GND.n111 236.048
R4038 GND.n3620 GND.n329 236.048
R4039 GND.n330 GND.n329 236.048
R4040 GND.n236 GND.n234 236.048
R4041 GND.n3925 GND.n236 236.048
R4042 GND.n255 GND.n254 236.048
R4043 GND.n3856 GND.n254 236.048
R4044 GND.n286 GND.n284 236.048
R4045 GND.n3763 GND.n286 236.048
R4046 GND.n305 GND.n304 236.048
R4047 GND.n3703 GND.n304 236.048
R4048 GND.n11 GND.n9 236.048
R4049 GND.n4282 GND.n11 236.048
R4050 GND.n525 GND.n520 236.048
R4051 GND.n522 GND.n520 236.048
R4052 GND.n655 GND.n654 236.048
R4053 GND.n2122 GND.n654 236.048
R4054 GND.n2995 GND.n2994 236.048
R4055 GND.n2996 GND.n2995 236.048
R4056 GND.n2477 GND.n2476 236.048
R4057 GND.n2844 GND.n2476 236.048
R4058 GND.n2776 GND.n2775 236.048
R4059 GND.n2777 GND.n2776 236.048
R4060 GND.n2893 GND.n2892 236.048
R4061 GND.n2951 GND.n2892 236.048
R4062 GND.n2984 GND.n2983 236.048
R4063 GND.n2983 GND.n2982 236.048
R4064 GND.n2361 GND.n2360 236.048
R4065 GND.n2419 GND.n2360 236.048
R4066 GND.n2449 GND.n2330 236.048
R4067 GND.n2449 GND.n2331 236.048
R4068 GND.n2234 GND.n2233 236.048
R4069 GND.n2292 GND.n2233 236.048
R4070 GND.n2322 GND.n2202 236.048
R4071 GND.n2322 GND.n2203 236.048
R4072 GND.n2556 GND.n2555 236.048
R4073 GND.n2614 GND.n2555 236.048
R4074 GND.n2644 GND.n2524 236.048
R4075 GND.n2644 GND.n2525 236.048
R4076 GND.n2677 GND.n2676 236.048
R4077 GND.n2735 GND.n2676 236.048
R4078 GND.n2768 GND.n2767 236.048
R4079 GND.n2767 GND.n2766 236.048
R4080 GND.n73 GND.n72 236.048
R4081 GND.n4190 GND.n72 236.048
R4082 GND.n52 GND.n51 236.048
R4083 GND.n4219 GND.n51 236.048
R4084 GND.n3143 GND.n563 236.048
R4085 GND.n564 GND.n563 236.048
R4086 GND.n3117 GND.n3116 236.048
R4087 GND.n3116 GND.n3115 236.048
R4088 GND.n3994 GND.n3993 236.048
R4089 GND.n3995 GND.n3994 236.048
R4090 GND.n3446 GND.n3445 227.064
R4091 GND.n3528 GND.n3527 227.064
R4092 GND.n3268 GND.n513 227.064
R4093 GND.n4258 GND.n4257 227.064
R4094 GND.t377 GND.n1909 217.311
R4095 GND.t696 GND.n1912 217.311
R4096 GND.n1822 GND.t589 215.714
R4097 GND.t96 GND.n1821 215.714
R4098 GND.n4235 GND.n4234 204.013
R4099 GND.n2992 GND.t741 203.526
R4100 GND.n2998 GND.t741 203.526
R4101 GND.n2999 GND.t424 203.526
R4102 GND.n3005 GND.t593 203.526
R4103 GND.n3006 GND.t393 203.526
R4104 GND.n3012 GND.t861 203.526
R4105 GND.n3014 GND.t265 203.526
R4106 GND.t265 GND.n3013 203.526
R4107 GND.n3013 GND.t872 203.526
R4108 GND.n3020 GND.t872 203.526
R4109 GND.t614 GND.n3021 203.526
R4110 GND.t402 GND.n639 203.526
R4111 GND.n481 GND.n480 192.982
R4112 GND.n474 GND.n473 192.982
R4113 GND.n460 GND.n459 192.982
R4114 GND.n3535 GND.n3534 192.982
R4115 GND.n3542 GND.n3541 192.982
R4116 GND.n3565 GND.n3564 192.982
R4117 GND.n3245 GND.n3244 192.982
R4118 GND.n3238 GND.n3237 192.982
R4119 GND.n3337 GND.n3336 192.982
R4120 GND.n3190 GND.n3189 192.982
R4121 GND.n4236 GND.n38 192.982
R4122 GND.n4251 GND.n4250 192.982
R4123 GND.n3590 GND.n3589 192.982
R4124 GND.n1906 GND.n1905 192.982
R4125 GND.n1939 GND.t328 190.261
R4126 GND.t373 GND.n1938 190.261
R4127 GND.n1758 GND.n1757 181.749
R4128 GND.n4206 GND.t673 179.623
R4129 GND.n1863 GND.t679 176.65
R4130 GND.n1868 GND.t203 176.65
R4131 GND.n1873 GND.t700 176.65
R4132 GND.n1878 GND.t283 176.65
R4133 GND.n1883 GND.t877 176.65
R4134 GND.n1888 GND.t463 176.65
R4135 GND.n1893 GND.t786 176.65
R4136 GND.n1894 GND.t73 176.65
R4137 GND.n2141 GND.n2140 176.091
R4138 GND.n1244 GND.n1242 176.091
R4139 GND.n1795 GND.n1794 174.518
R4140 GND.n1810 GND.n1809 174.518
R4141 GND.n1825 GND.n1824 174.518
R4142 GND.n1840 GND.n1839 174.518
R4143 GND.n1855 GND.n1854 174.518
R4144 GND.n1780 GND.n1779 174.518
R4145 GND.n1941 GND.n1935 174.518
R4146 GND.n3965 GND.n3963 173.012
R4147 GND.n3967 GND.n224 173.012
R4148 GND.n3972 GND.n220 173.012
R4149 GND.n3974 GND.n218 173.012
R4150 GND.n3979 GND.n215 173.012
R4151 GND.n3981 GND.n214 173.012
R4152 GND.n3986 GND.n211 173.012
R4153 GND.n3988 GND.n210 173.012
R4154 GND.n4010 GND.n198 173.012
R4155 GND.n4012 GND.n197 173.012
R4156 GND.n4017 GND.n193 173.012
R4157 GND.n4019 GND.n191 173.012
R4158 GND.n4024 GND.n187 173.012
R4159 GND.n4026 GND.n186 173.012
R4160 GND.n4031 GND.n183 173.012
R4161 GND.n4033 GND.n182 173.012
R4162 GND.n4038 GND.n179 173.012
R4163 GND.n4040 GND.n179 173.012
R4164 GND.n4060 GND.n167 173.012
R4165 GND.n4062 GND.n166 173.012
R4166 GND.n4067 GND.n162 173.012
R4167 GND.n4069 GND.n160 173.012
R4168 GND.n4074 GND.n157 173.012
R4169 GND.n4076 GND.n156 173.012
R4170 GND.n4081 GND.n153 173.012
R4171 GND.n4083 GND.n152 173.012
R4172 GND.n4088 GND.n149 173.012
R4173 GND.n4090 GND.n149 173.012
R4174 GND.n4105 GND.n140 173.012
R4175 GND.n4107 GND.n139 173.012
R4176 GND.n4112 GND.n135 173.012
R4177 GND.n4114 GND.n133 173.012
R4178 GND.n4119 GND.n129 173.012
R4179 GND.n4121 GND.n128 173.012
R4180 GND.n4126 GND.n125 173.012
R4181 GND.n4128 GND.n124 173.012
R4182 GND.n4133 GND.n121 173.012
R4183 GND.n4135 GND.n121 173.012
R4184 GND.n4155 GND.n108 173.012
R4185 GND.n4157 GND.n107 173.012
R4186 GND.n101 GND.n98 173.012
R4187 GND.n4164 GND.n97 173.012
R4188 GND.n90 GND.n89 173.012
R4189 GND.n87 GND.n86 173.012
R4190 GND.n3592 GND.n3588 173.012
R4191 GND.n3594 GND.n3588 173.012
R4192 GND.n4255 GND.n27 173.012
R4193 GND.n4253 GND.n28 173.012
R4194 GND.n4248 GND.n31 173.012
R4195 GND.n4246 GND.n33 173.012
R4196 GND.n4240 GND.n36 173.012
R4197 GND.n4238 GND.n37 173.012
R4198 GND.n3194 GND.n3193 173.012
R4199 GND.n546 GND.n545 173.012
R4200 GND.n3187 GND.n550 173.012
R4201 GND.n3185 GND.n550 173.012
R4202 GND.n3083 GND.n607 173.012
R4203 GND.n3084 GND.n3083 173.012
R4204 GND.n3036 GND.n3030 173.012
R4205 GND.n3042 GND.n3029 173.012
R4206 GND.n3046 GND.n2148 173.012
R4207 GND.n3047 GND.n3046 173.012
R4208 GND.n1611 GND.n1610 173.012
R4209 GND.n1616 GND.n1615 173.012
R4210 GND.n1597 GND.n1596 173.012
R4211 GND.n1602 GND.n1601 173.012
R4212 GND.n1589 GND.n1043 173.012
R4213 GND.n1590 GND.n1589 173.012
R4214 GND.n1789 GND.n1788 173.012
R4215 GND.n1804 GND.n1803 173.012
R4216 GND.n1819 GND.n1818 173.012
R4217 GND.n1834 GND.n1833 173.012
R4218 GND.n1849 GND.n1848 173.012
R4219 GND.n1774 GND.n1773 173.012
R4220 GND.n1275 GND.n1274 173.012
R4221 GND.n1275 GND.n1206 173.012
R4222 GND.n1268 GND.n1212 173.012
R4223 GND.n1266 GND.n1213 173.012
R4224 GND.n1261 GND.n1216 173.012
R4225 GND.n1259 GND.n1217 173.012
R4226 GND.n1254 GND.n1220 173.012
R4227 GND.n1252 GND.n1222 173.012
R4228 GND.n2067 GND.n695 173.012
R4229 GND.n2069 GND.n695 173.012
R4230 GND.n2074 GND.n692 173.012
R4231 GND.n2076 GND.n691 173.012
R4232 GND.n2081 GND.n688 173.012
R4233 GND.n2083 GND.n687 173.012
R4234 GND.n2088 GND.n683 173.012
R4235 GND.n2090 GND.n681 173.012
R4236 GND.n2095 GND.n678 173.012
R4237 GND.n2097 GND.n677 173.012
R4238 GND.n1354 GND.n1353 173.012
R4239 GND.n1354 GND.n1185 173.012
R4240 GND.n1347 GND.n1191 173.012
R4241 GND.n1345 GND.n1192 173.012
R4242 GND.n1340 GND.n1195 173.012
R4243 GND.n1338 GND.n1196 173.012
R4244 GND.n1333 GND.n1199 173.012
R4245 GND.n1331 GND.n1201 173.012
R4246 GND.n1325 GND.n1204 173.012
R4247 GND.n1323 GND.n1321 173.012
R4248 GND.n1984 GND.n826 173.012
R4249 GND.n1986 GND.n826 173.012
R4250 GND.n1991 GND.n823 173.012
R4251 GND.n1993 GND.n822 173.012
R4252 GND.n1998 GND.n819 173.012
R4253 GND.n2000 GND.n818 173.012
R4254 GND.n2005 GND.n814 173.012
R4255 GND.n2007 GND.n812 173.012
R4256 GND.n2012 GND.n809 173.012
R4257 GND.n2014 GND.n808 173.012
R4258 GND.n1753 GND.n1752 173.012
R4259 GND.n1748 GND.n1747 173.012
R4260 GND.n1709 GND.n880 173.012
R4261 GND.n1707 GND.n882 173.012
R4262 GND.n1715 GND.n876 173.012
R4263 GND.n1713 GND.n878 173.012
R4264 GND.n1720 GND.n1719 173.012
R4265 GND.n1719 GND.n874 173.012
R4266 GND.n1730 GND.n1729 173.012
R4267 GND.n1726 GND.n1725 173.012
R4268 GND.n1741 GND.n1740 173.012
R4269 GND.n1736 GND.n1735 173.012
R4270 GND.n1112 GND.n1092 173.012
R4271 GND.n1110 GND.n1107 173.012
R4272 GND.n1118 GND.n1088 173.012
R4273 GND.n1116 GND.n1090 173.012
R4274 GND.n1123 GND.n1122 173.012
R4275 GND.n1122 GND.n1085 173.012
R4276 GND.n1133 GND.n1074 173.012
R4277 GND.n1127 GND.n1075 173.012
R4278 GND.n1140 GND.n1139 173.012
R4279 GND.n1078 GND.n1072 173.012
R4280 GND.n1633 GND.n930 173.012
R4281 GND.n1631 GND.n932 173.012
R4282 GND.n1639 GND.n926 173.012
R4283 GND.n1637 GND.n928 173.012
R4284 GND.n1644 GND.n1643 173.012
R4285 GND.n1643 GND.n924 173.012
R4286 GND.n1654 GND.n1653 173.012
R4287 GND.n1650 GND.n1649 173.012
R4288 GND.n1665 GND.n1664 173.012
R4289 GND.n1660 GND.n1659 173.012
R4290 GND.n1625 GND.n1624 173.012
R4291 GND.n1625 GND.n933 173.012
R4292 GND.n1012 GND.n939 173.012
R4293 GND.n1010 GND.n940 173.012
R4294 GND.n1005 GND.n943 173.012
R4295 GND.n1003 GND.n944 173.012
R4296 GND.n998 GND.n947 173.012
R4297 GND.n996 GND.n949 173.012
R4298 GND.n990 GND.n952 173.012
R4299 GND.n988 GND.n986 173.012
R4300 GND.n1672 GND.n906 173.012
R4301 GND.n1674 GND.n906 173.012
R4302 GND.n1679 GND.n903 173.012
R4303 GND.n1681 GND.n902 173.012
R4304 GND.n1686 GND.n899 173.012
R4305 GND.n1688 GND.n898 173.012
R4306 GND.n893 GND.n890 173.012
R4307 GND.n1695 GND.n889 173.012
R4308 GND.n1699 GND.n887 173.012
R4309 GND.n1701 GND.n885 173.012
R4310 GND.n1565 GND.n1146 173.012
R4311 GND.n1563 GND.n1146 173.012
R4312 GND.n1558 GND.n1149 173.012
R4313 GND.n1556 GND.n1150 173.012
R4314 GND.n1551 GND.n1153 173.012
R4315 GND.n1549 GND.n1154 173.012
R4316 GND.n1544 GND.n1157 173.012
R4317 GND.n1542 GND.n1159 173.012
R4318 GND.n1536 GND.n1162 173.012
R4319 GND.n1534 GND.n1531 173.012
R4320 GND.n1506 GND.n1505 173.012
R4321 GND.n1506 GND.n1164 173.012
R4322 GND.n1498 GND.n1170 173.012
R4323 GND.n1496 GND.n1171 173.012
R4324 GND.n1491 GND.n1174 173.012
R4325 GND.n1489 GND.n1175 173.012
R4326 GND.n1484 GND.n1178 173.012
R4327 GND.n1482 GND.n1180 173.012
R4328 GND.n1476 GND.n1183 173.012
R4329 GND.n1474 GND.n1472 173.012
R4330 GND.n1946 GND.n848 173.012
R4331 GND.n1951 GND.n847 173.012
R4332 GND.n1955 GND.n845 173.012
R4333 GND.n1956 GND.n1955 173.012
R4334 GND.n1962 GND.n1961 173.012
R4335 GND.n1966 GND.n1965 173.012
R4336 GND.n1972 GND.n1971 173.012
R4337 GND.n1977 GND.n1976 173.012
R4338 GND.n1391 GND.n1390 173.012
R4339 GND.n1396 GND.n1395 173.012
R4340 GND.n1400 GND.n1379 173.012
R4341 GND.n1405 GND.n1378 173.012
R4342 GND.n1409 GND.n1376 173.012
R4343 GND.n1410 GND.n1409 173.012
R4344 GND.n1416 GND.n1415 173.012
R4345 GND.n1420 GND.n1419 173.012
R4346 GND.n1424 GND.n1360 173.012
R4347 GND.n1429 GND.n1359 173.012
R4348 GND.n2022 GND.n2021 173.012
R4349 GND.n2027 GND.n2026 173.012
R4350 GND.n796 GND.n789 173.012
R4351 GND.n2034 GND.n788 173.012
R4352 GND.n2038 GND.n786 173.012
R4353 GND.n2039 GND.n2038 173.012
R4354 GND.n2045 GND.n2044 173.012
R4355 GND.n2049 GND.n2048 173.012
R4356 GND.n2055 GND.n2054 173.012
R4357 GND.n2060 GND.n2059 173.012
R4358 GND.n772 GND.n771 173.012
R4359 GND.n760 GND.n759 173.012
R4360 GND.n765 GND.n764 173.012
R4361 GND.n756 GND.n755 173.012
R4362 GND.n751 GND.n750 173.012
R4363 GND.n751 GND.n711 173.012
R4364 GND.n743 GND.n742 173.012
R4365 GND.n738 GND.n737 173.012
R4366 GND.n731 GND.n730 173.012
R4367 GND.n725 GND.n724 173.012
R4368 GND.n3341 GND.n415 173.012
R4369 GND.n3339 GND.n416 173.012
R4370 GND.n3334 GND.n419 173.012
R4371 GND.n3332 GND.n3328 173.012
R4372 GND.n3233 GND.n3231 173.012
R4373 GND.n3235 GND.n3220 173.012
R4374 GND.n3240 GND.n3217 173.012
R4375 GND.n3242 GND.n3216 173.012
R4376 GND.n3248 GND.n3247 173.012
R4377 GND.n3248 GND.n3209 173.012
R4378 GND.n3313 GND.n3312 173.012
R4379 GND.n3301 GND.n3300 173.012
R4380 GND.n3306 GND.n3305 173.012
R4381 GND.n3298 GND.n3297 173.012
R4382 GND.n3291 GND.n3290 173.012
R4383 GND.n3290 GND.n501 173.012
R4384 GND.n3286 GND.n3285 173.012
R4385 GND.n3278 GND.n3277 173.012
R4386 GND.n3487 GND.n3486 173.012
R4387 GND.n3576 GND.n3575 173.012
R4388 GND.n3497 GND.n3477 173.012
R4389 GND.n3491 GND.n3478 173.012
R4390 GND.n3502 GND.n3501 173.012
R4391 GND.n3501 GND.n3474 173.012
R4392 GND.n3513 GND.n3512 173.012
R4393 GND.n3508 GND.n3507 173.012
R4394 GND.n3569 GND.n353 173.012
R4395 GND.n3567 GND.n354 173.012
R4396 GND.n3562 GND.n357 173.012
R4397 GND.n3560 GND.n3556 173.012
R4398 GND.n3546 GND.n3545 173.012
R4399 GND.n3452 GND.n3451 173.012
R4400 GND.n3539 GND.n366 173.012
R4401 GND.n3537 GND.n367 173.012
R4402 GND.n3532 GND.n370 173.012
R4403 GND.n3530 GND.n370 173.012
R4404 GND.n3449 GND.n3448 173.012
R4405 GND.n457 GND.n456 173.012
R4406 GND.n462 GND.n439 173.012
R4407 GND.n464 GND.n437 173.012
R4408 GND.n469 GND.n434 173.012
R4409 GND.n471 GND.n433 173.012
R4410 GND.n476 GND.n430 173.012
R4411 GND.n478 GND.n429 173.012
R4412 GND.n484 GND.n483 173.012
R4413 GND.n484 GND.n422 173.012
R4414 GND.n3383 GND.n3382 173.012
R4415 GND.n3379 GND.n3378 173.012
R4416 GND.n3389 GND.n3352 173.012
R4417 GND.n3389 GND.n3388 173.012
R4418 GND.n3437 GND.n3436 173.012
R4419 GND.n3442 GND.n3441 173.012
R4420 GND.n3427 GND.n3426 173.012
R4421 GND.n3431 GND.n3430 173.012
R4422 GND.n3419 GND.n395 173.012
R4423 GND.n3420 GND.n3419 173.012
R4424 GND.n3407 GND.n3406 173.012
R4425 GND.n3415 GND.n3414 173.012
R4426 GND.n3316 GND.n3315 173.012
R4427 GND.n3402 GND.n3401 173.012
R4428 GND.n3394 GND.n3393 173.012
R4429 GND.n3349 GND.n3348 173.012
R4430 GND.n3265 GND.n3264 173.012
R4431 GND.n532 GND.n531 173.012
R4432 GND.n4001 GND.n4000 173.012
R4433 GND.n4005 GND.n4004 173.012
R4434 GND.n4044 GND.n174 173.012
R4435 GND.n4050 GND.n173 173.012
R4436 GND.n4054 GND.n171 173.012
R4437 GND.n4055 GND.n4054 173.012
R4438 GND.n4096 GND.n4095 173.012
R4439 GND.n4100 GND.n4099 173.012
R4440 GND.n4139 GND.n116 173.012
R4441 GND.n4145 GND.n115 173.012
R4442 GND.n4149 GND.n112 173.012
R4443 GND.n4150 GND.n4149 173.012
R4444 GND.n3374 GND.n3364 173.012
R4445 GND.n3368 GND.n3365 173.012
R4446 GND.n3519 GND.n3518 173.012
R4447 GND.n3524 GND.n3523 173.012
R4448 GND.n3674 GND.n3673 173.012
R4449 GND.n3637 GND.n3636 173.012
R4450 GND.n3631 GND.n3630 173.012
R4451 GND.n3627 GND.n3626 173.012
R4452 GND.n3620 GND.n3619 173.012
R4453 GND.n3619 GND.n330 173.012
R4454 GND.n3615 GND.n3614 173.012
R4455 GND.n3607 GND.n3606 173.012
R4456 GND.n3602 GND.n3601 173.012
R4457 GND.n3579 GND.n3578 173.012
R4458 GND.n3910 GND.n3909 173.012
R4459 GND.n3905 GND.n3904 173.012
R4460 GND.n3920 GND.n3919 173.012
R4461 GND.n3916 GND.n3915 173.012
R4462 GND.n3926 GND.n234 173.012
R4463 GND.n3926 GND.n3925 173.012
R4464 GND.n3932 GND.n231 173.012
R4465 GND.n3930 GND.n233 173.012
R4466 GND.n3873 GND.n3872 173.012
R4467 GND.n3878 GND.n3877 173.012
R4468 GND.n3863 GND.n3862 173.012
R4469 GND.n3867 GND.n3866 173.012
R4470 GND.n3855 GND.n255 173.012
R4471 GND.n3856 GND.n3855 173.012
R4472 GND.n3843 GND.n3842 173.012
R4473 GND.n3851 GND.n3850 173.012
R4474 GND.n273 GND.n272 173.012
R4475 GND.n3838 GND.n3837 173.012
R4476 GND.n3748 GND.n3747 173.012
R4477 GND.n3827 GND.n3826 173.012
R4478 GND.n3758 GND.n3757 173.012
R4479 GND.n3754 GND.n3753 173.012
R4480 GND.n3764 GND.n284 173.012
R4481 GND.n3764 GND.n3763 173.012
R4482 GND.n3770 GND.n281 173.012
R4483 GND.n3768 GND.n283 173.012
R4484 GND.n3776 GND.n277 173.012
R4485 GND.n3774 GND.n279 173.012
R4486 GND.n3720 GND.n3719 173.012
R4487 GND.n3725 GND.n3724 173.012
R4488 GND.n3710 GND.n3709 173.012
R4489 GND.n3714 GND.n3713 173.012
R4490 GND.n3702 GND.n305 173.012
R4491 GND.n3703 GND.n3702 173.012
R4492 GND.n3690 GND.n3689 173.012
R4493 GND.n3698 GND.n3697 173.012
R4494 GND.n3641 GND.n3640 173.012
R4495 GND.n3685 GND.n3684 173.012
R4496 GND.n3936 GND.n229 173.012
R4497 GND.n3938 GND.n227 173.012
R4498 GND.n4267 GND.n4266 173.012
R4499 GND.n4262 GND.n4261 173.012
R4500 GND.n4277 GND.n4276 173.012
R4501 GND.n4273 GND.n4272 173.012
R4502 GND.n4283 GND.n9 173.012
R4503 GND.n4283 GND.n4282 173.012
R4504 GND.n4289 GND.n6 173.012
R4505 GND.n4287 GND.n8 173.012
R4506 GND.n4293 GND.n4 173.012
R4507 GND.n4295 GND.n2 173.012
R4508 GND.n3253 GND.n3252 173.012
R4509 GND.n3273 GND.n3272 173.012
R4510 GND.n525 GND.n524 173.012
R4511 GND.n524 GND.n522 173.012
R4512 GND.n2105 GND.n2104 173.012
R4513 GND.n2110 GND.n2109 173.012
R4514 GND.n665 GND.n658 173.012
R4515 GND.n2117 GND.n657 173.012
R4516 GND.n2121 GND.n655 173.012
R4517 GND.n2122 GND.n2121 173.012
R4518 GND.n2128 GND.n2127 173.012
R4519 GND.n2132 GND.n2131 173.012
R4520 GND.n2138 GND.n2137 173.012
R4521 GND.n1246 GND.n1225 173.012
R4522 GND.n3025 GND.n3024 173.012
R4523 GND.n2183 GND.n2182 173.012
R4524 GND.n3018 GND.n2156 173.012
R4525 GND.n3016 GND.n2158 173.012
R4526 GND.n3010 GND.n2161 173.012
R4527 GND.n3008 GND.n2162 173.012
R4528 GND.n3003 GND.n2165 173.012
R4529 GND.n3001 GND.n2166 173.012
R4530 GND.n2996 GND.n2169 173.012
R4531 GND.n2994 GND.n2169 173.012
R4532 GND.n2821 GND.n2820 173.012
R4533 GND.n2816 GND.n2813 173.012
R4534 GND.n2833 GND.n2481 173.012
R4535 GND.n2839 GND.n2480 173.012
R4536 GND.n2843 GND.n2477 173.012
R4537 GND.n2844 GND.n2843 173.012
R4538 GND.n2850 GND.n2849 173.012
R4539 GND.n2855 GND.n2854 173.012
R4540 GND.n2864 GND.n2459 173.012
R4541 GND.n2859 GND.n2460 173.012
R4542 GND.n2805 GND.n2802 173.012
R4543 GND.n2826 GND.n2800 173.012
R4544 GND.n2830 GND.n2493 173.012
R4545 GND.n2491 GND.n2490 173.012
R4546 GND.n2795 GND.n2794 173.012
R4547 GND.n2790 GND.n2789 173.012
R4548 GND.n2785 GND.n2784 173.012
R4549 GND.n2782 GND.n2498 173.012
R4550 GND.n2777 GND.n2506 173.012
R4551 GND.n2775 GND.n2506 173.012
R4552 GND.n2950 GND.n2893 173.012
R4553 GND.n2951 GND.n2950 173.012
R4554 GND.n2982 GND.n2175 173.012
R4555 GND.n2984 GND.n2175 173.012
R4556 GND.n2418 GND.n2361 173.012
R4557 GND.n2419 GND.n2418 173.012
R4558 GND.n2452 GND.n2331 173.012
R4559 GND.n2452 GND.n2330 173.012
R4560 GND.n2291 GND.n2234 173.012
R4561 GND.n2292 GND.n2291 173.012
R4562 GND.n2325 GND.n2203 173.012
R4563 GND.n2325 GND.n2202 173.012
R4564 GND.n2613 GND.n2556 173.012
R4565 GND.n2614 GND.n2613 173.012
R4566 GND.n2647 GND.n2525 173.012
R4567 GND.n2647 GND.n2524 173.012
R4568 GND.n2734 GND.n2677 173.012
R4569 GND.n2735 GND.n2734 173.012
R4570 GND.n2766 GND.n2509 173.012
R4571 GND.n2768 GND.n2509 173.012
R4572 GND.n1943 GND.n1761 173.012
R4573 GND.n1918 GND.n1857 173.012
R4574 GND.n1913 GND.n1901 173.012
R4575 GND.n4168 GND.n95 173.012
R4576 GND.n4170 GND.n93 173.012
R4577 GND.n1584 GND.n1583 173.012
R4578 GND.n1052 GND.n1051 173.012
R4579 GND.n4179 GND.n76 173.012
R4580 GND.n4185 GND.n75 173.012
R4581 GND.n4189 GND.n73 173.012
R4582 GND.n4190 GND.n4189 173.012
R4583 GND.n4198 GND.n4197 173.012
R4584 GND.n4202 GND.n4201 173.012
R4585 GND.n4208 GND.n55 173.012
R4586 GND.n4214 GND.n54 173.012
R4587 GND.n4218 GND.n52 173.012
R4588 GND.n4219 GND.n4218 173.012
R4589 GND.n4227 GND.n4226 173.012
R4590 GND.n4231 GND.n4230 173.012
R4591 GND.n3165 GND.n3164 173.012
R4592 GND.n3160 GND.n3159 173.012
R4593 GND.n3154 GND.n3153 173.012
R4594 GND.n3150 GND.n3149 173.012
R4595 GND.n3143 GND.n3142 173.012
R4596 GND.n3142 GND.n564 173.012
R4597 GND.n3138 GND.n3137 173.012
R4598 GND.n3130 GND.n3129 173.012
R4599 GND.n3125 GND.n3124 173.012
R4600 GND.n2517 GND.n2516 173.012
R4601 GND.n3115 GND.n579 173.012
R4602 GND.n3117 GND.n579 173.012
R4603 GND.n3993 GND.n207 173.012
R4604 GND.n3995 GND.n207 173.012
R4605 GND.n2987 GND.n2986 163.056
R4606 GND.n3050 GND.n634 163.056
R4607 GND.n2988 GND.n2172 163.056
R4608 GND.n3050 GND.n635 163.056
R4609 GND.n2206 GND.n2170 163.056
R4610 GND.n3050 GND.n636 163.056
R4611 GND.n3050 GND.n637 163.056
R4612 GND.n3050 GND.n638 163.056
R4613 GND.n3051 GND.n3050 163.056
R4614 GND.t821 GND.n82 152.346
R4615 GND.n3060 GND.n625 150.213
R4616 GND.n3054 GND.n628 150.213
R4617 GND.n3054 GND.n3053 150.213
R4618 GND.n3061 GND.n3060 150.213
R4619 GND.n3067 GND.n610 150.213
R4620 GND.n3071 GND.n3069 150.213
R4621 GND.n3072 GND.n3071 150.213
R4622 GND.n3066 GND.n610 150.213
R4623 GND.n3096 GND.n596 150.213
R4624 GND.n3090 GND.n599 150.213
R4625 GND.n3090 GND.n3089 150.213
R4626 GND.n3097 GND.n3096 150.213
R4627 GND.n3109 GND.n584 150.213
R4628 GND.n3103 GND.n587 150.213
R4629 GND.n3103 GND.n3102 150.213
R4630 GND.n3110 GND.n3109 150.213
R4631 GND.n2927 GND.n2911 150.213
R4632 GND.n2921 GND.n2918 150.213
R4633 GND.n2921 GND.n2920 150.213
R4634 GND.n2928 GND.n2927 150.213
R4635 GND.n2934 GND.n2896 150.213
R4636 GND.n2938 GND.n2936 150.213
R4637 GND.n2939 GND.n2938 150.213
R4638 GND.n2933 GND.n2896 150.213
R4639 GND.n2963 GND.n2882 150.213
R4640 GND.n2957 GND.n2885 150.213
R4641 GND.n2957 GND.n2956 150.213
R4642 GND.n2964 GND.n2963 150.213
R4643 GND.n2976 GND.n2180 150.213
R4644 GND.n2970 GND.n2873 150.213
R4645 GND.n2970 GND.n2969 150.213
R4646 GND.n2977 GND.n2976 150.213
R4647 GND.n2395 GND.n2379 150.213
R4648 GND.n2389 GND.n2386 150.213
R4649 GND.n2389 GND.n2388 150.213
R4650 GND.n2396 GND.n2395 150.213
R4651 GND.n2402 GND.n2364 150.213
R4652 GND.n2406 GND.n2404 150.213
R4653 GND.n2407 GND.n2406 150.213
R4654 GND.n2401 GND.n2364 150.213
R4655 GND.n2431 GND.n2350 150.213
R4656 GND.n2425 GND.n2353 150.213
R4657 GND.n2425 GND.n2424 150.213
R4658 GND.n2432 GND.n2431 150.213
R4659 GND.n2444 GND.n2338 150.213
R4660 GND.n2438 GND.n2341 150.213
R4661 GND.n2438 GND.n2437 150.213
R4662 GND.n2445 GND.n2444 150.213
R4663 GND.n2268 GND.n2252 150.213
R4664 GND.n2262 GND.n2259 150.213
R4665 GND.n2262 GND.n2261 150.213
R4666 GND.n2269 GND.n2268 150.213
R4667 GND.n2275 GND.n2237 150.213
R4668 GND.n2279 GND.n2277 150.213
R4669 GND.n2280 GND.n2279 150.213
R4670 GND.n2274 GND.n2237 150.213
R4671 GND.n2304 GND.n2223 150.213
R4672 GND.n2298 GND.n2226 150.213
R4673 GND.n2298 GND.n2297 150.213
R4674 GND.n2305 GND.n2304 150.213
R4675 GND.n2317 GND.n2211 150.213
R4676 GND.n2311 GND.n2214 150.213
R4677 GND.n2311 GND.n2310 150.213
R4678 GND.n2318 GND.n2317 150.213
R4679 GND.n2590 GND.n2574 150.213
R4680 GND.n2584 GND.n2581 150.213
R4681 GND.n2584 GND.n2583 150.213
R4682 GND.n2591 GND.n2590 150.213
R4683 GND.n2597 GND.n2559 150.213
R4684 GND.n2601 GND.n2599 150.213
R4685 GND.n2602 GND.n2601 150.213
R4686 GND.n2596 GND.n2559 150.213
R4687 GND.n2626 GND.n2545 150.213
R4688 GND.n2620 GND.n2548 150.213
R4689 GND.n2620 GND.n2619 150.213
R4690 GND.n2627 GND.n2626 150.213
R4691 GND.n2639 GND.n2533 150.213
R4692 GND.n2633 GND.n2536 150.213
R4693 GND.n2633 GND.n2632 150.213
R4694 GND.n2640 GND.n2639 150.213
R4695 GND.n2711 GND.n2695 150.213
R4696 GND.n2705 GND.n2702 150.213
R4697 GND.n2705 GND.n2704 150.213
R4698 GND.n2712 GND.n2711 150.213
R4699 GND.n2718 GND.n2680 150.213
R4700 GND.n2722 GND.n2720 150.213
R4701 GND.n2723 GND.n2722 150.213
R4702 GND.n2717 GND.n2680 150.213
R4703 GND.n2747 GND.n2666 150.213
R4704 GND.n2741 GND.n2669 150.213
R4705 GND.n2741 GND.n2740 150.213
R4706 GND.n2748 GND.n2747 150.213
R4707 GND.n2760 GND.n2514 150.213
R4708 GND.n2754 GND.n2657 150.213
R4709 GND.n2754 GND.n2753 150.213
R4710 GND.n2761 GND.n2760 150.213
R4711 GND.n2780 GND.n2779 147.843
R4712 GND.n2858 GND.n2857 147.843
R4713 GND.n2847 GND.n2846 147.843
R4714 GND.n2487 GND.n2486 147.843
R4715 GND.n2810 GND.n2809 147.843
R4716 GND.t505 GND.n4235 143.995
R4717 GND.n3680 GND.t469 137.369
R4718 GND.n3833 GND.t838 137.369
R4719 GND.n1777 GND.n841 127.168
R4720 GND.n1776 GND.n1758 127.168
R4721 GND.n1938 GND.n1936 124.918
R4722 GND.t377 GND.t694 119.632
R4723 GND.t696 GND.t781 119.632
R4724 GND.n3386 GND.n3385 119.019
R4725 GND.n529 GND.n527 119.019
R4726 GND.n4117 GND.n130 118.349
R4727 GND.n4022 GND.n188 118.349
R4728 GND.n3132 GND.n570 116.663
R4729 GND.n3135 GND.n3134 116.663
R4730 GND.n3147 GND.n3145 116.663
R4731 GND.n3157 GND.n3156 116.663
R4732 GND.n1580 GND.n1058 112.255
R4733 GND.n4223 GND.n47 112.255
R4734 GND.n4194 GND.n68 112.255
R4735 GND.n1807 GND.n841 106.32
R4736 GND.n1806 GND.n1758 106.32
R4737 GND.n1837 GND.n841 106.32
R4738 GND.n1836 GND.n1758 106.32
R4739 GND.n1792 GND.n841 106.32
R4740 GND.n1791 GND.n1758 106.32
R4741 GND.n1852 GND.n841 106.162
R4742 GND.n1851 GND.n1758 106.162
R4743 GND.n3963 GND.n225 105.082
R4744 GND.n225 GND.n224 105.082
R4745 GND.n3953 GND.n215 105.082
R4746 GND.n3953 GND.n214 105.082
R4747 GND.n3948 GND.n211 105.082
R4748 GND.n3948 GND.n210 105.082
R4749 GND.n3803 GND.n198 105.082
R4750 GND.n3803 GND.n197 105.082
R4751 GND.n3811 GND.n187 105.082
R4752 GND.n3811 GND.n186 105.082
R4753 GND.n3816 GND.n183 105.082
R4754 GND.n3816 GND.n182 105.082
R4755 GND.n3799 GND.n167 105.082
R4756 GND.n3799 GND.n166 105.082
R4757 GND.n3791 GND.n157 105.082
R4758 GND.n3791 GND.n156 105.082
R4759 GND.n3786 GND.n153 105.082
R4760 GND.n3786 GND.n152 105.082
R4761 GND.n3650 GND.n140 105.082
R4762 GND.n3650 GND.n139 105.082
R4763 GND.n3658 GND.n129 105.082
R4764 GND.n3658 GND.n128 105.082
R4765 GND.n3663 GND.n125 105.082
R4766 GND.n3663 GND.n124 105.082
R4767 GND.n3646 GND.n108 105.082
R4768 GND.n3646 GND.n107 105.082
R4769 GND.n4175 GND.n90 105.082
R4770 GND.n4175 GND.n86 105.082
R4771 GND.n3206 GND.n27 105.082
R4772 GND.n3206 GND.n28 105.082
R4773 GND.n3198 GND.n36 105.082
R4774 GND.n3198 GND.n37 105.082
R4775 GND.n3194 GND.n537 105.082
R4776 GND.n546 GND.n537 105.082
R4777 GND.n1788 GND.n1782 105.082
R4778 GND.n1803 GND.n1797 105.082
R4779 GND.n1818 GND.n1812 105.082
R4780 GND.n1833 GND.n1827 105.082
R4781 GND.n1848 GND.n1842 105.082
R4782 GND.n1773 GND.n1767 105.082
R4783 GND.n1229 GND.n1213 105.082
R4784 GND.n1229 GND.n1212 105.082
R4785 GND.n1234 GND.n1217 105.082
R4786 GND.n1234 GND.n1216 105.082
R4787 GND.n1296 GND.n691 105.082
R4788 GND.n1296 GND.n692 105.082
R4789 GND.n1291 GND.n687 105.082
R4790 GND.n1291 GND.n688 105.082
R4791 GND.n1283 GND.n677 105.082
R4792 GND.n1283 GND.n678 105.082
R4793 GND.n1306 GND.n1191 105.082
R4794 GND.n1306 GND.n1192 105.082
R4795 GND.n1311 GND.n1195 105.082
R4796 GND.n1311 GND.n1196 105.082
R4797 GND.n1321 GND.n1205 105.082
R4798 GND.n1205 GND.n1204 105.082
R4799 GND.n1447 GND.n822 105.082
R4800 GND.n1447 GND.n823 105.082
R4801 GND.n1442 GND.n818 105.082
R4802 GND.n1442 GND.n819 105.082
R4803 GND.n1434 GND.n808 105.082
R4804 GND.n1434 GND.n809 105.082
R4805 GND.n1752 GND.n854 105.082
R4806 GND.n1748 GND.n854 105.082
R4807 GND.n1709 GND.n1708 105.082
R4808 GND.n1708 GND.n1707 105.082
R4809 GND.n1715 GND.n1714 105.082
R4810 GND.n1714 GND.n1713 105.082
R4811 GND.n1740 GND.n862 105.082
R4812 GND.n1736 GND.n862 105.082
R4813 GND.n1112 GND.n1111 105.082
R4814 GND.n1111 GND.n1110 105.082
R4815 GND.n1118 GND.n1117 105.082
R4816 GND.n1117 GND.n1116 105.082
R4817 GND.n1139 GND.n1138 105.082
R4818 GND.n1138 GND.n1072 105.082
R4819 GND.n1633 GND.n1632 105.082
R4820 GND.n1632 GND.n1631 105.082
R4821 GND.n1639 GND.n1638 105.082
R4822 GND.n1638 GND.n1637 105.082
R4823 GND.n1664 GND.n912 105.082
R4824 GND.n1660 GND.n912 105.082
R4825 GND.n971 GND.n939 105.082
R4826 GND.n971 GND.n940 105.082
R4827 GND.n976 GND.n943 105.082
R4828 GND.n976 GND.n944 105.082
R4829 GND.n953 GND.n952 105.082
R4830 GND.n986 GND.n953 105.082
R4831 GND.n961 GND.n903 105.082
R4832 GND.n961 GND.n902 105.082
R4833 GND.n956 GND.n899 105.082
R4834 GND.n956 GND.n898 105.082
R4835 GND.n1700 GND.n1699 105.082
R4836 GND.n1701 GND.n1700 105.082
R4837 GND.n1516 GND.n1149 105.082
R4838 GND.n1516 GND.n1150 105.082
R4839 GND.n1521 GND.n1153 105.082
R4840 GND.n1521 GND.n1154 105.082
R4841 GND.n1163 GND.n1162 105.082
R4842 GND.n1531 GND.n1163 105.082
R4843 GND.n1457 GND.n1170 105.082
R4844 GND.n1457 GND.n1171 105.082
R4845 GND.n1462 GND.n1174 105.082
R4846 GND.n1462 GND.n1175 105.082
R4847 GND.n1184 GND.n1183 105.082
R4848 GND.n1472 GND.n1184 105.082
R4849 GND.n1951 GND.n1950 105.082
R4850 GND.n1950 GND.n848 105.082
R4851 GND.n1976 GND.n832 105.082
R4852 GND.n1972 GND.n832 105.082
R4853 GND.n1395 GND.n1385 105.082
R4854 GND.n1391 GND.n1385 105.082
R4855 GND.n1405 GND.n1404 105.082
R4856 GND.n1404 GND.n1379 105.082
R4857 GND.n1429 GND.n1428 105.082
R4858 GND.n1428 GND.n1360 105.082
R4859 GND.n2026 GND.n800 105.082
R4860 GND.n2022 GND.n800 105.082
R4861 GND.n2034 GND.n2033 105.082
R4862 GND.n2033 GND.n789 105.082
R4863 GND.n2059 GND.n701 105.082
R4864 GND.n2055 GND.n701 105.082
R4865 GND.n760 GND.n703 105.082
R4866 GND.n772 GND.n703 105.082
R4867 GND.n756 GND.n710 105.082
R4868 GND.n764 GND.n710 105.082
R4869 GND.n725 GND.n722 105.082
R4870 GND.n730 GND.n722 105.082
R4871 GND.n3322 GND.n415 105.082
R4872 GND.n3322 GND.n416 105.082
R4873 GND.n3231 GND.n3221 105.082
R4874 GND.n3221 GND.n3220 105.082
R4875 GND.n3224 GND.n3217 105.082
R4876 GND.n3224 GND.n3216 105.082
R4877 GND.n3301 GND.n489 105.082
R4878 GND.n3313 GND.n489 105.082
R4879 GND.n3277 GND.n503 105.082
R4880 GND.n3286 GND.n503 105.082
R4881 GND.n3486 GND.n346 105.082
R4882 GND.n3576 GND.n346 105.082
R4883 GND.n3512 GND.n3469 105.082
R4884 GND.n3508 GND.n3469 105.082
R4885 GND.n3550 GND.n353 105.082
R4886 GND.n3550 GND.n354 105.082
R4887 GND.n3546 GND.n360 105.082
R4888 GND.n3452 GND.n360 105.082
R4889 GND.n3456 GND.n366 105.082
R4890 GND.n3456 GND.n367 105.082
R4891 GND.n3449 GND.n377 105.082
R4892 GND.n456 GND.n377 105.082
R4893 GND.n448 GND.n434 105.082
R4894 GND.n448 GND.n433 105.082
R4895 GND.n443 GND.n430 105.082
R4896 GND.n443 GND.n429 105.082
R4897 GND.n3437 GND.n385 105.082
R4898 GND.n3441 GND.n385 105.082
R4899 GND.n3406 GND.n397 105.082
R4900 GND.n3415 GND.n397 105.082
R4901 GND.n3316 GND.n403 105.082
R4902 GND.n3402 GND.n403 105.082
R4903 GND.n3523 GND.n375 105.082
R4904 GND.n3519 GND.n375 105.082
R4905 GND.n3637 GND.n320 105.082
R4906 GND.n3673 GND.n320 105.082
R4907 GND.n3606 GND.n332 105.082
R4908 GND.n3615 GND.n332 105.082
R4909 GND.n3579 GND.n338 105.082
R4910 GND.n3602 GND.n338 105.082
R4911 GND.n3909 GND.n3901 105.082
R4912 GND.n3905 GND.n3901 105.082
R4913 GND.n3932 GND.n3931 105.082
R4914 GND.n3931 GND.n3930 105.082
R4915 GND.n3873 GND.n245 105.082
R4916 GND.n3877 GND.n245 105.082
R4917 GND.n3842 GND.n257 105.082
R4918 GND.n3851 GND.n257 105.082
R4919 GND.n273 GND.n263 105.082
R4920 GND.n3838 GND.n263 105.082
R4921 GND.n3747 GND.n270 105.082
R4922 GND.n3826 GND.n270 105.082
R4923 GND.n3770 GND.n3769 105.082
R4924 GND.n3769 GND.n3768 105.082
R4925 GND.n3776 GND.n3775 105.082
R4926 GND.n3775 GND.n3774 105.082
R4927 GND.n3720 GND.n295 105.082
R4928 GND.n3724 GND.n295 105.082
R4929 GND.n3689 GND.n307 105.082
R4930 GND.n3698 GND.n307 105.082
R4931 GND.n3641 GND.n313 105.082
R4932 GND.n3685 GND.n313 105.082
R4933 GND.n3938 GND.n3937 105.082
R4934 GND.n3937 GND.n3936 105.082
R4935 GND.n4266 GND.n22 105.082
R4936 GND.n4262 GND.n22 105.082
R4937 GND.n4289 GND.n4288 105.082
R4938 GND.n4288 GND.n4287 105.082
R4939 GND.n4295 GND.n4294 105.082
R4940 GND.n4294 GND.n4293 105.082
R4941 GND.n3253 GND.n509 105.082
R4942 GND.n3273 GND.n509 105.082
R4943 GND.n2109 GND.n669 105.082
R4944 GND.n2105 GND.n669 105.082
R4945 GND.n2117 GND.n2116 105.082
R4946 GND.n2116 GND.n658 105.082
R4947 GND.n2138 GND.n644 105.082
R4948 GND.n1226 GND.n1225 105.082
R4949 GND.n3025 GND.n2150 105.082
R4950 GND.n2183 GND.n2150 105.082
R4951 GND.n2190 GND.n2161 105.082
R4952 GND.n2190 GND.n2162 105.082
R4953 GND.n2195 GND.n2165 105.082
R4954 GND.n2195 GND.n2166 105.082
R4955 GND.n2816 GND.n2814 105.082
R4956 GND.n2820 GND.n2814 105.082
R4957 GND.n2854 GND.n2470 105.082
R4958 GND.n2850 GND.n2470 105.082
R4959 GND.n2864 GND.n2863 105.082
R4960 GND.n2863 GND.n2460 105.082
R4961 GND.n2826 GND.n2825 105.082
R4962 GND.n2825 GND.n2802 105.082
R4963 GND.n2789 GND.n2495 105.082
R4964 GND.n2795 GND.n2495 105.082
R4965 GND.n2498 GND.n2497 105.082
R4966 GND.n2785 GND.n2497 105.082
R4967 GND.n1762 GND.n1761 105.082
R4968 GND.n1918 GND.n1917 105.082
R4969 GND.n1917 GND.n1901 105.082
R4970 GND.n4169 GND.n4168 105.082
R4971 GND.n4170 GND.n4169 105.082
R4972 GND.n3160 GND.n554 105.082
R4973 GND.n3164 GND.n554 105.082
R4974 GND.n3129 GND.n566 105.082
R4975 GND.n3138 GND.n566 105.082
R4976 GND.n2517 GND.n572 105.082
R4977 GND.n3125 GND.n572 105.082
R4978 GND.t328 GND.t373 104.74
R4979 GND.n1958 GND.n841 88.201
R4980 GND.n2999 GND.n2998 86.184
R4981 GND.n3006 GND.n3005 86.184
R4982 GND.n3021 GND.n3020 86.184
R4983 GND.n4193 GND.n69 83.1314
R4984 GND.n4222 GND.n48 83.1314
R4985 GND.n2773 GND.n2772 73.9214
R4986 GND.n3050 GND.n633 73.9214
R4987 GND.n1351 GND.n1187 73.1255
R4988 GND.n1351 GND.t721 73.1255
R4989 GND.n1354 GND.n1186 73.1255
R4990 GND.t721 GND.n1186 73.1255
R4991 GND.n936 GND.n935 73.1255
R4992 GND.t641 GND.n936 73.1255
R4993 GND.n1625 GND.n934 73.1255
R4994 GND.t641 GND.n934 73.1255
R4995 GND.n1643 GND.n922 73.1255
R4996 GND.n922 GND.t844 73.1255
R4997 GND.n923 GND.n921 73.1255
R4998 GND.n921 GND.t844 73.1255
R4999 GND.n1673 GND.n905 73.1255
R5000 GND.n905 GND.t386 73.1255
R5001 GND.n906 GND.n904 73.1255
R5002 GND.n904 GND.t386 73.1255
R5003 GND.n1122 GND.n1083 73.1255
R5004 GND.n1083 GND.t451 73.1255
R5005 GND.n1084 GND.n1082 73.1255
R5006 GND.n1082 GND.t451 73.1255
R5007 GND.n1564 GND.n1145 73.1255
R5008 GND.n1145 GND.t406 73.1255
R5009 GND.n1146 GND.n1144 73.1255
R5010 GND.n1144 GND.t406 73.1255
R5011 GND.n1719 GND.n872 73.1255
R5012 GND.n872 GND.t11 73.1255
R5013 GND.n873 GND.n871 73.1255
R5014 GND.n871 GND.t11 73.1255
R5015 GND.n1167 GND.n1166 73.1255
R5016 GND.t751 GND.n1167 73.1255
R5017 GND.n1506 GND.n1165 73.1255
R5018 GND.t751 GND.n1165 73.1255
R5019 GND.n3389 GND.n3353 73.1255
R5020 GND.t618 GND.n3353 73.1255
R5021 GND.n3356 GND.n3354 73.1255
R5022 GND.t618 GND.n3356 73.1255
R5023 GND.n3419 GND.n393 73.1255
R5024 GND.n393 GND.t446 73.1255
R5025 GND.n394 GND.n392 73.1255
R5026 GND.n392 GND.t446 73.1255
R5027 GND.n426 GND.n424 73.1255
R5028 GND.t704 GND.n426 73.1255
R5029 GND.n484 GND.n423 73.1255
R5030 GND.t704 GND.n423 73.1255
R5031 GND.n3531 GND.n369 73.1255
R5032 GND.n369 GND.t30 73.1255
R5033 GND.n370 GND.n368 73.1255
R5034 GND.n368 GND.t30 73.1255
R5035 GND.n3501 GND.n3472 73.1255
R5036 GND.n3472 GND.t840 73.1255
R5037 GND.n3473 GND.n3471 73.1255
R5038 GND.n3471 GND.t840 73.1255
R5039 GND.n3702 GND.n303 73.1255
R5040 GND.n303 GND.t453 73.1255
R5041 GND.n304 GND.n302 73.1255
R5042 GND.n302 GND.t453 73.1255
R5043 GND.n3764 GND.n285 73.1255
R5044 GND.t224 GND.n285 73.1255
R5045 GND.n287 GND.n286 73.1255
R5046 GND.t224 GND.n287 73.1255
R5047 GND.n3855 GND.n253 73.1255
R5048 GND.n253 GND.t18 73.1255
R5049 GND.n254 GND.n252 73.1255
R5050 GND.n252 GND.t18 73.1255
R5051 GND.n3926 GND.n235 73.1255
R5052 GND.t457 GND.n235 73.1255
R5053 GND.n237 GND.n236 73.1255
R5054 GND.t457 GND.n237 73.1255
R5055 GND.n4283 GND.n10 73.1255
R5056 GND.t295 GND.n10 73.1255
R5057 GND.n12 GND.n11 73.1255
R5058 GND.t295 GND.n12 73.1255
R5059 GND.n3290 GND.n499 73.1255
R5060 GND.n499 GND.t459 73.1255
R5061 GND.n500 GND.n498 73.1255
R5062 GND.n498 GND.t459 73.1255
R5063 GND.n3213 GND.n3211 73.1255
R5064 GND.t335 GND.n3213 73.1255
R5065 GND.n3248 GND.n3210 73.1255
R5066 GND.t335 GND.n3210 73.1255
R5067 GND.n520 GND.n518 73.1255
R5068 GND.n518 GND.t355 73.1255
R5069 GND.n524 GND.n519 73.1255
R5070 GND.n519 GND.t355 73.1255
R5071 GND.n1272 GND.n1208 73.1255
R5072 GND.n1272 GND.t612 73.1255
R5073 GND.n1275 GND.n1207 73.1255
R5074 GND.t612 GND.n1207 73.1255
R5075 GND.n2776 GND.n2500 73.1255
R5076 GND.n2500 GND.t435 73.1255
R5077 GND.n2506 GND.n2499 73.1255
R5078 GND.n2499 GND.t435 73.1255
R5079 GND.n2843 GND.n2475 73.1255
R5080 GND.n2475 GND.t331 73.1255
R5081 GND.n2476 GND.n2474 73.1255
R5082 GND.n2474 GND.t331 73.1255
R5083 GND.n2983 GND.n2174 73.1255
R5084 GND.n2174 GND.t739 73.1255
R5085 GND.n2175 GND.n2173 73.1255
R5086 GND.n2173 GND.t739 73.1255
R5087 GND.n2950 GND.n2891 73.1255
R5088 GND.n2891 GND.t657 73.1255
R5089 GND.n2892 GND.n2890 73.1255
R5090 GND.n2890 GND.t657 73.1255
R5091 GND.n2450 GND.n2449 73.1255
R5092 GND.t735 GND.n2450 73.1255
R5093 GND.n2452 GND.n2451 73.1255
R5094 GND.n2451 GND.t735 73.1255
R5095 GND.n2418 GND.n2359 73.1255
R5096 GND.n2359 GND.t620 73.1255
R5097 GND.n2360 GND.n2358 73.1255
R5098 GND.n2358 GND.t620 73.1255
R5099 GND.n2323 GND.n2322 73.1255
R5100 GND.t849 GND.n2323 73.1255
R5101 GND.n2325 GND.n2324 73.1255
R5102 GND.n2324 GND.t849 73.1255
R5103 GND.n2291 GND.n2232 73.1255
R5104 GND.n2232 GND.t594 73.1255
R5105 GND.n2233 GND.n2231 73.1255
R5106 GND.n2231 GND.t594 73.1255
R5107 GND.n2645 GND.n2644 73.1255
R5108 GND.t737 GND.n2645 73.1255
R5109 GND.n2647 GND.n2646 73.1255
R5110 GND.n2646 GND.t737 73.1255
R5111 GND.n2613 GND.n2554 73.1255
R5112 GND.n2554 GND.t249 73.1255
R5113 GND.n2555 GND.n2553 73.1255
R5114 GND.n2553 GND.t249 73.1255
R5115 GND.n2767 GND.n2508 73.1255
R5116 GND.n2508 GND.t697 73.1255
R5117 GND.n2509 GND.n2507 73.1255
R5118 GND.n2507 GND.t697 73.1255
R5119 GND.n2734 GND.n2675 73.1255
R5120 GND.n2675 GND.t3 73.1255
R5121 GND.n2676 GND.n2674 73.1255
R5122 GND.n2674 GND.t3 73.1255
R5123 GND.n2995 GND.n2168 73.1255
R5124 GND.n2168 GND.t741 73.1255
R5125 GND.n2169 GND.n2167 73.1255
R5126 GND.n2167 GND.t741 73.1255
R5127 GND.n2121 GND.n653 73.1255
R5128 GND.n653 GND.t15 73.1255
R5129 GND.n654 GND.n652 73.1255
R5130 GND.n652 GND.t15 73.1255
R5131 GND.n2068 GND.n694 73.1255
R5132 GND.n694 GND.t798 73.1255
R5133 GND.n695 GND.n693 73.1255
R5134 GND.n693 GND.t798 73.1255
R5135 GND.n751 GND.n712 73.1255
R5136 GND.t455 GND.n712 73.1255
R5137 GND.n714 GND.n713 73.1255
R5138 GND.t455 GND.n714 73.1255
R5139 GND.n2038 GND.n784 73.1255
R5140 GND.n784 GND.t259 73.1255
R5141 GND.n785 GND.n783 73.1255
R5142 GND.n783 GND.t259 73.1255
R5143 GND.n1985 GND.n825 73.1255
R5144 GND.n825 GND.t23 73.1255
R5145 GND.n826 GND.n824 73.1255
R5146 GND.n824 GND.t23 73.1255
R5147 GND.n1409 GND.n1372 73.1255
R5148 GND.n1372 GND.t302 73.1255
R5149 GND.n1373 GND.n1371 73.1255
R5150 GND.n1371 GND.t302 73.1255
R5151 GND.n1955 GND.n843 73.1255
R5152 GND.t328 GND.n843 73.1255
R5153 GND.n844 GND.n842 73.1255
R5154 GND.t328 GND.n842 73.1255
R5155 GND.n1589 GND.n1041 73.1255
R5156 GND.n1041 GND.t726 73.1255
R5157 GND.n1042 GND.n1040 73.1255
R5158 GND.n1040 GND.t726 73.1255
R5159 GND.n3116 GND.n578 73.1255
R5160 GND.n578 GND.t851 73.1255
R5161 GND.n579 GND.n577 73.1255
R5162 GND.n577 GND.t851 73.1255
R5163 GND.n3083 GND.n605 73.1255
R5164 GND.n605 GND.t883 73.1255
R5165 GND.n606 GND.n604 73.1255
R5166 GND.n604 GND.t883 73.1255
R5167 GND.n3142 GND.n562 73.1255
R5168 GND.n562 GND.t793 73.1255
R5169 GND.n563 GND.n561 73.1255
R5170 GND.n561 GND.t793 73.1255
R5171 GND.n3186 GND.n542 73.1255
R5172 GND.n542 GND.t655 73.1255
R5173 GND.n550 GND.n541 73.1255
R5174 GND.n541 GND.t655 73.1255
R5175 GND.n3046 GND.n2146 73.1255
R5176 GND.n2146 GND.t644 73.1255
R5177 GND.n2147 GND.n2145 73.1255
R5178 GND.n2145 GND.t644 73.1255
R5179 GND.n4218 GND.n50 73.1255
R5180 GND.n50 GND.t757 73.1255
R5181 GND.n51 GND.n49 73.1255
R5182 GND.n49 GND.t757 73.1255
R5183 GND.n4189 GND.n71 73.1255
R5184 GND.n71 GND.t201 73.1255
R5185 GND.n72 GND.n70 73.1255
R5186 GND.n70 GND.t201 73.1255
R5187 GND.n3593 GND.n344 73.1255
R5188 GND.n344 GND.t83 73.1255
R5189 GND.n3588 GND.n343 73.1255
R5190 GND.n343 GND.t83 73.1255
R5191 GND.n3619 GND.n328 73.1255
R5192 GND.n328 GND.t13 73.1255
R5193 GND.n329 GND.n327 73.1255
R5194 GND.n327 GND.t13 73.1255
R5195 GND.n4134 GND.n120 73.1255
R5196 GND.n120 GND.t664 73.1255
R5197 GND.n121 GND.n119 73.1255
R5198 GND.n119 GND.t664 73.1255
R5199 GND.n4089 GND.n148 73.1255
R5200 GND.n148 GND.t0 73.1255
R5201 GND.n149 GND.n147 73.1255
R5202 GND.n147 GND.t0 73.1255
R5203 GND.n4039 GND.n178 73.1255
R5204 GND.n178 GND.t856 73.1255
R5205 GND.n179 GND.n177 73.1255
R5206 GND.n177 GND.t856 73.1255
R5207 GND.n4149 GND.n110 73.1255
R5208 GND.n110 GND.t215 73.1255
R5209 GND.n111 GND.n109 73.1255
R5210 GND.n109 GND.t215 73.1255
R5211 GND.n4054 GND.n169 73.1255
R5212 GND.n169 GND.t806 73.1255
R5213 GND.n170 GND.n168 73.1255
R5214 GND.n168 GND.t806 73.1255
R5215 GND.n3994 GND.n206 73.1255
R5216 GND.n206 GND.t91 73.1255
R5217 GND.n207 GND.n205 73.1255
R5218 GND.n205 GND.t91 73.1255
R5219 GND.n1909 GND.n841 71.34
R5220 GND.n1904 GND.n1758 71.34
R5221 GND.n1860 GND.t231 69.8913
R5222 GND.n1865 GND.t869 69.8913
R5223 GND.n1870 GND.t101 69.8913
R5224 GND.n1875 GND.t766 69.8913
R5225 GND.n1880 GND.t97 69.8913
R5226 GND.n1885 GND.t186 69.8913
R5227 GND.n1890 GND.t606 69.8913
R5228 GND.n1897 GND.t22 69.8913
R5229 GND.n1933 GND 68.0603
R5230 GND.t513 GND.n104 65.5144
R5231 GND.n1334 GND.n1333 65.0005
R5232 GND.n1335 GND.n1334 65.0005
R5233 GND.n1331 GND.n1330 65.0005
R5234 GND.n1330 GND.n1329 65.0005
R5235 GND.n1341 GND.n1340 65.0005
R5236 GND.n1342 GND.n1341 65.0005
R5237 GND.n1338 GND.n1337 65.0005
R5238 GND.n1337 GND.n1336 65.0005
R5239 GND.n1348 GND.n1347 65.0005
R5240 GND.n1349 GND.n1348 65.0005
R5241 GND.n1345 GND.n1344 65.0005
R5242 GND.n1344 GND.n1343 65.0005
R5243 GND.n1353 GND.n1352 65.0005
R5244 GND.n1352 GND.n805 65.0005
R5245 GND.n1188 GND.n1185 65.0005
R5246 GND.n1350 GND.n1188 65.0005
R5247 GND.n1326 GND.n1325 65.0005
R5248 GND.n1327 GND.n1326 65.0005
R5249 GND.n1323 GND.n1322 65.0005
R5250 GND.n1322 GND.n697 65.0005
R5251 GND.n991 GND.n990 65.0005
R5252 GND.n992 GND.n991 65.0005
R5253 GND.n988 GND.n987 65.0005
R5254 GND.n987 GND.n907 65.0005
R5255 GND.n999 GND.n998 65.0005
R5256 GND.n1000 GND.n999 65.0005
R5257 GND.n996 GND.n995 65.0005
R5258 GND.n995 GND.n994 65.0005
R5259 GND.n1006 GND.n1005 65.0005
R5260 GND.n1007 GND.n1006 65.0005
R5261 GND.n1003 GND.n1002 65.0005
R5262 GND.n1002 GND.n1001 65.0005
R5263 GND.n1013 GND.n1012 65.0005
R5264 GND.n1014 GND.n1013 65.0005
R5265 GND.n1010 GND.n1009 65.0005
R5266 GND.n1009 GND.n1008 65.0005
R5267 GND.n1624 GND.n1623 65.0005
R5268 GND.n1623 GND.n1622 65.0005
R5269 GND.n1015 GND.n933 65.0005
R5270 GND.n1016 GND.n1015 65.0005
R5271 GND.n1659 GND.n1658 65.0005
R5272 GND.n1658 GND.n1657 65.0005
R5273 GND.n1666 GND.n1665 65.0005
R5274 GND.n1667 GND.n1666 65.0005
R5275 GND.n1649 GND.n1648 65.0005
R5276 GND.n1648 GND.n1647 65.0005
R5277 GND.n1655 GND.n1654 65.0005
R5278 GND.n1656 GND.n1655 65.0005
R5279 GND.n1021 GND.n924 65.0005
R5280 GND.n1022 GND.n1021 65.0005
R5281 GND.n1645 GND.n1644 65.0005
R5282 GND.n1646 GND.n1645 65.0005
R5283 GND.n1025 GND.n928 65.0005
R5284 GND.n1026 GND.n1025 65.0005
R5285 GND.n1019 GND.n926 65.0005
R5286 GND.n1023 GND.n1019 65.0005
R5287 GND.n1029 GND.n932 65.0005
R5288 GND.n1030 GND.n1029 65.0005
R5289 GND.n1017 GND.n930 65.0005
R5290 GND.n1027 GND.n1017 65.0005
R5291 GND.n1062 GND.n887 65.0005
R5292 GND.n1065 GND.n1062 65.0005
R5293 GND.n1067 GND.n885 65.0005
R5294 GND.n1068 GND.n1067 65.0005
R5295 GND.n893 GND.n892 65.0005
R5296 GND.n1691 GND.n892 65.0005
R5297 GND.n891 GND.n889 65.0005
R5298 GND.n1064 GND.n891 65.0005
R5299 GND.n1686 GND.n1685 65.0005
R5300 GND.n1685 GND.n1684 65.0005
R5301 GND.n1689 GND.n1688 65.0005
R5302 GND.n1690 GND.n1689 65.0005
R5303 GND.n1679 GND.n1678 65.0005
R5304 GND.n1678 GND.n1677 65.0005
R5305 GND.n1682 GND.n1681 65.0005
R5306 GND.n1683 GND.n1682 65.0005
R5307 GND.n1672 GND.n1671 65.0005
R5308 GND.n1671 GND.n1670 65.0005
R5309 GND.n1675 GND.n1674 65.0005
R5310 GND.n1676 GND.n1675 65.0005
R5311 GND.n1079 GND.n1078 65.0005
R5312 GND.n1080 GND.n1079 65.0005
R5313 GND.n1141 GND.n1140 65.0005
R5314 GND.n1142 GND.n1141 65.0005
R5315 GND.n1127 GND.n1077 65.0005
R5316 GND.n1126 GND.n1077 65.0005
R5317 GND.n1076 GND.n1074 65.0005
R5318 GND.n1081 GND.n1076 65.0005
R5319 GND.n1096 GND.n1085 65.0005
R5320 GND.n1097 GND.n1096 65.0005
R5321 GND.n1124 GND.n1123 65.0005
R5322 GND.n1125 GND.n1124 65.0005
R5323 GND.n1102 GND.n1090 65.0005
R5324 GND.n1103 GND.n1102 65.0005
R5325 GND.n1099 GND.n1088 65.0005
R5326 GND.n1099 GND.n1098 65.0005
R5327 GND.n1107 GND.n1106 65.0005
R5328 GND.n1106 GND.n908 65.0005
R5329 GND.n1095 GND.n1092 65.0005
R5330 GND.n1104 GND.n1095 65.0005
R5331 GND.n1537 GND.n1536 65.0005
R5332 GND.n1538 GND.n1537 65.0005
R5333 GND.n1534 GND.n1533 65.0005
R5334 GND.n1533 GND.n1532 65.0005
R5335 GND.n1545 GND.n1544 65.0005
R5336 GND.n1546 GND.n1545 65.0005
R5337 GND.n1542 GND.n1541 65.0005
R5338 GND.n1541 GND.n1540 65.0005
R5339 GND.n1552 GND.n1551 65.0005
R5340 GND.n1553 GND.n1552 65.0005
R5341 GND.n1549 GND.n1548 65.0005
R5342 GND.n1548 GND.n1547 65.0005
R5343 GND.n1559 GND.n1558 65.0005
R5344 GND.n1560 GND.n1559 65.0005
R5345 GND.n1556 GND.n1555 65.0005
R5346 GND.n1555 GND.n1554 65.0005
R5347 GND.n1566 GND.n1565 65.0005
R5348 GND.n1567 GND.n1566 65.0005
R5349 GND.n1563 GND.n1562 65.0005
R5350 GND.n1562 GND.n1561 65.0005
R5351 GND.n1735 GND.n1734 65.0005
R5352 GND.n1734 GND.n1733 65.0005
R5353 GND.n1742 GND.n1741 65.0005
R5354 GND.n1743 GND.n1742 65.0005
R5355 GND.n1725 GND.n1724 65.0005
R5356 GND.n1724 GND.n1723 65.0005
R5357 GND.n1731 GND.n1730 65.0005
R5358 GND.n1732 GND.n1731 65.0005
R5359 GND.n1056 GND.n874 65.0005
R5360 GND.n1057 GND.n1056 65.0005
R5361 GND.n1721 GND.n1720 65.0005
R5362 GND.n1722 GND.n1721 65.0005
R5363 GND.n1574 GND.n878 65.0005
R5364 GND.n1574 GND.n1573 65.0005
R5365 GND.n1059 GND.n876 65.0005
R5366 GND.n1059 GND.n1058 65.0005
R5367 GND.n1060 GND.n882 65.0005
R5368 GND.n1569 GND.n1060 65.0005
R5369 GND.n1571 GND.n880 65.0005
R5370 GND.n1572 GND.n1571 65.0005
R5371 GND.n1477 GND.n1476 65.0005
R5372 GND.n1478 GND.n1477 65.0005
R5373 GND.n1474 GND.n1473 65.0005
R5374 GND.n1473 GND.n828 65.0005
R5375 GND.n1485 GND.n1484 65.0005
R5376 GND.n1486 GND.n1485 65.0005
R5377 GND.n1482 GND.n1481 65.0005
R5378 GND.n1481 GND.n1480 65.0005
R5379 GND.n1492 GND.n1491 65.0005
R5380 GND.n1493 GND.n1492 65.0005
R5381 GND.n1489 GND.n1488 65.0005
R5382 GND.n1488 GND.n1487 65.0005
R5383 GND.n1499 GND.n1498 65.0005
R5384 GND.n1500 GND.n1499 65.0005
R5385 GND.n1496 GND.n1495 65.0005
R5386 GND.n1495 GND.n1494 65.0005
R5387 GND.n1505 GND.n1504 65.0005
R5388 GND.n1504 GND.n1503 65.0005
R5389 GND.n1501 GND.n1164 65.0005
R5390 GND.n1502 GND.n1501 65.0005
R5391 GND.n1747 GND.n1746 65.0005
R5392 GND.n1746 GND.n1745 65.0005
R5393 GND.n1754 GND.n1753 65.0005
R5394 GND.n1755 GND.n1754 65.0005
R5395 GND.n1946 GND.n850 65.0005
R5396 GND.n1756 GND.n850 65.0005
R5397 GND.n3388 GND.n3387 65.0005
R5398 GND.n3387 GND.n3386 65.0005
R5399 GND.n3355 GND.n3352 65.0005
R5400 GND.n3355 GND.n381 65.0005
R5401 GND.n3378 GND.n3377 65.0005
R5402 GND.n3377 GND.n371 65.0005
R5403 GND.n3384 GND.n3383 65.0005
R5404 GND.n3385 GND.n3384 65.0005
R5405 GND.n3401 GND.n3400 65.0005
R5406 GND.n3400 GND.n401 65.0005
R5407 GND.n3315 GND.n406 65.0005
R5408 GND.n3398 GND.n406 65.0005
R5409 GND.n3414 GND.n3413 65.0005
R5410 GND.n3413 GND.n3412 65.0005
R5411 GND.n3408 GND.n3407 65.0005
R5412 GND.n3409 GND.n3408 65.0005
R5413 GND.n3421 GND.n3420 65.0005
R5414 GND.n3422 GND.n3421 65.0005
R5415 GND.n3410 GND.n395 65.0005
R5416 GND.n3411 GND.n3410 65.0005
R5417 GND.n3432 GND.n3431 65.0005
R5418 GND.n3433 GND.n3432 65.0005
R5419 GND.n3426 GND.n3425 65.0005
R5420 GND.n3425 GND.n3424 65.0005
R5421 GND.n3443 GND.n3442 65.0005
R5422 GND.n3444 GND.n3443 65.0005
R5423 GND.n3436 GND.n3435 65.0005
R5424 GND.n3435 GND.n3434 65.0005
R5425 GND.n483 GND.n482 65.0005
R5426 GND.n482 GND.n481 65.0005
R5427 GND.n425 GND.n422 65.0005
R5428 GND.n425 GND.n407 65.0005
R5429 GND.n476 GND.n475 65.0005
R5430 GND.n475 GND.n474 65.0005
R5431 GND.n479 GND.n478 65.0005
R5432 GND.n480 GND.n479 65.0005
R5433 GND.n469 GND.n468 65.0005
R5434 GND.n468 GND.n467 65.0005
R5435 GND.n472 GND.n471 65.0005
R5436 GND.n473 GND.n472 65.0005
R5437 GND.n462 GND.n461 65.0005
R5438 GND.n461 GND.n460 65.0005
R5439 GND.n465 GND.n464 65.0005
R5440 GND.n466 GND.n465 65.0005
R5441 GND.n3448 GND.n3447 65.0005
R5442 GND.n3447 GND.n3446 65.0005
R5443 GND.n458 GND.n457 65.0005
R5444 GND.n459 GND.n458 65.0005
R5445 GND.n3395 GND.n3394 65.0005
R5446 GND.n3396 GND.n3395 65.0005
R5447 GND.n3348 GND.n3347 65.0005
R5448 GND.n3347 GND.n3346 65.0005
R5449 GND.n3368 GND.n3367 65.0005
R5450 GND.n3367 GND.n342 65.0005
R5451 GND.n3366 GND.n3364 65.0005
R5452 GND.n3366 GND.n350 65.0005
R5453 GND.n3533 GND.n3532 65.0005
R5454 GND.n3534 GND.n3533 65.0005
R5455 GND.n3530 GND.n3529 65.0005
R5456 GND.n3529 GND.n3528 65.0005
R5457 GND.n3540 GND.n3539 65.0005
R5458 GND.n3541 GND.n3540 65.0005
R5459 GND.n3537 GND.n3536 65.0005
R5460 GND.n3536 GND.n3535 65.0005
R5461 GND.n3545 GND.n3544 65.0005
R5462 GND.n3544 GND.n69 65.0005
R5463 GND.n3451 GND.n363 65.0005
R5464 GND.n3542 GND.n363 65.0005
R5465 GND.n3563 GND.n3562 65.0005
R5466 GND.n3564 GND.n3563 65.0005
R5467 GND.n3560 GND.n3559 65.0005
R5468 GND.n3559 GND.n3558 65.0005
R5469 GND.n3570 GND.n3569 65.0005
R5470 GND.n3571 GND.n3570 65.0005
R5471 GND.n3567 GND.n3566 65.0005
R5472 GND.n3566 GND.n3565 65.0005
R5473 GND.n3507 GND.n3506 65.0005
R5474 GND.n3506 GND.n3505 65.0005
R5475 GND.n3514 GND.n3513 65.0005
R5476 GND.n3515 GND.n3514 65.0005
R5477 GND.n3481 GND.n3474 65.0005
R5478 GND.n3482 GND.n3481 65.0005
R5479 GND.n3503 GND.n3502 65.0005
R5480 GND.n3504 GND.n3503 65.0005
R5481 GND.n3491 GND.n3480 65.0005
R5482 GND.n3490 GND.n3480 65.0005
R5483 GND.n3479 GND.n3477 65.0005
R5484 GND.n3483 GND.n3479 65.0005
R5485 GND.n3575 GND.n3574 65.0005
R5486 GND.n3574 GND.n3573 65.0005
R5487 GND.n3488 GND.n3487 65.0005
R5488 GND.n3489 GND.n3488 65.0005
R5489 GND.n3518 GND.n3517 65.0005
R5490 GND.n3517 GND.n3516 65.0005
R5491 GND.n3525 GND.n3524 65.0005
R5492 GND.n3526 GND.n3525 65.0005
R5493 GND.n3684 GND.n3683 65.0005
R5494 GND.n3683 GND.n311 65.0005
R5495 GND.n3640 GND.n316 65.0005
R5496 GND.n3681 GND.n316 65.0005
R5497 GND.n3697 GND.n3696 65.0005
R5498 GND.n3696 GND.n3695 65.0005
R5499 GND.n3691 GND.n3690 65.0005
R5500 GND.n3692 GND.n3691 65.0005
R5501 GND.n3704 GND.n3703 65.0005
R5502 GND.n3705 GND.n3704 65.0005
R5503 GND.n3693 GND.n305 65.0005
R5504 GND.n3694 GND.n3693 65.0005
R5505 GND.n3715 GND.n3714 65.0005
R5506 GND.n3716 GND.n3715 65.0005
R5507 GND.n3709 GND.n3708 65.0005
R5508 GND.n3708 GND.n3707 65.0005
R5509 GND.n3726 GND.n3725 65.0005
R5510 GND.n3727 GND.n3726 65.0005
R5511 GND.n3719 GND.n3718 65.0005
R5512 GND.n3718 GND.n3717 65.0005
R5513 GND.n3731 GND.n279 65.0005
R5514 GND.n3732 GND.n3731 65.0005
R5515 GND.n290 GND.n277 65.0005
R5516 GND.n3729 GND.n290 65.0005
R5517 GND.n3735 GND.n283 65.0005
R5518 GND.n3736 GND.n3735 65.0005
R5519 GND.n288 GND.n281 65.0005
R5520 GND.n3733 GND.n288 65.0005
R5521 GND.n3763 GND.n3762 65.0005
R5522 GND.n3762 GND.n3761 65.0005
R5523 GND.n3737 GND.n284 65.0005
R5524 GND.n3738 GND.n3737 65.0005
R5525 GND.n3753 GND.n3752 65.0005
R5526 GND.n3752 GND.n3751 65.0005
R5527 GND.n3759 GND.n3758 65.0005
R5528 GND.n3760 GND.n3759 65.0005
R5529 GND.n3828 GND.n3827 65.0005
R5530 GND.n3829 GND.n3828 65.0005
R5531 GND.n3749 GND.n3748 65.0005
R5532 GND.n3750 GND.n3749 65.0005
R5533 GND.n3837 GND.n3836 65.0005
R5534 GND.n3836 GND.n261 65.0005
R5535 GND.n272 GND.n266 65.0005
R5536 GND.n3834 GND.n266 65.0005
R5537 GND.n3850 GND.n3849 65.0005
R5538 GND.n3849 GND.n3848 65.0005
R5539 GND.n3844 GND.n3843 65.0005
R5540 GND.n3845 GND.n3844 65.0005
R5541 GND.n3857 GND.n3856 65.0005
R5542 GND.n3858 GND.n3857 65.0005
R5543 GND.n3846 GND.n255 65.0005
R5544 GND.n3847 GND.n3846 65.0005
R5545 GND.n3868 GND.n3867 65.0005
R5546 GND.n3869 GND.n3868 65.0005
R5547 GND.n3862 GND.n3861 65.0005
R5548 GND.n3861 GND.n3860 65.0005
R5549 GND.n3879 GND.n3878 65.0005
R5550 GND.n3880 GND.n3879 65.0005
R5551 GND.n3872 GND.n3871 65.0005
R5552 GND.n3871 GND.n3870 65.0005
R5553 GND.n3888 GND.n233 65.0005
R5554 GND.n3889 GND.n3888 65.0005
R5555 GND.n238 GND.n231 65.0005
R5556 GND.n3886 GND.n238 65.0005
R5557 GND.n3925 GND.n3924 65.0005
R5558 GND.n3924 GND.n3923 65.0005
R5559 GND.n3890 GND.n234 65.0005
R5560 GND.n3891 GND.n3890 65.0005
R5561 GND.n3915 GND.n3914 65.0005
R5562 GND.n3914 GND.n3913 65.0005
R5563 GND.n3921 GND.n3920 65.0005
R5564 GND.n3922 GND.n3921 65.0005
R5565 GND.n3904 GND.n3903 65.0005
R5566 GND.n3911 GND.n3910 65.0005
R5567 GND.n3912 GND.n3911 65.0005
R5568 GND.n3884 GND.n229 65.0005
R5569 GND.n3885 GND.n3884 65.0005
R5570 GND.n240 GND.n227 65.0005
R5571 GND.n3882 GND.n240 65.0005
R5572 GND.n3170 GND.n8 65.0005
R5573 GND.n3174 GND.n3170 65.0005
R5574 GND.n3176 GND.n6 65.0005
R5575 GND.n3177 GND.n3176 65.0005
R5576 GND.n4282 GND.n4281 65.0005
R5577 GND.n4281 GND.n4280 65.0005
R5578 GND.n3172 GND.n9 65.0005
R5579 GND.n3173 GND.n3172 65.0005
R5580 GND.n4272 GND.n4271 65.0005
R5581 GND.n4271 GND.n4270 65.0005
R5582 GND.n4278 GND.n4277 65.0005
R5583 GND.n4279 GND.n4278 65.0005
R5584 GND.n4261 GND.n4260 65.0005
R5585 GND.n4260 GND.n4259 65.0005
R5586 GND.n4268 GND.n4267 65.0005
R5587 GND.n4269 GND.n4268 65.0005
R5588 GND.n3168 GND.n4 65.0005
R5589 GND.n3178 GND.n3168 65.0005
R5590 GND.n3180 GND.n2 65.0005
R5591 GND.n3181 GND.n3180 65.0005
R5592 GND.n3272 GND.n3271 65.0005
R5593 GND.n3271 GND.n507 65.0005
R5594 GND.n3252 GND.n512 65.0005
R5595 GND.n3269 GND.n512 65.0005
R5596 GND.n3285 GND.n3284 65.0005
R5597 GND.n3284 GND.n3283 65.0005
R5598 GND.n3279 GND.n3278 65.0005
R5599 GND.n3280 GND.n3279 65.0005
R5600 GND.n3292 GND.n3291 65.0005
R5601 GND.n3293 GND.n3292 65.0005
R5602 GND.n3281 GND.n501 65.0005
R5603 GND.n3282 GND.n3281 65.0005
R5604 GND.n3307 GND.n3306 65.0005
R5605 GND.n3308 GND.n3307 65.0005
R5606 GND.n3297 GND.n3296 65.0005
R5607 GND.n3296 GND.n3295 65.0005
R5608 GND.n3312 GND.n3311 65.0005
R5609 GND.n3311 GND.n412 65.0005
R5610 GND.n3300 GND.n492 65.0005
R5611 GND.n3309 GND.n492 65.0005
R5612 GND.n3247 GND.n3246 65.0005
R5613 GND.n3246 GND.n3245 65.0005
R5614 GND.n3212 GND.n3209 65.0005
R5615 GND.n3212 GND.n513 65.0005
R5616 GND.n3240 GND.n3239 65.0005
R5617 GND.n3239 GND.n3238 65.0005
R5618 GND.n3243 GND.n3242 65.0005
R5619 GND.n3244 GND.n3243 65.0005
R5620 GND.n3233 GND.n3232 65.0005
R5621 GND.n3232 GND.n48 65.0005
R5622 GND.n3236 GND.n3235 65.0005
R5623 GND.n3237 GND.n3236 65.0005
R5624 GND.n3335 GND.n3334 65.0005
R5625 GND.n3336 GND.n3335 65.0005
R5626 GND.n3332 GND.n3331 65.0005
R5627 GND.n3331 GND.n3330 65.0005
R5628 GND.n3342 GND.n3341 65.0005
R5629 GND.n3343 GND.n3342 65.0005
R5630 GND.n3339 GND.n3338 65.0005
R5631 GND.n3338 GND.n3337 65.0005
R5632 GND.n3266 GND.n3265 65.0005
R5633 GND.n3267 GND.n3266 65.0005
R5634 GND.n531 GND.n530 65.0005
R5635 GND.n530 GND.n529 65.0005
R5636 GND.n526 GND.n525 65.0005
R5637 GND.n527 GND.n526 65.0005
R5638 GND.n522 GND.n521 65.0005
R5639 GND.n521 GND.n24 65.0005
R5640 GND.n1247 GND.n1246 65.0005
R5641 GND.n1248 GND.n1247 65.0005
R5642 GND.n1244 GND.n1243 65.0005
R5643 GND.n1243 GND.n640 65.0005
R5644 GND.n1255 GND.n1254 65.0005
R5645 GND.n1256 GND.n1255 65.0005
R5646 GND.n1252 GND.n1251 65.0005
R5647 GND.n1251 GND.n1250 65.0005
R5648 GND.n1262 GND.n1261 65.0005
R5649 GND.n1263 GND.n1262 65.0005
R5650 GND.n1259 GND.n1258 65.0005
R5651 GND.n1258 GND.n1257 65.0005
R5652 GND.n1269 GND.n1268 65.0005
R5653 GND.n1270 GND.n1269 65.0005
R5654 GND.n1266 GND.n1265 65.0005
R5655 GND.n1265 GND.n1264 65.0005
R5656 GND.n1274 GND.n1273 65.0005
R5657 GND.n1273 GND.n674 65.0005
R5658 GND.n1209 GND.n1206 65.0005
R5659 GND.n1271 GND.n1209 65.0005
R5660 GND.n2778 GND.n2777 65.0005
R5661 GND.n2779 GND.n2778 65.0005
R5662 GND.n2775 GND.n2774 65.0005
R5663 GND.n2774 GND.n2773 65.0005
R5664 GND.n2784 GND.n2465 65.0005
R5665 GND.n2858 GND.n2465 65.0005
R5666 GND.n2782 GND.n2781 65.0005
R5667 GND.n2781 GND.n2780 65.0005
R5668 GND.n2794 GND.n2473 65.0005
R5669 GND.n2847 GND.n2473 65.0005
R5670 GND.n2790 GND.n2466 65.0005
R5671 GND.n2857 GND.n2466 65.0005
R5672 GND.n2493 GND.n2489 65.0005
R5673 GND.n2809 GND.n2489 65.0005
R5674 GND.n2491 GND.n2488 65.0005
R5675 GND.n2488 GND.n2487 65.0005
R5676 GND.n2805 GND.n2804 65.0005
R5677 GND.n2804 GND.n633 65.0005
R5678 GND.n2803 GND.n2800 65.0005
R5679 GND.n2810 GND.n2803 65.0005
R5680 GND.n2859 GND.n2462 65.0005
R5681 GND.n2858 GND.n2462 65.0005
R5682 GND.n2461 GND.n2459 65.0005
R5683 GND.n2780 GND.n2461 65.0005
R5684 GND.n2849 GND.n2848 65.0005
R5685 GND.n2848 GND.n2847 65.0005
R5686 GND.n2856 GND.n2855 65.0005
R5687 GND.n2857 GND.n2856 65.0005
R5688 GND.n2485 GND.n2477 65.0005
R5689 GND.n2486 GND.n2485 65.0005
R5690 GND.n2845 GND.n2844 65.0005
R5691 GND.n2846 GND.n2845 65.0005
R5692 GND.n2833 GND.n2483 65.0005
R5693 GND.n2809 GND.n2483 65.0005
R5694 GND.n2482 GND.n2480 65.0005
R5695 GND.n2487 GND.n2482 65.0005
R5696 GND.n2821 GND.n2812 65.0005
R5697 GND.n2812 GND.n633 65.0005
R5698 GND.n2813 GND.n2811 65.0005
R5699 GND.n2811 GND.n2810 65.0005
R5700 GND.n2982 GND.n2981 65.0005
R5701 GND.n2981 GND.n2980 65.0005
R5702 GND.n2985 GND.n2984 65.0005
R5703 GND.n2986 GND.n2985 65.0005
R5704 GND.n2877 GND.n2873 65.0005
R5705 GND.n2967 GND.n2877 65.0005
R5706 GND.n2180 GND.n2176 65.0005
R5707 GND.n2979 GND.n2176 65.0005
R5708 GND.n2889 GND.n2885 65.0005
R5709 GND.n2954 GND.n2889 65.0005
R5710 GND.n2882 GND.n2878 65.0005
R5711 GND.n2966 GND.n2878 65.0005
R5712 GND.n2936 GND.n2900 65.0005
R5713 GND.n2931 GND.n2900 65.0005
R5714 GND.n2934 GND.n2899 65.0005
R5715 GND.n2905 GND.n2899 65.0005
R5716 GND.n2918 GND.n2917 65.0005
R5717 GND.n2917 GND.n634 65.0005
R5718 GND.n2911 GND.n2907 65.0005
R5719 GND.n2930 GND.n2907 65.0005
R5720 GND.n2969 GND.n2968 65.0005
R5721 GND.n2968 GND.n2967 65.0005
R5722 GND.n2978 GND.n2977 65.0005
R5723 GND.n2979 GND.n2978 65.0005
R5724 GND.n2956 GND.n2955 65.0005
R5725 GND.n2955 GND.n2954 65.0005
R5726 GND.n2965 GND.n2964 65.0005
R5727 GND.n2966 GND.n2965 65.0005
R5728 GND.n2903 GND.n2893 65.0005
R5729 GND.n2904 GND.n2903 65.0005
R5730 GND.n2952 GND.n2951 65.0005
R5731 GND.n2953 GND.n2952 65.0005
R5732 GND.n2939 GND.n2932 65.0005
R5733 GND.n2932 GND.n2931 65.0005
R5734 GND.n2933 GND.n2906 65.0005
R5735 GND.n2906 GND.n2905 65.0005
R5736 GND.n2920 GND.n2919 65.0005
R5737 GND.n2919 GND.n634 65.0005
R5738 GND.n2929 GND.n2928 65.0005
R5739 GND.n2930 GND.n2929 65.0005
R5740 GND.n2333 GND.n2331 65.0005
R5741 GND.n2448 GND.n2333 65.0005
R5742 GND.n2332 GND.n2330 65.0005
R5743 GND.n2332 GND.n2172 65.0005
R5744 GND.n2345 GND.n2341 65.0005
R5745 GND.n2435 GND.n2345 65.0005
R5746 GND.n2338 GND.n2334 65.0005
R5747 GND.n2447 GND.n2334 65.0005
R5748 GND.n2357 GND.n2353 65.0005
R5749 GND.n2422 GND.n2357 65.0005
R5750 GND.n2350 GND.n2346 65.0005
R5751 GND.n2434 GND.n2346 65.0005
R5752 GND.n2404 GND.n2368 65.0005
R5753 GND.n2399 GND.n2368 65.0005
R5754 GND.n2402 GND.n2367 65.0005
R5755 GND.n2373 GND.n2367 65.0005
R5756 GND.n2386 GND.n2385 65.0005
R5757 GND.n2385 GND.n635 65.0005
R5758 GND.n2379 GND.n2375 65.0005
R5759 GND.n2398 GND.n2375 65.0005
R5760 GND.n2437 GND.n2436 65.0005
R5761 GND.n2436 GND.n2435 65.0005
R5762 GND.n2446 GND.n2445 65.0005
R5763 GND.n2447 GND.n2446 65.0005
R5764 GND.n2424 GND.n2423 65.0005
R5765 GND.n2423 GND.n2422 65.0005
R5766 GND.n2433 GND.n2432 65.0005
R5767 GND.n2434 GND.n2433 65.0005
R5768 GND.n2371 GND.n2361 65.0005
R5769 GND.n2372 GND.n2371 65.0005
R5770 GND.n2420 GND.n2419 65.0005
R5771 GND.n2421 GND.n2420 65.0005
R5772 GND.n2407 GND.n2400 65.0005
R5773 GND.n2400 GND.n2399 65.0005
R5774 GND.n2401 GND.n2374 65.0005
R5775 GND.n2374 GND.n2373 65.0005
R5776 GND.n2388 GND.n2387 65.0005
R5777 GND.n2387 GND.n635 65.0005
R5778 GND.n2397 GND.n2396 65.0005
R5779 GND.n2398 GND.n2397 65.0005
R5780 GND.n2205 GND.n2203 65.0005
R5781 GND.n2321 GND.n2205 65.0005
R5782 GND.n2204 GND.n2202 65.0005
R5783 GND.n2206 GND.n2204 65.0005
R5784 GND.n2218 GND.n2214 65.0005
R5785 GND.n2308 GND.n2218 65.0005
R5786 GND.n2211 GND.n2207 65.0005
R5787 GND.n2320 GND.n2207 65.0005
R5788 GND.n2230 GND.n2226 65.0005
R5789 GND.n2295 GND.n2230 65.0005
R5790 GND.n2223 GND.n2219 65.0005
R5791 GND.n2307 GND.n2219 65.0005
R5792 GND.n2277 GND.n2241 65.0005
R5793 GND.n2272 GND.n2241 65.0005
R5794 GND.n2275 GND.n2240 65.0005
R5795 GND.n2246 GND.n2240 65.0005
R5796 GND.n2259 GND.n2258 65.0005
R5797 GND.n2258 GND.n636 65.0005
R5798 GND.n2252 GND.n2248 65.0005
R5799 GND.n2271 GND.n2248 65.0005
R5800 GND.n2310 GND.n2309 65.0005
R5801 GND.n2309 GND.n2308 65.0005
R5802 GND.n2319 GND.n2318 65.0005
R5803 GND.n2320 GND.n2319 65.0005
R5804 GND.n2297 GND.n2296 65.0005
R5805 GND.n2296 GND.n2295 65.0005
R5806 GND.n2306 GND.n2305 65.0005
R5807 GND.n2307 GND.n2306 65.0005
R5808 GND.n2244 GND.n2234 65.0005
R5809 GND.n2245 GND.n2244 65.0005
R5810 GND.n2293 GND.n2292 65.0005
R5811 GND.n2294 GND.n2293 65.0005
R5812 GND.n2280 GND.n2273 65.0005
R5813 GND.n2273 GND.n2272 65.0005
R5814 GND.n2274 GND.n2247 65.0005
R5815 GND.n2247 GND.n2246 65.0005
R5816 GND.n2261 GND.n2260 65.0005
R5817 GND.n2260 GND.n636 65.0005
R5818 GND.n2270 GND.n2269 65.0005
R5819 GND.n2271 GND.n2270 65.0005
R5820 GND.n2527 GND.n2525 65.0005
R5821 GND.n2643 GND.n2527 65.0005
R5822 GND.n2526 GND.n2524 65.0005
R5823 GND.n2528 GND.n2526 65.0005
R5824 GND.n2540 GND.n2536 65.0005
R5825 GND.n2630 GND.n2540 65.0005
R5826 GND.n2533 GND.n2529 65.0005
R5827 GND.n2642 GND.n2529 65.0005
R5828 GND.n2552 GND.n2548 65.0005
R5829 GND.n2617 GND.n2552 65.0005
R5830 GND.n2545 GND.n2541 65.0005
R5831 GND.n2629 GND.n2541 65.0005
R5832 GND.n2599 GND.n2563 65.0005
R5833 GND.n2594 GND.n2563 65.0005
R5834 GND.n2597 GND.n2562 65.0005
R5835 GND.n2568 GND.n2562 65.0005
R5836 GND.n2581 GND.n2580 65.0005
R5837 GND.n2580 GND.n637 65.0005
R5838 GND.n2574 GND.n2570 65.0005
R5839 GND.n2593 GND.n2570 65.0005
R5840 GND.n2632 GND.n2631 65.0005
R5841 GND.n2631 GND.n2630 65.0005
R5842 GND.n2641 GND.n2640 65.0005
R5843 GND.n2642 GND.n2641 65.0005
R5844 GND.n2619 GND.n2618 65.0005
R5845 GND.n2618 GND.n2617 65.0005
R5846 GND.n2628 GND.n2627 65.0005
R5847 GND.n2629 GND.n2628 65.0005
R5848 GND.n2566 GND.n2556 65.0005
R5849 GND.n2567 GND.n2566 65.0005
R5850 GND.n2615 GND.n2614 65.0005
R5851 GND.n2616 GND.n2615 65.0005
R5852 GND.n2602 GND.n2595 65.0005
R5853 GND.n2595 GND.n2594 65.0005
R5854 GND.n2596 GND.n2569 65.0005
R5855 GND.n2569 GND.n2568 65.0005
R5856 GND.n2583 GND.n2582 65.0005
R5857 GND.n2582 GND.n637 65.0005
R5858 GND.n2592 GND.n2591 65.0005
R5859 GND.n2593 GND.n2592 65.0005
R5860 GND.n2766 GND.n2765 65.0005
R5861 GND.n2765 GND.n2764 65.0005
R5862 GND.n2769 GND.n2768 65.0005
R5863 GND.n2770 GND.n2769 65.0005
R5864 GND.n2661 GND.n2657 65.0005
R5865 GND.n2751 GND.n2661 65.0005
R5866 GND.n2514 GND.n2510 65.0005
R5867 GND.n2763 GND.n2510 65.0005
R5868 GND.n2673 GND.n2669 65.0005
R5869 GND.n2738 GND.n2673 65.0005
R5870 GND.n2666 GND.n2662 65.0005
R5871 GND.n2750 GND.n2662 65.0005
R5872 GND.n2720 GND.n2684 65.0005
R5873 GND.n2715 GND.n2684 65.0005
R5874 GND.n2718 GND.n2683 65.0005
R5875 GND.n2689 GND.n2683 65.0005
R5876 GND.n2702 GND.n2701 65.0005
R5877 GND.n2701 GND.n638 65.0005
R5878 GND.n2695 GND.n2691 65.0005
R5879 GND.n2714 GND.n2691 65.0005
R5880 GND.n2753 GND.n2752 65.0005
R5881 GND.n2752 GND.n2751 65.0005
R5882 GND.n2762 GND.n2761 65.0005
R5883 GND.n2763 GND.n2762 65.0005
R5884 GND.n2740 GND.n2739 65.0005
R5885 GND.n2739 GND.n2738 65.0005
R5886 GND.n2749 GND.n2748 65.0005
R5887 GND.n2750 GND.n2749 65.0005
R5888 GND.n2687 GND.n2677 65.0005
R5889 GND.n2688 GND.n2687 65.0005
R5890 GND.n2736 GND.n2735 65.0005
R5891 GND.n2737 GND.n2736 65.0005
R5892 GND.n2723 GND.n2716 65.0005
R5893 GND.n2716 GND.n2715 65.0005
R5894 GND.n2717 GND.n2690 65.0005
R5895 GND.n2690 GND.n2689 65.0005
R5896 GND.n2704 GND.n2703 65.0005
R5897 GND.n2703 GND.n638 65.0005
R5898 GND.n2713 GND.n2712 65.0005
R5899 GND.n2714 GND.n2713 65.0005
R5900 GND.n2997 GND.n2996 65.0005
R5901 GND.n2998 GND.n2997 65.0005
R5902 GND.n2994 GND.n2993 65.0005
R5903 GND.n2993 GND.n2992 65.0005
R5904 GND.n3004 GND.n3003 65.0005
R5905 GND.n3005 GND.n3004 65.0005
R5906 GND.n3001 GND.n3000 65.0005
R5907 GND.n3000 GND.n2999 65.0005
R5908 GND.n3011 GND.n3010 65.0005
R5909 GND.n3012 GND.n3011 65.0005
R5910 GND.n3008 GND.n3007 65.0005
R5911 GND.n3007 GND.n3006 65.0005
R5912 GND.n3019 GND.n3018 65.0005
R5913 GND.n3020 GND.n3019 65.0005
R5914 GND.n3016 GND.n3015 65.0005
R5915 GND.n3015 GND.n3014 65.0005
R5916 GND.n3024 GND.n3023 65.0005
R5917 GND.n3023 GND.n639 65.0005
R5918 GND.n2182 GND.n2153 65.0005
R5919 GND.n3021 GND.n2153 65.0005
R5920 GND.n2137 GND.n2136 65.0005
R5921 GND.n2136 GND.n2135 65.0005
R5922 GND.n2142 GND.n2141 65.0005
R5923 GND.n2143 GND.n2142 65.0005
R5924 GND.n2127 GND.n2126 65.0005
R5925 GND.n2126 GND.n2125 65.0005
R5926 GND.n2133 GND.n2132 65.0005
R5927 GND.n2134 GND.n2133 65.0005
R5928 GND.n659 GND.n655 65.0005
R5929 GND.n660 GND.n659 65.0005
R5930 GND.n2123 GND.n2122 65.0005
R5931 GND.n2124 GND.n2123 65.0005
R5932 GND.n2114 GND.n665 65.0005
R5933 GND.n2114 GND.n2113 65.0005
R5934 GND.n662 GND.n657 65.0005
R5935 GND.n662 GND.n661 65.0005
R5936 GND.n2104 GND.n2103 65.0005
R5937 GND.n2103 GND.n2102 65.0005
R5938 GND.n2111 GND.n2110 65.0005
R5939 GND.n2112 GND.n2111 65.0005
R5940 GND.n2095 GND.n2094 65.0005
R5941 GND.n2094 GND.n2093 65.0005
R5942 GND.n2098 GND.n2097 65.0005
R5943 GND.n2099 GND.n2098 65.0005
R5944 GND.n2088 GND.n2087 65.0005
R5945 GND.n2087 GND.n2086 65.0005
R5946 GND.n2091 GND.n2090 65.0005
R5947 GND.n2092 GND.n2091 65.0005
R5948 GND.n2081 GND.n2080 65.0005
R5949 GND.n2080 GND.n2079 65.0005
R5950 GND.n2084 GND.n2083 65.0005
R5951 GND.n2085 GND.n2084 65.0005
R5952 GND.n2074 GND.n2073 65.0005
R5953 GND.n2073 GND.n2072 65.0005
R5954 GND.n2077 GND.n2076 65.0005
R5955 GND.n2078 GND.n2077 65.0005
R5956 GND.n2067 GND.n2066 65.0005
R5957 GND.n2066 GND.n2065 65.0005
R5958 GND.n2070 GND.n2069 65.0005
R5959 GND.n2071 GND.n2070 65.0005
R5960 GND.n732 GND.n731 65.0005
R5961 GND.n733 GND.n732 65.0005
R5962 GND.n724 GND.n723 65.0005
R5963 GND.n723 GND.n673 65.0005
R5964 GND.n744 GND.n743 65.0005
R5965 GND.n745 GND.n744 65.0005
R5966 GND.n737 GND.n736 65.0005
R5967 GND.n736 GND.n735 65.0005
R5968 GND.n750 GND.n749 65.0005
R5969 GND.n749 GND.n748 65.0005
R5970 GND.n746 GND.n711 65.0005
R5971 GND.n747 GND.n746 65.0005
R5972 GND.n766 GND.n765 65.0005
R5973 GND.n767 GND.n766 65.0005
R5974 GND.n755 GND.n754 65.0005
R5975 GND.n754 GND.n47 65.0005
R5976 GND.n771 GND.n770 65.0005
R5977 GND.n770 GND.n696 65.0005
R5978 GND.n759 GND.n706 65.0005
R5979 GND.n768 GND.n706 65.0005
R5980 GND.n2054 GND.n2053 65.0005
R5981 GND.n2053 GND.n2052 65.0005
R5982 GND.n2061 GND.n2060 65.0005
R5983 GND.n2062 GND.n2061 65.0005
R5984 GND.n2044 GND.n2043 65.0005
R5985 GND.n2043 GND.n2042 65.0005
R5986 GND.n2050 GND.n2049 65.0005
R5987 GND.n2051 GND.n2050 65.0005
R5988 GND.n790 GND.n786 65.0005
R5989 GND.n791 GND.n790 65.0005
R5990 GND.n2040 GND.n2039 65.0005
R5991 GND.n2041 GND.n2040 65.0005
R5992 GND.n2031 GND.n796 65.0005
R5993 GND.n2031 GND.n2030 65.0005
R5994 GND.n793 GND.n788 65.0005
R5995 GND.n793 GND.n792 65.0005
R5996 GND.n2021 GND.n2020 65.0005
R5997 GND.n2020 GND.n2019 65.0005
R5998 GND.n2028 GND.n2027 65.0005
R5999 GND.n2029 GND.n2028 65.0005
R6000 GND.n2012 GND.n2011 65.0005
R6001 GND.n2011 GND.n2010 65.0005
R6002 GND.n2015 GND.n2014 65.0005
R6003 GND.n2016 GND.n2015 65.0005
R6004 GND.n2005 GND.n2004 65.0005
R6005 GND.n2004 GND.n2003 65.0005
R6006 GND.n2008 GND.n2007 65.0005
R6007 GND.n2009 GND.n2008 65.0005
R6008 GND.n1998 GND.n1997 65.0005
R6009 GND.n1997 GND.n1996 65.0005
R6010 GND.n2001 GND.n2000 65.0005
R6011 GND.n2002 GND.n2001 65.0005
R6012 GND.n1991 GND.n1990 65.0005
R6013 GND.n1990 GND.n1989 65.0005
R6014 GND.n1994 GND.n1993 65.0005
R6015 GND.n1995 GND.n1994 65.0005
R6016 GND.n1984 GND.n1983 65.0005
R6017 GND.n1983 GND.n1982 65.0005
R6018 GND.n1987 GND.n1986 65.0005
R6019 GND.n1988 GND.n1987 65.0005
R6020 GND.n1424 GND.n1362 65.0005
R6021 GND.n1423 GND.n1362 65.0005
R6022 GND.n1361 GND.n1359 65.0005
R6023 GND.n1361 GND.n804 65.0005
R6024 GND.n1415 GND.n1414 65.0005
R6025 GND.n1414 GND.n1413 65.0005
R6026 GND.n1421 GND.n1420 65.0005
R6027 GND.n1422 GND.n1421 65.0005
R6028 GND.n1376 GND.n1375 65.0005
R6029 GND.n1375 GND.n1374 65.0005
R6030 GND.n1411 GND.n1410 65.0005
R6031 GND.n1412 GND.n1411 65.0005
R6032 GND.n1400 GND.n1381 65.0005
R6033 GND.n1399 GND.n1381 65.0005
R6034 GND.n1380 GND.n1378 65.0005
R6035 GND.n1380 GND.n68 65.0005
R6036 GND.n1390 GND.n1389 65.0005
R6037 GND.n1389 GND.n827 65.0005
R6038 GND.n1397 GND.n1396 65.0005
R6039 GND.n1398 GND.n1397 65.0005
R6040 GND.n1971 GND.n1970 65.0005
R6041 GND.n1970 GND.n1969 65.0005
R6042 GND.n1978 GND.n1977 65.0005
R6043 GND.n1979 GND.n1978 65.0005
R6044 GND.n1961 GND.n1960 65.0005
R6045 GND.n1960 GND.n1959 65.0005
R6046 GND.n1967 GND.n1966 65.0005
R6047 GND.n1968 GND.n1967 65.0005
R6048 GND.n1957 GND.n1956 65.0005
R6049 GND.n1958 GND.n1957 65.0005
R6050 GND.n1775 GND.n1774 65.0005
R6051 GND.n1776 GND.n1775 65.0005
R6052 GND.n1779 GND.n1778 65.0005
R6053 GND.n1778 GND.n1777 65.0005
R6054 GND.n1805 GND.n1804 65.0005
R6055 GND.n1806 GND.n1805 65.0005
R6056 GND.n1809 GND.n1808 65.0005
R6057 GND.n1808 GND.n1807 65.0005
R6058 GND.n1835 GND.n1834 65.0005
R6059 GND.n1836 GND.n1835 65.0005
R6060 GND.n1839 GND.n1838 65.0005
R6061 GND.n1838 GND.n1837 65.0005
R6062 GND.n1850 GND.n1849 65.0005
R6063 GND.n1851 GND.n1850 65.0005
R6064 GND.n1854 GND.n1853 65.0005
R6065 GND.n1853 GND.n1852 65.0005
R6066 GND.n1820 GND.n1819 65.0005
R6067 GND.n1821 GND.n1820 65.0005
R6068 GND.n1824 GND.n1823 65.0005
R6069 GND.n1823 GND.n1822 65.0005
R6070 GND.n1790 GND.n1789 65.0005
R6071 GND.n1791 GND.n1790 65.0005
R6072 GND.n1794 GND.n1793 65.0005
R6073 GND.n1793 GND.n1792 65.0005
R6074 GND.n1937 GND.n845 65.0005
R6075 GND.n1938 GND.n1937 65.0005
R6076 GND.n849 GND.n847 65.0005
R6077 GND.n1936 GND.n849 65.0005
R6078 GND.n1944 GND.n1943 65.0005
R6079 GND.n1945 GND.n1944 65.0005
R6080 GND.n1941 GND.n1940 65.0005
R6081 GND.n1940 GND.n1939 65.0005
R6082 GND.n1911 GND.n95 65.0005
R6083 GND.n1912 GND.n1911 65.0005
R6084 GND.n1913 GND.n1903 65.0005
R6085 GND.n1904 GND.n1903 65.0005
R6086 GND.n1902 GND.n1857 65.0005
R6087 GND.n1909 GND.n1902 65.0005
R6088 GND.n1591 GND.n1590 65.0005
R6089 GND.n1592 GND.n1591 65.0005
R6090 GND.n1577 GND.n1043 65.0005
R6091 GND.n1578 GND.n1577 65.0005
R6092 GND.n1603 GND.n1602 65.0005
R6093 GND.n1604 GND.n1603 65.0005
R6094 GND.n1596 GND.n1595 65.0005
R6095 GND.n1595 GND.n1594 65.0005
R6096 GND.n1617 GND.n1616 65.0005
R6097 GND.n1618 GND.n1617 65.0005
R6098 GND.n1610 GND.n1609 65.0005
R6099 GND.n1609 GND.n1608 65.0005
R6100 GND.n1583 GND.n1582 65.0005
R6101 GND.n1582 GND.n1581 65.0005
R6102 GND.n1053 GND.n1052 65.0005
R6103 GND.n1054 GND.n1053 65.0005
R6104 GND.n3115 GND.n3114 65.0005
R6105 GND.n3114 GND.n3113 65.0005
R6106 GND.n3118 GND.n3117 65.0005
R6107 GND.n3119 GND.n3118 65.0005
R6108 GND.n591 GND.n587 65.0005
R6109 GND.n3100 GND.n591 65.0005
R6110 GND.n584 GND.n580 65.0005
R6111 GND.n3112 GND.n580 65.0005
R6112 GND.n603 GND.n599 65.0005
R6113 GND.n3087 GND.n603 65.0005
R6114 GND.n596 GND.n592 65.0005
R6115 GND.n3099 GND.n592 65.0005
R6116 GND.n3069 GND.n614 65.0005
R6117 GND.n3064 GND.n614 65.0005
R6118 GND.n3067 GND.n613 65.0005
R6119 GND.n619 GND.n613 65.0005
R6120 GND.n632 GND.n628 65.0005
R6121 GND.n3051 GND.n632 65.0005
R6122 GND.n625 GND.n621 65.0005
R6123 GND.n3063 GND.n621 65.0005
R6124 GND.n3102 GND.n3101 65.0005
R6125 GND.n3101 GND.n3100 65.0005
R6126 GND.n3111 GND.n3110 65.0005
R6127 GND.n3112 GND.n3111 65.0005
R6128 GND.n3089 GND.n3088 65.0005
R6129 GND.n3088 GND.n3087 65.0005
R6130 GND.n3098 GND.n3097 65.0005
R6131 GND.n3099 GND.n3098 65.0005
R6132 GND.n617 GND.n607 65.0005
R6133 GND.n618 GND.n617 65.0005
R6134 GND.n3085 GND.n3084 65.0005
R6135 GND.n3086 GND.n3085 65.0005
R6136 GND.n3072 GND.n3065 65.0005
R6137 GND.n3065 GND.n3064 65.0005
R6138 GND.n3066 GND.n620 65.0005
R6139 GND.n620 GND.n619 65.0005
R6140 GND.n3053 GND.n3052 65.0005
R6141 GND.n3052 GND.n3051 65.0005
R6142 GND.n3062 GND.n3061 65.0005
R6143 GND.n3063 GND.n3062 65.0005
R6144 GND.n3124 GND.n3123 65.0005
R6145 GND.n3123 GND.n570 65.0005
R6146 GND.n2516 GND.n575 65.0005
R6147 GND.n3121 GND.n575 65.0005
R6148 GND.n3137 GND.n3136 65.0005
R6149 GND.n3136 GND.n3135 65.0005
R6150 GND.n3131 GND.n3130 65.0005
R6151 GND.n3132 GND.n3131 65.0005
R6152 GND.n3144 GND.n3143 65.0005
R6153 GND.n3145 GND.n3144 65.0005
R6154 GND.n3133 GND.n564 65.0005
R6155 GND.n3134 GND.n3133 65.0005
R6156 GND.n3155 GND.n3154 65.0005
R6157 GND.n3156 GND.n3155 65.0005
R6158 GND.n3149 GND.n3148 65.0005
R6159 GND.n3148 GND.n3147 65.0005
R6160 GND.n3166 GND.n3165 65.0005
R6161 GND.n3167 GND.n3166 65.0005
R6162 GND.n3159 GND.n3158 65.0005
R6163 GND.n3158 GND.n3157 65.0005
R6164 GND.n3188 GND.n3187 65.0005
R6165 GND.n3189 GND.n3188 65.0005
R6166 GND.n3185 GND.n3184 65.0005
R6167 GND.n3184 GND.n3183 65.0005
R6168 GND.n3193 GND.n3192 65.0005
R6169 GND.n3192 GND.n38 65.0005
R6170 GND.n545 GND.n540 65.0005
R6171 GND.n3190 GND.n540 65.0005
R6172 GND.n4241 GND.n4240 65.0005
R6173 GND.n4242 GND.n4241 65.0005
R6174 GND.n4238 GND.n4237 65.0005
R6175 GND.n4237 GND.n4236 65.0005
R6176 GND.n4249 GND.n4248 65.0005
R6177 GND.n4250 GND.n4249 65.0005
R6178 GND.n4246 GND.n4245 65.0005
R6179 GND.n4245 GND.n4244 65.0005
R6180 GND.n4256 GND.n4255 65.0005
R6181 GND.n4257 GND.n4256 65.0005
R6182 GND.n4253 GND.n4252 65.0005
R6183 GND.n4252 GND.n4251 65.0005
R6184 GND.n3033 GND.n2148 65.0005
R6185 GND.n3034 GND.n3033 65.0005
R6186 GND.n3048 GND.n3047 65.0005
R6187 GND.n3049 GND.n3048 65.0005
R6188 GND.n3036 GND.n3032 65.0005
R6189 GND.n3032 GND.n39 65.0005
R6190 GND.n3031 GND.n3029 65.0005
R6191 GND.n3035 GND.n3031 65.0005
R6192 GND.n4226 GND.n4225 65.0005
R6193 GND.n4225 GND.n4224 65.0005
R6194 GND.n4232 GND.n4231 65.0005
R6195 GND.n4233 GND.n4232 65.0005
R6196 GND.n58 GND.n52 65.0005
R6197 GND.n59 GND.n58 65.0005
R6198 GND.n4220 GND.n4219 65.0005
R6199 GND.n4221 GND.n4220 65.0005
R6200 GND.n4208 GND.n57 65.0005
R6201 GND.n4207 GND.n57 65.0005
R6202 GND.n56 GND.n54 65.0005
R6203 GND.n60 GND.n56 65.0005
R6204 GND.n4197 GND.n4196 65.0005
R6205 GND.n4196 GND.n4195 65.0005
R6206 GND.n4203 GND.n4202 65.0005
R6207 GND.n4204 GND.n4203 65.0005
R6208 GND.n79 GND.n73 65.0005
R6209 GND.n80 GND.n79 65.0005
R6210 GND.n4191 GND.n4190 65.0005
R6211 GND.n4192 GND.n4191 65.0005
R6212 GND.n4179 GND.n78 65.0005
R6213 GND.n4178 GND.n78 65.0005
R6214 GND.n77 GND.n75 65.0005
R6215 GND.n81 GND.n77 65.0005
R6216 GND.n3592 GND.n3591 65.0005
R6217 GND.n3591 GND.n3590 65.0005
R6218 GND.n3595 GND.n3594 65.0005
R6219 GND.n3596 GND.n3595 65.0005
R6220 GND.n89 GND.n85 65.0005
R6221 GND.n1905 GND.n85 65.0005
R6222 GND.n87 GND.n84 65.0005
R6223 GND.n3589 GND.n84 65.0005
R6224 GND.n1907 GND.n93 65.0005
R6225 GND.n1907 GND.n1906 65.0005
R6226 GND.n3601 GND.n3600 65.0005
R6227 GND.n3600 GND.n336 65.0005
R6228 GND.n3578 GND.n341 65.0005
R6229 GND.n3598 GND.n341 65.0005
R6230 GND.n3614 GND.n3613 65.0005
R6231 GND.n3613 GND.n3612 65.0005
R6232 GND.n3608 GND.n3607 65.0005
R6233 GND.n3609 GND.n3608 65.0005
R6234 GND.n3621 GND.n3620 65.0005
R6235 GND.n3622 GND.n3621 65.0005
R6236 GND.n3610 GND.n330 65.0005
R6237 GND.n3611 GND.n3610 65.0005
R6238 GND.n3632 GND.n3631 65.0005
R6239 GND.n3633 GND.n3632 65.0005
R6240 GND.n3626 GND.n3625 65.0005
R6241 GND.n3625 GND.n3624 65.0005
R6242 GND.n3675 GND.n3674 65.0005
R6243 GND.n3676 GND.n3675 65.0005
R6244 GND.n3636 GND.n3635 65.0005
R6245 GND.n3635 GND.n3634 65.0005
R6246 GND.n101 GND.n100 65.0005
R6247 GND.n4160 GND.n100 65.0005
R6248 GND.n99 GND.n97 65.0005
R6249 GND.n1757 GND.n99 65.0005
R6250 GND.n4155 GND.n4154 65.0005
R6251 GND.n4154 GND.n4153 65.0005
R6252 GND.n4158 GND.n4157 65.0005
R6253 GND.n4159 GND.n4158 65.0005
R6254 GND.n4133 GND.n4132 65.0005
R6255 GND.n4132 GND.n4131 65.0005
R6256 GND.n4136 GND.n4135 65.0005
R6257 GND.n4137 GND.n4136 65.0005
R6258 GND.n4126 GND.n4125 65.0005
R6259 GND.n4125 GND.n4124 65.0005
R6260 GND.n4129 GND.n4128 65.0005
R6261 GND.n4130 GND.n4129 65.0005
R6262 GND.n4119 GND.n4118 65.0005
R6263 GND.n4118 GND.n4117 65.0005
R6264 GND.n4122 GND.n4121 65.0005
R6265 GND.n4123 GND.n4122 65.0005
R6266 GND.n4112 GND.n4111 65.0005
R6267 GND.n4111 GND.n4110 65.0005
R6268 GND.n4115 GND.n4114 65.0005
R6269 GND.n4116 GND.n4115 65.0005
R6270 GND.n4105 GND.n4104 65.0005
R6271 GND.n4104 GND.n4103 65.0005
R6272 GND.n4108 GND.n4107 65.0005
R6273 GND.n4109 GND.n4108 65.0005
R6274 GND.n4088 GND.n4087 65.0005
R6275 GND.n4087 GND.n4086 65.0005
R6276 GND.n4091 GND.n4090 65.0005
R6277 GND.n4092 GND.n4091 65.0005
R6278 GND.n4081 GND.n4080 65.0005
R6279 GND.n4080 GND.n4079 65.0005
R6280 GND.n4084 GND.n4083 65.0005
R6281 GND.n4085 GND.n4084 65.0005
R6282 GND.n4074 GND.n4073 65.0005
R6283 GND.n4073 GND.n4072 65.0005
R6284 GND.n4077 GND.n4076 65.0005
R6285 GND.n4078 GND.n4077 65.0005
R6286 GND.n4067 GND.n4066 65.0005
R6287 GND.n4066 GND.n4065 65.0005
R6288 GND.n4070 GND.n4069 65.0005
R6289 GND.n4071 GND.n4070 65.0005
R6290 GND.n4060 GND.n4059 65.0005
R6291 GND.n4059 GND.n4058 65.0005
R6292 GND.n4063 GND.n4062 65.0005
R6293 GND.n4064 GND.n4063 65.0005
R6294 GND.n4038 GND.n4037 65.0005
R6295 GND.n4037 GND.n4036 65.0005
R6296 GND.n4041 GND.n4040 65.0005
R6297 GND.n4042 GND.n4041 65.0005
R6298 GND.n4031 GND.n4030 65.0005
R6299 GND.n4030 GND.n4029 65.0005
R6300 GND.n4034 GND.n4033 65.0005
R6301 GND.n4035 GND.n4034 65.0005
R6302 GND.n4024 GND.n4023 65.0005
R6303 GND.n4023 GND.n4022 65.0005
R6304 GND.n4027 GND.n4026 65.0005
R6305 GND.n4028 GND.n4027 65.0005
R6306 GND.n4017 GND.n4016 65.0005
R6307 GND.n4016 GND.n4015 65.0005
R6308 GND.n4020 GND.n4019 65.0005
R6309 GND.n4021 GND.n4020 65.0005
R6310 GND.n4010 GND.n4009 65.0005
R6311 GND.n4009 GND.n4008 65.0005
R6312 GND.n4013 GND.n4012 65.0005
R6313 GND.n4014 GND.n4013 65.0005
R6314 GND.n3986 GND.n3985 65.0005
R6315 GND.n3985 GND.n3984 65.0005
R6316 GND.n3989 GND.n3988 65.0005
R6317 GND.n3990 GND.n3989 65.0005
R6318 GND.n3979 GND.n3978 65.0005
R6319 GND.n3978 GND.n3977 65.0005
R6320 GND.n3982 GND.n3981 65.0005
R6321 GND.n3983 GND.n3982 65.0005
R6322 GND.n3972 GND.n3971 65.0005
R6323 GND.n3971 GND.n3970 65.0005
R6324 GND.n3975 GND.n3974 65.0005
R6325 GND.n3976 GND.n3975 65.0005
R6326 GND.n3965 GND.n3964 65.0005
R6327 GND.n3968 GND.n3967 65.0005
R6328 GND.n3969 GND.n3968 65.0005
R6329 GND.n3677 GND.n112 65.0005
R6330 GND.n3678 GND.n3677 65.0005
R6331 GND.n4151 GND.n4150 65.0005
R6332 GND.n4152 GND.n4151 65.0005
R6333 GND.n4139 GND.n118 65.0005
R6334 GND.n4138 GND.n118 65.0005
R6335 GND.n117 GND.n115 65.0005
R6336 GND.n3679 GND.n117 65.0005
R6337 GND.n4095 GND.n4094 65.0005
R6338 GND.n4094 GND.n4093 65.0005
R6339 GND.n4101 GND.n4100 65.0005
R6340 GND.n4102 GND.n4101 65.0005
R6341 GND.n3830 GND.n171 65.0005
R6342 GND.n3831 GND.n3830 65.0005
R6343 GND.n4056 GND.n4055 65.0005
R6344 GND.n4057 GND.n4056 65.0005
R6345 GND.n4044 GND.n176 65.0005
R6346 GND.n4043 GND.n176 65.0005
R6347 GND.n175 GND.n173 65.0005
R6348 GND.n3832 GND.n175 65.0005
R6349 GND.n4000 GND.n3999 65.0005
R6350 GND.n3999 GND.n3998 65.0005
R6351 GND.n4006 GND.n4005 65.0005
R6352 GND.n4007 GND.n4006 65.0005
R6353 GND.n3993 GND.n3992 65.0005
R6354 GND.n3992 GND.n3991 65.0005
R6355 GND.n3996 GND.n3995 65.0005
R6356 GND.n3997 GND.n3996 65.0005
R6357 GND.n1939 GND.n841 62.4595
R6358 GND.n1945 GND.n1758 62.4595
R6359 GND.n4147 GND.t216 61.1579
R6360 GND.n145 GND.t70 61.1579
R6361 GND.n146 GND.t432 61.1579
R6362 GND.n4052 GND.t807 61.1579
R6363 GND.n203 GND.t79 61.1579
R6364 GND.n204 GND.t290 61.1579
R6365 GND.n3262 GND.t325 61.1579
R6366 GND.n3391 GND.t672 61.1579
R6367 GND.n3351 GND.t619 61.1579
R6368 GND.n3376 GND.t306 61.1579
R6369 GND.n3362 GND.t82 61.1579
R6370 GND.n3940 GND.t524 61.1579
R6371 GND.n3934 GND.t171 61.1579
R6372 GND.n3928 GND.t458 61.1579
R6373 GND.n3896 GND.t278 61.1579
R6374 GND.n3902 GND.t123 61.1579
R6375 GND.n275 GND.t579 61.1579
R6376 GND.n3840 GND.t121 61.1579
R6377 GND.n3853 GND.t19 61.1579
R6378 GND.n251 GND.t363 61.1579
R6379 GND.n246 GND.t814 61.1579
R6380 GND.n3778 GND.t547 61.1579
R6381 GND.n3772 GND.t149 61.1579
R6382 GND.n3766 GND.t225 61.1579
R6383 GND.n3743 GND.t228 61.1579
R6384 GND.n3745 GND.t103 61.1579
R6385 GND.n3643 GND.t534 61.1579
R6386 GND.n3687 GND.t834 61.1579
R6387 GND.n3700 GND.t454 61.1579
R6388 GND.n301 GND.t683 61.1579
R6389 GND.n296 GND.t165 61.1579
R6390 GND.n3581 GND.t486 61.1579
R6391 GND.n3604 GND.t117 61.1579
R6392 GND.n3617 GND.t14 61.1579
R6393 GND.n326 GND.t783 61.1579
R6394 GND.n321 GND.t179 61.1579
R6395 GND.n3465 GND.t510 61.1579
R6396 GND.n3470 GND.t147 61.1579
R6397 GND.n3475 GND.t841 61.1579
R6398 GND.n3499 GND.t247 61.1579
R6399 GND.n3484 GND.t145 61.1579
R6400 GND.n3318 GND.t571 61.1579
R6401 GND.n3404 GND.t828 61.1579
R6402 GND.n3417 GND.t447 61.1579
R6403 GND.n391 GND.t282 61.1579
R6404 GND.n386 GND.t163 61.1579
R6405 GND.n4297 GND.t530 61.1579
R6406 GND.n4291 GND.t816 61.1579
R6407 GND.n4285 GND.t296 61.1579
R6408 GND.n17 GND.t40 61.1579
R6409 GND.n23 GND.t119 61.1579
R6410 GND.n3255 GND.t545 61.1579
R6411 GND.n3275 GND.t151 61.1579
R6412 GND.n3288 GND.t460 61.1579
R6413 GND.n497 GND.t602 61.1579
R6414 GND.n3303 GND.t169 61.1579
R6415 GND.n523 GND.t356 61.1579
R6416 GND.n645 GND.t141 61.1579
R6417 GND.n650 GND.t347 61.1579
R6418 GND.n2119 GND.t16 61.1579
R6419 GND.n671 GND.t824 61.1579
R6420 GND.n672 GND.t502 61.1579
R6421 GND.n728 GND.t113 61.1579
R6422 GND.n740 GND.t344 61.1579
R6423 GND.n753 GND.t456 61.1579
R6424 GND.n762 GND.t143 61.1579
R6425 GND.n774 GND.t516 61.1579
R6426 GND.n776 GND.t830 61.1579
R6427 GND.n781 GND.t34 61.1579
R6428 GND.n2036 GND.t260 61.1579
R6429 GND.n802 GND.t131 61.1579
R6430 GND.n803 GND.t559 61.1579
R6431 GND.n1368 GND.t157 61.1579
R6432 GND.n1369 GND.t233 61.1579
R6433 GND.n1407 GND.t303 61.1579
R6434 GND.n1387 GND.t109 61.1579
R6435 GND.n1388 GND.t488 61.1579
R6436 GND.n834 GND.t822 61.1579
R6437 GND.n839 GND.t184 61.1579
R6438 GND.n1953 GND.t329 61.1579
R6439 GND.n856 GND.t161 61.1579
R6440 GND.n857 GND.t536 61.1579
R6441 GND.n864 GND.t139 61.1579
R6442 GND.n869 GND.t309 61.1579
R6443 GND.n1717 GND.t12 61.1579
R6444 GND.n1711 GND.t137 61.1579
R6445 GND.n1705 GND.t549 61.1579
R6446 GND.n1135 GND.t111 61.1579
R6447 GND.n1086 GND.t812 61.1579
R6448 GND.n1120 GND.t452 61.1579
R6449 GND.n1114 GND.t177 61.1579
R6450 GND.n1108 GND.t573 61.1579
R6451 GND.n914 GND.t492 61.1579
R6452 GND.n919 GND.t371 61.1579
R6453 GND.n1641 GND.t845 61.1579
R6454 GND.n1635 GND.t522 61.1579
R6455 GND.n1629 GND.t155 61.1579
R6456 GND.n1627 GND.t642 61.1579
R6457 GND.n969 GND.t563 61.1579
R6458 GND.n974 GND.t127 61.1579
R6459 GND.n979 GND.t860 61.1579
R6460 GND.n982 GND.t167 61.1579
R6461 GND.n966 GND.t387 61.1579
R6462 GND.n964 GND.t175 61.1579
R6463 GND.n959 GND.t526 61.1579
R6464 GND.n954 GND.t871 61.1579
R6465 GND.n1697 GND.t500 61.1579
R6466 GND.n1512 GND.t407 61.1579
R6467 GND.n1514 GND.t832 61.1579
R6468 GND.n1519 GND.t581 61.1579
R6469 GND.n1524 GND.t312 61.1579
R6470 GND.n1527 GND.t575 61.1579
R6471 GND.n1508 GND.t752 61.1579
R6472 GND.n1455 GND.t115 61.1579
R6473 GND.n1460 GND.t551 61.1579
R6474 GND.n1465 GND.t788 61.1579
R6475 GND.n1468 GND.t520 61.1579
R6476 GND.n1452 GND.t24 61.1579
R6477 GND.n1450 GND.t173 61.1579
R6478 GND.n1445 GND.t480 61.1579
R6479 GND.n1440 GND.t690 61.1579
R6480 GND.n1437 GND.t557 61.1579
R6481 GND.n1356 GND.t722 61.1579
R6482 GND.n1304 GND.t826 61.1579
R6483 GND.n1309 GND.t490 61.1579
R6484 GND.n1314 GND.t411 61.1579
R6485 GND.n1317 GND.t512 61.1579
R6486 GND.n1301 GND.t799 61.1579
R6487 GND.n1299 GND.t135 61.1579
R6488 GND.n1294 GND.t567 61.1579
R6489 GND.n1289 GND.t257 61.1579
R6490 GND.n1286 GND.t498 61.1579
R6491 GND.n1277 GND.t613 61.1579
R6492 GND.n1227 GND.t159 61.1579
R6493 GND.n1232 GND.t518 61.1579
R6494 GND.n1237 GND.t65 61.1579
R6495 GND.n1240 GND.t569 61.1579
R6496 GND.n2866 GND.t8 61.1579
R6497 GND.n2472 GND.t541 61.1579
R6498 GND.n2478 GND.t332 61.1579
R6499 GND.n2841 GND.t675 61.1579
R6500 GND.n2815 GND.t496 61.1579
R6501 GND.n2828 GND.t771 61.1579
R6502 GND.n2797 GND.t804 61.1579
R6503 GND.n2787 GND.t468 61.1579
R6504 GND.n2504 GND.t426 61.1579
R6505 GND.n2502 GND.t436 61.1579
R6506 GND.n2872 GND.t543 61.1579
R6507 GND.n2872 GND.t748 61.1579
R6508 GND.n2884 GND.t238 61.1579
R6509 GND.n2884 GND.t275 61.1579
R6510 GND.n2894 GND.t658 61.1579
R6511 GND.n2948 GND.t853 61.1579
R6512 GND.n2948 GND.t790 61.1579
R6513 GND.n2913 GND.t761 61.1579
R6514 GND.n2913 GND.t385 61.1579
R6515 GND.n2870 GND.t740 61.1579
R6516 GND.n2340 GND.t240 61.1579
R6517 GND.n2340 GND.t719 61.1579
R6518 GND.n2352 GND.t750 61.1579
R6519 GND.n2352 GND.t763 61.1579
R6520 GND.n2362 GND.t621 61.1579
R6521 GND.n2416 GND.t367 61.1579
R6522 GND.n2416 GND.t636 61.1579
R6523 GND.n2381 GND.t639 61.1579
R6524 GND.n2381 GND.t236 61.1579
R6525 GND.n2454 GND.t736 61.1579
R6526 GND.n2213 GND.t390 61.1579
R6527 GND.n2213 GND.t396 61.1579
R6528 GND.n2225 GND.t716 61.1579
R6529 GND.n2225 GND.t428 61.1579
R6530 GND.n2235 GND.t595 61.1579
R6531 GND.n2289 GND.t597 61.1579
R6532 GND.n2289 GND.t320 61.1579
R6533 GND.n2254 GND.t723 61.1579
R6534 GND.n2254 GND.t652 61.1579
R6535 GND.n2327 GND.t850 61.1579
R6536 GND.n2535 GND.t242 61.1579
R6537 GND.n2535 GND.t680 61.1579
R6538 GND.n2547 GND.t274 61.1579
R6539 GND.n2547 GND.t653 61.1579
R6540 GND.n2557 GND.t250 61.1579
R6541 GND.n2611 GND.t608 61.1579
R6542 GND.n2611 GND.t873 61.1579
R6543 GND.n2576 GND.t663 61.1579
R6544 GND.n2576 GND.t6 61.1579
R6545 GND.n2649 GND.t738 61.1579
R6546 GND.n2656 GND.t650 61.1579
R6547 GND.n2656 GND.t772 61.1579
R6548 GND.n2668 GND.t28 61.1579
R6549 GND.n2668 GND.t399 61.1579
R6550 GND.n2678 GND.t4 61.1579
R6551 GND.n2732 GND.t632 61.1579
R6552 GND.n2732 GND.t669 61.1579
R6553 GND.n2697 GND.t681 61.1579
R6554 GND.n2697 GND.t423 61.1579
R6555 GND.n2654 GND.t698 61.1579
R6556 GND.n45 GND.t847 61.1579
R6557 GND.n4216 GND.t758 61.1579
R6558 GND.n65 GND.t744 61.1579
R6559 GND.n66 GND.t718 61.1579
R6560 GND.n4187 GND.t202 61.1579
R6561 GND.n1044 GND.t863 61.1579
R6562 GND.n1586 GND.t747 61.1579
R6563 GND.n1587 GND.t727 61.1579
R6564 GND.n1599 GND.t334 61.1579
R6565 GND.n1613 GND.t401 61.1579
R6566 GND.n3044 GND.t645 61.1579
R6567 GND.n3027 GND.t59 61.1579
R6568 GND.n2185 GND.t615 61.1579
R6569 GND.n2188 GND.t266 61.1579
R6570 GND.n2193 GND.t394 61.1579
R6571 GND.n2198 GND.t425 61.1579
R6572 GND.n2200 GND.t742 61.1579
R6573 GND.n2519 GND.t837 61.1579
R6574 GND.n3127 GND.t398 61.1579
R6575 GND.n3140 GND.t794 61.1579
R6576 GND.n560 GND.t253 61.1579
R6577 GND.n555 GND.t421 61.1579
R6578 GND.n586 GND.t764 61.1579
R6579 GND.n586 GND.t271 61.1579
R6580 GND.n598 GND.t854 61.1579
R6581 GND.n598 GND.t339 61.1579
R6582 GND.n608 GND.t884 61.1579
R6583 GND.n3081 GND.t341 61.1579
R6584 GND.n3081 GND.t616 61.1579
R6585 GND.n627 GND.t192 61.1579
R6586 GND.n627 GND.t10 61.1579
R6587 GND.n2521 GND.t852 61.1579
R6588 GND.n3959 GND.t577 61.1579
R6589 GND.n3956 GND.t264 61.1579
R6590 GND.n3951 GND.t528 61.1579
R6591 GND.n3946 GND.t133 61.1579
R6592 GND.n3944 GND.t92 61.1579
R6593 GND.n3806 GND.t508 61.1579
R6594 GND.n3809 GND.t445 61.1579
R6595 GND.n3814 GND.t476 61.1579
R6596 GND.n3819 GND.t818 61.1579
R6597 GND.n3821 GND.t857 61.1579
R6598 GND.n3797 GND.t494 61.1579
R6599 GND.n3794 GND.t625 61.1579
R6600 GND.n3789 GND.t555 61.1579
R6601 GND.n3784 GND.t105 61.1579
R6602 GND.n3782 GND.t1 61.1579
R6603 GND.n3653 GND.t538 61.1579
R6604 GND.n3656 GND.t430 61.1579
R6605 GND.n3661 GND.t478 61.1579
R6606 GND.n3666 GND.t125 61.1579
R6607 GND.n3668 GND.t665 61.1579
R6608 GND.n3644 GND.t514 61.1579
R6609 GND.n4166 GND.t630 61.1579
R6610 GND.n4172 GND.t482 61.1579
R6611 GND.n3586 GND.t181 61.1579
R6612 GND.n3585 GND.t84 61.1579
R6613 GND.n3553 GND.t565 61.1579
R6614 GND.n3548 GND.t245 61.1579
R6615 GND.n3454 GND.t561 61.1579
R6616 GND.n3459 GND.t153 61.1579
R6617 GND.n3461 GND.t31 61.1579
R6618 GND.n454 GND.t540 61.1579
R6619 GND.n451 GND.t314 61.1579
R6620 GND.n446 GND.t504 61.1579
R6621 GND.n441 GND.t820 61.1579
R6622 GND.n486 GND.t705 61.1579
R6623 GND.n3325 GND.t532 61.1579
R6624 GND.n421 GND.t785 61.1579
R6625 GND.n3227 GND.t553 61.1579
R6626 GND.n3222 GND.t107 61.1579
R6627 GND.n3250 GND.t336 61.1579
R6628 GND.n3204 GND.t484 61.1579
R6629 GND.n3201 GND.t667 61.1579
R6630 GND.n3196 GND.t506 61.1579
R6631 GND.n548 GND.t129 61.1579
R6632 GND.n544 GND.t656 61.1579
R6633 GND GND.t374 61.1525
R6634 GND GND.t205 61.1525
R6635 GND GND.t702 61.1525
R6636 GND GND.t317 61.1525
R6637 GND GND.t590 61.1525
R6638 GND GND.t48 61.1525
R6639 GND GND.t778 61.1525
R6640 GND.n1856 GND.t695 61.1525
R6641 GND.n3445 GND.n381 59.5094
R6642 GND.n3527 GND.n371 59.5094
R6643 GND.n3346 GND.n3344 59.5094
R6644 GND.n3397 GND.n3396 59.5094
R6645 GND.n3572 GND.n350 59.5094
R6646 GND.n3597 GND.n342 59.5094
R6647 GND.n4258 GND.n24 59.5094
R6648 GND.n3268 GND.n3267 59.5094
R6649 GND.n1931 GND 58.3538
R6650 GND.n3059 GND.n626 57.536
R6651 GND.n3055 GND.n626 57.536
R6652 GND.n3095 GND.n597 57.536
R6653 GND.n3091 GND.n597 57.536
R6654 GND.n3108 GND.n585 57.536
R6655 GND.n3104 GND.n585 57.536
R6656 GND.n2926 GND.n2912 57.536
R6657 GND.n2922 GND.n2912 57.536
R6658 GND.n2962 GND.n2883 57.536
R6659 GND.n2958 GND.n2883 57.536
R6660 GND.n2975 GND.n2181 57.536
R6661 GND.n2971 GND.n2181 57.536
R6662 GND.n2394 GND.n2380 57.536
R6663 GND.n2390 GND.n2380 57.536
R6664 GND.n2430 GND.n2351 57.536
R6665 GND.n2426 GND.n2351 57.536
R6666 GND.n2443 GND.n2339 57.536
R6667 GND.n2439 GND.n2339 57.536
R6668 GND.n2267 GND.n2253 57.536
R6669 GND.n2263 GND.n2253 57.536
R6670 GND.n2303 GND.n2224 57.536
R6671 GND.n2299 GND.n2224 57.536
R6672 GND.n2316 GND.n2212 57.536
R6673 GND.n2312 GND.n2212 57.536
R6674 GND.n2589 GND.n2575 57.536
R6675 GND.n2585 GND.n2575 57.536
R6676 GND.n2625 GND.n2546 57.536
R6677 GND.n2621 GND.n2546 57.536
R6678 GND.n2638 GND.n2534 57.536
R6679 GND.n2634 GND.n2534 57.536
R6680 GND.n2710 GND.n2696 57.536
R6681 GND.n2706 GND.n2696 57.536
R6682 GND.n2746 GND.n2667 57.536
R6683 GND.n2742 GND.n2667 57.536
R6684 GND.n2759 GND.n2515 57.536
R6685 GND.n2755 GND.n2515 57.536
R6686 GND.n1580 GND.n1579 54.9156
R6687 GND.n1606 GND.n1605 54.9156
R6688 GND.n4223 GND.n4222 54.9156
R6689 GND.n4206 GND.n4205 54.9156
R6690 GND.n4194 GND.n4193 54.9156
R6691 GND.n220 GND.n219 52.5417
R6692 GND.n219 GND.n218 52.5417
R6693 GND.n193 GND.n192 52.5417
R6694 GND.n192 GND.n191 52.5417
R6695 GND.n162 GND.n161 52.5417
R6696 GND.n161 GND.n160 52.5417
R6697 GND.n135 GND.n134 52.5417
R6698 GND.n134 GND.n133 52.5417
R6699 GND.n4163 GND.n98 52.5417
R6700 GND.n4164 GND.n4163 52.5417
R6701 GND.n32 GND.n31 52.5417
R6702 GND.n33 GND.n32 52.5417
R6703 GND.n3042 GND.n3041 52.5417
R6704 GND.n3041 GND.n3030 52.5417
R6705 GND.n1611 GND.n1034 52.5417
R6706 GND.n1615 GND.n1034 52.5417
R6707 GND.n1597 GND.n1039 52.5417
R6708 GND.n1601 GND.n1039 52.5417
R6709 GND.n1222 GND.n1221 52.5417
R6710 GND.n1221 GND.n1220 52.5417
R6711 GND.n682 GND.n681 52.5417
R6712 GND.n683 GND.n682 52.5417
R6713 GND.n1200 GND.n1199 52.5417
R6714 GND.n1201 GND.n1200 52.5417
R6715 GND.n813 GND.n812 52.5417
R6716 GND.n814 GND.n813 52.5417
R6717 GND.n1729 GND.n868 52.5417
R6718 GND.n1726 GND.n868 52.5417
R6719 GND.n1133 GND.n1132 52.5417
R6720 GND.n1132 GND.n1075 52.5417
R6721 GND.n1653 GND.n918 52.5417
R6722 GND.n1650 GND.n918 52.5417
R6723 GND.n948 GND.n947 52.5417
R6724 GND.n949 GND.n948 52.5417
R6725 GND.n1694 GND.n890 52.5417
R6726 GND.n1695 GND.n1694 52.5417
R6727 GND.n1158 GND.n1157 52.5417
R6728 GND.n1159 GND.n1158 52.5417
R6729 GND.n1179 GND.n1178 52.5417
R6730 GND.n1180 GND.n1179 52.5417
R6731 GND.n1965 GND.n838 52.5417
R6732 GND.n1962 GND.n838 52.5417
R6733 GND.n1419 GND.n1366 52.5417
R6734 GND.n1416 GND.n1366 52.5417
R6735 GND.n2048 GND.n780 52.5417
R6736 GND.n2045 GND.n780 52.5417
R6737 GND.n738 GND.n718 52.5417
R6738 GND.n742 GND.n718 52.5417
R6739 GND.n420 GND.n419 52.5417
R6740 GND.n3328 GND.n420 52.5417
R6741 GND.n3298 GND.n496 52.5417
R6742 GND.n3305 GND.n496 52.5417
R6743 GND.n3497 GND.n3496 52.5417
R6744 GND.n3496 GND.n3478 52.5417
R6745 GND.n358 GND.n357 52.5417
R6746 GND.n3556 GND.n358 52.5417
R6747 GND.n439 GND.n438 52.5417
R6748 GND.n438 GND.n437 52.5417
R6749 GND.n3382 GND.n3361 52.5417
R6750 GND.n3379 GND.n3361 52.5417
R6751 GND.n3427 GND.n390 52.5417
R6752 GND.n3430 GND.n390 52.5417
R6753 GND.n3349 GND.n411 52.5417
R6754 GND.n3393 GND.n411 52.5417
R6755 GND.n532 GND.n517 52.5417
R6756 GND.n3264 GND.n517 52.5417
R6757 GND.n4004 GND.n202 52.5417
R6758 GND.n4001 GND.n202 52.5417
R6759 GND.n4050 GND.n4049 52.5417
R6760 GND.n4049 GND.n174 52.5417
R6761 GND.n4099 GND.n144 52.5417
R6762 GND.n4096 GND.n144 52.5417
R6763 GND.n4145 GND.n4144 52.5417
R6764 GND.n4144 GND.n116 52.5417
R6765 GND.n3374 GND.n3373 52.5417
R6766 GND.n3373 GND.n3365 52.5417
R6767 GND.n3627 GND.n325 52.5417
R6768 GND.n3630 GND.n325 52.5417
R6769 GND.n3919 GND.n3895 52.5417
R6770 GND.n3916 GND.n3895 52.5417
R6771 GND.n3863 GND.n250 52.5417
R6772 GND.n3866 GND.n250 52.5417
R6773 GND.n3757 GND.n3742 52.5417
R6774 GND.n3754 GND.n3742 52.5417
R6775 GND.n3710 GND.n300 52.5417
R6776 GND.n3713 GND.n300 52.5417
R6777 GND.n4276 GND.n16 52.5417
R6778 GND.n4273 GND.n16 52.5417
R6779 GND.n2131 GND.n649 52.5417
R6780 GND.n2128 GND.n649 52.5417
R6781 GND.n2157 GND.n2156 52.5417
R6782 GND.n2158 GND.n2157 52.5417
R6783 GND.n2839 GND.n2838 52.5417
R6784 GND.n2838 GND.n2481 52.5417
R6785 GND.n2831 GND.n2490 52.5417
R6786 GND.n2831 GND.n2830 52.5417
R6787 GND.n1051 GND.n1046 52.5417
R6788 GND.n1584 GND.n1046 52.5417
R6789 GND.n4185 GND.n4184 52.5417
R6790 GND.n4184 GND.n76 52.5417
R6791 GND.n4201 GND.n64 52.5417
R6792 GND.n4198 GND.n64 52.5417
R6793 GND.n4214 GND.n4213 52.5417
R6794 GND.n4213 GND.n55 52.5417
R6795 GND.n4230 GND.n43 52.5417
R6796 GND.n4227 GND.n43 52.5417
R6797 GND.n3150 GND.n559 52.5417
R6798 GND.n3153 GND.n559 52.5417
R6799 GND.n3050 GND.n3049 52.3938
R6800 GND.n1929 GND 48.6472
R6801 GND.n1822 GND.n841 45.6728
R6802 GND.n1821 GND.n1758 45.6728
R6803 GND.t25 GND.n1054 45.3202
R6804 GND.n1055 GND.t25 45.3202
R6805 GND.t746 GND.n1055 45.3202
R6806 GND.n1581 GND.t746 45.3202
R6807 GND.n1578 GND.t726 45.3202
R6808 GND.n1592 GND.t726 45.3202
R6809 GND.n1594 GND.t416 45.3202
R6810 GND.t416 GND.n1593 45.3202
R6811 GND.n1593 GND.t333 45.3202
R6812 GND.n1604 GND.t333 45.3202
R6813 GND.n1608 GND.t795 45.3202
R6814 GND.t795 GND.n1607 45.3202
R6815 GND.n1607 GND.t400 45.3202
R6816 GND.n1618 GND.t400 45.3202
R6817 GND.n3049 GND.t644 45.3202
R6818 GND.n3034 GND.t644 45.3202
R6819 GND.t379 GND.n3035 45.3202
R6820 GND.n3039 GND.t379 45.3202
R6821 GND.n3039 GND.t58 45.3202
R6822 GND.t58 GND.n39 45.3202
R6823 GND.n4233 GND.t874 45.3202
R6824 GND.n46 GND.t874 45.3202
R6825 GND.t846 GND.n46 45.3202
R6826 GND.n4224 GND.t846 45.3202
R6827 GND.n4221 GND.t757 45.3202
R6828 GND.n59 GND.t757 45.3202
R6829 GND.t294 GND.n60 45.3202
R6830 GND.n4211 GND.t294 45.3202
R6831 GND.n4211 GND.t743 45.3202
R6832 GND.t743 GND.n4207 45.3202
R6833 GND.n4204 GND.t801 45.3202
R6834 GND.n67 GND.t801 45.3202
R6835 GND.t717 GND.n67 45.3202
R6836 GND.n4195 GND.t717 45.3202
R6837 GND.n4192 GND.t201 45.3202
R6838 GND.n80 GND.t201 45.3202
R6839 GND.t418 GND.n81 45.3202
R6840 GND.n4182 GND.t418 45.3202
R6841 GND.n4182 GND.t862 45.3202
R6842 GND.t862 GND.n4178 45.3202
R6843 GND.n3050 GND.n639 43.0923
R6844 GND.n1332 GND.n1198 34.4123
R6845 GND.n1328 GND.n1198 34.4123
R6846 GND.n1200 GND.n1197 34.4123
R6847 GND.n1328 GND.n1197 34.4123
R6848 GND.n997 GND.n946 34.4123
R6849 GND.n993 GND.n946 34.4123
R6850 GND.n948 GND.n945 34.4123
R6851 GND.n993 GND.n945 34.4123
R6852 GND.n918 GND.n916 34.4123
R6853 GND.n920 GND.n916 34.4123
R6854 GND.n917 GND.n915 34.4123
R6855 GND.n920 GND.n915 34.4123
R6856 GND.n895 GND.n894 34.4123
R6857 GND.n1692 GND.n895 34.4123
R6858 GND.n1694 GND.n1693 34.4123
R6859 GND.n1693 GND.n1692 34.4123
R6860 GND.n1132 GND.n1131 34.4123
R6861 GND.n1131 GND.n1130 34.4123
R6862 GND.n1129 GND.n1128 34.4123
R6863 GND.n1130 GND.n1129 34.4123
R6864 GND.n1543 GND.n1156 34.4123
R6865 GND.n1539 GND.n1156 34.4123
R6866 GND.n1158 GND.n1155 34.4123
R6867 GND.n1539 GND.n1155 34.4123
R6868 GND.n868 GND.n866 34.4123
R6869 GND.n870 GND.n866 34.4123
R6870 GND.n867 GND.n865 34.4123
R6871 GND.n870 GND.n865 34.4123
R6872 GND.n1483 GND.n1177 34.4123
R6873 GND.n1479 GND.n1177 34.4123
R6874 GND.n1179 GND.n1176 34.4123
R6875 GND.n1479 GND.n1176 34.4123
R6876 GND.n3361 GND.n3359 34.4123
R6877 GND.n3359 GND.n3358 34.4123
R6878 GND.n3360 GND.n3357 34.4123
R6879 GND.n3358 GND.n3357 34.4123
R6880 GND.n390 GND.n388 34.4123
R6881 GND.n3423 GND.n388 34.4123
R6882 GND.n389 GND.n387 34.4123
R6883 GND.n3423 GND.n387 34.4123
R6884 GND.n463 GND.n436 34.4123
R6885 GND.n440 GND.n436 34.4123
R6886 GND.n438 GND.n435 34.4123
R6887 GND.n440 GND.n435 34.4123
R6888 GND.n411 GND.n409 34.4123
R6889 GND.n3345 GND.n409 34.4123
R6890 GND.n410 GND.n408 34.4123
R6891 GND.n3345 GND.n408 34.4123
R6892 GND.n3373 GND.n3372 34.4123
R6893 GND.n3372 GND.n3371 34.4123
R6894 GND.n3370 GND.n3369 34.4123
R6895 GND.n3371 GND.n3370 34.4123
R6896 GND.n3561 GND.n356 34.4123
R6897 GND.n3557 GND.n356 34.4123
R6898 GND.n358 GND.n355 34.4123
R6899 GND.n3557 GND.n355 34.4123
R6900 GND.n3496 GND.n3495 34.4123
R6901 GND.n3495 GND.n3494 34.4123
R6902 GND.n3493 GND.n3492 34.4123
R6903 GND.n3494 GND.n3493 34.4123
R6904 GND.n300 GND.n298 34.4123
R6905 GND.n3706 GND.n298 34.4123
R6906 GND.n299 GND.n297 34.4123
R6907 GND.n3706 GND.n297 34.4123
R6908 GND.n3742 GND.n3740 34.4123
R6909 GND.n3744 GND.n3740 34.4123
R6910 GND.n3741 GND.n3739 34.4123
R6911 GND.n3744 GND.n3739 34.4123
R6912 GND.n250 GND.n248 34.4123
R6913 GND.n3859 GND.n248 34.4123
R6914 GND.n249 GND.n247 34.4123
R6915 GND.n3859 GND.n247 34.4123
R6916 GND.n3895 GND.n3893 34.4123
R6917 GND.n3897 GND.n3893 34.4123
R6918 GND.n3894 GND.n3892 34.4123
R6919 GND.n3897 GND.n3892 34.4123
R6920 GND.n16 GND.n14 34.4123
R6921 GND.n18 GND.n14 34.4123
R6922 GND.n15 GND.n13 34.4123
R6923 GND.n18 GND.n13 34.4123
R6924 GND.n496 GND.n494 34.4123
R6925 GND.n3294 GND.n494 34.4123
R6926 GND.n495 GND.n493 34.4123
R6927 GND.n3294 GND.n493 34.4123
R6928 GND.n3333 GND.n418 34.4123
R6929 GND.n3329 GND.n418 34.4123
R6930 GND.n420 GND.n417 34.4123
R6931 GND.n3329 GND.n417 34.4123
R6932 GND.n517 GND.n515 34.4123
R6933 GND.n528 GND.n515 34.4123
R6934 GND.n516 GND.n514 34.4123
R6935 GND.n528 GND.n514 34.4123
R6936 GND.n1253 GND.n1219 34.4123
R6937 GND.n1249 GND.n1219 34.4123
R6938 GND.n1221 GND.n1218 34.4123
R6939 GND.n1249 GND.n1218 34.4123
R6940 GND.n2492 GND.n2484 34.4123
R6941 GND.n2836 GND.n2484 34.4123
R6942 GND.n2832 GND.n2831 34.4123
R6943 GND.n2836 GND.n2832 34.4123
R6944 GND.n2838 GND.n2837 34.4123
R6945 GND.n2837 GND.n2836 34.4123
R6946 GND.n2835 GND.n2834 34.4123
R6947 GND.n2836 GND.n2835 34.4123
R6948 GND.n2935 GND.n2902 34.4123
R6949 GND.n2942 GND.n2902 34.4123
R6950 GND.n2944 GND.n2943 34.4123
R6951 GND.n2943 GND.n2942 34.4123
R6952 GND.n2901 GND.n2897 34.4123
R6953 GND.n2942 GND.n2901 34.4123
R6954 GND.n2941 GND.n2940 34.4123
R6955 GND.n2942 GND.n2941 34.4123
R6956 GND.n2403 GND.n2370 34.4123
R6957 GND.n2410 GND.n2370 34.4123
R6958 GND.n2412 GND.n2411 34.4123
R6959 GND.n2411 GND.n2410 34.4123
R6960 GND.n2369 GND.n2365 34.4123
R6961 GND.n2410 GND.n2369 34.4123
R6962 GND.n2409 GND.n2408 34.4123
R6963 GND.n2410 GND.n2409 34.4123
R6964 GND.n2276 GND.n2243 34.4123
R6965 GND.n2283 GND.n2243 34.4123
R6966 GND.n2285 GND.n2284 34.4123
R6967 GND.n2284 GND.n2283 34.4123
R6968 GND.n2242 GND.n2238 34.4123
R6969 GND.n2283 GND.n2242 34.4123
R6970 GND.n2282 GND.n2281 34.4123
R6971 GND.n2283 GND.n2282 34.4123
R6972 GND.n2598 GND.n2565 34.4123
R6973 GND.n2605 GND.n2565 34.4123
R6974 GND.n2607 GND.n2606 34.4123
R6975 GND.n2606 GND.n2605 34.4123
R6976 GND.n2564 GND.n2560 34.4123
R6977 GND.n2605 GND.n2564 34.4123
R6978 GND.n2604 GND.n2603 34.4123
R6979 GND.n2605 GND.n2604 34.4123
R6980 GND.n2719 GND.n2686 34.4123
R6981 GND.n2726 GND.n2686 34.4123
R6982 GND.n2728 GND.n2727 34.4123
R6983 GND.n2727 GND.n2726 34.4123
R6984 GND.n2685 GND.n2681 34.4123
R6985 GND.n2726 GND.n2685 34.4123
R6986 GND.n2725 GND.n2724 34.4123
R6987 GND.n2726 GND.n2725 34.4123
R6988 GND.n3017 GND.n2155 34.4123
R6989 GND.n3013 GND.n2155 34.4123
R6990 GND.n2157 GND.n2154 34.4123
R6991 GND.n3013 GND.n2154 34.4123
R6992 GND.n649 GND.n647 34.4123
R6993 GND.n651 GND.n647 34.4123
R6994 GND.n648 GND.n646 34.4123
R6995 GND.n651 GND.n646 34.4123
R6996 GND.n2089 GND.n680 34.4123
R6997 GND.n684 GND.n680 34.4123
R6998 GND.n682 GND.n679 34.4123
R6999 GND.n684 GND.n679 34.4123
R7000 GND.n718 GND.n716 34.4123
R7001 GND.n734 GND.n716 34.4123
R7002 GND.n717 GND.n715 34.4123
R7003 GND.n734 GND.n715 34.4123
R7004 GND.n780 GND.n778 34.4123
R7005 GND.n782 GND.n778 34.4123
R7006 GND.n779 GND.n777 34.4123
R7007 GND.n782 GND.n777 34.4123
R7008 GND.n2006 GND.n811 34.4123
R7009 GND.n815 GND.n811 34.4123
R7010 GND.n813 GND.n810 34.4123
R7011 GND.n815 GND.n810 34.4123
R7012 GND.n1366 GND.n1364 34.4123
R7013 GND.n1370 GND.n1364 34.4123
R7014 GND.n1365 GND.n1363 34.4123
R7015 GND.n1370 GND.n1363 34.4123
R7016 GND.n838 GND.n836 34.4123
R7017 GND.n840 GND.n836 34.4123
R7018 GND.n837 GND.n835 34.4123
R7019 GND.n840 GND.n835 34.4123
R7020 GND.n1039 GND.n1037 34.4123
R7021 GND.n1593 GND.n1037 34.4123
R7022 GND.n1038 GND.n1036 34.4123
R7023 GND.n1593 GND.n1036 34.4123
R7024 GND.n1034 GND.n1032 34.4123
R7025 GND.n1607 GND.n1032 34.4123
R7026 GND.n1033 GND.n1031 34.4123
R7027 GND.n1607 GND.n1031 34.4123
R7028 GND.n1049 GND.n1046 34.4123
R7029 GND.n1055 GND.n1049 34.4123
R7030 GND.n1048 GND.n1047 34.4123
R7031 GND.n1055 GND.n1048 34.4123
R7032 GND.n3068 GND.n616 34.4123
R7033 GND.n3075 GND.n616 34.4123
R7034 GND.n3077 GND.n3076 34.4123
R7035 GND.n3076 GND.n3075 34.4123
R7036 GND.n615 GND.n611 34.4123
R7037 GND.n3075 GND.n615 34.4123
R7038 GND.n3074 GND.n3073 34.4123
R7039 GND.n3075 GND.n3074 34.4123
R7040 GND.n559 GND.n557 34.4123
R7041 GND.n3146 GND.n557 34.4123
R7042 GND.n558 GND.n556 34.4123
R7043 GND.n3146 GND.n556 34.4123
R7044 GND.n4247 GND.n30 34.4123
R7045 GND.n4243 GND.n30 34.4123
R7046 GND.n32 GND.n29 34.4123
R7047 GND.n4243 GND.n29 34.4123
R7048 GND.n3041 GND.n3040 34.4123
R7049 GND.n3040 GND.n3039 34.4123
R7050 GND.n3038 GND.n3037 34.4123
R7051 GND.n3039 GND.n3038 34.4123
R7052 GND.n43 GND.n41 34.4123
R7053 GND.n46 GND.n41 34.4123
R7054 GND.n42 GND.n40 34.4123
R7055 GND.n46 GND.n40 34.4123
R7056 GND.n4213 GND.n4212 34.4123
R7057 GND.n4212 GND.n4211 34.4123
R7058 GND.n4210 GND.n4209 34.4123
R7059 GND.n4211 GND.n4210 34.4123
R7060 GND.n64 GND.n62 34.4123
R7061 GND.n67 GND.n62 34.4123
R7062 GND.n63 GND.n61 34.4123
R7063 GND.n67 GND.n61 34.4123
R7064 GND.n4184 GND.n4183 34.4123
R7065 GND.n4183 GND.n4182 34.4123
R7066 GND.n4181 GND.n4180 34.4123
R7067 GND.n4182 GND.n4181 34.4123
R7068 GND.n325 GND.n323 34.4123
R7069 GND.n3623 GND.n323 34.4123
R7070 GND.n324 GND.n322 34.4123
R7071 GND.n3623 GND.n322 34.4123
R7072 GND.n103 GND.n102 34.4123
R7073 GND.n4161 GND.n103 34.4123
R7074 GND.n4163 GND.n4162 34.4123
R7075 GND.n4162 GND.n4161 34.4123
R7076 GND.n4113 GND.n132 34.4123
R7077 GND.n136 GND.n132 34.4123
R7078 GND.n134 GND.n131 34.4123
R7079 GND.n136 GND.n131 34.4123
R7080 GND.n4068 GND.n159 34.4123
R7081 GND.n163 GND.n159 34.4123
R7082 GND.n161 GND.n158 34.4123
R7083 GND.n163 GND.n158 34.4123
R7084 GND.n4018 GND.n190 34.4123
R7085 GND.n194 GND.n190 34.4123
R7086 GND.n192 GND.n189 34.4123
R7087 GND.n194 GND.n189 34.4123
R7088 GND.n3973 GND.n217 34.4123
R7089 GND.n221 GND.n217 34.4123
R7090 GND.n219 GND.n216 34.4123
R7091 GND.n221 GND.n216 34.4123
R7092 GND.n4144 GND.n4143 34.4123
R7093 GND.n4143 GND.n4142 34.4123
R7094 GND.n4141 GND.n4140 34.4123
R7095 GND.n4142 GND.n4141 34.4123
R7096 GND.n144 GND.n142 34.4123
R7097 GND.n3728 GND.n142 34.4123
R7098 GND.n143 GND.n141 34.4123
R7099 GND.n3728 GND.n141 34.4123
R7100 GND.n4049 GND.n4048 34.4123
R7101 GND.n4048 GND.n4047 34.4123
R7102 GND.n4046 GND.n4045 34.4123
R7103 GND.n4047 GND.n4046 34.4123
R7104 GND.n202 GND.n200 34.4123
R7105 GND.n3881 GND.n200 34.4123
R7106 GND.n201 GND.n199 34.4123
R7107 GND.n3881 GND.n199 34.4123
R7108 GND.n3259 GND.n535 33.6641
R7109 GND.n3078 GND.n611 29.7417
R7110 GND.n612 GND.n611 29.7417
R7111 GND.n3078 GND.n3077 29.7417
R7112 GND.n3077 GND.n612 29.7417
R7113 GND.n2945 GND.n2897 29.7417
R7114 GND.n2898 GND.n2897 29.7417
R7115 GND.n2945 GND.n2944 29.7417
R7116 GND.n2944 GND.n2898 29.7417
R7117 GND.n2413 GND.n2365 29.7417
R7118 GND.n2366 GND.n2365 29.7417
R7119 GND.n2413 GND.n2412 29.7417
R7120 GND.n2412 GND.n2366 29.7417
R7121 GND.n2286 GND.n2238 29.7417
R7122 GND.n2239 GND.n2238 29.7417
R7123 GND.n2286 GND.n2285 29.7417
R7124 GND.n2285 GND.n2239 29.7417
R7125 GND.n2608 GND.n2560 29.7417
R7126 GND.n2561 GND.n2560 29.7417
R7127 GND.n2608 GND.n2607 29.7417
R7128 GND.n2607 GND.n2561 29.7417
R7129 GND.n2729 GND.n2681 29.7417
R7130 GND.n2682 GND.n2681 29.7417
R7131 GND.n2729 GND.n2728 29.7417
R7132 GND.n2728 GND.n2682 29.7417
R7133 GND.n1927 GND 29.2342
R7134 GND.n1050 GND.n104 27.4581
R7135 GND.n4177 GND.n82 27.4581
R7136 GND.n4098 GND 26.3103
R7137 GND.n4053 GND 26.3103
R7138 GND.n4003 GND 26.3103
R7139 GND.n3350 GND 26.3103
R7140 GND GND.n3390 26.3103
R7141 GND GND.n3375 26.3103
R7142 GND.n4217 GND 26.3103
R7143 GND.n4200 GND 26.3103
R7144 GND.n4188 GND 26.3103
R7145 GND.n1045 GND 26.3103
R7146 GND.n1588 GND 26.3103
R7147 GND.n1612 GND 26.3103
R7148 GND GND.n44 24.8229
R7149 GND.n1339 GND.n1194 22.5005
R7150 GND.t659 GND.n1194 22.5005
R7151 GND.n1311 GND.n1193 22.5005
R7152 GND.t659 GND.n1193 22.5005
R7153 GND.n1346 GND.n1190 22.5005
R7154 GND.t720 GND.n1190 22.5005
R7155 GND.n1306 GND.n1189 22.5005
R7156 GND.t720 GND.n1189 22.5005
R7157 GND.n1205 GND.n1202 22.5005
R7158 GND.t626 GND.n1202 22.5005
R7159 GND.n1324 GND.n1203 22.5005
R7160 GND.n1203 GND.t626 22.5005
R7161 GND.n989 GND.n951 22.5005
R7162 GND.n951 GND.t41 22.5005
R7163 GND.n953 GND.n950 22.5005
R7164 GND.t41 GND.n950 22.5005
R7165 GND.n1004 GND.n942 22.5005
R7166 GND.t760 GND.n942 22.5005
R7167 GND.n976 GND.n941 22.5005
R7168 GND.t760 GND.n941 22.5005
R7169 GND.n1011 GND.n938 22.5005
R7170 GND.t676 GND.n938 22.5005
R7171 GND.n971 GND.n937 22.5005
R7172 GND.t676 GND.n937 22.5005
R7173 GND.n912 GND.n910 22.5005
R7174 GND.t464 GND.n910 22.5005
R7175 GND.n911 GND.n909 22.5005
R7176 GND.t464 GND.n909 22.5005
R7177 GND.n1638 GND.n927 22.5005
R7178 GND.t732 GND.n927 22.5005
R7179 GND.n1024 GND.n1020 22.5005
R7180 GND.n1024 GND.t732 22.5005
R7181 GND.n1632 GND.n931 22.5005
R7182 GND.t213 GND.n931 22.5005
R7183 GND.n1028 GND.n1018 22.5005
R7184 GND.n1028 GND.t213 22.5005
R7185 GND.n1066 GND.n1063 22.5005
R7186 GND.n1066 GND.t471 22.5005
R7187 GND.n1700 GND.n886 22.5005
R7188 GND.t471 GND.n886 22.5005
R7189 GND.n1687 GND.n897 22.5005
R7190 GND.t214 GND.n897 22.5005
R7191 GND.n956 GND.n896 22.5005
R7192 GND.t214 GND.n896 22.5005
R7193 GND.n1680 GND.n901 22.5005
R7194 GND.t762 GND.n901 22.5005
R7195 GND.n961 GND.n900 22.5005
R7196 GND.t762 GND.n900 22.5005
R7197 GND.n1138 GND.n1070 22.5005
R7198 GND.t691 GND.n1070 22.5005
R7199 GND.n1071 GND.n1069 22.5005
R7200 GND.t691 GND.n1069 22.5005
R7201 GND.n1117 GND.n1089 22.5005
R7202 GND.n1089 GND.t712 22.5005
R7203 GND.n1101 GND.n1100 22.5005
R7204 GND.n1101 GND.t712 22.5005
R7205 GND.n1111 GND.n1093 22.5005
R7206 GND.t466 GND.n1093 22.5005
R7207 GND.n1105 GND.n1094 22.5005
R7208 GND.n1105 GND.t466 22.5005
R7209 GND.n1535 GND.n1161 22.5005
R7210 GND.t276 GND.n1161 22.5005
R7211 GND.n1163 GND.n1160 22.5005
R7212 GND.t276 GND.n1160 22.5005
R7213 GND.n1550 GND.n1152 22.5005
R7214 GND.t93 GND.n1152 22.5005
R7215 GND.n1521 GND.n1151 22.5005
R7216 GND.t93 GND.n1151 22.5005
R7217 GND.n1557 GND.n1148 22.5005
R7218 GND.t797 GND.n1148 22.5005
R7219 GND.n1516 GND.n1147 22.5005
R7220 GND.t797 GND.n1147 22.5005
R7221 GND.n862 GND.n860 22.5005
R7222 GND.t88 GND.n860 22.5005
R7223 GND.n861 GND.n859 22.5005
R7224 GND.t88 GND.n859 22.5005
R7225 GND.n1714 GND.n877 22.5005
R7226 GND.t219 GND.n877 22.5005
R7227 GND.n1576 GND.n1575 22.5005
R7228 GND.t219 GND.n1576 22.5005
R7229 GND.n1708 GND.n881 22.5005
R7230 GND.t864 GND.n881 22.5005
R7231 GND.n1570 GND.n1061 22.5005
R7232 GND.n1570 GND.t864 22.5005
R7233 GND.n1475 GND.n1182 22.5005
R7234 GND.n1182 GND.t280 22.5005
R7235 GND.n1184 GND.n1181 22.5005
R7236 GND.t280 GND.n1181 22.5005
R7237 GND.n1490 GND.n1173 22.5005
R7238 GND.t866 GND.n1173 22.5005
R7239 GND.n1462 GND.n1172 22.5005
R7240 GND.t866 GND.n1172 22.5005
R7241 GND.n1497 GND.n1169 22.5005
R7242 GND.t638 GND.n1169 22.5005
R7243 GND.n1457 GND.n1168 22.5005
R7244 GND.t638 GND.n1168 22.5005
R7245 GND.n854 GND.n852 22.5005
R7246 GND.t767 GND.n852 22.5005
R7247 GND.n853 GND.n851 22.5005
R7248 GND.t767 GND.n851 22.5005
R7249 GND.n3399 GND.n403 22.5005
R7250 GND.n3399 GND.t441 22.5005
R7251 GND.n405 GND.n404 22.5005
R7252 GND.t441 GND.n405 22.5005
R7253 GND.n400 GND.n397 22.5005
R7254 GND.t182 GND.n400 22.5005
R7255 GND.n399 GND.n398 22.5005
R7256 GND.t182 GND.n399 22.5005
R7257 GND.n385 GND.n383 22.5005
R7258 GND.t745 GND.n383 22.5005
R7259 GND.n384 GND.n382 22.5005
R7260 GND.t745 GND.n382 22.5005
R7261 GND.n477 GND.n428 22.5005
R7262 GND.t670 GND.n428 22.5005
R7263 GND.n443 GND.n427 22.5005
R7264 GND.t670 GND.n427 22.5005
R7265 GND.n470 GND.n432 22.5005
R7266 GND.n432 GND.t354 22.5005
R7267 GND.n448 GND.n431 22.5005
R7268 GND.n431 GND.t354 22.5005
R7269 GND.n380 GND.n378 22.5005
R7270 GND.t582 GND.n380 22.5005
R7271 GND.n379 GND.n377 22.5005
R7272 GND.t582 GND.n379 22.5005
R7273 GND.n3538 GND.n365 22.5005
R7274 GND.t26 GND.n365 22.5005
R7275 GND.n3456 GND.n364 22.5005
R7276 GND.t26 GND.n364 22.5005
R7277 GND.n3543 GND.n361 22.5005
R7278 GND.n3543 GND.t617 22.5005
R7279 GND.n362 GND.n360 22.5005
R7280 GND.t617 GND.n362 22.5005
R7281 GND.n3568 GND.n352 22.5005
R7282 GND.t197 GND.n352 22.5005
R7283 GND.n3550 GND.n351 22.5005
R7284 GND.t197 GND.n351 22.5005
R7285 GND.n3469 GND.n3467 22.5005
R7286 GND.t710 GND.n3467 22.5005
R7287 GND.n3468 GND.n3466 22.5005
R7288 GND.t710 GND.n3466 22.5005
R7289 GND.n349 GND.n346 22.5005
R7290 GND.t775 GND.n349 22.5005
R7291 GND.n348 GND.n347 22.5005
R7292 GND.t775 GND.n348 22.5005
R7293 GND.n375 GND.n373 22.5005
R7294 GND.t731 GND.n373 22.5005
R7295 GND.n374 GND.n372 22.5005
R7296 GND.t731 GND.n372 22.5005
R7297 GND.n3682 GND.n313 22.5005
R7298 GND.n3682 GND.t623 22.5005
R7299 GND.n315 GND.n314 22.5005
R7300 GND.t623 GND.n315 22.5005
R7301 GND.n310 GND.n307 22.5005
R7302 GND.t770 GND.n310 22.5005
R7303 GND.n309 GND.n308 22.5005
R7304 GND.t770 GND.n309 22.5005
R7305 GND.n295 GND.n293 22.5005
R7306 GND.t769 GND.n293 22.5005
R7307 GND.n294 GND.n292 22.5005
R7308 GND.t769 GND.n292 22.5005
R7309 GND.n3775 GND.n278 22.5005
R7310 GND.t258 GND.n278 22.5005
R7311 GND.n3730 GND.n291 22.5005
R7312 GND.n3730 GND.t258 22.5005
R7313 GND.n3769 GND.n282 22.5005
R7314 GND.t634 GND.n282 22.5005
R7315 GND.n3734 GND.n289 22.5005
R7316 GND.n3734 GND.t634 22.5005
R7317 GND.n270 GND.n268 22.5005
R7318 GND.t217 GND.n268 22.5005
R7319 GND.n269 GND.n267 22.5005
R7320 GND.t217 GND.n267 22.5005
R7321 GND.n3835 GND.n263 22.5005
R7322 GND.n3835 GND.t809 22.5005
R7323 GND.n265 GND.n264 22.5005
R7324 GND.t809 GND.n265 22.5005
R7325 GND.n260 GND.n257 22.5005
R7326 GND.t591 GND.n260 22.5005
R7327 GND.n259 GND.n258 22.5005
R7328 GND.t591 GND.n259 22.5005
R7329 GND.n245 GND.n243 22.5005
R7330 GND.t220 GND.n243 22.5005
R7331 GND.n244 GND.n242 22.5005
R7332 GND.t220 GND.n242 22.5005
R7333 GND.n3931 GND.n232 22.5005
R7334 GND.t759 GND.n232 22.5005
R7335 GND.n3887 GND.n239 22.5005
R7336 GND.n3887 GND.t759 22.5005
R7337 GND.n3901 GND.n3899 22.5005
R7338 GND.t71 GND.n3899 22.5005
R7339 GND.n3900 GND.n3898 22.5005
R7340 GND.t71 GND.n3898 22.5005
R7341 GND.n3937 GND.n228 22.5005
R7342 GND.t191 GND.n228 22.5005
R7343 GND.n3883 GND.n241 22.5005
R7344 GND.n3883 GND.t191 22.5005
R7345 GND.n4288 GND.n7 22.5005
R7346 GND.t190 GND.n7 22.5005
R7347 GND.n3175 GND.n3171 22.5005
R7348 GND.n3175 GND.t190 22.5005
R7349 GND.n22 GND.n20 22.5005
R7350 GND.t218 GND.n20 22.5005
R7351 GND.n21 GND.n19 22.5005
R7352 GND.t218 GND.n19 22.5005
R7353 GND.n4294 GND.n3 22.5005
R7354 GND.t611 GND.n3 22.5005
R7355 GND.n3179 GND.n3169 22.5005
R7356 GND.n3179 GND.t611 22.5005
R7357 GND.n3270 GND.n509 22.5005
R7358 GND.n3270 GND.t867 22.5005
R7359 GND.n511 GND.n510 22.5005
R7360 GND.t867 GND.n511 22.5005
R7361 GND.n506 GND.n503 22.5005
R7362 GND.t287 GND.n506 22.5005
R7363 GND.n505 GND.n504 22.5005
R7364 GND.t287 GND.n505 22.5005
R7365 GND.n3310 GND.n489 22.5005
R7366 GND.n3310 GND.t647 22.5005
R7367 GND.n491 GND.n490 22.5005
R7368 GND.t647 GND.n491 22.5005
R7369 GND.n3241 GND.n3215 22.5005
R7370 GND.t357 GND.n3215 22.5005
R7371 GND.n3224 GND.n3214 22.5005
R7372 GND.t357 GND.n3214 22.5005
R7373 GND.n3234 GND.n3219 22.5005
R7374 GND.n3219 GND.t756 22.5005
R7375 GND.n3221 GND.n3218 22.5005
R7376 GND.t756 GND.n3218 22.5005
R7377 GND.n3340 GND.n414 22.5005
R7378 GND.t707 GND.n414 22.5005
R7379 GND.n3322 GND.n413 22.5005
R7380 GND.t707 GND.n413 22.5005
R7381 GND.n1245 GND.n1224 22.5005
R7382 GND.n1224 GND.t211 22.5005
R7383 GND.n1226 GND.n1223 22.5005
R7384 GND.t211 GND.n1223 22.5005
R7385 GND.n1260 GND.n1215 22.5005
R7386 GND.t286 GND.n1215 22.5005
R7387 GND.n1234 GND.n1214 22.5005
R7388 GND.t286 GND.n1214 22.5005
R7389 GND.n1267 GND.n1211 22.5005
R7390 GND.t395 GND.n1211 22.5005
R7391 GND.n1229 GND.n1210 22.5005
R7392 GND.t395 GND.n1210 22.5005
R7393 GND.n2783 GND.n2464 22.5005
R7394 GND.t648 GND.n2464 22.5005
R7395 GND.n2497 GND.n2463 22.5005
R7396 GND.t648 GND.n2463 22.5005
R7397 GND.n2793 GND.n2792 22.5005
R7398 GND.n2792 GND.t434 22.5005
R7399 GND.n2791 GND.n2495 22.5005
R7400 GND.t434 GND.n2791 22.5005
R7401 GND.n2807 GND.n2806 22.5005
R7402 GND.t353 GND.n2807 22.5005
R7403 GND.n2825 GND.n2824 22.5005
R7404 GND.n2824 GND.t353 22.5005
R7405 GND.n2863 GND.n2862 22.5005
R7406 GND.n2862 GND.t648 22.5005
R7407 GND.n2861 GND.n2860 22.5005
R7408 GND.t648 GND.n2861 22.5005
R7409 GND.n2470 GND.n2468 22.5005
R7410 GND.t434 GND.n2468 22.5005
R7411 GND.n2469 GND.n2467 22.5005
R7412 GND.t434 GND.n2467 22.5005
R7413 GND.n2814 GND.n2808 22.5005
R7414 GND.t353 GND.n2808 22.5005
R7415 GND.n2823 GND.n2822 22.5005
R7416 GND.t353 GND.n2823 22.5005
R7417 GND.n2876 GND.n2875 22.5005
R7418 GND.n2876 GND.t438 22.5005
R7419 GND.n2874 GND.n2181 22.5005
R7420 GND.t438 GND.n2874 22.5005
R7421 GND.n2888 GND.n2887 22.5005
R7422 GND.n2888 GND.t465 22.5005
R7423 GND.n2886 GND.n2883 22.5005
R7424 GND.t465 GND.n2886 22.5005
R7425 GND.n2916 GND.n2914 22.5005
R7426 GND.n2916 GND.t365 22.5005
R7427 GND.n2915 GND.n2912 22.5005
R7428 GND.t365 GND.n2915 22.5005
R7429 GND.n2181 GND.n2178 22.5005
R7430 GND.t438 GND.n2178 22.5005
R7431 GND.n2179 GND.n2177 22.5005
R7432 GND.t438 GND.n2177 22.5005
R7433 GND.n2883 GND.n2880 22.5005
R7434 GND.t465 GND.n2880 22.5005
R7435 GND.n2881 GND.n2879 22.5005
R7436 GND.t465 GND.n2879 22.5005
R7437 GND.n2912 GND.n2909 22.5005
R7438 GND.t365 GND.n2909 22.5005
R7439 GND.n2910 GND.n2908 22.5005
R7440 GND.t365 GND.n2908 22.5005
R7441 GND.n2344 GND.n2343 22.5005
R7442 GND.n2344 GND.t95 22.5005
R7443 GND.n2342 GND.n2339 22.5005
R7444 GND.t95 GND.n2342 22.5005
R7445 GND.n2356 GND.n2355 22.5005
R7446 GND.n2356 GND.t713 22.5005
R7447 GND.n2354 GND.n2351 22.5005
R7448 GND.t713 GND.n2354 22.5005
R7449 GND.n2384 GND.n2382 22.5005
R7450 GND.n2384 GND.t350 22.5005
R7451 GND.n2383 GND.n2380 22.5005
R7452 GND.t350 GND.n2383 22.5005
R7453 GND.n2339 GND.n2336 22.5005
R7454 GND.t95 GND.n2336 22.5005
R7455 GND.n2337 GND.n2335 22.5005
R7456 GND.t95 GND.n2335 22.5005
R7457 GND.n2351 GND.n2348 22.5005
R7458 GND.t713 GND.n2348 22.5005
R7459 GND.n2349 GND.n2347 22.5005
R7460 GND.t713 GND.n2347 22.5005
R7461 GND.n2380 GND.n2377 22.5005
R7462 GND.t350 GND.n2377 22.5005
R7463 GND.n2378 GND.n2376 22.5005
R7464 GND.t350 GND.n2376 22.5005
R7465 GND.n2217 GND.n2216 22.5005
R7466 GND.n2217 GND.t383 22.5005
R7467 GND.n2215 GND.n2212 22.5005
R7468 GND.t383 GND.n2215 22.5005
R7469 GND.n2229 GND.n2228 22.5005
R7470 GND.n2229 GND.t87 22.5005
R7471 GND.n2227 GND.n2224 22.5005
R7472 GND.t87 GND.n2227 22.5005
R7473 GND.n2257 GND.n2255 22.5005
R7474 GND.n2257 GND.t55 22.5005
R7475 GND.n2256 GND.n2253 22.5005
R7476 GND.t55 GND.n2256 22.5005
R7477 GND.n2212 GND.n2209 22.5005
R7478 GND.t383 GND.n2209 22.5005
R7479 GND.n2210 GND.n2208 22.5005
R7480 GND.t383 GND.n2208 22.5005
R7481 GND.n2224 GND.n2221 22.5005
R7482 GND.t87 GND.n2221 22.5005
R7483 GND.n2222 GND.n2220 22.5005
R7484 GND.t87 GND.n2220 22.5005
R7485 GND.n2253 GND.n2250 22.5005
R7486 GND.t55 GND.n2250 22.5005
R7487 GND.n2251 GND.n2249 22.5005
R7488 GND.t55 GND.n2249 22.5005
R7489 GND.n2539 GND.n2538 22.5005
R7490 GND.n2539 GND.t437 22.5005
R7491 GND.n2537 GND.n2534 22.5005
R7492 GND.t437 GND.n2537 22.5005
R7493 GND.n2551 GND.n2550 22.5005
R7494 GND.n2551 GND.t711 22.5005
R7495 GND.n2549 GND.n2546 22.5005
R7496 GND.t711 GND.n2549 22.5005
R7497 GND.n2579 GND.n2577 22.5005
R7498 GND.n2579 GND.t725 22.5005
R7499 GND.n2578 GND.n2575 22.5005
R7500 GND.t725 GND.n2578 22.5005
R7501 GND.n2534 GND.n2531 22.5005
R7502 GND.t437 GND.n2531 22.5005
R7503 GND.n2532 GND.n2530 22.5005
R7504 GND.t437 GND.n2530 22.5005
R7505 GND.n2546 GND.n2543 22.5005
R7506 GND.t711 GND.n2543 22.5005
R7507 GND.n2544 GND.n2542 22.5005
R7508 GND.t711 GND.n2542 22.5005
R7509 GND.n2575 GND.n2572 22.5005
R7510 GND.t725 GND.n2572 22.5005
R7511 GND.n2573 GND.n2571 22.5005
R7512 GND.t725 GND.n2571 22.5005
R7513 GND.n2660 GND.n2659 22.5005
R7514 GND.n2660 GND.t633 22.5005
R7515 GND.n2658 GND.n2515 22.5005
R7516 GND.t633 GND.n2658 22.5005
R7517 GND.n2672 GND.n2671 22.5005
R7518 GND.n2672 GND.t75 22.5005
R7519 GND.n2670 GND.n2667 22.5005
R7520 GND.t75 GND.n2670 22.5005
R7521 GND.n2700 GND.n2698 22.5005
R7522 GND.n2700 GND.t470 22.5005
R7523 GND.n2699 GND.n2696 22.5005
R7524 GND.t470 GND.n2699 22.5005
R7525 GND.n2515 GND.n2512 22.5005
R7526 GND.t633 GND.n2512 22.5005
R7527 GND.n2513 GND.n2511 22.5005
R7528 GND.t633 GND.n2511 22.5005
R7529 GND.n2667 GND.n2664 22.5005
R7530 GND.t75 GND.n2664 22.5005
R7531 GND.n2665 GND.n2663 22.5005
R7532 GND.t75 GND.n2663 22.5005
R7533 GND.n2696 GND.n2693 22.5005
R7534 GND.t470 GND.n2693 22.5005
R7535 GND.n2694 GND.n2692 22.5005
R7536 GND.t470 GND.n2692 22.5005
R7537 GND.n3002 GND.n2164 22.5005
R7538 GND.t439 GND.n2164 22.5005
R7539 GND.n2195 GND.n2163 22.5005
R7540 GND.t439 GND.n2163 22.5005
R7541 GND.n3009 GND.n2160 22.5005
R7542 GND.t57 GND.n2160 22.5005
R7543 GND.n2190 GND.n2159 22.5005
R7544 GND.t57 GND.n2159 22.5005
R7545 GND.n3022 GND.n2151 22.5005
R7546 GND.n3022 GND.t442 22.5005
R7547 GND.n2152 GND.n2150 22.5005
R7548 GND.t442 GND.n2152 22.5005
R7549 GND.n644 GND.n642 22.5005
R7550 GND.t660 GND.n642 22.5005
R7551 GND.n643 GND.n641 22.5005
R7552 GND.t660 GND.n641 22.5005
R7553 GND.n2116 GND.n2115 22.5005
R7554 GND.n2115 GND.t774 22.5005
R7555 GND.n664 GND.n663 22.5005
R7556 GND.n663 GND.t774 22.5005
R7557 GND.n669 GND.n667 22.5005
R7558 GND.t345 GND.n667 22.5005
R7559 GND.n668 GND.n666 22.5005
R7560 GND.t345 GND.n666 22.5005
R7561 GND.n2096 GND.n676 22.5005
R7562 GND.t474 GND.n676 22.5005
R7563 GND.n1283 GND.n675 22.5005
R7564 GND.t474 GND.n675 22.5005
R7565 GND.n2082 GND.n686 22.5005
R7566 GND.t198 GND.n686 22.5005
R7567 GND.n1291 GND.n685 22.5005
R7568 GND.t198 GND.n685 22.5005
R7569 GND.n2075 GND.n690 22.5005
R7570 GND.t800 GND.n690 22.5005
R7571 GND.n1296 GND.n689 22.5005
R7572 GND.t800 GND.n689 22.5005
R7573 GND.n722 GND.n720 22.5005
R7574 GND.n720 GND.t730 22.5005
R7575 GND.n721 GND.n719 22.5005
R7576 GND.t730 GND.n719 22.5005
R7577 GND.n710 GND.n708 22.5005
R7578 GND.n708 GND.t635 22.5005
R7579 GND.n709 GND.n707 22.5005
R7580 GND.t635 GND.n707 22.5005
R7581 GND.n769 GND.n703 22.5005
R7582 GND.n769 GND.t433 22.5005
R7583 GND.n705 GND.n704 22.5005
R7584 GND.t433 GND.n705 22.5005
R7585 GND.n701 GND.n699 22.5005
R7586 GND.t440 GND.n699 22.5005
R7587 GND.n700 GND.n698 22.5005
R7588 GND.t440 GND.n698 22.5005
R7589 GND.n2033 GND.n2032 22.5005
R7590 GND.n2032 GND.t404 22.5005
R7591 GND.n795 GND.n794 22.5005
R7592 GND.n794 GND.t404 22.5005
R7593 GND.n800 GND.n798 22.5005
R7594 GND.t780 GND.n798 22.5005
R7595 GND.n799 GND.n797 22.5005
R7596 GND.t780 GND.n797 22.5005
R7597 GND.n2013 GND.n807 22.5005
R7598 GND.t38 GND.n807 22.5005
R7599 GND.n1434 GND.n806 22.5005
R7600 GND.t38 GND.n806 22.5005
R7601 GND.n1999 GND.n817 22.5005
R7602 GND.t321 GND.n817 22.5005
R7603 GND.n1442 GND.n816 22.5005
R7604 GND.t321 GND.n816 22.5005
R7605 GND.n1992 GND.n821 22.5005
R7606 GND.t692 GND.n821 22.5005
R7607 GND.n1447 GND.n820 22.5005
R7608 GND.t692 GND.n820 22.5005
R7609 GND.n1428 GND.n1427 22.5005
R7610 GND.n1427 GND.t221 22.5005
R7611 GND.n1426 GND.n1425 22.5005
R7612 GND.t221 GND.n1426 22.5005
R7613 GND.n1404 GND.n1403 22.5005
R7614 GND.n1403 GND.t56 22.5005
R7615 GND.n1402 GND.n1401 22.5005
R7616 GND.t56 GND.n1402 22.5005
R7617 GND.n1385 GND.n1383 22.5005
R7618 GND.n1383 GND.t472 22.5005
R7619 GND.n1384 GND.n1382 22.5005
R7620 GND.t472 GND.n1382 22.5005
R7621 GND.n832 GND.n830 22.5005
R7622 GND.n830 GND.t604 22.5005
R7623 GND.n831 GND.n829 22.5005
R7624 GND.t604 GND.n829 22.5005
R7625 GND.n1770 GND.n1768 22.5005
R7626 GND.t206 GND.n1770 22.5005
R7627 GND.n1769 GND.n1767 22.5005
R7628 GND.t206 GND.n1769 22.5005
R7629 GND.n1800 GND.n1798 22.5005
R7630 GND.t318 GND.n1800 22.5005
R7631 GND.n1799 GND.n1797 22.5005
R7632 GND.t318 GND.n1799 22.5005
R7633 GND.n1830 GND.n1828 22.5005
R7634 GND.t49 GND.n1830 22.5005
R7635 GND.n1829 GND.n1827 22.5005
R7636 GND.t49 GND.n1829 22.5005
R7637 GND.n1845 GND.n1843 22.5005
R7638 GND.t779 GND.n1845 22.5005
R7639 GND.n1844 GND.n1842 22.5005
R7640 GND.t779 GND.n1844 22.5005
R7641 GND.n1815 GND.n1813 22.5005
R7642 GND.t876 GND.n1815 22.5005
R7643 GND.n1814 GND.n1812 22.5005
R7644 GND.t876 GND.n1814 22.5005
R7645 GND.n1785 GND.n1783 22.5005
R7646 GND.t703 GND.n1785 22.5005
R7647 GND.n1784 GND.n1782 22.5005
R7648 GND.t703 GND.n1784 22.5005
R7649 GND.n1950 GND.n1949 22.5005
R7650 GND.n1949 GND.t685 22.5005
R7651 GND.n1948 GND.n1947 22.5005
R7652 GND.t685 GND.n1948 22.5005
R7653 GND.n1762 GND.n1759 22.5005
R7654 GND.t678 GND.n1759 22.5005
R7655 GND.n1942 GND.n1760 22.5005
R7656 GND.t678 GND.n1760 22.5005
R7657 GND.n1910 GND.n1908 22.5005
R7658 GND.n1910 GND.t377 22.5005
R7659 GND.n4169 GND.n94 22.5005
R7660 GND.t377 GND.n94 22.5005
R7661 GND.n1917 GND.n1916 22.5005
R7662 GND.n1916 GND.t696 22.5005
R7663 GND.n1915 GND.n1914 22.5005
R7664 GND.t696 GND.n1915 22.5005
R7665 GND.n590 GND.n589 22.5005
R7666 GND.n590 GND.t699 22.5005
R7667 GND.n588 GND.n585 22.5005
R7668 GND.t699 GND.n588 22.5005
R7669 GND.n602 GND.n601 22.5005
R7670 GND.n602 GND.t255 22.5005
R7671 GND.n600 GND.n597 22.5005
R7672 GND.t255 GND.n600 22.5005
R7673 GND.n631 GND.n630 22.5005
R7674 GND.n631 GND.t462 22.5005
R7675 GND.n629 GND.n626 22.5005
R7676 GND.t462 GND.n629 22.5005
R7677 GND.n585 GND.n582 22.5005
R7678 GND.t699 GND.n582 22.5005
R7679 GND.n583 GND.n581 22.5005
R7680 GND.t699 GND.n581 22.5005
R7681 GND.n597 GND.n594 22.5005
R7682 GND.t255 GND.n594 22.5005
R7683 GND.n595 GND.n593 22.5005
R7684 GND.t255 GND.n593 22.5005
R7685 GND.n626 GND.n623 22.5005
R7686 GND.t462 GND.n623 22.5005
R7687 GND.n624 GND.n622 22.5005
R7688 GND.t462 GND.n622 22.5005
R7689 GND.n3122 GND.n572 22.5005
R7690 GND.n3122 GND.t865 22.5005
R7691 GND.n574 GND.n573 22.5005
R7692 GND.t865 GND.n574 22.5005
R7693 GND.n569 GND.n566 22.5005
R7694 GND.t89 GND.n569 22.5005
R7695 GND.n568 GND.n567 22.5005
R7696 GND.t89 GND.n568 22.5005
R7697 GND.n554 GND.n552 22.5005
R7698 GND.t687 GND.n552 22.5005
R7699 GND.n553 GND.n551 22.5005
R7700 GND.t687 GND.n551 22.5005
R7701 GND.n3191 GND.n538 22.5005
R7702 GND.n3191 GND.t654 22.5005
R7703 GND.n539 GND.n537 22.5005
R7704 GND.t654 GND.n539 22.5005
R7705 GND.n4239 GND.n35 22.5005
R7706 GND.t610 GND.n35 22.5005
R7707 GND.n3198 GND.n34 22.5005
R7708 GND.t610 GND.n34 22.5005
R7709 GND.n4254 GND.n26 22.5005
R7710 GND.t361 GND.n26 22.5005
R7711 GND.n3206 GND.n25 22.5005
R7712 GND.t361 GND.n25 22.5005
R7713 GND.n88 GND.n83 22.5005
R7714 GND.t80 GND.n83 22.5005
R7715 GND.n4176 GND.n4175 22.5005
R7716 GND.t80 GND.n4176 22.5005
R7717 GND.n3599 GND.n338 22.5005
R7718 GND.n3599 GND.t755 22.5005
R7719 GND.n340 GND.n339 22.5005
R7720 GND.t755 GND.n340 22.5005
R7721 GND.n335 GND.n332 22.5005
R7722 GND.t733 GND.n335 22.5005
R7723 GND.n334 GND.n333 22.5005
R7724 GND.t733 GND.n334 22.5005
R7725 GND.n320 GND.n318 22.5005
R7726 GND.t94 GND.n318 22.5005
R7727 GND.n319 GND.n317 22.5005
R7728 GND.t94 GND.n317 22.5005
R7729 GND.n4156 GND.n106 22.5005
R7730 GND.t643 GND.n106 22.5005
R7731 GND.n3646 GND.n105 22.5005
R7732 GND.t643 GND.n105 22.5005
R7733 GND.n4127 GND.n123 22.5005
R7734 GND.t662 GND.n123 22.5005
R7735 GND.n3663 GND.n122 22.5005
R7736 GND.t662 GND.n122 22.5005
R7737 GND.n4120 GND.n127 22.5005
R7738 GND.t36 GND.n127 22.5005
R7739 GND.n3658 GND.n126 22.5005
R7740 GND.t36 GND.n126 22.5005
R7741 GND.n4106 GND.n138 22.5005
R7742 GND.t880 GND.n138 22.5005
R7743 GND.n3650 GND.n137 22.5005
R7744 GND.t880 GND.n137 22.5005
R7745 GND.n4082 GND.n151 22.5005
R7746 GND.t98 GND.n151 22.5005
R7747 GND.n3786 GND.n150 22.5005
R7748 GND.t98 GND.n150 22.5005
R7749 GND.n4075 GND.n155 22.5005
R7750 GND.t408 GND.n155 22.5005
R7751 GND.n3791 GND.n154 22.5005
R7752 GND.t408 GND.n154 22.5005
R7753 GND.n4061 GND.n165 22.5005
R7754 GND.t734 GND.n165 22.5005
R7755 GND.n3799 GND.n164 22.5005
R7756 GND.t734 GND.n164 22.5005
R7757 GND.n4032 GND.n181 22.5005
R7758 GND.t855 GND.n181 22.5005
R7759 GND.n3816 GND.n180 22.5005
R7760 GND.t855 GND.n180 22.5005
R7761 GND.n4025 GND.n185 22.5005
R7762 GND.t839 GND.n185 22.5005
R7763 GND.n3811 GND.n184 22.5005
R7764 GND.t839 GND.n184 22.5005
R7765 GND.n4011 GND.n196 22.5005
R7766 GND.t352 GND.n196 22.5005
R7767 GND.n3803 GND.n195 22.5005
R7768 GND.t352 GND.n195 22.5005
R7769 GND.n3987 GND.n209 22.5005
R7770 GND.t291 GND.n209 22.5005
R7771 GND.n3948 GND.n208 22.5005
R7772 GND.t291 GND.n208 22.5005
R7773 GND.n3980 GND.n213 22.5005
R7774 GND.t45 GND.n213 22.5005
R7775 GND.n3953 GND.n212 22.5005
R7776 GND.t45 GND.n212 22.5005
R7777 GND.n3966 GND.n223 22.5005
R7778 GND.t473 GND.n223 22.5005
R7779 GND.n225 GND.n222 22.5005
R7780 GND.t473 GND.n222 22.5005
R7781 GND.t678 GND.t768 20.1796
R7782 GND.t685 GND.t230 20.1796
R7783 GND.n1925 GND 19.5277
R7784 GND GND.n1927 19.2885
R7785 GND.n1594 GND.n1592 19.1913
R7786 GND.n3035 GND.n3034 19.1913
R7787 GND.n60 GND.n59 19.1913
R7788 GND.n81 GND.n80 19.1913
R7789 GND.n968 GND.n913 18.6076
R7790 GND.n1704 GND.n1703 18.6076
R7791 GND.n1510 GND.n863 18.6076
R7792 GND.n1454 GND.n833 18.6076
R7793 GND.n1432 GND.n1431 18.6076
R7794 GND.n1303 GND.n775 18.6076
R7795 GND.n3942 GND.n3941 18.6076
R7796 GND.n3824 GND.n3823 18.6076
R7797 GND.n3780 GND.n3779 18.6076
R7798 GND.n3671 GND.n3670 18.6076
R7799 GND.n3583 GND.n3582 18.6076
R7800 GND.n3464 GND.n3463 18.6076
R7801 GND.n3320 GND.n3319 18.6076
R7802 GND.n3257 GND.n3256 18.6076
R7803 GND.n1920 GND.n113 17.3253
R7804 GND.n2501 GND 17.1782
R7805 GND.n2869 GND 17.1782
R7806 GND.n2455 GND 17.1782
R7807 GND.n2328 GND 17.1782
R7808 GND.n2650 GND 17.1782
R7809 GND.n2653 GND 17.1782
R7810 GND.n2201 GND 17.1782
R7811 GND.n2522 GND 17.1782
R7812 GND.n3943 GND 17.1782
R7813 GND.n3822 GND 17.1782
R7814 GND.n3781 GND 17.1782
R7815 GND.n3669 GND 17.1782
R7816 GND.n3584 GND 17.1782
R7817 GND.n3462 GND 17.1782
R7818 GND.n487 GND 17.1782
R7819 GND.n3251 GND 17.1782
R7820 GND.n543 GND 17.1782
R7821 GND.n4148 GND.n113 15.8782
R7822 GND.n3055 GND.n3054 13.8976
R7823 GND.n3060 GND.n3059 13.8976
R7824 GND.n3070 GND.n612 13.8976
R7825 GND.n3071 GND.n3070 13.8976
R7826 GND.n3079 GND.n610 13.8976
R7827 GND.n3079 GND.n3078 13.8976
R7828 GND.n3091 GND.n3090 13.8976
R7829 GND.n3096 GND.n3095 13.8976
R7830 GND.n3104 GND.n3103 13.8976
R7831 GND.n3109 GND.n3108 13.8976
R7832 GND.n2922 GND.n2921 13.8976
R7833 GND.n2927 GND.n2926 13.8976
R7834 GND.n2937 GND.n2898 13.8976
R7835 GND.n2938 GND.n2937 13.8976
R7836 GND.n2946 GND.n2896 13.8976
R7837 GND.n2946 GND.n2945 13.8976
R7838 GND.n2958 GND.n2957 13.8976
R7839 GND.n2963 GND.n2962 13.8976
R7840 GND.n2971 GND.n2970 13.8976
R7841 GND.n2976 GND.n2975 13.8976
R7842 GND.n2390 GND.n2389 13.8976
R7843 GND.n2395 GND.n2394 13.8976
R7844 GND.n2405 GND.n2366 13.8976
R7845 GND.n2406 GND.n2405 13.8976
R7846 GND.n2414 GND.n2364 13.8976
R7847 GND.n2414 GND.n2413 13.8976
R7848 GND.n2426 GND.n2425 13.8976
R7849 GND.n2431 GND.n2430 13.8976
R7850 GND.n2439 GND.n2438 13.8976
R7851 GND.n2444 GND.n2443 13.8976
R7852 GND.n2263 GND.n2262 13.8976
R7853 GND.n2268 GND.n2267 13.8976
R7854 GND.n2278 GND.n2239 13.8976
R7855 GND.n2279 GND.n2278 13.8976
R7856 GND.n2287 GND.n2237 13.8976
R7857 GND.n2287 GND.n2286 13.8976
R7858 GND.n2299 GND.n2298 13.8976
R7859 GND.n2304 GND.n2303 13.8976
R7860 GND.n2312 GND.n2311 13.8976
R7861 GND.n2317 GND.n2316 13.8976
R7862 GND.n2585 GND.n2584 13.8976
R7863 GND.n2590 GND.n2589 13.8976
R7864 GND.n2600 GND.n2561 13.8976
R7865 GND.n2601 GND.n2600 13.8976
R7866 GND.n2609 GND.n2559 13.8976
R7867 GND.n2609 GND.n2608 13.8976
R7868 GND.n2621 GND.n2620 13.8976
R7869 GND.n2626 GND.n2625 13.8976
R7870 GND.n2634 GND.n2633 13.8976
R7871 GND.n2639 GND.n2638 13.8976
R7872 GND.n2706 GND.n2705 13.8976
R7873 GND.n2711 GND.n2710 13.8976
R7874 GND.n2721 GND.n2682 13.8976
R7875 GND.n2722 GND.n2721 13.8976
R7876 GND.n2730 GND.n2680 13.8976
R7877 GND.n2730 GND.n2729 13.8976
R7878 GND.n2742 GND.n2741 13.8976
R7879 GND.n2747 GND.n2746 13.8976
R7880 GND.n2755 GND.n2754 13.8976
R7881 GND.n2760 GND.n2759 13.8976
R7882 GND.n2523 GND.n2519 13.2764
R7883 GND.n2329 GND.n2201 10.7601
R7884 GND.n1281 GND.n1280 10.6976
R7885 GND GND.n4297 10.5092
R7886 GND.n2867 GND.n2866 10.4893
R7887 GND GND.n113 10.3837
R7888 GND.n1923 GND 9.81028
R7889 GND.n1280 GND.n44 9.62522
R7890 GND GND.n1923 9.59289
R7891 GND GND.n1931 9.58202
R7892 GND GND.n1929 9.58202
R7893 GND GND.n1925 9.58202
R7894 GND GND.n1921 9.53583
R7895 GND GND.n1933 8.38365
R7896 GND.n1860 GND.n1765 8.32958
R7897 GND.n1898 GND.n1897 8.32958
R7898 GND.n3259 GND.n3258 8.16273
R7899 GND.n543 GND.n0 7.9965
R7900 GND.n2501 GND.n2457 7.973
R7901 GND.n2869 GND.n2868 7.973
R7902 GND.n2456 GND.n2455 7.973
R7903 GND.n2329 GND.n2328 7.973
R7904 GND.n2651 GND.n2650 7.973
R7905 GND.n2653 GND.n2652 7.973
R7906 GND.n2523 GND.n2522 7.973
R7907 GND.n1869 GND.n1781 7.9105
R7908 GND.n1874 GND.n1796 7.9105
R7909 GND.n1879 GND.n1811 7.9105
R7910 GND.n1884 GND.n1826 7.9105
R7911 GND.n1889 GND.n1841 7.9105
R7912 GND.n1864 GND.n1766 7.9105
R7913 GND.n3260 GND.n3259 7.9105
R7914 GND.n1280 GND.n1279 7.9105
R7915 GND.n2058 GND.n775 7.0005
R7916 GND.n1431 GND.n1430 7.0005
R7917 GND.n1975 GND.n833 7.0005
R7918 GND.n1739 GND.n863 7.0005
R7919 GND.n1704 GND.n883 7.0005
R7920 GND.n1663 GND.n913 7.0005
R7921 GND.n985 GND.n968 7.0005
R7922 GND.n1703 GND.n1702 7.0005
R7923 GND.n1530 GND.n1510 7.0005
R7924 GND.n1471 GND.n1454 7.0005
R7925 GND.n1433 GND.n1432 7.0005
R7926 GND.n1320 GND.n1303 7.0005
R7927 GND.n1282 GND.n1281 7.0005
R7928 GND.n3941 GND 5.98963
R7929 GND GND.n3824 5.98963
R7930 GND.n3779 GND 5.98963
R7931 GND GND.n3671 5.98963
R7932 GND.n3582 GND 5.98963
R7933 GND.n3464 GND 5.98963
R7934 GND.n3319 GND 5.98963
R7935 GND.n3256 GND 5.98963
R7936 GND.n3942 GND 5.98963
R7937 GND.n3823 GND 5.98963
R7938 GND.n3780 GND 5.98963
R7939 GND.n3670 GND 5.98963
R7940 GND.n3583 GND 5.98963
R7941 GND.n3463 GND 5.98963
R7942 GND GND.n3320 5.98963
R7943 GND.n1879 GND.n1878 4.47177
R7944 GND.n3258 GND 4.35376
R7945 GND.n1279 GND.n535 4.15267
R7946 GND GND.n978 3.03311
R7947 GND.n955 GND 3.03311
R7948 GND GND.n1523 3.03311
R7949 GND GND.n1464 3.03311
R7950 GND.n1441 GND 3.03311
R7951 GND GND.n1313 3.03311
R7952 GND.n1290 GND 3.03311
R7953 GND GND.n1236 3.03311
R7954 GND.n726 GND.n535 2.79941
R7955 GND.n2456 GND.n2329 2.7876
R7956 GND.n2868 GND.n2456 2.7876
R7957 GND.n2868 GND.n2867 2.7876
R7958 GND.n2652 GND.n2457 2.7876
R7959 GND.n2652 GND.n2651 2.7876
R7960 GND.n2651 GND.n2523 2.7876
R7961 GND.n4298 GND.n0 2.7406
R7962 GND.n4229 GND.n44 2.6816
R7963 GND.n3941 GND.n3940 2.5793
R7964 GND.n3824 GND.n275 2.5793
R7965 GND.n3779 GND.n3778 2.5793
R7966 GND.n3671 GND.n3643 2.5793
R7967 GND.n3582 GND.n3581 2.5793
R7968 GND.n3465 GND.n3464 2.5793
R7969 GND.n3319 GND.n3318 2.5793
R7970 GND.n3256 GND.n3255 2.5793
R7971 GND.n0 GND 2.49506
R7972 GND.n2797 GND 2.42713
R7973 GND GND.n2188 2.42713
R7974 GND.n3956 GND 2.42713
R7975 GND GND.n3809 2.42713
R7976 GND.n3794 GND 2.42713
R7977 GND GND.n3656 2.42713
R7978 GND GND.n4166 2.42713
R7979 GND.n3548 GND 2.42713
R7980 GND.n451 GND 2.42713
R7981 GND GND.n421 2.42713
R7982 GND.n3201 GND 2.42713
R7983 GND.n1859 GND 2.32659
R7984 GND.n1279 GND 2.17441
R7985 GND.n775 GND 2.17441
R7986 GND.n1431 GND 2.17441
R7987 GND GND.n833 2.17441
R7988 GND.n863 GND 2.17441
R7989 GND GND.n1704 2.17441
R7990 GND GND.n913 2.17441
R7991 GND.n524 GND.n523 2.15648
R7992 GND.n3045 GND 1.74454
R7993 GND.n2140 GND.n2139 1.71489
R7994 GND.n1242 GND.n1241 1.71489
R7995 GND.n1889 GND.n1888 1.67683
R7996 GND.n1884 GND.n1883 1.6737
R7997 GND.n1874 GND.n1873 1.6737
R7998 GND.n1869 GND.n1868 1.67363
R7999 GND.n4146 GND.n114 1.66898
R8000 GND.n4098 GND.n4097 1.66898
R8001 GND.n4051 GND.n172 1.66898
R8002 GND.n4003 GND.n4002 1.66898
R8003 GND.n3392 GND.n3350 1.66898
R8004 GND.n3381 GND.n3380 1.66898
R8005 GND.n3375 GND.n3363 1.66898
R8006 GND.n3939 GND.n226 1.66898
R8007 GND.n3935 GND.n226 1.66898
R8008 GND.n3933 GND.n230 1.66898
R8009 GND.n3929 GND.n230 1.66898
R8010 GND.n3918 GND.n3917 1.66898
R8011 GND.n3908 GND.n3907 1.66898
R8012 GND.n3907 GND.n3906 1.66898
R8013 GND.n274 GND.n262 1.66898
R8014 GND.n3839 GND.n262 1.66898
R8015 GND.n3841 GND.n256 1.66898
R8016 GND.n3852 GND.n256 1.66898
R8017 GND.n3865 GND.n3864 1.66898
R8018 GND.n3875 GND.n3874 1.66898
R8019 GND.n3876 GND.n3875 1.66898
R8020 GND.n3777 GND.n276 1.66898
R8021 GND.n3773 GND.n276 1.66898
R8022 GND.n3771 GND.n280 1.66898
R8023 GND.n3767 GND.n280 1.66898
R8024 GND.n3756 GND.n3755 1.66898
R8025 GND.n3746 GND.n271 1.66898
R8026 GND.n3825 GND.n271 1.66898
R8027 GND.n3642 GND.n312 1.66898
R8028 GND.n3686 GND.n312 1.66898
R8029 GND.n3688 GND.n306 1.66898
R8030 GND.n3699 GND.n306 1.66898
R8031 GND.n3712 GND.n3711 1.66898
R8032 GND.n3722 GND.n3721 1.66898
R8033 GND.n3723 GND.n3722 1.66898
R8034 GND.n3580 GND.n337 1.66898
R8035 GND.n3603 GND.n337 1.66898
R8036 GND.n3605 GND.n331 1.66898
R8037 GND.n3616 GND.n331 1.66898
R8038 GND.n3629 GND.n3628 1.66898
R8039 GND.n3639 GND.n3638 1.66898
R8040 GND.n3672 GND.n3639 1.66898
R8041 GND.n3522 GND.n3521 1.66898
R8042 GND.n3521 GND.n3520 1.66898
R8043 GND.n3511 GND.n3510 1.66898
R8044 GND.n3510 GND.n3509 1.66898
R8045 GND.n3498 GND.n3476 1.66898
R8046 GND.n3485 GND.n345 1.66898
R8047 GND.n3577 GND.n345 1.66898
R8048 GND.n3317 GND.n402 1.66898
R8049 GND.n3403 GND.n402 1.66898
R8050 GND.n3405 GND.n396 1.66898
R8051 GND.n3416 GND.n396 1.66898
R8052 GND.n3429 GND.n3428 1.66898
R8053 GND.n3439 GND.n3438 1.66898
R8054 GND.n3440 GND.n3439 1.66898
R8055 GND.n4296 GND.n1 1.66898
R8056 GND.n4292 GND.n1 1.66898
R8057 GND.n4290 GND.n5 1.66898
R8058 GND.n4286 GND.n5 1.66898
R8059 GND.n4275 GND.n4274 1.66898
R8060 GND.n4265 GND.n4264 1.66898
R8061 GND.n4264 GND.n4263 1.66898
R8062 GND.n3254 GND.n508 1.66898
R8063 GND.n3274 GND.n508 1.66898
R8064 GND.n3276 GND.n502 1.66898
R8065 GND.n3287 GND.n502 1.66898
R8066 GND.n3304 GND.n3299 1.66898
R8067 GND.n3302 GND.n488 1.66898
R8068 GND.n3314 GND.n488 1.66898
R8069 GND.n2130 GND.n2129 1.66898
R8070 GND.n2118 GND.n656 1.66898
R8071 GND.n670 GND.n656 1.66898
R8072 GND.n2108 GND.n2107 1.66898
R8073 GND.n2107 GND.n2106 1.66898
R8074 GND.n727 GND.n726 1.66898
R8075 GND.n729 GND.n727 1.66898
R8076 GND.n741 GND.n739 1.66898
R8077 GND.n758 GND.n757 1.66898
R8078 GND.n763 GND.n758 1.66898
R8079 GND.n761 GND.n702 1.66898
R8080 GND.n773 GND.n702 1.66898
R8081 GND.n2058 GND.n2057 1.66898
R8082 GND.n2057 GND.n2056 1.66898
R8083 GND.n2047 GND.n2046 1.66898
R8084 GND.n2035 GND.n787 1.66898
R8085 GND.n801 GND.n787 1.66898
R8086 GND.n2025 GND.n2024 1.66898
R8087 GND.n2024 GND.n2023 1.66898
R8088 GND.n1430 GND.n1358 1.66898
R8089 GND.n1367 GND.n1358 1.66898
R8090 GND.n1418 GND.n1417 1.66898
R8091 GND.n1406 GND.n1377 1.66898
R8092 GND.n1386 GND.n1377 1.66898
R8093 GND.n1394 GND.n1393 1.66898
R8094 GND.n1393 GND.n1392 1.66898
R8095 GND.n1975 GND.n1974 1.66898
R8096 GND.n1974 GND.n1973 1.66898
R8097 GND.n1964 GND.n1963 1.66898
R8098 GND.n1952 GND.n846 1.66898
R8099 GND.n855 GND.n846 1.66898
R8100 GND.n1751 GND.n1750 1.66898
R8101 GND.n1750 GND.n1749 1.66898
R8102 GND.n1739 GND.n1738 1.66898
R8103 GND.n1738 GND.n1737 1.66898
R8104 GND.n1728 GND.n1727 1.66898
R8105 GND.n1716 GND.n875 1.66898
R8106 GND.n1712 GND.n875 1.66898
R8107 GND.n1710 GND.n879 1.66898
R8108 GND.n1706 GND.n879 1.66898
R8109 GND.n1137 GND.n883 1.66898
R8110 GND.n1137 GND.n1136 1.66898
R8111 GND.n1134 GND.n1073 1.66898
R8112 GND.n1119 GND.n1087 1.66898
R8113 GND.n1115 GND.n1087 1.66898
R8114 GND.n1113 GND.n1091 1.66898
R8115 GND.n1109 GND.n1091 1.66898
R8116 GND.n1663 GND.n1662 1.66898
R8117 GND.n1662 GND.n1661 1.66898
R8118 GND.n1652 GND.n1651 1.66898
R8119 GND.n1640 GND.n925 1.66898
R8120 GND.n1636 GND.n925 1.66898
R8121 GND.n1634 GND.n929 1.66898
R8122 GND.n1630 GND.n929 1.66898
R8123 GND.n985 GND.n984 1.66898
R8124 GND.n984 GND.n983 1.66898
R8125 GND.n981 GND.n980 1.66898
R8126 GND.n978 GND.n977 1.66898
R8127 GND.n977 GND.n975 1.66898
R8128 GND.n973 GND.n972 1.66898
R8129 GND.n972 GND.n970 1.66898
R8130 GND.n1702 GND.n884 1.66898
R8131 GND.n1698 GND.n884 1.66898
R8132 GND.n1696 GND.n888 1.66898
R8133 GND.n957 GND.n955 1.66898
R8134 GND.n958 GND.n957 1.66898
R8135 GND.n962 GND.n960 1.66898
R8136 GND.n963 GND.n962 1.66898
R8137 GND.n1530 GND.n1529 1.66898
R8138 GND.n1529 GND.n1528 1.66898
R8139 GND.n1526 GND.n1525 1.66898
R8140 GND.n1523 GND.n1522 1.66898
R8141 GND.n1522 GND.n1520 1.66898
R8142 GND.n1518 GND.n1517 1.66898
R8143 GND.n1517 GND.n1515 1.66898
R8144 GND.n1471 GND.n1470 1.66898
R8145 GND.n1470 GND.n1469 1.66898
R8146 GND.n1467 GND.n1466 1.66898
R8147 GND.n1464 GND.n1463 1.66898
R8148 GND.n1463 GND.n1461 1.66898
R8149 GND.n1459 GND.n1458 1.66898
R8150 GND.n1458 GND.n1456 1.66898
R8151 GND.n1435 GND.n1433 1.66898
R8152 GND.n1436 GND.n1435 1.66898
R8153 GND.n1439 GND.n1438 1.66898
R8154 GND.n1443 GND.n1441 1.66898
R8155 GND.n1444 GND.n1443 1.66898
R8156 GND.n1448 GND.n1446 1.66898
R8157 GND.n1449 GND.n1448 1.66898
R8158 GND.n1320 GND.n1319 1.66898
R8159 GND.n1319 GND.n1318 1.66898
R8160 GND.n1316 GND.n1315 1.66898
R8161 GND.n1313 GND.n1312 1.66898
R8162 GND.n1312 GND.n1310 1.66898
R8163 GND.n1308 GND.n1307 1.66898
R8164 GND.n1307 GND.n1305 1.66898
R8165 GND.n1284 GND.n1282 1.66898
R8166 GND.n1285 GND.n1284 1.66898
R8167 GND.n1288 GND.n1287 1.66898
R8168 GND.n1292 GND.n1290 1.66898
R8169 GND.n1293 GND.n1292 1.66898
R8170 GND.n1297 GND.n1295 1.66898
R8171 GND.n1298 GND.n1297 1.66898
R8172 GND.n1239 GND.n1238 1.66898
R8173 GND.n1236 GND.n1235 1.66898
R8174 GND.n1235 GND.n1233 1.66898
R8175 GND.n1231 GND.n1230 1.66898
R8176 GND.n1230 GND.n1228 1.66898
R8177 GND.n2865 GND.n2458 1.66898
R8178 GND.n2471 GND.n2458 1.66898
R8179 GND.n2853 GND.n2852 1.66898
R8180 GND.n2852 GND.n2851 1.66898
R8181 GND.n2840 GND.n2479 1.66898
R8182 GND.n2818 GND.n2817 1.66898
R8183 GND.n2819 GND.n2818 1.66898
R8184 GND.n2503 GND.n2496 1.66898
R8185 GND.n2786 GND.n2496 1.66898
R8186 GND.n2788 GND.n2494 1.66898
R8187 GND.n2796 GND.n2494 1.66898
R8188 GND.n2829 GND.n2798 1.66898
R8189 GND.n2827 GND.n2799 1.66898
R8190 GND.n2801 GND.n2799 1.66898
R8191 GND.n2974 GND.n2973 1.66898
R8192 GND.n2973 GND.n2972 1.66898
R8193 GND.n2961 GND.n2960 1.66898
R8194 GND.n2960 GND.n2959 1.66898
R8195 GND.n2947 GND.n2895 1.66898
R8196 GND.n2925 GND.n2924 1.66898
R8197 GND.n2924 GND.n2923 1.66898
R8198 GND.n2442 GND.n2441 1.66898
R8199 GND.n2441 GND.n2440 1.66898
R8200 GND.n2429 GND.n2428 1.66898
R8201 GND.n2428 GND.n2427 1.66898
R8202 GND.n2415 GND.n2363 1.66898
R8203 GND.n2393 GND.n2392 1.66898
R8204 GND.n2392 GND.n2391 1.66898
R8205 GND.n2315 GND.n2314 1.66898
R8206 GND.n2314 GND.n2313 1.66898
R8207 GND.n2302 GND.n2301 1.66898
R8208 GND.n2301 GND.n2300 1.66898
R8209 GND.n2288 GND.n2236 1.66898
R8210 GND.n2266 GND.n2265 1.66898
R8211 GND.n2265 GND.n2264 1.66898
R8212 GND.n2637 GND.n2636 1.66898
R8213 GND.n2636 GND.n2635 1.66898
R8214 GND.n2624 GND.n2623 1.66898
R8215 GND.n2623 GND.n2622 1.66898
R8216 GND.n2610 GND.n2558 1.66898
R8217 GND.n2588 GND.n2587 1.66898
R8218 GND.n2587 GND.n2586 1.66898
R8219 GND.n2758 GND.n2757 1.66898
R8220 GND.n2757 GND.n2756 1.66898
R8221 GND.n2745 GND.n2744 1.66898
R8222 GND.n2744 GND.n2743 1.66898
R8223 GND.n2731 GND.n2679 1.66898
R8224 GND.n2709 GND.n2708 1.66898
R8225 GND.n2708 GND.n2707 1.66898
R8226 GND.n4229 GND.n4228 1.66898
R8227 GND.n4215 GND.n53 1.66898
R8228 GND.n4200 GND.n4199 1.66898
R8229 GND.n4186 GND.n74 1.66898
R8230 GND.n1585 GND.n1045 1.66898
R8231 GND.n1600 GND.n1598 1.66898
R8232 GND.n1614 GND.n1612 1.66898
R8233 GND.n3043 GND.n3028 1.66898
R8234 GND.n2197 GND.n2196 1.66898
R8235 GND.n2196 GND.n2194 1.66898
R8236 GND.n2192 GND.n2191 1.66898
R8237 GND.n2191 GND.n2189 1.66898
R8238 GND.n2187 GND.n2186 1.66898
R8239 GND.n2184 GND.n2149 1.66898
R8240 GND.n3026 GND.n2149 1.66898
R8241 GND.n2518 GND.n571 1.66898
R8242 GND.n3126 GND.n571 1.66898
R8243 GND.n3128 GND.n565 1.66898
R8244 GND.n3139 GND.n565 1.66898
R8245 GND.n3152 GND.n3151 1.66898
R8246 GND.n3162 GND.n3161 1.66898
R8247 GND.n3163 GND.n3162 1.66898
R8248 GND.n3107 GND.n3106 1.66898
R8249 GND.n3106 GND.n3105 1.66898
R8250 GND.n3094 GND.n3093 1.66898
R8251 GND.n3093 GND.n3092 1.66898
R8252 GND.n3080 GND.n609 1.66898
R8253 GND.n3058 GND.n3057 1.66898
R8254 GND.n3057 GND.n3056 1.66898
R8255 GND.n3949 GND.n3947 1.66898
R8256 GND.n3950 GND.n3949 1.66898
R8257 GND.n3954 GND.n3952 1.66898
R8258 GND.n3955 GND.n3954 1.66898
R8259 GND.n3958 GND.n3957 1.66898
R8260 GND.n3961 GND.n3960 1.66898
R8261 GND.n3962 GND.n3961 1.66898
R8262 GND.n3818 GND.n3817 1.66898
R8263 GND.n3817 GND.n3815 1.66898
R8264 GND.n3813 GND.n3812 1.66898
R8265 GND.n3812 GND.n3810 1.66898
R8266 GND.n3808 GND.n3807 1.66898
R8267 GND.n3805 GND.n3804 1.66898
R8268 GND.n3804 GND.n3802 1.66898
R8269 GND.n3787 GND.n3785 1.66898
R8270 GND.n3788 GND.n3787 1.66898
R8271 GND.n3792 GND.n3790 1.66898
R8272 GND.n3793 GND.n3792 1.66898
R8273 GND.n3796 GND.n3795 1.66898
R8274 GND.n3800 GND.n3798 1.66898
R8275 GND.n3801 GND.n3800 1.66898
R8276 GND.n3665 GND.n3664 1.66898
R8277 GND.n3664 GND.n3662 1.66898
R8278 GND.n3660 GND.n3659 1.66898
R8279 GND.n3659 GND.n3657 1.66898
R8280 GND.n3655 GND.n3654 1.66898
R8281 GND.n3652 GND.n3651 1.66898
R8282 GND.n3651 GND.n3649 1.66898
R8283 GND.n4174 GND.n91 1.66898
R8284 GND.n4174 GND.n4173 1.66898
R8285 GND.n4171 GND.n92 1.66898
R8286 GND.n4167 GND.n92 1.66898
R8287 GND.n4165 GND.n96 1.66898
R8288 GND.n3647 GND.n3645 1.66898
R8289 GND.n3648 GND.n3647 1.66898
R8290 GND.n3458 GND.n3457 1.66898
R8291 GND.n3457 GND.n3455 1.66898
R8292 GND.n3453 GND.n359 1.66898
R8293 GND.n3547 GND.n359 1.66898
R8294 GND.n3555 GND.n3554 1.66898
R8295 GND.n3552 GND.n3551 1.66898
R8296 GND.n3551 GND.n3549 1.66898
R8297 GND.n444 GND.n442 1.66898
R8298 GND.n445 GND.n444 1.66898
R8299 GND.n449 GND.n447 1.66898
R8300 GND.n450 GND.n449 1.66898
R8301 GND.n453 GND.n452 1.66898
R8302 GND.n455 GND.n376 1.66898
R8303 GND.n3450 GND.n376 1.66898
R8304 GND.n3225 GND.n3223 1.66898
R8305 GND.n3226 GND.n3225 1.66898
R8306 GND.n3229 GND.n3228 1.66898
R8307 GND.n3230 GND.n3229 1.66898
R8308 GND.n3327 GND.n3326 1.66898
R8309 GND.n3324 GND.n3323 1.66898
R8310 GND.n3323 GND.n3321 1.66898
R8311 GND.n547 GND.n536 1.66898
R8312 GND.n3195 GND.n536 1.66898
R8313 GND.n3199 GND.n3197 1.66898
R8314 GND.n3200 GND.n3199 1.66898
R8315 GND.n3203 GND.n3202 1.66898
R8316 GND.n3207 GND.n3205 1.66898
R8317 GND.n3208 GND.n3207 1.66898
R8318 GND.n534 GND 1.66083
R8319 GND.n2867 GND.n2457 1.65255
R8320 GND.n3258 GND.n3257 1.58746
R8321 GND.n1788 GND.n1787 1.5505
R8322 GND.n1803 GND.n1802 1.5505
R8323 GND.n1818 GND.n1817 1.5505
R8324 GND.n1833 GND.n1832 1.5505
R8325 GND.n1848 GND.n1847 1.5505
R8326 GND.n1773 GND.n1772 1.5505
R8327 GND.n4149 GND.n4148 1.5505
R8328 GND.n4146 GND.n4145 1.5505
R8329 GND.n116 GND.n114 1.5505
R8330 GND.n4099 GND.n4098 1.5505
R8331 GND.n4097 GND.n4096 1.5505
R8332 GND.n4054 GND.n4053 1.5505
R8333 GND.n4051 GND.n4050 1.5505
R8334 GND.n174 GND.n172 1.5505
R8335 GND.n4004 GND.n4003 1.5505
R8336 GND.n4002 GND.n4001 1.5505
R8337 GND.n3264 GND.n3263 1.5505
R8338 GND.n3350 GND.n3349 1.5505
R8339 GND.n3393 GND.n3392 1.5505
R8340 GND.n3390 GND.n3389 1.5505
R8341 GND.n3382 GND.n3381 1.5505
R8342 GND.n3380 GND.n3379 1.5505
R8343 GND.n3375 GND.n3374 1.5505
R8344 GND.n3365 GND.n3363 1.5505
R8345 GND.n3939 GND.n3938 1.5505
R8346 GND.n3937 GND.n226 1.5505
R8347 GND.n3936 GND.n3935 1.5505
R8348 GND.n3933 GND.n3932 1.5505
R8349 GND.n3931 GND.n230 1.5505
R8350 GND.n3930 GND.n3929 1.5505
R8351 GND.n3927 GND.n3926 1.5505
R8352 GND.n3919 GND.n3918 1.5505
R8353 GND.n3917 GND.n3916 1.5505
R8354 GND.n3909 GND.n3908 1.5505
R8355 GND.n3907 GND.n3901 1.5505
R8356 GND.n3906 GND.n3905 1.5505
R8357 GND.n274 GND.n273 1.5505
R8358 GND.n263 GND.n262 1.5505
R8359 GND.n3839 GND.n3838 1.5505
R8360 GND.n3842 GND.n3841 1.5505
R8361 GND.n257 GND.n256 1.5505
R8362 GND.n3852 GND.n3851 1.5505
R8363 GND.n3855 GND.n3854 1.5505
R8364 GND.n3864 GND.n3863 1.5505
R8365 GND.n3866 GND.n3865 1.5505
R8366 GND.n3874 GND.n3873 1.5505
R8367 GND.n3875 GND.n245 1.5505
R8368 GND.n3877 GND.n3876 1.5505
R8369 GND.n3777 GND.n3776 1.5505
R8370 GND.n3775 GND.n276 1.5505
R8371 GND.n3774 GND.n3773 1.5505
R8372 GND.n3771 GND.n3770 1.5505
R8373 GND.n3769 GND.n280 1.5505
R8374 GND.n3768 GND.n3767 1.5505
R8375 GND.n3765 GND.n3764 1.5505
R8376 GND.n3757 GND.n3756 1.5505
R8377 GND.n3755 GND.n3754 1.5505
R8378 GND.n3747 GND.n3746 1.5505
R8379 GND.n271 GND.n270 1.5505
R8380 GND.n3826 GND.n3825 1.5505
R8381 GND.n3642 GND.n3641 1.5505
R8382 GND.n313 GND.n312 1.5505
R8383 GND.n3686 GND.n3685 1.5505
R8384 GND.n3689 GND.n3688 1.5505
R8385 GND.n307 GND.n306 1.5505
R8386 GND.n3699 GND.n3698 1.5505
R8387 GND.n3702 GND.n3701 1.5505
R8388 GND.n3711 GND.n3710 1.5505
R8389 GND.n3713 GND.n3712 1.5505
R8390 GND.n3721 GND.n3720 1.5505
R8391 GND.n3722 GND.n295 1.5505
R8392 GND.n3724 GND.n3723 1.5505
R8393 GND.n3580 GND.n3579 1.5505
R8394 GND.n338 GND.n337 1.5505
R8395 GND.n3603 GND.n3602 1.5505
R8396 GND.n3606 GND.n3605 1.5505
R8397 GND.n332 GND.n331 1.5505
R8398 GND.n3616 GND.n3615 1.5505
R8399 GND.n3619 GND.n3618 1.5505
R8400 GND.n3628 GND.n3627 1.5505
R8401 GND.n3630 GND.n3629 1.5505
R8402 GND.n3638 GND.n3637 1.5505
R8403 GND.n3639 GND.n320 1.5505
R8404 GND.n3673 GND.n3672 1.5505
R8405 GND.n3523 GND.n3522 1.5505
R8406 GND.n3521 GND.n375 1.5505
R8407 GND.n3520 GND.n3519 1.5505
R8408 GND.n3512 GND.n3511 1.5505
R8409 GND.n3510 GND.n3469 1.5505
R8410 GND.n3509 GND.n3508 1.5505
R8411 GND.n3501 GND.n3500 1.5505
R8412 GND.n3498 GND.n3497 1.5505
R8413 GND.n3478 GND.n3476 1.5505
R8414 GND.n3486 GND.n3485 1.5505
R8415 GND.n346 GND.n345 1.5505
R8416 GND.n3577 GND.n3576 1.5505
R8417 GND.n3317 GND.n3316 1.5505
R8418 GND.n403 GND.n402 1.5505
R8419 GND.n3403 GND.n3402 1.5505
R8420 GND.n3406 GND.n3405 1.5505
R8421 GND.n397 GND.n396 1.5505
R8422 GND.n3416 GND.n3415 1.5505
R8423 GND.n3419 GND.n3418 1.5505
R8424 GND.n3428 GND.n3427 1.5505
R8425 GND.n3430 GND.n3429 1.5505
R8426 GND.n3438 GND.n3437 1.5505
R8427 GND.n3439 GND.n385 1.5505
R8428 GND.n3441 GND.n3440 1.5505
R8429 GND.n4296 GND.n4295 1.5505
R8430 GND.n4294 GND.n1 1.5505
R8431 GND.n4293 GND.n4292 1.5505
R8432 GND.n4290 GND.n4289 1.5505
R8433 GND.n4288 GND.n5 1.5505
R8434 GND.n4287 GND.n4286 1.5505
R8435 GND.n4284 GND.n4283 1.5505
R8436 GND.n4276 GND.n4275 1.5505
R8437 GND.n4274 GND.n4273 1.5505
R8438 GND.n4266 GND.n4265 1.5505
R8439 GND.n4264 GND.n22 1.5505
R8440 GND.n4263 GND.n4262 1.5505
R8441 GND.n3277 GND.n3276 1.5505
R8442 GND.n503 GND.n502 1.5505
R8443 GND.n3287 GND.n3286 1.5505
R8444 GND.n3290 GND.n3289 1.5505
R8445 GND.n3299 GND.n3298 1.5505
R8446 GND.n3305 GND.n3304 1.5505
R8447 GND.n3302 GND.n3301 1.5505
R8448 GND.n489 GND.n488 1.5505
R8449 GND.n3314 GND.n3313 1.5505
R8450 GND.n3254 GND.n3253 1.5505
R8451 GND.n509 GND.n508 1.5505
R8452 GND.n3274 GND.n3273 1.5505
R8453 GND.n533 GND.n532 1.5505
R8454 GND.n2139 GND.n2138 1.5505
R8455 GND.n2131 GND.n2130 1.5505
R8456 GND.n2129 GND.n2128 1.5505
R8457 GND.n2121 GND.n2120 1.5505
R8458 GND.n2118 GND.n2117 1.5505
R8459 GND.n2116 GND.n656 1.5505
R8460 GND.n670 GND.n658 1.5505
R8461 GND.n2109 GND.n2108 1.5505
R8462 GND.n2107 GND.n669 1.5505
R8463 GND.n2106 GND.n2105 1.5505
R8464 GND.n726 GND.n725 1.5505
R8465 GND.n727 GND.n722 1.5505
R8466 GND.n730 GND.n729 1.5505
R8467 GND.n739 GND.n738 1.5505
R8468 GND.n742 GND.n741 1.5505
R8469 GND.n752 GND.n751 1.5505
R8470 GND.n757 GND.n756 1.5505
R8471 GND.n758 GND.n710 1.5505
R8472 GND.n764 GND.n763 1.5505
R8473 GND.n761 GND.n760 1.5505
R8474 GND.n703 GND.n702 1.5505
R8475 GND.n773 GND.n772 1.5505
R8476 GND.n2059 GND.n2058 1.5505
R8477 GND.n2057 GND.n701 1.5505
R8478 GND.n2056 GND.n2055 1.5505
R8479 GND.n2048 GND.n2047 1.5505
R8480 GND.n2046 GND.n2045 1.5505
R8481 GND.n2038 GND.n2037 1.5505
R8482 GND.n2035 GND.n2034 1.5505
R8483 GND.n2033 GND.n787 1.5505
R8484 GND.n801 GND.n789 1.5505
R8485 GND.n2026 GND.n2025 1.5505
R8486 GND.n2024 GND.n800 1.5505
R8487 GND.n2023 GND.n2022 1.5505
R8488 GND.n1430 GND.n1429 1.5505
R8489 GND.n1428 GND.n1358 1.5505
R8490 GND.n1367 GND.n1360 1.5505
R8491 GND.n1419 GND.n1418 1.5505
R8492 GND.n1417 GND.n1416 1.5505
R8493 GND.n1409 GND.n1408 1.5505
R8494 GND.n1406 GND.n1405 1.5505
R8495 GND.n1404 GND.n1377 1.5505
R8496 GND.n1386 GND.n1379 1.5505
R8497 GND.n1395 GND.n1394 1.5505
R8498 GND.n1393 GND.n1385 1.5505
R8499 GND.n1392 GND.n1391 1.5505
R8500 GND.n1976 GND.n1975 1.5505
R8501 GND.n1974 GND.n832 1.5505
R8502 GND.n1973 GND.n1972 1.5505
R8503 GND.n1965 GND.n1964 1.5505
R8504 GND.n1963 GND.n1962 1.5505
R8505 GND.n1955 GND.n1954 1.5505
R8506 GND.n1952 GND.n1951 1.5505
R8507 GND.n1950 GND.n846 1.5505
R8508 GND.n855 GND.n848 1.5505
R8509 GND.n1752 GND.n1751 1.5505
R8510 GND.n1750 GND.n854 1.5505
R8511 GND.n1749 GND.n1748 1.5505
R8512 GND.n1740 GND.n1739 1.5505
R8513 GND.n1738 GND.n862 1.5505
R8514 GND.n1737 GND.n1736 1.5505
R8515 GND.n1729 GND.n1728 1.5505
R8516 GND.n1727 GND.n1726 1.5505
R8517 GND.n1719 GND.n1718 1.5505
R8518 GND.n1716 GND.n1715 1.5505
R8519 GND.n1714 GND.n875 1.5505
R8520 GND.n1713 GND.n1712 1.5505
R8521 GND.n1710 GND.n1709 1.5505
R8522 GND.n1708 GND.n879 1.5505
R8523 GND.n1707 GND.n1706 1.5505
R8524 GND.n1139 GND.n883 1.5505
R8525 GND.n1138 GND.n1137 1.5505
R8526 GND.n1136 GND.n1072 1.5505
R8527 GND.n1134 GND.n1133 1.5505
R8528 GND.n1075 GND.n1073 1.5505
R8529 GND.n1122 GND.n1121 1.5505
R8530 GND.n1119 GND.n1118 1.5505
R8531 GND.n1117 GND.n1087 1.5505
R8532 GND.n1116 GND.n1115 1.5505
R8533 GND.n1113 GND.n1112 1.5505
R8534 GND.n1111 GND.n1091 1.5505
R8535 GND.n1110 GND.n1109 1.5505
R8536 GND.n1664 GND.n1663 1.5505
R8537 GND.n1662 GND.n912 1.5505
R8538 GND.n1661 GND.n1660 1.5505
R8539 GND.n1653 GND.n1652 1.5505
R8540 GND.n1651 GND.n1650 1.5505
R8541 GND.n1643 GND.n1642 1.5505
R8542 GND.n1640 GND.n1639 1.5505
R8543 GND.n1638 GND.n925 1.5505
R8544 GND.n1637 GND.n1636 1.5505
R8545 GND.n1634 GND.n1633 1.5505
R8546 GND.n1632 GND.n929 1.5505
R8547 GND.n1631 GND.n1630 1.5505
R8548 GND.n986 GND.n985 1.5505
R8549 GND.n984 GND.n953 1.5505
R8550 GND.n983 GND.n952 1.5505
R8551 GND.n981 GND.n949 1.5505
R8552 GND.n980 GND.n947 1.5505
R8553 GND.n978 GND.n944 1.5505
R8554 GND.n977 GND.n976 1.5505
R8555 GND.n975 GND.n943 1.5505
R8556 GND.n973 GND.n940 1.5505
R8557 GND.n972 GND.n971 1.5505
R8558 GND.n970 GND.n939 1.5505
R8559 GND.n1626 GND.n1625 1.5505
R8560 GND.n1702 GND.n1701 1.5505
R8561 GND.n1700 GND.n884 1.5505
R8562 GND.n1699 GND.n1698 1.5505
R8563 GND.n1696 GND.n1695 1.5505
R8564 GND.n890 GND.n888 1.5505
R8565 GND.n955 GND.n898 1.5505
R8566 GND.n957 GND.n956 1.5505
R8567 GND.n958 GND.n899 1.5505
R8568 GND.n960 GND.n902 1.5505
R8569 GND.n962 GND.n961 1.5505
R8570 GND.n963 GND.n903 1.5505
R8571 GND.n965 GND.n906 1.5505
R8572 GND.n1531 GND.n1530 1.5505
R8573 GND.n1529 GND.n1163 1.5505
R8574 GND.n1528 GND.n1162 1.5505
R8575 GND.n1526 GND.n1159 1.5505
R8576 GND.n1525 GND.n1157 1.5505
R8577 GND.n1523 GND.n1154 1.5505
R8578 GND.n1522 GND.n1521 1.5505
R8579 GND.n1520 GND.n1153 1.5505
R8580 GND.n1518 GND.n1150 1.5505
R8581 GND.n1517 GND.n1516 1.5505
R8582 GND.n1515 GND.n1149 1.5505
R8583 GND.n1513 GND.n1146 1.5505
R8584 GND.n1472 GND.n1471 1.5505
R8585 GND.n1470 GND.n1184 1.5505
R8586 GND.n1469 GND.n1183 1.5505
R8587 GND.n1467 GND.n1180 1.5505
R8588 GND.n1466 GND.n1178 1.5505
R8589 GND.n1464 GND.n1175 1.5505
R8590 GND.n1463 GND.n1462 1.5505
R8591 GND.n1461 GND.n1174 1.5505
R8592 GND.n1459 GND.n1171 1.5505
R8593 GND.n1458 GND.n1457 1.5505
R8594 GND.n1456 GND.n1170 1.5505
R8595 GND.n1507 GND.n1506 1.5505
R8596 GND.n1433 GND.n808 1.5505
R8597 GND.n1435 GND.n1434 1.5505
R8598 GND.n1436 GND.n809 1.5505
R8599 GND.n1438 GND.n812 1.5505
R8600 GND.n1439 GND.n814 1.5505
R8601 GND.n1441 GND.n818 1.5505
R8602 GND.n1443 GND.n1442 1.5505
R8603 GND.n1444 GND.n819 1.5505
R8604 GND.n1446 GND.n822 1.5505
R8605 GND.n1448 GND.n1447 1.5505
R8606 GND.n1449 GND.n823 1.5505
R8607 GND.n1451 GND.n826 1.5505
R8608 GND.n1321 GND.n1320 1.5505
R8609 GND.n1319 GND.n1205 1.5505
R8610 GND.n1318 GND.n1204 1.5505
R8611 GND.n1316 GND.n1201 1.5505
R8612 GND.n1315 GND.n1199 1.5505
R8613 GND.n1313 GND.n1196 1.5505
R8614 GND.n1312 GND.n1311 1.5505
R8615 GND.n1310 GND.n1195 1.5505
R8616 GND.n1308 GND.n1192 1.5505
R8617 GND.n1307 GND.n1306 1.5505
R8618 GND.n1305 GND.n1191 1.5505
R8619 GND.n1355 GND.n1354 1.5505
R8620 GND.n1282 GND.n677 1.5505
R8621 GND.n1284 GND.n1283 1.5505
R8622 GND.n1285 GND.n678 1.5505
R8623 GND.n1287 GND.n681 1.5505
R8624 GND.n1288 GND.n683 1.5505
R8625 GND.n1290 GND.n687 1.5505
R8626 GND.n1292 GND.n1291 1.5505
R8627 GND.n1293 GND.n688 1.5505
R8628 GND.n1295 GND.n691 1.5505
R8629 GND.n1297 GND.n1296 1.5505
R8630 GND.n1298 GND.n692 1.5505
R8631 GND.n1300 GND.n695 1.5505
R8632 GND.n1239 GND.n1222 1.5505
R8633 GND.n1238 GND.n1220 1.5505
R8634 GND.n1236 GND.n1217 1.5505
R8635 GND.n1235 GND.n1234 1.5505
R8636 GND.n1233 GND.n1216 1.5505
R8637 GND.n1231 GND.n1213 1.5505
R8638 GND.n1230 GND.n1229 1.5505
R8639 GND.n1228 GND.n1212 1.5505
R8640 GND.n1276 GND.n1275 1.5505
R8641 GND.n1241 GND.n1225 1.5505
R8642 GND.n2854 GND.n2853 1.5505
R8643 GND.n2852 GND.n2470 1.5505
R8644 GND.n2851 GND.n2850 1.5505
R8645 GND.n2843 GND.n2842 1.5505
R8646 GND.n2840 GND.n2839 1.5505
R8647 GND.n2481 GND.n2479 1.5505
R8648 GND.n2817 GND.n2816 1.5505
R8649 GND.n2818 GND.n2814 1.5505
R8650 GND.n2820 GND.n2819 1.5505
R8651 GND.n2865 GND.n2864 1.5505
R8652 GND.n2863 GND.n2458 1.5505
R8653 GND.n2471 GND.n2460 1.5505
R8654 GND.n2503 GND.n2498 1.5505
R8655 GND.n2497 GND.n2496 1.5505
R8656 GND.n2786 GND.n2785 1.5505
R8657 GND.n2789 GND.n2788 1.5505
R8658 GND.n2495 GND.n2494 1.5505
R8659 GND.n2796 GND.n2795 1.5505
R8660 GND.n2798 GND.n2490 1.5505
R8661 GND.n2830 GND.n2829 1.5505
R8662 GND.n2827 GND.n2826 1.5505
R8663 GND.n2825 GND.n2799 1.5505
R8664 GND.n2802 GND.n2801 1.5505
R8665 GND.n2506 GND.n2505 1.5505
R8666 GND.n2975 GND.n2974 1.5505
R8667 GND.n2973 GND.n2181 1.5505
R8668 GND.n2972 GND.n2971 1.5505
R8669 GND.n2962 GND.n2961 1.5505
R8670 GND.n2960 GND.n2883 1.5505
R8671 GND.n2959 GND.n2958 1.5505
R8672 GND.n2950 GND.n2949 1.5505
R8673 GND.n2947 GND.n2946 1.5505
R8674 GND.n2937 GND.n2895 1.5505
R8675 GND.n2926 GND.n2925 1.5505
R8676 GND.n2924 GND.n2912 1.5505
R8677 GND.n2923 GND.n2922 1.5505
R8678 GND.n2871 GND.n2175 1.5505
R8679 GND.n2443 GND.n2442 1.5505
R8680 GND.n2441 GND.n2339 1.5505
R8681 GND.n2440 GND.n2439 1.5505
R8682 GND.n2430 GND.n2429 1.5505
R8683 GND.n2428 GND.n2351 1.5505
R8684 GND.n2427 GND.n2426 1.5505
R8685 GND.n2418 GND.n2417 1.5505
R8686 GND.n2415 GND.n2414 1.5505
R8687 GND.n2405 GND.n2363 1.5505
R8688 GND.n2394 GND.n2393 1.5505
R8689 GND.n2392 GND.n2380 1.5505
R8690 GND.n2391 GND.n2390 1.5505
R8691 GND.n2453 GND.n2452 1.5505
R8692 GND.n2316 GND.n2315 1.5505
R8693 GND.n2314 GND.n2212 1.5505
R8694 GND.n2313 GND.n2312 1.5505
R8695 GND.n2303 GND.n2302 1.5505
R8696 GND.n2301 GND.n2224 1.5505
R8697 GND.n2300 GND.n2299 1.5505
R8698 GND.n2291 GND.n2290 1.5505
R8699 GND.n2288 GND.n2287 1.5505
R8700 GND.n2278 GND.n2236 1.5505
R8701 GND.n2267 GND.n2266 1.5505
R8702 GND.n2265 GND.n2253 1.5505
R8703 GND.n2264 GND.n2263 1.5505
R8704 GND.n2326 GND.n2325 1.5505
R8705 GND.n2638 GND.n2637 1.5505
R8706 GND.n2636 GND.n2534 1.5505
R8707 GND.n2635 GND.n2634 1.5505
R8708 GND.n2625 GND.n2624 1.5505
R8709 GND.n2623 GND.n2546 1.5505
R8710 GND.n2622 GND.n2621 1.5505
R8711 GND.n2613 GND.n2612 1.5505
R8712 GND.n2610 GND.n2609 1.5505
R8713 GND.n2600 GND.n2558 1.5505
R8714 GND.n2589 GND.n2588 1.5505
R8715 GND.n2587 GND.n2575 1.5505
R8716 GND.n2586 GND.n2585 1.5505
R8717 GND.n2648 GND.n2647 1.5505
R8718 GND.n2759 GND.n2758 1.5505
R8719 GND.n2757 GND.n2515 1.5505
R8720 GND.n2756 GND.n2755 1.5505
R8721 GND.n2746 GND.n2745 1.5505
R8722 GND.n2744 GND.n2667 1.5505
R8723 GND.n2743 GND.n2742 1.5505
R8724 GND.n2734 GND.n2733 1.5505
R8725 GND.n2731 GND.n2730 1.5505
R8726 GND.n2721 GND.n2679 1.5505
R8727 GND.n2710 GND.n2709 1.5505
R8728 GND.n2708 GND.n2696 1.5505
R8729 GND.n2707 GND.n2706 1.5505
R8730 GND.n2655 GND.n2509 1.5505
R8731 GND.n1763 GND.n1761 1.5505
R8732 GND.n1919 GND.n1918 1.5505
R8733 GND.n1917 GND.n1858 1.5505
R8734 GND.n1901 GND.n1900 1.5505
R8735 GND.n4230 GND.n4229 1.5505
R8736 GND.n4228 GND.n4227 1.5505
R8737 GND.n4218 GND.n4217 1.5505
R8738 GND.n4215 GND.n4214 1.5505
R8739 GND.n55 GND.n53 1.5505
R8740 GND.n4201 GND.n4200 1.5505
R8741 GND.n4199 GND.n4198 1.5505
R8742 GND.n4189 GND.n4188 1.5505
R8743 GND.n4186 GND.n4185 1.5505
R8744 GND.n76 GND.n74 1.5505
R8745 GND.n1051 GND.n1045 1.5505
R8746 GND.n1585 GND.n1584 1.5505
R8747 GND.n1589 GND.n1588 1.5505
R8748 GND.n1598 GND.n1597 1.5505
R8749 GND.n1601 GND.n1600 1.5505
R8750 GND.n1612 GND.n1611 1.5505
R8751 GND.n1615 GND.n1614 1.5505
R8752 GND.n3046 GND.n3045 1.5505
R8753 GND.n3043 GND.n3042 1.5505
R8754 GND.n3030 GND.n3028 1.5505
R8755 GND.n2199 GND.n2169 1.5505
R8756 GND.n2197 GND.n2166 1.5505
R8757 GND.n2196 GND.n2195 1.5505
R8758 GND.n2194 GND.n2165 1.5505
R8759 GND.n2192 GND.n2162 1.5505
R8760 GND.n2191 GND.n2190 1.5505
R8761 GND.n2189 GND.n2161 1.5505
R8762 GND.n2187 GND.n2158 1.5505
R8763 GND.n2186 GND.n2156 1.5505
R8764 GND.n2184 GND.n2183 1.5505
R8765 GND.n2150 GND.n2149 1.5505
R8766 GND.n3026 GND.n3025 1.5505
R8767 GND.n2518 GND.n2517 1.5505
R8768 GND.n572 GND.n571 1.5505
R8769 GND.n3126 GND.n3125 1.5505
R8770 GND.n3129 GND.n3128 1.5505
R8771 GND.n566 GND.n565 1.5505
R8772 GND.n3139 GND.n3138 1.5505
R8773 GND.n3142 GND.n3141 1.5505
R8774 GND.n3151 GND.n3150 1.5505
R8775 GND.n3153 GND.n3152 1.5505
R8776 GND.n3161 GND.n3160 1.5505
R8777 GND.n3162 GND.n554 1.5505
R8778 GND.n3164 GND.n3163 1.5505
R8779 GND.n3108 GND.n3107 1.5505
R8780 GND.n3106 GND.n585 1.5505
R8781 GND.n3105 GND.n3104 1.5505
R8782 GND.n3095 GND.n3094 1.5505
R8783 GND.n3093 GND.n597 1.5505
R8784 GND.n3092 GND.n3091 1.5505
R8785 GND.n3083 GND.n3082 1.5505
R8786 GND.n3080 GND.n3079 1.5505
R8787 GND.n3070 GND.n609 1.5505
R8788 GND.n3059 GND.n3058 1.5505
R8789 GND.n3057 GND.n626 1.5505
R8790 GND.n3056 GND.n3055 1.5505
R8791 GND.n2520 GND.n579 1.5505
R8792 GND.n3945 GND.n207 1.5505
R8793 GND.n3947 GND.n210 1.5505
R8794 GND.n3949 GND.n3948 1.5505
R8795 GND.n3950 GND.n211 1.5505
R8796 GND.n3952 GND.n214 1.5505
R8797 GND.n3954 GND.n3953 1.5505
R8798 GND.n3955 GND.n215 1.5505
R8799 GND.n3957 GND.n218 1.5505
R8800 GND.n3958 GND.n220 1.5505
R8801 GND.n3960 GND.n224 1.5505
R8802 GND.n3961 GND.n225 1.5505
R8803 GND.n3963 GND.n3962 1.5505
R8804 GND.n3820 GND.n179 1.5505
R8805 GND.n3818 GND.n182 1.5505
R8806 GND.n3817 GND.n3816 1.5505
R8807 GND.n3815 GND.n183 1.5505
R8808 GND.n3813 GND.n186 1.5505
R8809 GND.n3812 GND.n3811 1.5505
R8810 GND.n3810 GND.n187 1.5505
R8811 GND.n3808 GND.n191 1.5505
R8812 GND.n3807 GND.n193 1.5505
R8813 GND.n3805 GND.n197 1.5505
R8814 GND.n3804 GND.n3803 1.5505
R8815 GND.n3802 GND.n198 1.5505
R8816 GND.n3783 GND.n149 1.5505
R8817 GND.n3785 GND.n152 1.5505
R8818 GND.n3787 GND.n3786 1.5505
R8819 GND.n3788 GND.n153 1.5505
R8820 GND.n3790 GND.n156 1.5505
R8821 GND.n3792 GND.n3791 1.5505
R8822 GND.n3793 GND.n157 1.5505
R8823 GND.n3795 GND.n160 1.5505
R8824 GND.n3796 GND.n162 1.5505
R8825 GND.n3798 GND.n166 1.5505
R8826 GND.n3800 GND.n3799 1.5505
R8827 GND.n3801 GND.n167 1.5505
R8828 GND.n3667 GND.n121 1.5505
R8829 GND.n3665 GND.n124 1.5505
R8830 GND.n3664 GND.n3663 1.5505
R8831 GND.n3662 GND.n125 1.5505
R8832 GND.n3660 GND.n128 1.5505
R8833 GND.n3659 GND.n3658 1.5505
R8834 GND.n3657 GND.n129 1.5505
R8835 GND.n3655 GND.n133 1.5505
R8836 GND.n3654 GND.n135 1.5505
R8837 GND.n3652 GND.n139 1.5505
R8838 GND.n3651 GND.n3650 1.5505
R8839 GND.n3649 GND.n140 1.5505
R8840 GND.n3588 GND.n3587 1.5505
R8841 GND.n91 GND.n86 1.5505
R8842 GND.n4175 GND.n4174 1.5505
R8843 GND.n4173 GND.n90 1.5505
R8844 GND.n4171 GND.n4170 1.5505
R8845 GND.n4169 GND.n92 1.5505
R8846 GND.n4168 GND.n4167 1.5505
R8847 GND.n4165 GND.n4164 1.5505
R8848 GND.n98 GND.n96 1.5505
R8849 GND.n3645 GND.n107 1.5505
R8850 GND.n3647 GND.n3646 1.5505
R8851 GND.n3648 GND.n108 1.5505
R8852 GND.n3460 GND.n370 1.5505
R8853 GND.n3458 GND.n367 1.5505
R8854 GND.n3457 GND.n3456 1.5505
R8855 GND.n3455 GND.n366 1.5505
R8856 GND.n3453 GND.n3452 1.5505
R8857 GND.n360 GND.n359 1.5505
R8858 GND.n3547 GND.n3546 1.5505
R8859 GND.n3556 GND.n3555 1.5505
R8860 GND.n3554 GND.n357 1.5505
R8861 GND.n3552 GND.n354 1.5505
R8862 GND.n3551 GND.n3550 1.5505
R8863 GND.n3549 GND.n353 1.5505
R8864 GND.n485 GND.n484 1.5505
R8865 GND.n442 GND.n429 1.5505
R8866 GND.n444 GND.n443 1.5505
R8867 GND.n445 GND.n430 1.5505
R8868 GND.n447 GND.n433 1.5505
R8869 GND.n449 GND.n448 1.5505
R8870 GND.n450 GND.n434 1.5505
R8871 GND.n452 GND.n437 1.5505
R8872 GND.n453 GND.n439 1.5505
R8873 GND.n456 GND.n455 1.5505
R8874 GND.n377 GND.n376 1.5505
R8875 GND.n3450 GND.n3449 1.5505
R8876 GND.n3249 GND.n3248 1.5505
R8877 GND.n3223 GND.n3216 1.5505
R8878 GND.n3225 GND.n3224 1.5505
R8879 GND.n3226 GND.n3217 1.5505
R8880 GND.n3228 GND.n3220 1.5505
R8881 GND.n3229 GND.n3221 1.5505
R8882 GND.n3231 GND.n3230 1.5505
R8883 GND.n3328 GND.n3327 1.5505
R8884 GND.n3326 GND.n419 1.5505
R8885 GND.n3324 GND.n416 1.5505
R8886 GND.n3323 GND.n3322 1.5505
R8887 GND.n3321 GND.n415 1.5505
R8888 GND.n550 GND.n549 1.5505
R8889 GND.n547 GND.n546 1.5505
R8890 GND.n537 GND.n536 1.5505
R8891 GND.n3195 GND.n3194 1.5505
R8892 GND.n3197 GND.n37 1.5505
R8893 GND.n3199 GND.n3198 1.5505
R8894 GND.n3200 GND.n36 1.5505
R8895 GND.n3202 GND.n33 1.5505
R8896 GND.n3203 GND.n31 1.5505
R8897 GND.n3205 GND.n28 1.5505
R8898 GND.n3207 GND.n3206 1.5505
R8899 GND.n3208 GND.n27 1.5505
R8900 GND.n1764 GND 1.54738
R8901 GND.n1786 GND 1.54738
R8902 GND.n1801 GND 1.54738
R8903 GND.n1816 GND 1.54738
R8904 GND.n1831 GND 1.54738
R8905 GND.n1846 GND 1.54738
R8906 GND.n1899 GND 1.54738
R8907 GND.n1771 GND 1.54738
R8908 GND.n1935 GND.n1762 1.50658
R8909 GND.n1780 GND.n1767 1.50658
R8910 GND.n1795 GND.n1782 1.50658
R8911 GND.n1810 GND.n1797 1.50658
R8912 GND.n1825 GND.n1812 1.50658
R8913 GND.n1840 GND.n1827 1.50658
R8914 GND.n1855 GND.n1842 1.50658
R8915 GND.n2140 GND.n644 1.48372
R8916 GND.n1242 GND.n1226 1.48372
R8917 GND.n1864 GND.n1863 1.32825
R8918 GND.n1764 GND.n1763 1.1418
R8919 GND.n1787 GND.n1786 1.1418
R8920 GND.n1802 GND.n1801 1.1418
R8921 GND.n1817 GND.n1816 1.1418
R8922 GND.n1832 GND.n1831 1.1418
R8923 GND.n1847 GND.n1846 1.1418
R8924 GND.n1900 GND.n1899 1.1418
R8925 GND.n1772 GND.n1771 1.1418
R8926 GND.n1920 GND.n1919 1.11191
R8927 GND.n3261 GND 1.06886
R8928 GND.n1858 GND.n1856 1.06843
R8929 GND.n534 GND.n533 1.01952
R8930 GND.n1763 GND 1.01137
R8931 GND.n1787 GND 1.01137
R8932 GND.n1802 GND 1.01137
R8933 GND.n1817 GND 1.01137
R8934 GND.n1832 GND 1.01137
R8935 GND.n1847 GND 1.01137
R8936 GND.n1900 GND 1.01137
R8937 GND.n1772 GND 1.01137
R8938 GND GND.n4146 1.01137
R8939 GND GND.n4051 1.01137
R8940 GND.n3381 GND 1.01137
R8941 GND.n3935 GND 1.01137
R8942 GND.n3929 GND 1.01137
R8943 GND.n3927 GND 1.01137
R8944 GND.n3917 GND 1.01137
R8945 GND.n3906 GND 1.01137
R8946 GND GND.n3839 1.01137
R8947 GND GND.n3852 1.01137
R8948 GND.n3854 GND 1.01137
R8949 GND.n3865 GND 1.01137
R8950 GND.n3876 GND 1.01137
R8951 GND.n3773 GND 1.01137
R8952 GND.n3767 GND 1.01137
R8953 GND.n3765 GND 1.01137
R8954 GND.n3755 GND 1.01137
R8955 GND.n3825 GND 1.01137
R8956 GND GND.n3686 1.01137
R8957 GND GND.n3699 1.01137
R8958 GND.n3701 GND 1.01137
R8959 GND.n3712 GND 1.01137
R8960 GND.n3723 GND 1.01137
R8961 GND GND.n3603 1.01137
R8962 GND GND.n3616 1.01137
R8963 GND.n3618 GND 1.01137
R8964 GND.n3629 GND 1.01137
R8965 GND.n3672 GND 1.01137
R8966 GND.n3520 GND 1.01137
R8967 GND.n3509 GND 1.01137
R8968 GND.n3500 GND 1.01137
R8969 GND GND.n3476 1.01137
R8970 GND GND.n3577 1.01137
R8971 GND GND.n3403 1.01137
R8972 GND GND.n3416 1.01137
R8973 GND.n3418 GND 1.01137
R8974 GND.n3429 GND 1.01137
R8975 GND.n3440 GND 1.01137
R8976 GND.n4292 GND 1.01137
R8977 GND.n4286 GND 1.01137
R8978 GND.n4284 GND 1.01137
R8979 GND.n4274 GND 1.01137
R8980 GND.n4263 GND 1.01137
R8981 GND GND.n3274 1.01137
R8982 GND GND.n3287 1.01137
R8983 GND.n3289 GND 1.01137
R8984 GND.n3304 GND 1.01137
R8985 GND GND.n3314 1.01137
R8986 GND.n533 GND 1.01137
R8987 GND.n2130 GND 1.01137
R8988 GND.n2120 GND 1.01137
R8989 GND GND.n2118 1.01137
R8990 GND.n2108 GND 1.01137
R8991 GND.n739 GND 1.01137
R8992 GND.n752 GND 1.01137
R8993 GND.n757 GND 1.01137
R8994 GND GND.n761 1.01137
R8995 GND.n2047 GND 1.01137
R8996 GND.n2037 GND 1.01137
R8997 GND GND.n2035 1.01137
R8998 GND.n2025 GND 1.01137
R8999 GND.n1418 GND 1.01137
R9000 GND.n1408 GND 1.01137
R9001 GND GND.n1406 1.01137
R9002 GND.n1394 GND 1.01137
R9003 GND.n1964 GND 1.01137
R9004 GND.n1954 GND 1.01137
R9005 GND GND.n1952 1.01137
R9006 GND.n1751 GND 1.01137
R9007 GND.n1728 GND 1.01137
R9008 GND.n1718 GND 1.01137
R9009 GND GND.n1716 1.01137
R9010 GND GND.n1710 1.01137
R9011 GND GND.n1134 1.01137
R9012 GND.n1121 GND 1.01137
R9013 GND GND.n1119 1.01137
R9014 GND GND.n1113 1.01137
R9015 GND.n1652 GND 1.01137
R9016 GND.n1642 GND 1.01137
R9017 GND GND.n1640 1.01137
R9018 GND GND.n1634 1.01137
R9019 GND GND.n981 1.01137
R9020 GND GND.n973 1.01137
R9021 GND.n1626 GND 1.01137
R9022 GND GND.n1696 1.01137
R9023 GND.n960 GND 1.01137
R9024 GND.n965 GND 1.01137
R9025 GND GND.n1526 1.01137
R9026 GND GND.n1518 1.01137
R9027 GND GND.n1513 1.01137
R9028 GND GND.n1467 1.01137
R9029 GND GND.n1459 1.01137
R9030 GND.n1507 GND 1.01137
R9031 GND.n1438 GND 1.01137
R9032 GND.n1446 GND 1.01137
R9033 GND.n1451 GND 1.01137
R9034 GND GND.n1316 1.01137
R9035 GND GND.n1308 1.01137
R9036 GND.n1355 GND 1.01137
R9037 GND.n1287 GND 1.01137
R9038 GND.n1295 GND 1.01137
R9039 GND.n1300 GND 1.01137
R9040 GND GND.n1239 1.01137
R9041 GND GND.n1231 1.01137
R9042 GND.n1276 GND 1.01137
R9043 GND GND.n2471 1.01137
R9044 GND.n2851 GND 1.01137
R9045 GND.n2842 GND 1.01137
R9046 GND GND.n2479 1.01137
R9047 GND.n2819 GND 1.01137
R9048 GND.n2505 GND 1.01137
R9049 GND GND.n2786 1.01137
R9050 GND GND.n2796 1.01137
R9051 GND.n2829 GND 1.01137
R9052 GND.n2801 GND 1.01137
R9053 GND GND.n2871 1.01137
R9054 GND.n2972 GND 1.01137
R9055 GND.n2959 GND 1.01137
R9056 GND.n2949 GND 1.01137
R9057 GND GND.n2895 1.01137
R9058 GND.n2923 GND 1.01137
R9059 GND.n2453 GND 1.01137
R9060 GND.n2440 GND 1.01137
R9061 GND.n2427 GND 1.01137
R9062 GND.n2417 GND 1.01137
R9063 GND GND.n2363 1.01137
R9064 GND.n2391 GND 1.01137
R9065 GND.n2326 GND 1.01137
R9066 GND.n2313 GND 1.01137
R9067 GND.n2300 GND 1.01137
R9068 GND.n2290 GND 1.01137
R9069 GND GND.n2236 1.01137
R9070 GND.n2264 GND 1.01137
R9071 GND.n2648 GND 1.01137
R9072 GND.n2635 GND 1.01137
R9073 GND.n2622 GND 1.01137
R9074 GND.n2612 GND 1.01137
R9075 GND GND.n2558 1.01137
R9076 GND.n2586 GND 1.01137
R9077 GND GND.n2655 1.01137
R9078 GND.n2756 GND 1.01137
R9079 GND.n2743 GND 1.01137
R9080 GND.n2733 GND 1.01137
R9081 GND GND.n2679 1.01137
R9082 GND.n2707 GND 1.01137
R9083 GND GND.n4215 1.01137
R9084 GND GND.n4186 1.01137
R9085 GND.n1598 GND 1.01137
R9086 GND GND.n3043 1.01137
R9087 GND.n2199 GND 1.01137
R9088 GND.n2194 GND 1.01137
R9089 GND.n2189 GND 1.01137
R9090 GND.n2186 GND 1.01137
R9091 GND GND.n3026 1.01137
R9092 GND GND.n3126 1.01137
R9093 GND GND.n3139 1.01137
R9094 GND.n3141 GND 1.01137
R9095 GND.n3152 GND 1.01137
R9096 GND.n3163 GND 1.01137
R9097 GND.n2520 GND 1.01137
R9098 GND.n3105 GND 1.01137
R9099 GND.n3092 GND 1.01137
R9100 GND.n3082 GND 1.01137
R9101 GND GND.n609 1.01137
R9102 GND.n3056 GND 1.01137
R9103 GND GND.n3945 1.01137
R9104 GND GND.n3950 1.01137
R9105 GND GND.n3955 1.01137
R9106 GND GND.n3958 1.01137
R9107 GND.n3962 GND 1.01137
R9108 GND.n3820 GND 1.01137
R9109 GND.n3815 GND 1.01137
R9110 GND.n3810 GND 1.01137
R9111 GND.n3807 GND 1.01137
R9112 GND.n3802 GND 1.01137
R9113 GND GND.n3783 1.01137
R9114 GND GND.n3788 1.01137
R9115 GND GND.n3793 1.01137
R9116 GND GND.n3796 1.01137
R9117 GND GND.n3801 1.01137
R9118 GND.n3667 GND 1.01137
R9119 GND.n3662 GND 1.01137
R9120 GND.n3657 GND 1.01137
R9121 GND.n3654 GND 1.01137
R9122 GND.n3649 GND 1.01137
R9123 GND.n3587 GND 1.01137
R9124 GND.n4173 GND 1.01137
R9125 GND.n4167 GND 1.01137
R9126 GND GND.n96 1.01137
R9127 GND GND.n3648 1.01137
R9128 GND.n3460 GND 1.01137
R9129 GND.n3455 GND 1.01137
R9130 GND GND.n3547 1.01137
R9131 GND.n3554 GND 1.01137
R9132 GND.n3549 GND 1.01137
R9133 GND.n485 GND 1.01137
R9134 GND GND.n445 1.01137
R9135 GND GND.n450 1.01137
R9136 GND GND.n453 1.01137
R9137 GND GND.n3450 1.01137
R9138 GND.n3249 GND 1.01137
R9139 GND GND.n3226 1.01137
R9140 GND.n3230 GND 1.01137
R9141 GND.n3326 GND 1.01137
R9142 GND.n3321 GND 1.01137
R9143 GND.n549 GND 1.01137
R9144 GND GND.n3195 1.01137
R9145 GND GND.n3200 1.01137
R9146 GND GND.n3203 1.01137
R9147 GND GND.n3208 1.01137
R9148 GND.n1862 GND.n1861 0.645183
R9149 GND.n1896 GND.n1895 0.645183
R9150 GND.n1892 GND.n1891 0.645183
R9151 GND.n1887 GND.n1886 0.645183
R9152 GND.n1882 GND.n1881 0.645183
R9153 GND.n1877 GND.n1876 0.645183
R9154 GND.n1872 GND.n1871 0.645183
R9155 GND.n1867 GND.n1866 0.645183
R9156 GND.n4148 GND.n4147 0.606478
R9157 GND.n145 GND.n114 0.606478
R9158 GND.n4097 GND.n146 0.606478
R9159 GND.n4053 GND.n4052 0.606478
R9160 GND.n203 GND.n172 0.606478
R9161 GND.n4002 GND.n204 0.606478
R9162 GND.n3263 GND.n3262 0.606478
R9163 GND.n3392 GND.n3391 0.606478
R9164 GND.n3390 GND.n3351 0.606478
R9165 GND.n3380 GND.n3376 0.606478
R9166 GND.n3363 GND.n3362 0.606478
R9167 GND.n3940 GND.n3939 0.606478
R9168 GND.n3934 GND.n3933 0.606478
R9169 GND.n3928 GND.n3927 0.606478
R9170 GND.n3918 GND.n3896 0.606478
R9171 GND.n3908 GND.n3902 0.606478
R9172 GND.n275 GND.n274 0.606478
R9173 GND.n3841 GND.n3840 0.606478
R9174 GND.n3854 GND.n3853 0.606478
R9175 GND.n3864 GND.n251 0.606478
R9176 GND.n3874 GND.n246 0.606478
R9177 GND.n3778 GND.n3777 0.606478
R9178 GND.n3772 GND.n3771 0.606478
R9179 GND.n3766 GND.n3765 0.606478
R9180 GND.n3756 GND.n3743 0.606478
R9181 GND.n3746 GND.n3745 0.606478
R9182 GND.n3643 GND.n3642 0.606478
R9183 GND.n3688 GND.n3687 0.606478
R9184 GND.n3701 GND.n3700 0.606478
R9185 GND.n3711 GND.n301 0.606478
R9186 GND.n3721 GND.n296 0.606478
R9187 GND.n3581 GND.n3580 0.606478
R9188 GND.n3605 GND.n3604 0.606478
R9189 GND.n3618 GND.n3617 0.606478
R9190 GND.n3628 GND.n326 0.606478
R9191 GND.n3638 GND.n321 0.606478
R9192 GND.n3522 GND.n3465 0.606478
R9193 GND.n3511 GND.n3470 0.606478
R9194 GND.n3500 GND.n3475 0.606478
R9195 GND.n3499 GND.n3498 0.606478
R9196 GND.n3485 GND.n3484 0.606478
R9197 GND.n3318 GND.n3317 0.606478
R9198 GND.n3405 GND.n3404 0.606478
R9199 GND.n3418 GND.n3417 0.606478
R9200 GND.n3428 GND.n391 0.606478
R9201 GND.n3438 GND.n386 0.606478
R9202 GND.n4297 GND.n4296 0.606478
R9203 GND.n4291 GND.n4290 0.606478
R9204 GND.n4285 GND.n4284 0.606478
R9205 GND.n4275 GND.n17 0.606478
R9206 GND.n4265 GND.n23 0.606478
R9207 GND.n3255 GND.n3254 0.606478
R9208 GND.n3276 GND.n3275 0.606478
R9209 GND.n3289 GND.n3288 0.606478
R9210 GND.n3299 GND.n497 0.606478
R9211 GND.n3303 GND.n3302 0.606478
R9212 GND.n2139 GND.n645 0.606478
R9213 GND.n2129 GND.n650 0.606478
R9214 GND.n2120 GND.n2119 0.606478
R9215 GND.n671 GND.n670 0.606478
R9216 GND.n2106 GND.n672 0.606478
R9217 GND.n729 GND.n728 0.606478
R9218 GND.n741 GND.n740 0.606478
R9219 GND.n753 GND.n752 0.606478
R9220 GND.n763 GND.n762 0.606478
R9221 GND.n774 GND.n773 0.606478
R9222 GND.n2056 GND.n776 0.606478
R9223 GND.n2046 GND.n781 0.606478
R9224 GND.n2037 GND.n2036 0.606478
R9225 GND.n802 GND.n801 0.606478
R9226 GND.n2023 GND.n803 0.606478
R9227 GND.n1368 GND.n1367 0.606478
R9228 GND.n1417 GND.n1369 0.606478
R9229 GND.n1408 GND.n1407 0.606478
R9230 GND.n1387 GND.n1386 0.606478
R9231 GND.n1392 GND.n1388 0.606478
R9232 GND.n1973 GND.n834 0.606478
R9233 GND.n1963 GND.n839 0.606478
R9234 GND.n1954 GND.n1953 0.606478
R9235 GND.n856 GND.n855 0.606478
R9236 GND.n1749 GND.n857 0.606478
R9237 GND.n1737 GND.n864 0.606478
R9238 GND.n1727 GND.n869 0.606478
R9239 GND.n1718 GND.n1717 0.606478
R9240 GND.n1712 GND.n1711 0.606478
R9241 GND.n1706 GND.n1705 0.606478
R9242 GND.n1136 GND.n1135 0.606478
R9243 GND.n1086 GND.n1073 0.606478
R9244 GND.n1121 GND.n1120 0.606478
R9245 GND.n1115 GND.n1114 0.606478
R9246 GND.n1109 GND.n1108 0.606478
R9247 GND.n1661 GND.n914 0.606478
R9248 GND.n1651 GND.n919 0.606478
R9249 GND.n1642 GND.n1641 0.606478
R9250 GND.n1636 GND.n1635 0.606478
R9251 GND.n1630 GND.n1629 0.606478
R9252 GND.n983 GND.n982 0.606478
R9253 GND.n980 GND.n979 0.606478
R9254 GND.n975 GND.n974 0.606478
R9255 GND.n970 GND.n969 0.606478
R9256 GND.n1627 GND.n1626 0.606478
R9257 GND.n1698 GND.n1697 0.606478
R9258 GND.n954 GND.n888 0.606478
R9259 GND.n959 GND.n958 0.606478
R9260 GND.n964 GND.n963 0.606478
R9261 GND.n966 GND.n965 0.606478
R9262 GND.n1528 GND.n1527 0.606478
R9263 GND.n1525 GND.n1524 0.606478
R9264 GND.n1520 GND.n1519 0.606478
R9265 GND.n1515 GND.n1514 0.606478
R9266 GND.n1513 GND.n1512 0.606478
R9267 GND.n1469 GND.n1468 0.606478
R9268 GND.n1466 GND.n1465 0.606478
R9269 GND.n1461 GND.n1460 0.606478
R9270 GND.n1456 GND.n1455 0.606478
R9271 GND.n1508 GND.n1507 0.606478
R9272 GND.n1437 GND.n1436 0.606478
R9273 GND.n1440 GND.n1439 0.606478
R9274 GND.n1445 GND.n1444 0.606478
R9275 GND.n1450 GND.n1449 0.606478
R9276 GND.n1452 GND.n1451 0.606478
R9277 GND.n1318 GND.n1317 0.606478
R9278 GND.n1315 GND.n1314 0.606478
R9279 GND.n1310 GND.n1309 0.606478
R9280 GND.n1305 GND.n1304 0.606478
R9281 GND.n1356 GND.n1355 0.606478
R9282 GND.n1286 GND.n1285 0.606478
R9283 GND.n1289 GND.n1288 0.606478
R9284 GND.n1294 GND.n1293 0.606478
R9285 GND.n1299 GND.n1298 0.606478
R9286 GND.n1301 GND.n1300 0.606478
R9287 GND.n1241 GND.n1240 0.606478
R9288 GND.n1238 GND.n1237 0.606478
R9289 GND.n1233 GND.n1232 0.606478
R9290 GND.n1228 GND.n1227 0.606478
R9291 GND.n1277 GND.n1276 0.606478
R9292 GND.n2866 GND.n2865 0.606478
R9293 GND.n2853 GND.n2472 0.606478
R9294 GND.n2842 GND.n2478 0.606478
R9295 GND.n2841 GND.n2840 0.606478
R9296 GND.n2817 GND.n2815 0.606478
R9297 GND.n2505 GND.n2502 0.606478
R9298 GND.n2504 GND.n2503 0.606478
R9299 GND.n2788 GND.n2787 0.606478
R9300 GND.n2798 GND.n2797 0.606478
R9301 GND.n2828 GND.n2827 0.606478
R9302 GND.n2871 GND.n2870 0.606478
R9303 GND.n2974 GND.n2872 0.606478
R9304 GND.n2961 GND.n2884 0.606478
R9305 GND.n2949 GND.n2894 0.606478
R9306 GND.n2948 GND.n2947 0.606478
R9307 GND.n2925 GND.n2913 0.606478
R9308 GND.n2454 GND.n2453 0.606478
R9309 GND.n2442 GND.n2340 0.606478
R9310 GND.n2429 GND.n2352 0.606478
R9311 GND.n2417 GND.n2362 0.606478
R9312 GND.n2416 GND.n2415 0.606478
R9313 GND.n2393 GND.n2381 0.606478
R9314 GND.n2327 GND.n2326 0.606478
R9315 GND.n2315 GND.n2213 0.606478
R9316 GND.n2302 GND.n2225 0.606478
R9317 GND.n2290 GND.n2235 0.606478
R9318 GND.n2289 GND.n2288 0.606478
R9319 GND.n2266 GND.n2254 0.606478
R9320 GND.n2649 GND.n2648 0.606478
R9321 GND.n2637 GND.n2535 0.606478
R9322 GND.n2624 GND.n2547 0.606478
R9323 GND.n2612 GND.n2557 0.606478
R9324 GND.n2611 GND.n2610 0.606478
R9325 GND.n2588 GND.n2576 0.606478
R9326 GND.n2655 GND.n2654 0.606478
R9327 GND.n2758 GND.n2656 0.606478
R9328 GND.n2745 GND.n2668 0.606478
R9329 GND.n2733 GND.n2678 0.606478
R9330 GND.n2732 GND.n2731 0.606478
R9331 GND.n2709 GND.n2697 0.606478
R9332 GND.n4228 GND.n45 0.606478
R9333 GND.n4217 GND.n4216 0.606478
R9334 GND.n65 GND.n53 0.606478
R9335 GND.n4199 GND.n66 0.606478
R9336 GND.n4188 GND.n4187 0.606478
R9337 GND.n1044 GND.n74 0.606478
R9338 GND.n1586 GND.n1585 0.606478
R9339 GND.n1588 GND.n1587 0.606478
R9340 GND.n1600 GND.n1599 0.606478
R9341 GND.n1614 GND.n1613 0.606478
R9342 GND.n3045 GND.n3044 0.606478
R9343 GND.n3028 GND.n3027 0.606478
R9344 GND.n2200 GND.n2199 0.606478
R9345 GND.n2198 GND.n2197 0.606478
R9346 GND.n2193 GND.n2192 0.606478
R9347 GND.n2188 GND.n2187 0.606478
R9348 GND.n2185 GND.n2184 0.606478
R9349 GND.n2519 GND.n2518 0.606478
R9350 GND.n3128 GND.n3127 0.606478
R9351 GND.n3141 GND.n3140 0.606478
R9352 GND.n3151 GND.n560 0.606478
R9353 GND.n3161 GND.n555 0.606478
R9354 GND.n2521 GND.n2520 0.606478
R9355 GND.n3107 GND.n586 0.606478
R9356 GND.n3094 GND.n598 0.606478
R9357 GND.n3082 GND.n608 0.606478
R9358 GND.n3081 GND.n3080 0.606478
R9359 GND.n3058 GND.n627 0.606478
R9360 GND.n3945 GND.n3944 0.606478
R9361 GND.n3947 GND.n3946 0.606478
R9362 GND.n3952 GND.n3951 0.606478
R9363 GND.n3957 GND.n3956 0.606478
R9364 GND.n3960 GND.n3959 0.606478
R9365 GND.n3821 GND.n3820 0.606478
R9366 GND.n3819 GND.n3818 0.606478
R9367 GND.n3814 GND.n3813 0.606478
R9368 GND.n3809 GND.n3808 0.606478
R9369 GND.n3806 GND.n3805 0.606478
R9370 GND.n3783 GND.n3782 0.606478
R9371 GND.n3785 GND.n3784 0.606478
R9372 GND.n3790 GND.n3789 0.606478
R9373 GND.n3795 GND.n3794 0.606478
R9374 GND.n3798 GND.n3797 0.606478
R9375 GND.n3668 GND.n3667 0.606478
R9376 GND.n3666 GND.n3665 0.606478
R9377 GND.n3661 GND.n3660 0.606478
R9378 GND.n3656 GND.n3655 0.606478
R9379 GND.n3653 GND.n3652 0.606478
R9380 GND.n3587 GND.n3585 0.606478
R9381 GND.n3586 GND.n91 0.606478
R9382 GND.n4172 GND.n4171 0.606478
R9383 GND.n4166 GND.n4165 0.606478
R9384 GND.n3645 GND.n3644 0.606478
R9385 GND.n3461 GND.n3460 0.606478
R9386 GND.n3459 GND.n3458 0.606478
R9387 GND.n3454 GND.n3453 0.606478
R9388 GND.n3555 GND.n3548 0.606478
R9389 GND.n3553 GND.n3552 0.606478
R9390 GND.n486 GND.n485 0.606478
R9391 GND.n442 GND.n441 0.606478
R9392 GND.n447 GND.n446 0.606478
R9393 GND.n452 GND.n451 0.606478
R9394 GND.n455 GND.n454 0.606478
R9395 GND.n3250 GND.n3249 0.606478
R9396 GND.n3223 GND.n3222 0.606478
R9397 GND.n3228 GND.n3227 0.606478
R9398 GND.n3327 GND.n421 0.606478
R9399 GND.n3325 GND.n3324 0.606478
R9400 GND.n549 GND.n544 0.606478
R9401 GND.n548 GND.n547 0.606478
R9402 GND.n3197 GND.n3196 0.606478
R9403 GND.n3202 GND.n3201 0.606478
R9404 GND.n3205 GND.n3204 0.606478
R9405 GND.n1919 GND.n1856 0.601043
R9406 GND.n1861 GND 0.590136
R9407 GND.n1895 GND 0.590136
R9408 GND.n1891 GND 0.590136
R9409 GND.n1886 GND 0.590136
R9410 GND.n1881 GND 0.590136
R9411 GND.n1876 GND 0.590136
R9412 GND.n1871 GND 0.590136
R9413 GND.n1866 GND 0.590136
R9414 GND.n1894 GND.n1893 0.547267
R9415 GND.n2502 GND.n2501 0.495065
R9416 GND.n2870 GND.n2869 0.495065
R9417 GND.n2455 GND.n2454 0.495065
R9418 GND.n2328 GND.n2327 0.495065
R9419 GND.n2650 GND.n2649 0.495065
R9420 GND.n2654 GND.n2653 0.495065
R9421 GND.n2201 GND.n2200 0.495065
R9422 GND.n2522 GND.n2521 0.495065
R9423 GND.n3944 GND.n3943 0.495065
R9424 GND.n3822 GND.n3821 0.495065
R9425 GND.n3782 GND.n3781 0.495065
R9426 GND.n3669 GND.n3668 0.495065
R9427 GND.n3585 GND.n3584 0.495065
R9428 GND.n3462 GND.n3461 0.495065
R9429 GND.n487 GND.n486 0.495065
R9430 GND.n3251 GND.n3250 0.495065
R9431 GND.n544 GND.n543 0.495065
R9432 GND.n3263 GND.n3261 0.476043
R9433 GND.n1890 GND.n1889 0.419583
R9434 GND.n1885 GND.n1884 0.419583
R9435 GND.n1880 GND.n1879 0.419583
R9436 GND.n1875 GND.n1874 0.419583
R9437 GND.n1870 GND.n1869 0.419583
R9438 GND.n1865 GND.n1864 0.419583
R9439 GND.n4147 GND 0.405391
R9440 GND GND.n145 0.405391
R9441 GND GND.n146 0.405391
R9442 GND.n4052 GND 0.405391
R9443 GND GND.n203 0.405391
R9444 GND.n204 GND 0.405391
R9445 GND.n3262 GND 0.405391
R9446 GND.n3391 GND 0.405391
R9447 GND GND.n3351 0.405391
R9448 GND.n3376 GND 0.405391
R9449 GND.n3362 GND 0.405391
R9450 GND GND.n3934 0.405391
R9451 GND GND.n3928 0.405391
R9452 GND.n3896 GND 0.405391
R9453 GND.n3902 GND 0.405391
R9454 GND.n3840 GND 0.405391
R9455 GND.n3853 GND 0.405391
R9456 GND GND.n251 0.405391
R9457 GND GND.n246 0.405391
R9458 GND GND.n3772 0.405391
R9459 GND GND.n3766 0.405391
R9460 GND.n3743 GND 0.405391
R9461 GND.n3745 GND 0.405391
R9462 GND.n3687 GND 0.405391
R9463 GND.n3700 GND 0.405391
R9464 GND GND.n301 0.405391
R9465 GND GND.n296 0.405391
R9466 GND.n3604 GND 0.405391
R9467 GND.n3617 GND 0.405391
R9468 GND GND.n326 0.405391
R9469 GND GND.n321 0.405391
R9470 GND.n3470 GND 0.405391
R9471 GND.n3475 GND 0.405391
R9472 GND GND.n3499 0.405391
R9473 GND.n3484 GND 0.405391
R9474 GND.n3404 GND 0.405391
R9475 GND.n3417 GND 0.405391
R9476 GND GND.n391 0.405391
R9477 GND GND.n386 0.405391
R9478 GND GND.n4291 0.405391
R9479 GND GND.n4285 0.405391
R9480 GND.n17 GND 0.405391
R9481 GND.n23 GND 0.405391
R9482 GND.n3275 GND 0.405391
R9483 GND.n3288 GND 0.405391
R9484 GND GND.n497 0.405391
R9485 GND GND.n3303 0.405391
R9486 GND.n523 GND 0.405391
R9487 GND GND.n645 0.405391
R9488 GND GND.n650 0.405391
R9489 GND.n2119 GND 0.405391
R9490 GND GND.n671 0.405391
R9491 GND GND.n672 0.405391
R9492 GND.n728 GND 0.405391
R9493 GND.n740 GND 0.405391
R9494 GND GND.n753 0.405391
R9495 GND.n762 GND 0.405391
R9496 GND GND.n774 0.405391
R9497 GND GND.n776 0.405391
R9498 GND GND.n781 0.405391
R9499 GND.n2036 GND 0.405391
R9500 GND GND.n802 0.405391
R9501 GND GND.n803 0.405391
R9502 GND GND.n1368 0.405391
R9503 GND GND.n1369 0.405391
R9504 GND.n1407 GND 0.405391
R9505 GND GND.n1387 0.405391
R9506 GND.n1388 GND 0.405391
R9507 GND GND.n834 0.405391
R9508 GND GND.n839 0.405391
R9509 GND.n1953 GND 0.405391
R9510 GND GND.n856 0.405391
R9511 GND GND.n857 0.405391
R9512 GND GND.n864 0.405391
R9513 GND GND.n869 0.405391
R9514 GND.n1717 GND 0.405391
R9515 GND.n1711 GND 0.405391
R9516 GND.n1705 GND 0.405391
R9517 GND.n1135 GND 0.405391
R9518 GND GND.n1086 0.405391
R9519 GND.n1120 GND 0.405391
R9520 GND.n1114 GND 0.405391
R9521 GND.n1108 GND 0.405391
R9522 GND GND.n914 0.405391
R9523 GND GND.n919 0.405391
R9524 GND.n1641 GND 0.405391
R9525 GND.n1635 GND 0.405391
R9526 GND.n1629 GND 0.405391
R9527 GND.n982 GND 0.405391
R9528 GND.n979 GND 0.405391
R9529 GND.n974 GND 0.405391
R9530 GND.n969 GND 0.405391
R9531 GND GND.n1627 0.405391
R9532 GND.n1697 GND 0.405391
R9533 GND GND.n954 0.405391
R9534 GND GND.n959 0.405391
R9535 GND GND.n964 0.405391
R9536 GND GND.n966 0.405391
R9537 GND.n1527 GND 0.405391
R9538 GND.n1524 GND 0.405391
R9539 GND.n1519 GND 0.405391
R9540 GND.n1514 GND 0.405391
R9541 GND.n1512 GND 0.405391
R9542 GND.n1468 GND 0.405391
R9543 GND.n1465 GND 0.405391
R9544 GND.n1460 GND 0.405391
R9545 GND.n1455 GND 0.405391
R9546 GND GND.n1508 0.405391
R9547 GND GND.n1437 0.405391
R9548 GND GND.n1440 0.405391
R9549 GND GND.n1445 0.405391
R9550 GND GND.n1450 0.405391
R9551 GND GND.n1452 0.405391
R9552 GND.n1317 GND 0.405391
R9553 GND.n1314 GND 0.405391
R9554 GND.n1309 GND 0.405391
R9555 GND.n1304 GND 0.405391
R9556 GND GND.n1356 0.405391
R9557 GND GND.n1286 0.405391
R9558 GND GND.n1289 0.405391
R9559 GND GND.n1294 0.405391
R9560 GND GND.n1299 0.405391
R9561 GND GND.n1301 0.405391
R9562 GND.n1240 GND 0.405391
R9563 GND.n1237 GND 0.405391
R9564 GND.n1232 GND 0.405391
R9565 GND.n1227 GND 0.405391
R9566 GND GND.n1277 0.405391
R9567 GND.n2472 GND 0.405391
R9568 GND.n2478 GND 0.405391
R9569 GND GND.n2841 0.405391
R9570 GND.n2815 GND 0.405391
R9571 GND GND.n2504 0.405391
R9572 GND.n2787 GND 0.405391
R9573 GND GND.n2828 0.405391
R9574 GND.n2872 GND 0.405391
R9575 GND.n2884 GND 0.405391
R9576 GND.n2894 GND 0.405391
R9577 GND GND.n2948 0.405391
R9578 GND.n2913 GND 0.405391
R9579 GND.n2340 GND 0.405391
R9580 GND.n2352 GND 0.405391
R9581 GND.n2362 GND 0.405391
R9582 GND GND.n2416 0.405391
R9583 GND.n2381 GND 0.405391
R9584 GND.n2213 GND 0.405391
R9585 GND.n2225 GND 0.405391
R9586 GND.n2235 GND 0.405391
R9587 GND GND.n2289 0.405391
R9588 GND.n2254 GND 0.405391
R9589 GND.n2535 GND 0.405391
R9590 GND.n2547 GND 0.405391
R9591 GND.n2557 GND 0.405391
R9592 GND GND.n2611 0.405391
R9593 GND.n2576 GND 0.405391
R9594 GND.n2656 GND 0.405391
R9595 GND.n2668 GND 0.405391
R9596 GND.n2678 GND 0.405391
R9597 GND GND.n2732 0.405391
R9598 GND.n2697 GND 0.405391
R9599 GND GND.n45 0.405391
R9600 GND.n4216 GND 0.405391
R9601 GND GND.n65 0.405391
R9602 GND GND.n66 0.405391
R9603 GND.n4187 GND 0.405391
R9604 GND GND.n1044 0.405391
R9605 GND GND.n1586 0.405391
R9606 GND.n1587 GND 0.405391
R9607 GND.n1599 GND 0.405391
R9608 GND.n1613 GND 0.405391
R9609 GND.n3044 GND 0.405391
R9610 GND.n3027 GND 0.405391
R9611 GND GND.n2198 0.405391
R9612 GND GND.n2193 0.405391
R9613 GND GND.n2185 0.405391
R9614 GND.n3127 GND 0.405391
R9615 GND.n3140 GND 0.405391
R9616 GND GND.n560 0.405391
R9617 GND GND.n555 0.405391
R9618 GND GND.n586 0.405391
R9619 GND.n598 GND 0.405391
R9620 GND.n608 GND 0.405391
R9621 GND GND.n3081 0.405391
R9622 GND.n627 GND 0.405391
R9623 GND.n3946 GND 0.405391
R9624 GND.n3951 GND 0.405391
R9625 GND.n3959 GND 0.405391
R9626 GND GND.n3819 0.405391
R9627 GND GND.n3814 0.405391
R9628 GND GND.n3806 0.405391
R9629 GND.n3784 GND 0.405391
R9630 GND.n3789 GND 0.405391
R9631 GND.n3797 GND 0.405391
R9632 GND GND.n3666 0.405391
R9633 GND GND.n3661 0.405391
R9634 GND GND.n3653 0.405391
R9635 GND GND.n3586 0.405391
R9636 GND GND.n4172 0.405391
R9637 GND.n3644 GND 0.405391
R9638 GND GND.n3459 0.405391
R9639 GND GND.n3454 0.405391
R9640 GND GND.n3553 0.405391
R9641 GND.n441 GND 0.405391
R9642 GND.n446 GND 0.405391
R9643 GND.n454 GND 0.405391
R9644 GND.n3222 GND 0.405391
R9645 GND.n3227 GND 0.405391
R9646 GND GND.n3325 0.405391
R9647 GND GND.n548 0.405391
R9648 GND.n3196 GND 0.405391
R9649 GND.n3204 GND 0.405391
R9650 GND.n1859 GND.n1858 0.353761
R9651 GND.n1921 GND 0.149957
R9652 GND.n1628 GND 0.0901739
R9653 GND.n967 GND 0.0901739
R9654 GND GND.n1511 0.0901739
R9655 GND.n1509 GND 0.0901739
R9656 GND.n1453 GND 0.0901739
R9657 GND.n1357 GND 0.0901739
R9658 GND.n1302 GND 0.0901739
R9659 GND.n1278 GND 0.0901739
R9660 GND.n1934 GND.n1765 0.063
R9661 GND.n1765 GND.n1764 0.063
R9662 GND.n1930 GND.n1781 0.063
R9663 GND.n1786 GND.n1781 0.063
R9664 GND.n1928 GND.n1796 0.063
R9665 GND.n1801 GND.n1796 0.063
R9666 GND.n1926 GND.n1811 0.063
R9667 GND.n1816 GND.n1811 0.063
R9668 GND.n1924 GND.n1826 0.063
R9669 GND.n1831 GND.n1826 0.063
R9670 GND.n1922 GND.n1841 0.063
R9671 GND.n1846 GND.n1841 0.063
R9672 GND.n1898 GND.n1859 0.063
R9673 GND.n1899 GND.n1898 0.063
R9674 GND.n1932 GND.n1766 0.063
R9675 GND.n1771 GND.n1766 0.063
R9676 GND.n3260 GND.n534 0.063
R9677 GND.n3261 GND.n3260 0.063
R9678 GND.n1921 GND.n1920 0.063
R9679 GND.n3943 GND.n3942 0.063
R9680 GND.n3823 GND.n3822 0.063
R9681 GND.n3781 GND.n3780 0.063
R9682 GND.n3670 GND.n3669 0.063
R9683 GND.n3584 GND.n3583 0.063
R9684 GND.n3463 GND.n3462 0.063
R9685 GND.n3320 GND.n487 0.063
R9686 GND.n3257 GND.n3251 0.063
R9687 GND.n968 GND 0.0454219
R9688 GND.n1703 GND 0.0454219
R9689 GND.n1510 GND 0.0454219
R9690 GND.n1454 GND 0.0454219
R9691 GND.n1432 GND 0.0454219
R9692 GND.n1303 GND 0.0454219
R9693 GND.n1281 GND 0.0454219
R9694 GND.n1920 GND 0.0454219
R9695 GND.n1628 GND 0.0249565
R9696 GND.n967 GND 0.0249565
R9697 GND.n1511 GND 0.0249565
R9698 GND.n1509 GND 0.0249565
R9699 GND.n1453 GND 0.0249565
R9700 GND.n1357 GND 0.0249565
R9701 GND.n1302 GND 0.0249565
R9702 GND.n1278 GND 0.0249565
R9703 GND.n1861 GND.n1860 0.024
R9704 GND.n1895 GND.n1894 0.024
R9705 GND.n1891 GND.n1890 0.024
R9706 GND.n1886 GND.n1885 0.024
R9707 GND.n1881 GND.n1880 0.024
R9708 GND.n1876 GND.n1875 0.024
R9709 GND.n1871 GND.n1870 0.024
R9710 GND.n1866 GND.n1865 0.024
R9711 GND.n1935 GND.n1934 0.0232079
R9712 GND.n1932 GND.n1780 0.0232079
R9713 GND.n1930 GND.n1795 0.0232079
R9714 GND.n1928 GND.n1810 0.0232079
R9715 GND.n1926 GND.n1825 0.0232079
R9716 GND.n1924 GND.n1840 0.0232079
R9717 GND.n1922 GND.n1855 0.0232079
R9718 GND.n1863 GND 0.0204394
R9719 GND.n1897 GND 0.0204394
R9720 GND.n1893 GND 0.0204394
R9721 GND.n1888 GND 0.0204394
R9722 GND.n1883 GND 0.0204394
R9723 GND.n1878 GND 0.0204394
R9724 GND.n1873 GND 0.0204394
R9725 GND.n1868 GND 0.0204394
R9726 GND GND.n1628 0.0180781
R9727 GND GND.n967 0.0180781
R9728 GND.n1511 GND 0.0180781
R9729 GND GND.n1509 0.0180781
R9730 GND GND.n1453 0.0180781
R9731 GND GND.n1357 0.0180781
R9732 GND GND.n1302 0.0180781
R9733 GND GND.n1278 0.0180781
R9734 GND.n1862 GND 0.00441667
R9735 GND.n1896 GND 0.00441667
R9736 GND.n1892 GND 0.00441667
R9737 GND.n1887 GND 0.00441667
R9738 GND.n1882 GND 0.00441667
R9739 GND.n1877 GND 0.00441667
R9740 GND.n1872 GND 0.00441667
R9741 GND.n1867 GND 0.00441667
R9742 GND GND.n4298 0.00441667
R9743 GND GND.n1862 0.00406061
R9744 GND GND.n1896 0.00406061
R9745 GND GND.n1892 0.00406061
R9746 GND GND.n1887 0.00406061
R9747 GND GND.n1882 0.00406061
R9748 GND GND.n1877 0.00406061
R9749 GND GND.n1872 0.00406061
R9750 GND GND.n1867 0.00406061
R9751 GND.n4298 GND 0.00406061
R9752 GND.n1934 GND 0.00287997
R9753 GND.n1933 GND.n1932 0.00287997
R9754 GND.n1932 GND 0.00287997
R9755 GND.n1931 GND.n1930 0.00287997
R9756 GND.n1930 GND 0.00287997
R9757 GND.n1929 GND.n1928 0.00287997
R9758 GND.n1928 GND 0.00287997
R9759 GND.n1927 GND.n1926 0.00287997
R9760 GND.n1926 GND 0.00287997
R9761 GND.n1925 GND.n1924 0.00287997
R9762 GND.n1924 GND 0.00287997
R9763 GND.n1923 GND.n1922 0.00287997
R9764 GND.n1922 GND 0.00287997
R9765 CLK.n244 CLK.t23 158.207
R9766 CLK.n231 CLK.t8 158.207
R9767 CLK.n218 CLK.t59 158.207
R9768 CLK.n205 CLK.t2 158.207
R9769 CLK.n192 CLK.t93 158.207
R9770 CLK.n179 CLK.t22 158.207
R9771 CLK.n166 CLK.t5 158.207
R9772 CLK.n154 CLK.t102 158.207
R9773 CLK.n104 CLK.t13 158.207
R9774 CLK.n91 CLK.t80 158.207
R9775 CLK.n78 CLK.t51 158.207
R9776 CLK.n65 CLK.t114 158.207
R9777 CLK.n52 CLK.t84 158.207
R9778 CLK.n39 CLK.t54 158.207
R9779 CLK.n27 CLK.t117 158.207
R9780 CLK.n15 CLK.t27 158.207
R9781 CLK.n3 CLK.t95 158.207
R9782 CLK CLK.t100 158.202
R9783 CLK CLK.t72 158.202
R9784 CLK CLK.t15 158.202
R9785 CLK CLK.t62 158.202
R9786 CLK CLK.t37 158.202
R9787 CLK CLK.t97 158.202
R9788 CLK CLK.t69 158.202
R9789 CLK CLK.t45 158.202
R9790 CLK CLK.t83 158.202
R9791 CLK CLK.t30 158.202
R9792 CLK CLK.t16 158.202
R9793 CLK CLK.t63 158.202
R9794 CLK CLK.t38 158.202
R9795 CLK CLK.t19 158.202
R9796 CLK CLK.t70 158.202
R9797 CLK CLK.t113 158.202
R9798 CLK CLK.t42 158.202
R9799 CLK.n246 CLK.t39 150.293
R9800 CLK.t100 CLK.n249 150.293
R9801 CLK.n233 CLK.t26 150.293
R9802 CLK.t72 CLK.n236 150.293
R9803 CLK.n220 CLK.t108 150.293
R9804 CLK.t15 CLK.n223 150.293
R9805 CLK.n207 CLK.t75 150.293
R9806 CLK.t62 CLK.n210 150.293
R9807 CLK.n194 CLK.t47 150.293
R9808 CLK.t37 CLK.n197 150.293
R9809 CLK.n181 CLK.t111 150.293
R9810 CLK.t97 CLK.n184 150.293
R9811 CLK.n168 CLK.t78 150.293
R9812 CLK.t69 CLK.n171 150.293
R9813 CLK.n156 CLK.t17 150.293
R9814 CLK.t45 CLK.n159 150.293
R9815 CLK.n128 CLK.t44 150.293
R9816 CLK.n131 CLK.t87 150.293
R9817 CLK.n134 CLK.t34 150.293
R9818 CLK.n125 CLK.t18 150.293
R9819 CLK.n106 CLK.t31 150.293
R9820 CLK.t83 CLK.n109 150.293
R9821 CLK.n93 CLK.t52 150.293
R9822 CLK.t30 CLK.n96 150.293
R9823 CLK.n80 CLK.t25 150.293
R9824 CLK.t16 CLK.n83 150.293
R9825 CLK.n67 CLK.t11 150.293
R9826 CLK.t63 CLK.n70 150.293
R9827 CLK.n54 CLK.t55 150.293
R9828 CLK.t38 CLK.n57 150.293
R9829 CLK.n41 CLK.t28 150.293
R9830 CLK.t19 CLK.n44 150.293
R9831 CLK.n29 CLK.t88 150.293
R9832 CLK.t70 CLK.n32 150.293
R9833 CLK.n17 CLK.t57 150.293
R9834 CLK.t113 CLK.n20 150.293
R9835 CLK.n5 CLK.t33 150.293
R9836 CLK.t42 CLK.n8 150.293
R9837 CLK.t23 CLK.n243 150.273
R9838 CLK.t8 CLK.n230 150.273
R9839 CLK.t59 CLK.n217 150.273
R9840 CLK.t2 CLK.n204 150.273
R9841 CLK.t93 CLK.n191 150.273
R9842 CLK.t22 CLK.n178 150.273
R9843 CLK.t5 CLK.n165 150.273
R9844 CLK.t102 CLK.n153 150.273
R9845 CLK.n123 CLK.t105 150.273
R9846 CLK.n119 CLK.t77 150.273
R9847 CLK.n141 CLK.t74 150.273
R9848 CLK.n146 CLK.t110 150.273
R9849 CLK.t13 CLK.n103 150.273
R9850 CLK.t80 CLK.n90 150.273
R9851 CLK.t51 CLK.n77 150.273
R9852 CLK.t114 CLK.n64 150.273
R9853 CLK.t84 CLK.n51 150.273
R9854 CLK.t54 CLK.n38 150.273
R9855 CLK.t117 CLK.n26 150.273
R9856 CLK.t27 CLK.n14 150.273
R9857 CLK.t95 CLK.n2 150.273
R9858 CLK.n241 CLK.t40 73.6406
R9859 CLK.n228 CLK.t98 73.6406
R9860 CLK.n215 CLK.t29 73.6406
R9861 CLK.n202 CLK.t89 73.6406
R9862 CLK.n189 CLK.t60 73.6406
R9863 CLK.n176 CLK.t35 73.6406
R9864 CLK.n163 CLK.t96 73.6406
R9865 CLK.n151 CLK.t68 73.6406
R9866 CLK.n101 CLK.t20 73.6406
R9867 CLK.n88 CLK.t91 73.6406
R9868 CLK.n75 CLK.t65 73.6406
R9869 CLK.n62 CLK.t41 73.6406
R9870 CLK.n49 CLK.t99 73.6406
R9871 CLK.n36 CLK.t71 73.6406
R9872 CLK.n24 CLK.t9 73.6406
R9873 CLK.n12 CLK.t46 73.6406
R9874 CLK.n0 CLK.t64 73.6406
R9875 CLK.n248 CLK.t58 73.6304
R9876 CLK.n247 CLK.t107 73.6304
R9877 CLK.n235 CLK.t1 73.6304
R9878 CLK.n234 CLK.t94 73.6304
R9879 CLK.n222 CLK.t53 73.6304
R9880 CLK.n221 CLK.t67 73.6304
R9881 CLK.n209 CLK.t116 73.6304
R9882 CLK.n208 CLK.t6 73.6304
R9883 CLK.n196 CLK.t85 73.6304
R9884 CLK.n195 CLK.t103 73.6304
R9885 CLK.n183 CLK.t56 73.6304
R9886 CLK.n182 CLK.t24 73.6304
R9887 CLK.n170 CLK.t0 73.6304
R9888 CLK.n169 CLK.t10 73.6304
R9889 CLK.n158 CLK.t90 73.6304
R9890 CLK.n157 CLK.t106 73.6304
R9891 CLK.n129 CLK.t81 73.6304
R9892 CLK.n132 CLK.t48 73.6304
R9893 CLK.n120 CLK.t21 73.6304
R9894 CLK.n116 CLK.t3 73.6304
R9895 CLK.n138 CLK.t115 73.6304
R9896 CLK.n143 CLK.t61 73.6304
R9897 CLK.n135 CLK.t43 73.6304
R9898 CLK.n126 CLK.t49 73.6304
R9899 CLK.n108 CLK.t50 73.6304
R9900 CLK.n107 CLK.t104 73.6304
R9901 CLK.n95 CLK.t12 73.6304
R9902 CLK.n94 CLK.t32 73.6304
R9903 CLK.n82 CLK.t109 73.6304
R9904 CLK.n81 CLK.t92 73.6304
R9905 CLK.n69 CLK.t76 73.6304
R9906 CLK.n68 CLK.t66 73.6304
R9907 CLK.n56 CLK.t14 73.6304
R9908 CLK.n55 CLK.t4 73.6304
R9909 CLK.n43 CLK.t112 73.6304
R9910 CLK.n42 CLK.t101 73.6304
R9911 CLK.n31 CLK.t36 73.6304
R9912 CLK.n30 CLK.t73 73.6304
R9913 CLK.n19 CLK.t79 73.6304
R9914 CLK.n18 CLK.t7 73.6304
R9915 CLK.n7 CLK.t86 73.6304
R9916 CLK.n6 CLK.t82 73.6304
R9917 CLK.n124 CLK.n119 64.4516
R9918 CLK.n147 CLK.n142 59.9516
R9919 CLK.n133 CLK.n130 59.9516
R9920 CLK.n136 CLK.n135 54.8429
R9921 CLK.n142 CLK.n137 37.8646
R9922 CLK.n127 CLK.n126 34.5521
R9923 CLK.n137 CLK.n136 30.474
R9924 CLK.n130 CLK.n127 29.8239
R9925 CLK.n148 CLK.n115 23.654
R9926 CLK.n137 CLK.n124 22.0114
R9927 CLK.n248 CLK.n247 16.332
R9928 CLK.n235 CLK.n234 16.332
R9929 CLK.n222 CLK.n221 16.332
R9930 CLK.n209 CLK.n208 16.332
R9931 CLK.n196 CLK.n195 16.332
R9932 CLK.n183 CLK.n182 16.332
R9933 CLK.n170 CLK.n169 16.332
R9934 CLK.n158 CLK.n157 16.332
R9935 CLK.n108 CLK.n107 16.332
R9936 CLK.n95 CLK.n94 16.332
R9937 CLK.n82 CLK.n81 16.332
R9938 CLK.n69 CLK.n68 16.332
R9939 CLK.n56 CLK.n55 16.332
R9940 CLK.n43 CLK.n42 16.332
R9941 CLK.n31 CLK.n30 16.332
R9942 CLK.n19 CLK.n18 16.332
R9943 CLK.n7 CLK.n6 16.332
R9944 CLK.n175 CLK.n162 12.0538
R9945 CLK.n48 CLK.n35 12.0538
R9946 CLK.n136 CLK.n133 9.53311
R9947 CLK.n149 CLK.n11 9.40927
R9948 CLK.n188 CLK.n175 8.6438
R9949 CLK.n201 CLK.n188 8.6438
R9950 CLK.n214 CLK.n201 8.6438
R9951 CLK.n227 CLK.n214 8.6438
R9952 CLK.n240 CLK.n227 8.6438
R9953 CLK.n253 CLK.n240 8.6438
R9954 CLK.n61 CLK.n48 8.6438
R9955 CLK.n74 CLK.n61 8.6438
R9956 CLK.n87 CLK.n74 8.6438
R9957 CLK.n100 CLK.n87 8.6438
R9958 CLK.n113 CLK.n100 8.6438
R9959 CLK.n114 CLK.n23 6.21797
R9960 CLK.n115 CLK.n114 6.0284
R9961 CLK.n149 CLK.n148 5.92422
R9962 CLK.n114 CLK.n113 5.83163
R9963 CLK.n148 CLK.n147 4.90235
R9964 CLK.n124 CLK.n123 4.5005
R9965 CLK.n147 CLK.n146 4.5005
R9966 CLK.n142 CLK.n141 4.5005
R9967 CLK.n133 CLK.n132 4.5005
R9968 CLK.n130 CLK.n129 4.5005
R9969 CLK.n175 CLK.n174 3.4105
R9970 CLK.n188 CLK.n187 3.4105
R9971 CLK.n201 CLK.n200 3.4105
R9972 CLK.n214 CLK.n213 3.4105
R9973 CLK.n227 CLK.n226 3.4105
R9974 CLK.n240 CLK.n239 3.4105
R9975 CLK.n48 CLK.n47 3.4105
R9976 CLK.n61 CLK.n60 3.4105
R9977 CLK.n74 CLK.n73 3.4105
R9978 CLK.n87 CLK.n86 3.4105
R9979 CLK.n100 CLK.n99 3.4105
R9980 CLK.n113 CLK.n112 3.4105
R9981 CLK.n127 CLK.n115 3.4105
R9982 CLK.n253 CLK.n252 3.4105
R9983 CLK.n254 CLK.n150 2.59333
R9984 CLK.n150 CLK 2.35833
R9985 CLK.n242 CLK.n241 1.19615
R9986 CLK.n229 CLK.n228 1.19615
R9987 CLK.n216 CLK.n215 1.19615
R9988 CLK.n203 CLK.n202 1.19615
R9989 CLK.n190 CLK.n189 1.19615
R9990 CLK.n177 CLK.n176 1.19615
R9991 CLK.n164 CLK.n163 1.19615
R9992 CLK.n152 CLK.n151 1.19615
R9993 CLK.n102 CLK.n101 1.19615
R9994 CLK.n89 CLK.n88 1.19615
R9995 CLK.n76 CLK.n75 1.19615
R9996 CLK.n63 CLK.n62 1.19615
R9997 CLK.n50 CLK.n49 1.19615
R9998 CLK.n37 CLK.n36 1.19615
R9999 CLK.n25 CLK.n24 1.19615
R10000 CLK.n13 CLK.n12 1.19615
R10001 CLK.n1 CLK.n0 1.19615
R10002 CLK.n247 CLK.n246 1.1717
R10003 CLK.n249 CLK.n248 1.1717
R10004 CLK.n234 CLK.n233 1.1717
R10005 CLK.n236 CLK.n235 1.1717
R10006 CLK.n221 CLK.n220 1.1717
R10007 CLK.n223 CLK.n222 1.1717
R10008 CLK.n208 CLK.n207 1.1717
R10009 CLK.n210 CLK.n209 1.1717
R10010 CLK.n195 CLK.n194 1.1717
R10011 CLK.n197 CLK.n196 1.1717
R10012 CLK.n182 CLK.n181 1.1717
R10013 CLK.n184 CLK.n183 1.1717
R10014 CLK.n169 CLK.n168 1.1717
R10015 CLK.n171 CLK.n170 1.1717
R10016 CLK.n157 CLK.n156 1.1717
R10017 CLK.n159 CLK.n158 1.1717
R10018 CLK.n129 CLK.n128 1.1717
R10019 CLK.n132 CLK.n131 1.1717
R10020 CLK.n122 CLK.n121 1.1717
R10021 CLK.n118 CLK.n117 1.1717
R10022 CLK.n140 CLK.n139 1.1717
R10023 CLK.n145 CLK.n144 1.1717
R10024 CLK.n135 CLK.n134 1.1717
R10025 CLK.n126 CLK.n125 1.1717
R10026 CLK.n107 CLK.n106 1.1717
R10027 CLK.n109 CLK.n108 1.1717
R10028 CLK.n94 CLK.n93 1.1717
R10029 CLK.n96 CLK.n95 1.1717
R10030 CLK.n81 CLK.n80 1.1717
R10031 CLK.n83 CLK.n82 1.1717
R10032 CLK.n68 CLK.n67 1.1717
R10033 CLK.n70 CLK.n69 1.1717
R10034 CLK.n55 CLK.n54 1.1717
R10035 CLK.n57 CLK.n56 1.1717
R10036 CLK.n42 CLK.n41 1.1717
R10037 CLK.n44 CLK.n43 1.1717
R10038 CLK.n30 CLK.n29 1.1717
R10039 CLK.n32 CLK.n31 1.1717
R10040 CLK.n18 CLK.n17 1.1717
R10041 CLK.n20 CLK.n19 1.1717
R10042 CLK.n6 CLK.n5 1.1717
R10043 CLK.n8 CLK.n7 1.1717
R10044 CLK.n122 CLK 0.932141
R10045 CLK.n118 CLK 0.932141
R10046 CLK.n140 CLK 0.932141
R10047 CLK.n145 CLK 0.932141
R10048 CLK.n249 CLK 0.447191
R10049 CLK.n236 CLK 0.447191
R10050 CLK.n223 CLK 0.447191
R10051 CLK.n210 CLK 0.447191
R10052 CLK.n197 CLK 0.447191
R10053 CLK.n184 CLK 0.447191
R10054 CLK.n171 CLK 0.447191
R10055 CLK.n159 CLK 0.447191
R10056 CLK.n128 CLK 0.447191
R10057 CLK.n131 CLK 0.447191
R10058 CLK.n134 CLK 0.447191
R10059 CLK.n125 CLK 0.447191
R10060 CLK.n109 CLK 0.447191
R10061 CLK.n96 CLK 0.447191
R10062 CLK.n83 CLK 0.447191
R10063 CLK.n70 CLK 0.447191
R10064 CLK.n57 CLK 0.447191
R10065 CLK.n44 CLK 0.447191
R10066 CLK.n32 CLK 0.447191
R10067 CLK.n20 CLK 0.447191
R10068 CLK.n8 CLK 0.447191
R10069 CLK.n246 CLK 0.436162
R10070 CLK.n233 CLK 0.436162
R10071 CLK.n220 CLK 0.436162
R10072 CLK.n207 CLK 0.436162
R10073 CLK.n194 CLK 0.436162
R10074 CLK.n181 CLK 0.436162
R10075 CLK.n168 CLK 0.436162
R10076 CLK.n156 CLK 0.436162
R10077 CLK.n106 CLK 0.436162
R10078 CLK.n93 CLK 0.436162
R10079 CLK.n80 CLK 0.436162
R10080 CLK.n67 CLK 0.436162
R10081 CLK.n54 CLK 0.436162
R10082 CLK.n41 CLK 0.436162
R10083 CLK.n29 CLK 0.436162
R10084 CLK.n17 CLK 0.436162
R10085 CLK.n5 CLK 0.436162
R10086 CLK.n244 CLK 0.321667
R10087 CLK.n231 CLK 0.321667
R10088 CLK.n218 CLK 0.321667
R10089 CLK.n205 CLK 0.321667
R10090 CLK.n192 CLK 0.321667
R10091 CLK.n179 CLK 0.321667
R10092 CLK.n166 CLK 0.321667
R10093 CLK.n154 CLK 0.321667
R10094 CLK.n104 CLK 0.321667
R10095 CLK.n91 CLK 0.321667
R10096 CLK.n78 CLK 0.321667
R10097 CLK.n65 CLK 0.321667
R10098 CLK.n52 CLK 0.321667
R10099 CLK.n39 CLK 0.321667
R10100 CLK.n27 CLK 0.321667
R10101 CLK.n15 CLK 0.321667
R10102 CLK.n3 CLK 0.321667
R10103 CLK.n241 CLK 0.217464
R10104 CLK.n228 CLK 0.217464
R10105 CLK.n215 CLK 0.217464
R10106 CLK.n202 CLK 0.217464
R10107 CLK.n189 CLK 0.217464
R10108 CLK.n176 CLK 0.217464
R10109 CLK.n163 CLK 0.217464
R10110 CLK.n151 CLK 0.217464
R10111 CLK.n101 CLK 0.217464
R10112 CLK.n88 CLK 0.217464
R10113 CLK.n75 CLK 0.217464
R10114 CLK.n62 CLK 0.217464
R10115 CLK.n49 CLK 0.217464
R10116 CLK.n36 CLK 0.217464
R10117 CLK.n24 CLK 0.217464
R10118 CLK.n12 CLK 0.217464
R10119 CLK.n0 CLK 0.217464
R10120 CLK.n245 CLK 0.208867
R10121 CLK.n232 CLK 0.208867
R10122 CLK.n219 CLK 0.208867
R10123 CLK.n206 CLK 0.208867
R10124 CLK.n193 CLK 0.208867
R10125 CLK.n180 CLK 0.208867
R10126 CLK.n167 CLK 0.208867
R10127 CLK.n155 CLK 0.208867
R10128 CLK.n105 CLK 0.208867
R10129 CLK.n92 CLK 0.208867
R10130 CLK.n79 CLK 0.208867
R10131 CLK.n66 CLK 0.208867
R10132 CLK.n53 CLK 0.208867
R10133 CLK.n40 CLK 0.208867
R10134 CLK.n28 CLK 0.208867
R10135 CLK.n16 CLK 0.208867
R10136 CLK.n4 CLK 0.208867
R10137 CLK.n248 CLK 0.149957
R10138 CLK.n235 CLK 0.149957
R10139 CLK.n222 CLK 0.149957
R10140 CLK.n209 CLK 0.149957
R10141 CLK.n196 CLK 0.149957
R10142 CLK.n183 CLK 0.149957
R10143 CLK.n170 CLK 0.149957
R10144 CLK.n158 CLK 0.149957
R10145 CLK.n129 CLK 0.149957
R10146 CLK.n132 CLK 0.149957
R10147 CLK.n135 CLK 0.149957
R10148 CLK.n126 CLK 0.149957
R10149 CLK.n108 CLK 0.149957
R10150 CLK.n95 CLK 0.149957
R10151 CLK.n82 CLK 0.149957
R10152 CLK.n69 CLK 0.149957
R10153 CLK.n56 CLK 0.149957
R10154 CLK.n43 CLK 0.149957
R10155 CLK.n31 CLK 0.149957
R10156 CLK.n19 CLK 0.149957
R10157 CLK.n7 CLK 0.149957
R10158 CLK.n245 CLK.n244 0.145417
R10159 CLK.n251 CLK.n250 0.145417
R10160 CLK.n232 CLK.n231 0.145417
R10161 CLK.n238 CLK.n237 0.145417
R10162 CLK.n219 CLK.n218 0.145417
R10163 CLK.n225 CLK.n224 0.145417
R10164 CLK.n206 CLK.n205 0.145417
R10165 CLK.n212 CLK.n211 0.145417
R10166 CLK.n193 CLK.n192 0.145417
R10167 CLK.n199 CLK.n198 0.145417
R10168 CLK.n180 CLK.n179 0.145417
R10169 CLK.n186 CLK.n185 0.145417
R10170 CLK.n167 CLK.n166 0.145417
R10171 CLK.n173 CLK.n172 0.145417
R10172 CLK.n155 CLK.n154 0.145417
R10173 CLK.n161 CLK.n160 0.145417
R10174 CLK.n105 CLK.n104 0.145417
R10175 CLK.n111 CLK.n110 0.145417
R10176 CLK.n92 CLK.n91 0.145417
R10177 CLK.n98 CLK.n97 0.145417
R10178 CLK.n79 CLK.n78 0.145417
R10179 CLK.n85 CLK.n84 0.145417
R10180 CLK.n66 CLK.n65 0.145417
R10181 CLK.n72 CLK.n71 0.145417
R10182 CLK.n53 CLK.n52 0.145417
R10183 CLK.n59 CLK.n58 0.145417
R10184 CLK.n40 CLK.n39 0.145417
R10185 CLK.n46 CLK.n45 0.145417
R10186 CLK.n28 CLK.n27 0.145417
R10187 CLK.n34 CLK.n33 0.145417
R10188 CLK.n16 CLK.n15 0.145417
R10189 CLK.n22 CLK.n21 0.145417
R10190 CLK.n4 CLK.n3 0.145417
R10191 CLK.n10 CLK.n9 0.145417
R10192 CLK.n242 CLK 0.1255
R10193 CLK.n229 CLK 0.1255
R10194 CLK.n216 CLK 0.1255
R10195 CLK.n203 CLK 0.1255
R10196 CLK.n190 CLK 0.1255
R10197 CLK.n177 CLK 0.1255
R10198 CLK.n164 CLK 0.1255
R10199 CLK.n152 CLK 0.1255
R10200 CLK.n121 CLK 0.1255
R10201 CLK.n117 CLK 0.1255
R10202 CLK.n139 CLK 0.1255
R10203 CLK.n144 CLK 0.1255
R10204 CLK.n102 CLK 0.1255
R10205 CLK.n89 CLK 0.1255
R10206 CLK.n76 CLK 0.1255
R10207 CLK.n63 CLK 0.1255
R10208 CLK.n50 CLK 0.1255
R10209 CLK.n37 CLK 0.1255
R10210 CLK.n25 CLK 0.1255
R10211 CLK.n13 CLK 0.1255
R10212 CLK.n1 CLK 0.1255
R10213 CLK.n251 CLK 0.118
R10214 CLK.n238 CLK 0.118
R10215 CLK.n225 CLK 0.118
R10216 CLK.n212 CLK 0.118
R10217 CLK.n199 CLK 0.118
R10218 CLK.n186 CLK 0.118
R10219 CLK.n173 CLK 0.118
R10220 CLK.n161 CLK 0.118
R10221 CLK.n111 CLK 0.118
R10222 CLK.n98 CLK 0.118
R10223 CLK.n85 CLK 0.118
R10224 CLK.n72 CLK 0.118
R10225 CLK.n59 CLK 0.118
R10226 CLK.n46 CLK 0.118
R10227 CLK.n34 CLK 0.118
R10228 CLK.n22 CLK 0.118
R10229 CLK.n10 CLK 0.118
R10230 CLK.n247 CLK 0.117348
R10231 CLK.n234 CLK 0.117348
R10232 CLK.n221 CLK 0.117348
R10233 CLK.n208 CLK 0.117348
R10234 CLK.n195 CLK 0.117348
R10235 CLK.n182 CLK 0.117348
R10236 CLK.n169 CLK 0.117348
R10237 CLK.n157 CLK 0.117348
R10238 CLK.n107 CLK 0.117348
R10239 CLK.n94 CLK 0.117348
R10240 CLK.n81 CLK 0.117348
R10241 CLK.n68 CLK 0.117348
R10242 CLK.n55 CLK 0.117348
R10243 CLK.n42 CLK 0.117348
R10244 CLK.n30 CLK 0.117348
R10245 CLK.n18 CLK 0.117348
R10246 CLK.n6 CLK 0.117348
R10247 CLK.n123 CLK.n122 0.063
R10248 CLK.n119 CLK.n118 0.063
R10249 CLK.n141 CLK.n140 0.063
R10250 CLK.n146 CLK.n145 0.063
R10251 CLK.n247 CLK 0.0454219
R10252 CLK.n248 CLK 0.0454219
R10253 CLK.n234 CLK 0.0454219
R10254 CLK.n235 CLK 0.0454219
R10255 CLK.n221 CLK 0.0454219
R10256 CLK.n222 CLK 0.0454219
R10257 CLK.n208 CLK 0.0454219
R10258 CLK.n209 CLK 0.0454219
R10259 CLK.n195 CLK 0.0454219
R10260 CLK.n196 CLK 0.0454219
R10261 CLK.n182 CLK 0.0454219
R10262 CLK.n183 CLK 0.0454219
R10263 CLK.n169 CLK 0.0454219
R10264 CLK.n170 CLK 0.0454219
R10265 CLK.n157 CLK 0.0454219
R10266 CLK.n158 CLK 0.0454219
R10267 CLK.n129 CLK 0.0454219
R10268 CLK.n132 CLK 0.0454219
R10269 CLK.n135 CLK 0.0454219
R10270 CLK.n126 CLK 0.0454219
R10271 CLK.n107 CLK 0.0454219
R10272 CLK.n108 CLK 0.0454219
R10273 CLK.n94 CLK 0.0454219
R10274 CLK.n95 CLK 0.0454219
R10275 CLK.n81 CLK 0.0454219
R10276 CLK.n82 CLK 0.0454219
R10277 CLK.n68 CLK 0.0454219
R10278 CLK.n69 CLK 0.0454219
R10279 CLK.n55 CLK 0.0454219
R10280 CLK.n56 CLK 0.0454219
R10281 CLK.n42 CLK 0.0454219
R10282 CLK.n43 CLK 0.0454219
R10283 CLK.n30 CLK 0.0454219
R10284 CLK.n31 CLK 0.0454219
R10285 CLK.n18 CLK 0.0454219
R10286 CLK.n19 CLK 0.0454219
R10287 CLK.n6 CLK 0.0454219
R10288 CLK.n7 CLK 0.0454219
R10289 CLK.n252 CLK.n245 0.024
R10290 CLK.n252 CLK.n251 0.024
R10291 CLK.n239 CLK.n232 0.024
R10292 CLK.n239 CLK.n238 0.024
R10293 CLK.n226 CLK.n219 0.024
R10294 CLK.n226 CLK.n225 0.024
R10295 CLK.n213 CLK.n206 0.024
R10296 CLK.n213 CLK.n212 0.024
R10297 CLK.n200 CLK.n193 0.024
R10298 CLK.n200 CLK.n199 0.024
R10299 CLK.n187 CLK.n180 0.024
R10300 CLK.n187 CLK.n186 0.024
R10301 CLK.n174 CLK.n167 0.024
R10302 CLK.n174 CLK.n173 0.024
R10303 CLK.n162 CLK.n155 0.024
R10304 CLK.n162 CLK.n161 0.024
R10305 CLK.n112 CLK.n105 0.024
R10306 CLK.n112 CLK.n111 0.024
R10307 CLK.n99 CLK.n92 0.024
R10308 CLK.n99 CLK.n98 0.024
R10309 CLK.n86 CLK.n79 0.024
R10310 CLK.n86 CLK.n85 0.024
R10311 CLK.n73 CLK.n66 0.024
R10312 CLK.n73 CLK.n72 0.024
R10313 CLK.n60 CLK.n53 0.024
R10314 CLK.n60 CLK.n59 0.024
R10315 CLK.n47 CLK.n40 0.024
R10316 CLK.n47 CLK.n46 0.024
R10317 CLK.n35 CLK.n28 0.024
R10318 CLK.n35 CLK.n34 0.024
R10319 CLK.n23 CLK.n16 0.024
R10320 CLK.n23 CLK.n22 0.024
R10321 CLK.n11 CLK.n4 0.024
R10322 CLK.n11 CLK.n10 0.024
R10323 CLK.n150 CLK.n149 0.024
R10324 CLK CLK.n253 0.0232879
R10325 CLK.n243 CLK.n242 0.0216397
R10326 CLK.n243 CLK 0.0216397
R10327 CLK.n230 CLK.n229 0.0216397
R10328 CLK.n230 CLK 0.0216397
R10329 CLK.n217 CLK.n216 0.0216397
R10330 CLK.n217 CLK 0.0216397
R10331 CLK.n204 CLK.n203 0.0216397
R10332 CLK.n204 CLK 0.0216397
R10333 CLK.n191 CLK.n190 0.0216397
R10334 CLK.n191 CLK 0.0216397
R10335 CLK.n178 CLK.n177 0.0216397
R10336 CLK.n178 CLK 0.0216397
R10337 CLK.n165 CLK.n164 0.0216397
R10338 CLK.n165 CLK 0.0216397
R10339 CLK.n153 CLK.n152 0.0216397
R10340 CLK.n153 CLK 0.0216397
R10341 CLK.n103 CLK.n102 0.0216397
R10342 CLK.n103 CLK 0.0216397
R10343 CLK.n90 CLK.n89 0.0216397
R10344 CLK.n90 CLK 0.0216397
R10345 CLK.n77 CLK.n76 0.0216397
R10346 CLK.n77 CLK 0.0216397
R10347 CLK.n64 CLK.n63 0.0216397
R10348 CLK.n64 CLK 0.0216397
R10349 CLK.n51 CLK.n50 0.0216397
R10350 CLK.n51 CLK 0.0216397
R10351 CLK.n38 CLK.n37 0.0216397
R10352 CLK.n38 CLK 0.0216397
R10353 CLK.n26 CLK.n25 0.0216397
R10354 CLK.n26 CLK 0.0216397
R10355 CLK.n14 CLK.n13 0.0216397
R10356 CLK.n14 CLK 0.0216397
R10357 CLK.n2 CLK.n1 0.0216397
R10358 CLK.n2 CLK 0.0216397
R10359 CLK.n121 CLK.n120 0.0107679
R10360 CLK.n120 CLK 0.0107679
R10361 CLK.n117 CLK.n116 0.0107679
R10362 CLK.n116 CLK 0.0107679
R10363 CLK.n139 CLK.n138 0.0107679
R10364 CLK.n138 CLK 0.0107679
R10365 CLK.n144 CLK.n143 0.0107679
R10366 CLK.n143 CLK 0.0107679
R10367 CLK.n250 CLK 0.00441667
R10368 CLK.n237 CLK 0.00441667
R10369 CLK.n224 CLK 0.00441667
R10370 CLK.n211 CLK 0.00441667
R10371 CLK.n198 CLK 0.00441667
R10372 CLK.n185 CLK 0.00441667
R10373 CLK.n172 CLK 0.00441667
R10374 CLK.n160 CLK 0.00441667
R10375 CLK.n110 CLK 0.00441667
R10376 CLK.n97 CLK 0.00441667
R10377 CLK.n84 CLK 0.00441667
R10378 CLK.n71 CLK 0.00441667
R10379 CLK.n58 CLK 0.00441667
R10380 CLK.n45 CLK 0.00441667
R10381 CLK.n33 CLK 0.00441667
R10382 CLK.n21 CLK 0.00441667
R10383 CLK.n9 CLK 0.00441667
R10384 CLK.n250 CLK 0.00406061
R10385 CLK.n237 CLK 0.00406061
R10386 CLK.n224 CLK 0.00406061
R10387 CLK.n211 CLK 0.00406061
R10388 CLK.n198 CLK 0.00406061
R10389 CLK.n185 CLK 0.00406061
R10390 CLK.n172 CLK 0.00406061
R10391 CLK.n160 CLK 0.00406061
R10392 CLK.n110 CLK 0.00406061
R10393 CLK.n97 CLK 0.00406061
R10394 CLK.n84 CLK 0.00406061
R10395 CLK.n71 CLK 0.00406061
R10396 CLK.n58 CLK 0.00406061
R10397 CLK.n45 CLK 0.00406061
R10398 CLK.n33 CLK 0.00406061
R10399 CLK.n21 CLK 0.00406061
R10400 CLK.n9 CLK 0.00406061
R10401 CLK.n254 CLK 0.00128333
R10402 CLK.n254 CLK 0.00121212
R10403 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 169.46
R10404 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 168.089
R10405 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 167.809
R10406 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 150.293
R10407 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 73.6304
R10408 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 60.4568
R10409 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 12.0358
R10410 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 11.4489
R10411 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.981478
R10412 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 0.788543
R10413 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.769522
R10414 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 0.720633
R10415 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 0.682565
R10416 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.580578
R10417 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 0.55213
R10418 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 0.470609
R10419 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.447191
R10420 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.428234
R10421 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.1255
R10422 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.1255
R10423 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 0.063
R10424 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 0.063
R10425 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.063
R10426 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 0.063
R10427 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 0.063
R10428 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 0.0435206
R10429 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 0.0107679
R10430 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.0107679
R10431 Nand_Gate_4.A.n33 Nand_Gate_4.A.t1 169.46
R10432 Nand_Gate_4.A.n35 Nand_Gate_4.A.t3 167.809
R10433 Nand_Gate_4.A.n33 Nand_Gate_4.A.t0 167.809
R10434 Nand_Gate_4.A Nand_Gate_4.A.t4 158.585
R10435 Nand_Gate_4.A.n21 Nand_Gate_4.A.t8 150.293
R10436 Nand_Gate_4.A.t4 Nand_Gate_4.A.n2 150.293
R10437 Nand_Gate_4.A.n14 Nand_Gate_4.A.t7 150.273
R10438 Nand_Gate_4.A.n8 Nand_Gate_4.A.t11 150.273
R10439 Nand_Gate_4.A.n12 Nand_Gate_4.A.t9 73.6406
R10440 Nand_Gate_4.A.n6 Nand_Gate_4.A.t5 73.6406
R10441 Nand_Gate_4.A.n23 Nand_Gate_4.A.t6 73.6304
R10442 Nand_Gate_4.A.n0 Nand_Gate_4.A.t10 73.6304
R10443 Nand_Gate_4.A.n4 Nand_Gate_4.A.t2 60.3809
R10444 Nand_Gate_4.A.n27 Nand_Gate_4.A.n26 14.3097
R10445 Nand_Gate_4.A.n34 Nand_Gate_4.A.n33 11.4489
R10446 Nand_Gate_4.A.n36 Nand_Gate_4.A.n35 8.21389
R10447 Nand_Gate_4.A.n18 Nand_Gate_4.A.n11 8.1418
R10448 Nand_Gate_4.A.n29 Nand_Gate_4.A.n28 5.61191
R10449 Nand_Gate_4.A.n29 Nand_Gate_4.A 5.35402
R10450 Nand_Gate_4.A.n30 Nand_Gate_4.A.n29 4.563
R10451 Nand_Gate_4.A.n18 Nand_Gate_4.A.n17 4.5005
R10452 Nand_Gate_4.A.n28 Nand_Gate_4.A 1.83746
R10453 Nand_Gate_4.A.n20 Nand_Gate_4.A.n19 1.62007
R10454 Nand_Gate_4.A.n2 Nand_Gate_4.A.n1 1.19615
R10455 Nand_Gate_4.A.n5 Nand_Gate_4.A 1.08746
R10456 Nand_Gate_4.A.n20 Nand_Gate_4.A 1.01739
R10457 Nand_Gate_4.A.n13 Nand_Gate_4.A 0.851043
R10458 Nand_Gate_4.A.n7 Nand_Gate_4.A 0.851043
R10459 Nand_Gate_4.A.n4 Nand_Gate_4.A 0.848156
R10460 Nand_Gate_4.A.n32 Nand_Gate_4.A.n31 0.788543
R10461 Nand_Gate_4.A.n22 Nand_Gate_4.A 0.769522
R10462 Nand_Gate_4.A.n5 Nand_Gate_4.A.n4 0.682565
R10463 Nand_Gate_4.A.n31 Nand_Gate_4.A 0.65675
R10464 Nand_Gate_4.A.n22 Nand_Gate_4.A.n21 0.55213
R10465 Nand_Gate_4.A.n16 Nand_Gate_4.A.n15 0.55213
R10466 Nand_Gate_4.A.n10 Nand_Gate_4.A.n9 0.55213
R10467 Nand_Gate_4.A.n16 Nand_Gate_4.A 0.486828
R10468 Nand_Gate_4.A.n10 Nand_Gate_4.A 0.486828
R10469 Nand_Gate_4.A.n25 Nand_Gate_4.A.n24 0.470609
R10470 Nand_Gate_4.A.n13 Nand_Gate_4.A.n12 0.470609
R10471 Nand_Gate_4.A.n7 Nand_Gate_4.A.n6 0.470609
R10472 Nand_Gate_4.A.n21 Nand_Gate_4.A 0.447191
R10473 Nand_Gate_4.A.n2 Nand_Gate_4.A 0.447191
R10474 Nand_Gate_4.A.n25 Nand_Gate_4.A 0.428234
R10475 Nand_Gate_4.A.n36 Nand_Gate_4.A.n3 0.425067
R10476 Nand_Gate_4.A Nand_Gate_4.A.n36 0.39003
R10477 Nand_Gate_4.A.n35 Nand_Gate_4.A.n34 0.280391
R10478 Nand_Gate_4.A.n34 Nand_Gate_4.A.n32 0.262643
R10479 Nand_Gate_4.A.n12 Nand_Gate_4.A 0.217464
R10480 Nand_Gate_4.A.n6 Nand_Gate_4.A 0.217464
R10481 Nand_Gate_4.A.n24 Nand_Gate_4.A 0.1255
R10482 Nand_Gate_4.A.n15 Nand_Gate_4.A 0.1255
R10483 Nand_Gate_4.A.n9 Nand_Gate_4.A 0.1255
R10484 Nand_Gate_4.A.n32 Nand_Gate_4.A 0.1255
R10485 Nand_Gate_4.A.n1 Nand_Gate_4.A 0.1255
R10486 Nand_Gate_4.A.n26 Nand_Gate_4.A.n22 0.063
R10487 Nand_Gate_4.A.n26 Nand_Gate_4.A.n25 0.063
R10488 Nand_Gate_4.A.n17 Nand_Gate_4.A.n13 0.063
R10489 Nand_Gate_4.A.n17 Nand_Gate_4.A.n16 0.063
R10490 Nand_Gate_4.A.n11 Nand_Gate_4.A.n7 0.063
R10491 Nand_Gate_4.A.n11 Nand_Gate_4.A.n10 0.063
R10492 Nand_Gate_4.A.n28 Nand_Gate_4.A.n27 0.063
R10493 Nand_Gate_4.A.n27 Nand_Gate_4.A.n20 0.063
R10494 Nand_Gate_4.A.n30 Nand_Gate_4.A.n5 0.063
R10495 Nand_Gate_4.A.n31 Nand_Gate_4.A.n30 0.063
R10496 Nand_Gate_4.A.n32 Nand_Gate_4.A 0.063
R10497 Nand_Gate_4.A Nand_Gate_4.A.n18 0.0512812
R10498 Nand_Gate_4.A.n15 Nand_Gate_4.A.n14 0.0216397
R10499 Nand_Gate_4.A.n14 Nand_Gate_4.A 0.0216397
R10500 Nand_Gate_4.A.n9 Nand_Gate_4.A.n8 0.0216397
R10501 Nand_Gate_4.A.n8 Nand_Gate_4.A 0.0216397
R10502 Nand_Gate_4.A.n19 Nand_Gate_4.A 0.0168043
R10503 Nand_Gate_4.A.n19 Nand_Gate_4.A 0.0122188
R10504 Nand_Gate_4.A.n24 Nand_Gate_4.A.n23 0.0107679
R10505 Nand_Gate_4.A.n23 Nand_Gate_4.A 0.0107679
R10506 Nand_Gate_4.A.n1 Nand_Gate_4.A.n0 0.0107679
R10507 Nand_Gate_4.A.n0 Nand_Gate_4.A 0.0107679
R10508 Nand_Gate_4.A.n3 Nand_Gate_4.A 0.00441667
R10509 Nand_Gate_4.A.n3 Nand_Gate_4.A 0.00406061
R10510 VDD.n311 VDD.n310 55259.3
R10511 VDD.n311 VDD.n309 49126.7
R10512 VDD.n317 VDD.n310 32898.4
R10513 VDD.n318 VDD.n317 29988.1
R10514 VDD.n319 VDD.n318 29374.8
R10515 VDD.n313 VDD.n312 27016.6
R10516 VDD.n319 VDD.n309 25484.7
R10517 VDD.n312 VDD.n306 24146.4
R10518 VDD.n316 VDD.n313 16939.4
R10519 VDD.n316 VDD.n308 15719.7
R10520 VDD.n320 VDD.n308 15072.6
R10521 VDD.n320 VDD.n306 13411.9
R10522 VDD.n338 VDD.n289 12650.1
R10523 VDD.n292 VDD.n289 12650.1
R10524 VDD.n338 VDD.n290 12650.1
R10525 VDD.n330 VDD.n299 10684.6
R10526 VDD.n335 VDD.n294 10684.6
R10527 VDD.n335 VDD.n295 10684.6
R10528 VDD.n303 VDD.n302 10167.6
R10529 VDD.n302 VDD.n300 10167.6
R10530 VDD.n314 VDD.n305 6073.28
R10531 VDD.n322 VDD.n305 5168.82
R10532 VDD.n315 VDD.n314 4059.29
R10533 VDD.n315 VDD.n307 3849.04
R10534 VDD.n321 VDD.n307 3690.92
R10535 VDD.n322 VDD.n321 2993.95
R10536 VDD.n291 VDD.n288 2427.48
R10537 VDD.n291 VDD.n287 2427.48
R10538 VDD.n339 VDD.n288 2349.78
R10539 VDD.n339 VDD.n287 2349.78
R10540 VDD.n293 VDD.n292 2128.85
R10541 VDD.n334 VDD.n333 2051.01
R10542 VDD.n331 VDD.n298 2051.01
R10543 VDD.n334 VDD.n296 1973.31
R10544 VDD.n327 VDD.n298 1973.31
R10545 VDD.n326 VDD.n297 1952
R10546 VDD.n332 VDD.n297 1952
R10547 VDD.n7646 VDD.n7633 1084.97
R10548 VDD.n7646 VDD.n7634 1084.97
R10549 VDD.n7653 VDD.n7634 1084.97
R10550 VDD.n7653 VDD.n7633 1084.97
R10551 VDD.n7656 VDD.n7623 1084.97
R10552 VDD.n7656 VDD.n7624 1084.97
R10553 VDD.n7663 VDD.n7624 1084.97
R10554 VDD.n7663 VDD.n7623 1084.97
R10555 VDD.n7666 VDD.n7612 1084.97
R10556 VDD.n7666 VDD.n7613 1084.97
R10557 VDD.n7673 VDD.n7613 1084.97
R10558 VDD.n7673 VDD.n7612 1084.97
R10559 VDD.n7676 VDD.n7599 1084.97
R10560 VDD.n7676 VDD.n7600 1084.97
R10561 VDD.n7683 VDD.n7600 1084.97
R10562 VDD.n7683 VDD.n7599 1084.97
R10563 VDD.n7686 VDD.n7587 1084.97
R10564 VDD.n7686 VDD.n7588 1084.97
R10565 VDD.n7693 VDD.n7588 1084.97
R10566 VDD.n7693 VDD.n7587 1084.97
R10567 VDD.n7703 VDD.n7571 1084.97
R10568 VDD.n7703 VDD.n7572 1084.97
R10569 VDD.n7710 VDD.n7572 1084.97
R10570 VDD.n7710 VDD.n7571 1084.97
R10571 VDD.n7713 VDD.n7562 1084.97
R10572 VDD.n7713 VDD.n7563 1084.97
R10573 VDD.n7720 VDD.n7563 1084.97
R10574 VDD.n7720 VDD.n7562 1084.97
R10575 VDD.n7728 VDD.n7724 1084.97
R10576 VDD.n7724 VDD.n3 1084.97
R10577 VDD.n7723 VDD.n3 1084.97
R10578 VDD.n7728 VDD.n7723 1084.97
R10579 VDD.n7554 VDD.n8 1084.97
R10580 VDD.n7554 VDD.n9 1084.97
R10581 VDD.n7547 VDD.n9 1084.97
R10582 VDD.n7547 VDD.n8 1084.97
R10583 VDD.n7544 VDD.n17 1084.97
R10584 VDD.n7544 VDD.n18 1084.97
R10585 VDD.n7537 VDD.n18 1084.97
R10586 VDD.n7537 VDD.n17 1084.97
R10587 VDD.n7534 VDD.n30 1084.97
R10588 VDD.n7534 VDD.n31 1084.97
R10589 VDD.n7527 VDD.n31 1084.97
R10590 VDD.n7527 VDD.n30 1084.97
R10591 VDD.n7649 VDD.n7648 1084.97
R10592 VDD.n7648 VDD.n7642 1084.97
R10593 VDD.n7642 VDD.n7632 1084.97
R10594 VDD.n7649 VDD.n7632 1084.97
R10595 VDD.n7659 VDD.n7658 1084.97
R10596 VDD.n7658 VDD.n7629 1084.97
R10597 VDD.n7629 VDD.n7622 1084.97
R10598 VDD.n7659 VDD.n7622 1084.97
R10599 VDD.n7669 VDD.n7668 1084.97
R10600 VDD.n7668 VDD.n7619 1084.97
R10601 VDD.n7619 VDD.n7611 1084.97
R10602 VDD.n7669 VDD.n7611 1084.97
R10603 VDD.n7679 VDD.n7678 1084.97
R10604 VDD.n7678 VDD.n7608 1084.97
R10605 VDD.n7608 VDD.n7598 1084.97
R10606 VDD.n7679 VDD.n7598 1084.97
R10607 VDD.n7689 VDD.n7688 1084.97
R10608 VDD.n7688 VDD.n7595 1084.97
R10609 VDD.n7595 VDD.n7586 1084.97
R10610 VDD.n7689 VDD.n7586 1084.97
R10611 VDD.n7696 VDD.n7583 1084.97
R10612 VDD.n7696 VDD.n7584 1084.97
R10613 VDD.n7700 VDD.n7584 1084.97
R10614 VDD.n7700 VDD.n7583 1084.97
R10615 VDD.n7706 VDD.n7705 1084.97
R10616 VDD.n7705 VDD.n7580 1084.97
R10617 VDD.n7580 VDD.n7570 1084.97
R10618 VDD.n7706 VDD.n7570 1084.97
R10619 VDD.n7716 VDD.n7715 1084.97
R10620 VDD.n7715 VDD.n7567 1084.97
R10621 VDD.n7567 VDD.n7561 1084.97
R10622 VDD.n7716 VDD.n7561 1084.97
R10623 VDD.n7729 VDD.n6 1084.97
R10624 VDD.n7560 VDD.n6 1084.97
R10625 VDD.n7560 VDD.n5 1084.97
R10626 VDD.n7729 VDD.n5 1084.97
R10627 VDD.n7550 VDD.n7 1084.97
R10628 VDD.n13 VDD.n7 1084.97
R10629 VDD.n7549 VDD.n13 1084.97
R10630 VDD.n7550 VDD.n7549 1084.97
R10631 VDD.n7540 VDD.n16 1084.97
R10632 VDD.n26 VDD.n16 1084.97
R10633 VDD.n7539 VDD.n26 1084.97
R10634 VDD.n7540 VDD.n7539 1084.97
R10635 VDD.n7530 VDD.n29 1084.97
R10636 VDD.n36 VDD.n29 1084.97
R10637 VDD.n7529 VDD.n36 1084.97
R10638 VDD.n7530 VDD.n7529 1084.97
R10639 VDD.n43 VDD.n39 1084.97
R10640 VDD.n7524 VDD.n39 1084.97
R10641 VDD.n7524 VDD.n40 1084.97
R10642 VDD.n1779 VDD.n1766 1084.97
R10643 VDD.n1779 VDD.n1767 1084.97
R10644 VDD.n1786 VDD.n1767 1084.97
R10645 VDD.n1786 VDD.n1766 1084.97
R10646 VDD.n1789 VDD.n1756 1084.97
R10647 VDD.n1789 VDD.n1757 1084.97
R10648 VDD.n1796 VDD.n1757 1084.97
R10649 VDD.n1796 VDD.n1756 1084.97
R10650 VDD.n1799 VDD.n1745 1084.97
R10651 VDD.n1799 VDD.n1746 1084.97
R10652 VDD.n1806 VDD.n1746 1084.97
R10653 VDD.n1806 VDD.n1745 1084.97
R10654 VDD.n1809 VDD.n1732 1084.97
R10655 VDD.n1809 VDD.n1733 1084.97
R10656 VDD.n1816 VDD.n1733 1084.97
R10657 VDD.n1816 VDD.n1732 1084.97
R10658 VDD.n1819 VDD.n1720 1084.97
R10659 VDD.n1819 VDD.n1721 1084.97
R10660 VDD.n1826 VDD.n1721 1084.97
R10661 VDD.n1826 VDD.n1720 1084.97
R10662 VDD.n1836 VDD.n1704 1084.97
R10663 VDD.n1836 VDD.n1705 1084.97
R10664 VDD.n1843 VDD.n1705 1084.97
R10665 VDD.n1843 VDD.n1704 1084.97
R10666 VDD.n1846 VDD.n1694 1084.97
R10667 VDD.n1846 VDD.n1695 1084.97
R10668 VDD.n1853 VDD.n1695 1084.97
R10669 VDD.n1853 VDD.n1694 1084.97
R10670 VDD.n1856 VDD.n1683 1084.97
R10671 VDD.n1856 VDD.n1684 1084.97
R10672 VDD.n1863 VDD.n1684 1084.97
R10673 VDD.n1863 VDD.n1683 1084.97
R10674 VDD.n1866 VDD.n1670 1084.97
R10675 VDD.n1866 VDD.n1671 1084.97
R10676 VDD.n1873 VDD.n1671 1084.97
R10677 VDD.n1873 VDD.n1670 1084.97
R10678 VDD.n1876 VDD.n1660 1084.97
R10679 VDD.n1876 VDD.n1661 1084.97
R10680 VDD.n1883 VDD.n1661 1084.97
R10681 VDD.n1883 VDD.n1660 1084.97
R10682 VDD.n1886 VDD.n1649 1084.97
R10683 VDD.n1886 VDD.n1650 1084.97
R10684 VDD.n1893 VDD.n1650 1084.97
R10685 VDD.n1893 VDD.n1649 1084.97
R10686 VDD.n1782 VDD.n1781 1084.97
R10687 VDD.n1781 VDD.n1775 1084.97
R10688 VDD.n1775 VDD.n1765 1084.97
R10689 VDD.n1782 VDD.n1765 1084.97
R10690 VDD.n1792 VDD.n1791 1084.97
R10691 VDD.n1791 VDD.n1762 1084.97
R10692 VDD.n1762 VDD.n1755 1084.97
R10693 VDD.n1792 VDD.n1755 1084.97
R10694 VDD.n1802 VDD.n1801 1084.97
R10695 VDD.n1801 VDD.n1752 1084.97
R10696 VDD.n1752 VDD.n1744 1084.97
R10697 VDD.n1802 VDD.n1744 1084.97
R10698 VDD.n1812 VDD.n1811 1084.97
R10699 VDD.n1811 VDD.n1741 1084.97
R10700 VDD.n1741 VDD.n1731 1084.97
R10701 VDD.n1812 VDD.n1731 1084.97
R10702 VDD.n1822 VDD.n1821 1084.97
R10703 VDD.n1821 VDD.n1728 1084.97
R10704 VDD.n1728 VDD.n1719 1084.97
R10705 VDD.n1822 VDD.n1719 1084.97
R10706 VDD.n1829 VDD.n1716 1084.97
R10707 VDD.n1829 VDD.n1717 1084.97
R10708 VDD.n1833 VDD.n1717 1084.97
R10709 VDD.n1833 VDD.n1716 1084.97
R10710 VDD.n1839 VDD.n1838 1084.97
R10711 VDD.n1838 VDD.n1713 1084.97
R10712 VDD.n1713 VDD.n1703 1084.97
R10713 VDD.n1839 VDD.n1703 1084.97
R10714 VDD.n1849 VDD.n1848 1084.97
R10715 VDD.n1848 VDD.n1700 1084.97
R10716 VDD.n1700 VDD.n1693 1084.97
R10717 VDD.n1849 VDD.n1693 1084.97
R10718 VDD.n1859 VDD.n1858 1084.97
R10719 VDD.n1858 VDD.n1690 1084.97
R10720 VDD.n1690 VDD.n1682 1084.97
R10721 VDD.n1859 VDD.n1682 1084.97
R10722 VDD.n1869 VDD.n1868 1084.97
R10723 VDD.n1868 VDD.n1679 1084.97
R10724 VDD.n1679 VDD.n1669 1084.97
R10725 VDD.n1869 VDD.n1669 1084.97
R10726 VDD.n1879 VDD.n1878 1084.97
R10727 VDD.n1878 VDD.n1666 1084.97
R10728 VDD.n1666 VDD.n1659 1084.97
R10729 VDD.n1879 VDD.n1659 1084.97
R10730 VDD.n1889 VDD.n1888 1084.97
R10731 VDD.n1888 VDD.n1656 1084.97
R10732 VDD.n1656 VDD.n1648 1084.97
R10733 VDD.n1889 VDD.n1648 1084.97
R10734 VDD.n1646 VDD.n1645 1084.97
R10735 VDD.n1896 VDD.n1645 1084.97
R10736 VDD.n1896 VDD.n1643 1084.97
R10737 VDD.n1519 VDD.n1506 1084.97
R10738 VDD.n1519 VDD.n1507 1084.97
R10739 VDD.n1526 VDD.n1507 1084.97
R10740 VDD.n1526 VDD.n1506 1084.97
R10741 VDD.n1529 VDD.n1496 1084.97
R10742 VDD.n1529 VDD.n1497 1084.97
R10743 VDD.n1536 VDD.n1497 1084.97
R10744 VDD.n1536 VDD.n1496 1084.97
R10745 VDD.n1539 VDD.n1485 1084.97
R10746 VDD.n1539 VDD.n1486 1084.97
R10747 VDD.n1546 VDD.n1486 1084.97
R10748 VDD.n1546 VDD.n1485 1084.97
R10749 VDD.n1549 VDD.n1472 1084.97
R10750 VDD.n1549 VDD.n1473 1084.97
R10751 VDD.n1556 VDD.n1473 1084.97
R10752 VDD.n1556 VDD.n1472 1084.97
R10753 VDD.n1559 VDD.n1460 1084.97
R10754 VDD.n1559 VDD.n1461 1084.97
R10755 VDD.n1566 VDD.n1461 1084.97
R10756 VDD.n1566 VDD.n1460 1084.97
R10757 VDD.n1576 VDD.n1444 1084.97
R10758 VDD.n1576 VDD.n1445 1084.97
R10759 VDD.n1583 VDD.n1445 1084.97
R10760 VDD.n1583 VDD.n1444 1084.97
R10761 VDD.n1586 VDD.n1434 1084.97
R10762 VDD.n1586 VDD.n1435 1084.97
R10763 VDD.n1593 VDD.n1435 1084.97
R10764 VDD.n1593 VDD.n1434 1084.97
R10765 VDD.n1596 VDD.n1423 1084.97
R10766 VDD.n1596 VDD.n1424 1084.97
R10767 VDD.n1603 VDD.n1424 1084.97
R10768 VDD.n1603 VDD.n1423 1084.97
R10769 VDD.n1606 VDD.n1410 1084.97
R10770 VDD.n1606 VDD.n1411 1084.97
R10771 VDD.n1613 VDD.n1411 1084.97
R10772 VDD.n1613 VDD.n1410 1084.97
R10773 VDD.n1616 VDD.n1400 1084.97
R10774 VDD.n1616 VDD.n1401 1084.97
R10775 VDD.n1623 VDD.n1401 1084.97
R10776 VDD.n1623 VDD.n1400 1084.97
R10777 VDD.n1626 VDD.n1389 1084.97
R10778 VDD.n1626 VDD.n1390 1084.97
R10779 VDD.n1633 VDD.n1390 1084.97
R10780 VDD.n1633 VDD.n1389 1084.97
R10781 VDD.n1522 VDD.n1521 1084.97
R10782 VDD.n1521 VDD.n1515 1084.97
R10783 VDD.n1515 VDD.n1505 1084.97
R10784 VDD.n1522 VDD.n1505 1084.97
R10785 VDD.n1532 VDD.n1531 1084.97
R10786 VDD.n1531 VDD.n1502 1084.97
R10787 VDD.n1502 VDD.n1495 1084.97
R10788 VDD.n1532 VDD.n1495 1084.97
R10789 VDD.n1542 VDD.n1541 1084.97
R10790 VDD.n1541 VDD.n1492 1084.97
R10791 VDD.n1492 VDD.n1484 1084.97
R10792 VDD.n1542 VDD.n1484 1084.97
R10793 VDD.n1552 VDD.n1551 1084.97
R10794 VDD.n1551 VDD.n1481 1084.97
R10795 VDD.n1481 VDD.n1471 1084.97
R10796 VDD.n1552 VDD.n1471 1084.97
R10797 VDD.n1562 VDD.n1561 1084.97
R10798 VDD.n1561 VDD.n1468 1084.97
R10799 VDD.n1468 VDD.n1459 1084.97
R10800 VDD.n1562 VDD.n1459 1084.97
R10801 VDD.n1569 VDD.n1456 1084.97
R10802 VDD.n1569 VDD.n1457 1084.97
R10803 VDD.n1573 VDD.n1457 1084.97
R10804 VDD.n1573 VDD.n1456 1084.97
R10805 VDD.n1579 VDD.n1578 1084.97
R10806 VDD.n1578 VDD.n1453 1084.97
R10807 VDD.n1453 VDD.n1443 1084.97
R10808 VDD.n1579 VDD.n1443 1084.97
R10809 VDD.n1589 VDD.n1588 1084.97
R10810 VDD.n1588 VDD.n1440 1084.97
R10811 VDD.n1440 VDD.n1433 1084.97
R10812 VDD.n1589 VDD.n1433 1084.97
R10813 VDD.n1599 VDD.n1598 1084.97
R10814 VDD.n1598 VDD.n1430 1084.97
R10815 VDD.n1430 VDD.n1422 1084.97
R10816 VDD.n1599 VDD.n1422 1084.97
R10817 VDD.n1609 VDD.n1608 1084.97
R10818 VDD.n1608 VDD.n1419 1084.97
R10819 VDD.n1419 VDD.n1409 1084.97
R10820 VDD.n1609 VDD.n1409 1084.97
R10821 VDD.n1619 VDD.n1618 1084.97
R10822 VDD.n1618 VDD.n1406 1084.97
R10823 VDD.n1406 VDD.n1399 1084.97
R10824 VDD.n1619 VDD.n1399 1084.97
R10825 VDD.n1629 VDD.n1628 1084.97
R10826 VDD.n1628 VDD.n1396 1084.97
R10827 VDD.n1396 VDD.n1388 1084.97
R10828 VDD.n1629 VDD.n1388 1084.97
R10829 VDD.n1386 VDD.n1385 1084.97
R10830 VDD.n1636 VDD.n1385 1084.97
R10831 VDD.n1636 VDD.n1383 1084.97
R10832 VDD.n1259 VDD.n1246 1084.97
R10833 VDD.n1259 VDD.n1247 1084.97
R10834 VDD.n1266 VDD.n1247 1084.97
R10835 VDD.n1266 VDD.n1246 1084.97
R10836 VDD.n1269 VDD.n1236 1084.97
R10837 VDD.n1269 VDD.n1237 1084.97
R10838 VDD.n1276 VDD.n1237 1084.97
R10839 VDD.n1276 VDD.n1236 1084.97
R10840 VDD.n1279 VDD.n1225 1084.97
R10841 VDD.n1279 VDD.n1226 1084.97
R10842 VDD.n1286 VDD.n1226 1084.97
R10843 VDD.n1286 VDD.n1225 1084.97
R10844 VDD.n1289 VDD.n1212 1084.97
R10845 VDD.n1289 VDD.n1213 1084.97
R10846 VDD.n1296 VDD.n1213 1084.97
R10847 VDD.n1296 VDD.n1212 1084.97
R10848 VDD.n1299 VDD.n1200 1084.97
R10849 VDD.n1299 VDD.n1201 1084.97
R10850 VDD.n1306 VDD.n1201 1084.97
R10851 VDD.n1306 VDD.n1200 1084.97
R10852 VDD.n1316 VDD.n1184 1084.97
R10853 VDD.n1316 VDD.n1185 1084.97
R10854 VDD.n1323 VDD.n1185 1084.97
R10855 VDD.n1323 VDD.n1184 1084.97
R10856 VDD.n1326 VDD.n1174 1084.97
R10857 VDD.n1326 VDD.n1175 1084.97
R10858 VDD.n1333 VDD.n1175 1084.97
R10859 VDD.n1333 VDD.n1174 1084.97
R10860 VDD.n1336 VDD.n1163 1084.97
R10861 VDD.n1336 VDD.n1164 1084.97
R10862 VDD.n1343 VDD.n1164 1084.97
R10863 VDD.n1343 VDD.n1163 1084.97
R10864 VDD.n1346 VDD.n1150 1084.97
R10865 VDD.n1346 VDD.n1151 1084.97
R10866 VDD.n1353 VDD.n1151 1084.97
R10867 VDD.n1353 VDD.n1150 1084.97
R10868 VDD.n1356 VDD.n1140 1084.97
R10869 VDD.n1356 VDD.n1141 1084.97
R10870 VDD.n1363 VDD.n1141 1084.97
R10871 VDD.n1363 VDD.n1140 1084.97
R10872 VDD.n1366 VDD.n1129 1084.97
R10873 VDD.n1366 VDD.n1130 1084.97
R10874 VDD.n1373 VDD.n1130 1084.97
R10875 VDD.n1373 VDD.n1129 1084.97
R10876 VDD.n1262 VDD.n1261 1084.97
R10877 VDD.n1261 VDD.n1255 1084.97
R10878 VDD.n1255 VDD.n1245 1084.97
R10879 VDD.n1262 VDD.n1245 1084.97
R10880 VDD.n1272 VDD.n1271 1084.97
R10881 VDD.n1271 VDD.n1242 1084.97
R10882 VDD.n1242 VDD.n1235 1084.97
R10883 VDD.n1272 VDD.n1235 1084.97
R10884 VDD.n1282 VDD.n1281 1084.97
R10885 VDD.n1281 VDD.n1232 1084.97
R10886 VDD.n1232 VDD.n1224 1084.97
R10887 VDD.n1282 VDD.n1224 1084.97
R10888 VDD.n1292 VDD.n1291 1084.97
R10889 VDD.n1291 VDD.n1221 1084.97
R10890 VDD.n1221 VDD.n1211 1084.97
R10891 VDD.n1292 VDD.n1211 1084.97
R10892 VDD.n1302 VDD.n1301 1084.97
R10893 VDD.n1301 VDD.n1208 1084.97
R10894 VDD.n1208 VDD.n1199 1084.97
R10895 VDD.n1302 VDD.n1199 1084.97
R10896 VDD.n1309 VDD.n1196 1084.97
R10897 VDD.n1309 VDD.n1197 1084.97
R10898 VDD.n1313 VDD.n1197 1084.97
R10899 VDD.n1313 VDD.n1196 1084.97
R10900 VDD.n1319 VDD.n1318 1084.97
R10901 VDD.n1318 VDD.n1193 1084.97
R10902 VDD.n1193 VDD.n1183 1084.97
R10903 VDD.n1319 VDD.n1183 1084.97
R10904 VDD.n1329 VDD.n1328 1084.97
R10905 VDD.n1328 VDD.n1180 1084.97
R10906 VDD.n1180 VDD.n1173 1084.97
R10907 VDD.n1329 VDD.n1173 1084.97
R10908 VDD.n1339 VDD.n1338 1084.97
R10909 VDD.n1338 VDD.n1170 1084.97
R10910 VDD.n1170 VDD.n1162 1084.97
R10911 VDD.n1339 VDD.n1162 1084.97
R10912 VDD.n1349 VDD.n1348 1084.97
R10913 VDD.n1348 VDD.n1159 1084.97
R10914 VDD.n1159 VDD.n1149 1084.97
R10915 VDD.n1349 VDD.n1149 1084.97
R10916 VDD.n1359 VDD.n1358 1084.97
R10917 VDD.n1358 VDD.n1146 1084.97
R10918 VDD.n1146 VDD.n1139 1084.97
R10919 VDD.n1359 VDD.n1139 1084.97
R10920 VDD.n1369 VDD.n1368 1084.97
R10921 VDD.n1368 VDD.n1136 1084.97
R10922 VDD.n1136 VDD.n1128 1084.97
R10923 VDD.n1369 VDD.n1128 1084.97
R10924 VDD.n1126 VDD.n1125 1084.97
R10925 VDD.n1376 VDD.n1125 1084.97
R10926 VDD.n1376 VDD.n1123 1084.97
R10927 VDD.n999 VDD.n986 1084.97
R10928 VDD.n999 VDD.n987 1084.97
R10929 VDD.n1006 VDD.n987 1084.97
R10930 VDD.n1006 VDD.n986 1084.97
R10931 VDD.n1009 VDD.n976 1084.97
R10932 VDD.n1009 VDD.n977 1084.97
R10933 VDD.n1016 VDD.n977 1084.97
R10934 VDD.n1016 VDD.n976 1084.97
R10935 VDD.n1019 VDD.n965 1084.97
R10936 VDD.n1019 VDD.n966 1084.97
R10937 VDD.n1026 VDD.n966 1084.97
R10938 VDD.n1026 VDD.n965 1084.97
R10939 VDD.n1029 VDD.n952 1084.97
R10940 VDD.n1029 VDD.n953 1084.97
R10941 VDD.n1036 VDD.n953 1084.97
R10942 VDD.n1036 VDD.n952 1084.97
R10943 VDD.n1039 VDD.n940 1084.97
R10944 VDD.n1039 VDD.n941 1084.97
R10945 VDD.n1046 VDD.n941 1084.97
R10946 VDD.n1046 VDD.n940 1084.97
R10947 VDD.n1056 VDD.n924 1084.97
R10948 VDD.n1056 VDD.n925 1084.97
R10949 VDD.n1063 VDD.n925 1084.97
R10950 VDD.n1063 VDD.n924 1084.97
R10951 VDD.n1066 VDD.n914 1084.97
R10952 VDD.n1066 VDD.n915 1084.97
R10953 VDD.n1073 VDD.n915 1084.97
R10954 VDD.n1073 VDD.n914 1084.97
R10955 VDD.n1076 VDD.n903 1084.97
R10956 VDD.n1076 VDD.n904 1084.97
R10957 VDD.n1083 VDD.n904 1084.97
R10958 VDD.n1083 VDD.n903 1084.97
R10959 VDD.n1086 VDD.n890 1084.97
R10960 VDD.n1086 VDD.n891 1084.97
R10961 VDD.n1093 VDD.n891 1084.97
R10962 VDD.n1093 VDD.n890 1084.97
R10963 VDD.n1096 VDD.n880 1084.97
R10964 VDD.n1096 VDD.n881 1084.97
R10965 VDD.n1103 VDD.n881 1084.97
R10966 VDD.n1103 VDD.n880 1084.97
R10967 VDD.n1106 VDD.n869 1084.97
R10968 VDD.n1106 VDD.n870 1084.97
R10969 VDD.n1113 VDD.n870 1084.97
R10970 VDD.n1113 VDD.n869 1084.97
R10971 VDD.n1002 VDD.n1001 1084.97
R10972 VDD.n1001 VDD.n995 1084.97
R10973 VDD.n995 VDD.n985 1084.97
R10974 VDD.n1002 VDD.n985 1084.97
R10975 VDD.n1012 VDD.n1011 1084.97
R10976 VDD.n1011 VDD.n982 1084.97
R10977 VDD.n982 VDD.n975 1084.97
R10978 VDD.n1012 VDD.n975 1084.97
R10979 VDD.n1022 VDD.n1021 1084.97
R10980 VDD.n1021 VDD.n972 1084.97
R10981 VDD.n972 VDD.n964 1084.97
R10982 VDD.n1022 VDD.n964 1084.97
R10983 VDD.n1032 VDD.n1031 1084.97
R10984 VDD.n1031 VDD.n961 1084.97
R10985 VDD.n961 VDD.n951 1084.97
R10986 VDD.n1032 VDD.n951 1084.97
R10987 VDD.n1042 VDD.n1041 1084.97
R10988 VDD.n1041 VDD.n948 1084.97
R10989 VDD.n948 VDD.n939 1084.97
R10990 VDD.n1042 VDD.n939 1084.97
R10991 VDD.n1049 VDD.n936 1084.97
R10992 VDD.n1049 VDD.n937 1084.97
R10993 VDD.n1053 VDD.n937 1084.97
R10994 VDD.n1053 VDD.n936 1084.97
R10995 VDD.n1059 VDD.n1058 1084.97
R10996 VDD.n1058 VDD.n933 1084.97
R10997 VDD.n933 VDD.n923 1084.97
R10998 VDD.n1059 VDD.n923 1084.97
R10999 VDD.n1069 VDD.n1068 1084.97
R11000 VDD.n1068 VDD.n920 1084.97
R11001 VDD.n920 VDD.n913 1084.97
R11002 VDD.n1069 VDD.n913 1084.97
R11003 VDD.n1079 VDD.n1078 1084.97
R11004 VDD.n1078 VDD.n910 1084.97
R11005 VDD.n910 VDD.n902 1084.97
R11006 VDD.n1079 VDD.n902 1084.97
R11007 VDD.n1089 VDD.n1088 1084.97
R11008 VDD.n1088 VDD.n899 1084.97
R11009 VDD.n899 VDD.n889 1084.97
R11010 VDD.n1089 VDD.n889 1084.97
R11011 VDD.n1099 VDD.n1098 1084.97
R11012 VDD.n1098 VDD.n886 1084.97
R11013 VDD.n886 VDD.n879 1084.97
R11014 VDD.n1099 VDD.n879 1084.97
R11015 VDD.n1109 VDD.n1108 1084.97
R11016 VDD.n1108 VDD.n876 1084.97
R11017 VDD.n876 VDD.n868 1084.97
R11018 VDD.n1109 VDD.n868 1084.97
R11019 VDD.n866 VDD.n865 1084.97
R11020 VDD.n1116 VDD.n865 1084.97
R11021 VDD.n1116 VDD.n863 1084.97
R11022 VDD.n739 VDD.n726 1084.97
R11023 VDD.n739 VDD.n727 1084.97
R11024 VDD.n746 VDD.n727 1084.97
R11025 VDD.n746 VDD.n726 1084.97
R11026 VDD.n749 VDD.n716 1084.97
R11027 VDD.n749 VDD.n717 1084.97
R11028 VDD.n756 VDD.n717 1084.97
R11029 VDD.n756 VDD.n716 1084.97
R11030 VDD.n759 VDD.n705 1084.97
R11031 VDD.n759 VDD.n706 1084.97
R11032 VDD.n766 VDD.n706 1084.97
R11033 VDD.n766 VDD.n705 1084.97
R11034 VDD.n769 VDD.n692 1084.97
R11035 VDD.n769 VDD.n693 1084.97
R11036 VDD.n776 VDD.n693 1084.97
R11037 VDD.n776 VDD.n692 1084.97
R11038 VDD.n779 VDD.n680 1084.97
R11039 VDD.n779 VDD.n681 1084.97
R11040 VDD.n786 VDD.n681 1084.97
R11041 VDD.n786 VDD.n680 1084.97
R11042 VDD.n796 VDD.n664 1084.97
R11043 VDD.n796 VDD.n665 1084.97
R11044 VDD.n803 VDD.n665 1084.97
R11045 VDD.n803 VDD.n664 1084.97
R11046 VDD.n806 VDD.n654 1084.97
R11047 VDD.n806 VDD.n655 1084.97
R11048 VDD.n813 VDD.n655 1084.97
R11049 VDD.n813 VDD.n654 1084.97
R11050 VDD.n816 VDD.n643 1084.97
R11051 VDD.n816 VDD.n644 1084.97
R11052 VDD.n823 VDD.n644 1084.97
R11053 VDD.n823 VDD.n643 1084.97
R11054 VDD.n826 VDD.n630 1084.97
R11055 VDD.n826 VDD.n631 1084.97
R11056 VDD.n833 VDD.n631 1084.97
R11057 VDD.n833 VDD.n630 1084.97
R11058 VDD.n836 VDD.n620 1084.97
R11059 VDD.n836 VDD.n621 1084.97
R11060 VDD.n843 VDD.n621 1084.97
R11061 VDD.n843 VDD.n620 1084.97
R11062 VDD.n846 VDD.n609 1084.97
R11063 VDD.n846 VDD.n610 1084.97
R11064 VDD.n853 VDD.n610 1084.97
R11065 VDD.n853 VDD.n609 1084.97
R11066 VDD.n742 VDD.n741 1084.97
R11067 VDD.n741 VDD.n735 1084.97
R11068 VDD.n735 VDD.n725 1084.97
R11069 VDD.n742 VDD.n725 1084.97
R11070 VDD.n752 VDD.n751 1084.97
R11071 VDD.n751 VDD.n722 1084.97
R11072 VDD.n722 VDD.n715 1084.97
R11073 VDD.n752 VDD.n715 1084.97
R11074 VDD.n762 VDD.n761 1084.97
R11075 VDD.n761 VDD.n712 1084.97
R11076 VDD.n712 VDD.n704 1084.97
R11077 VDD.n762 VDD.n704 1084.97
R11078 VDD.n772 VDD.n771 1084.97
R11079 VDD.n771 VDD.n701 1084.97
R11080 VDD.n701 VDD.n691 1084.97
R11081 VDD.n772 VDD.n691 1084.97
R11082 VDD.n782 VDD.n781 1084.97
R11083 VDD.n781 VDD.n688 1084.97
R11084 VDD.n688 VDD.n679 1084.97
R11085 VDD.n782 VDD.n679 1084.97
R11086 VDD.n789 VDD.n676 1084.97
R11087 VDD.n789 VDD.n677 1084.97
R11088 VDD.n793 VDD.n677 1084.97
R11089 VDD.n793 VDD.n676 1084.97
R11090 VDD.n799 VDD.n798 1084.97
R11091 VDD.n798 VDD.n673 1084.97
R11092 VDD.n673 VDD.n663 1084.97
R11093 VDD.n799 VDD.n663 1084.97
R11094 VDD.n809 VDD.n808 1084.97
R11095 VDD.n808 VDD.n660 1084.97
R11096 VDD.n660 VDD.n653 1084.97
R11097 VDD.n809 VDD.n653 1084.97
R11098 VDD.n819 VDD.n818 1084.97
R11099 VDD.n818 VDD.n650 1084.97
R11100 VDD.n650 VDD.n642 1084.97
R11101 VDD.n819 VDD.n642 1084.97
R11102 VDD.n829 VDD.n828 1084.97
R11103 VDD.n828 VDD.n639 1084.97
R11104 VDD.n639 VDD.n629 1084.97
R11105 VDD.n829 VDD.n629 1084.97
R11106 VDD.n839 VDD.n838 1084.97
R11107 VDD.n838 VDD.n626 1084.97
R11108 VDD.n626 VDD.n619 1084.97
R11109 VDD.n839 VDD.n619 1084.97
R11110 VDD.n849 VDD.n848 1084.97
R11111 VDD.n848 VDD.n616 1084.97
R11112 VDD.n616 VDD.n608 1084.97
R11113 VDD.n849 VDD.n608 1084.97
R11114 VDD.n606 VDD.n605 1084.97
R11115 VDD.n856 VDD.n605 1084.97
R11116 VDD.n856 VDD.n603 1084.97
R11117 VDD.n479 VDD.n466 1084.97
R11118 VDD.n479 VDD.n467 1084.97
R11119 VDD.n486 VDD.n467 1084.97
R11120 VDD.n486 VDD.n466 1084.97
R11121 VDD.n489 VDD.n456 1084.97
R11122 VDD.n489 VDD.n457 1084.97
R11123 VDD.n496 VDD.n457 1084.97
R11124 VDD.n496 VDD.n456 1084.97
R11125 VDD.n499 VDD.n445 1084.97
R11126 VDD.n499 VDD.n446 1084.97
R11127 VDD.n506 VDD.n446 1084.97
R11128 VDD.n506 VDD.n445 1084.97
R11129 VDD.n509 VDD.n432 1084.97
R11130 VDD.n509 VDD.n433 1084.97
R11131 VDD.n516 VDD.n433 1084.97
R11132 VDD.n516 VDD.n432 1084.97
R11133 VDD.n519 VDD.n420 1084.97
R11134 VDD.n519 VDD.n421 1084.97
R11135 VDD.n526 VDD.n421 1084.97
R11136 VDD.n526 VDD.n420 1084.97
R11137 VDD.n536 VDD.n404 1084.97
R11138 VDD.n536 VDD.n405 1084.97
R11139 VDD.n543 VDD.n405 1084.97
R11140 VDD.n543 VDD.n404 1084.97
R11141 VDD.n546 VDD.n394 1084.97
R11142 VDD.n546 VDD.n395 1084.97
R11143 VDD.n553 VDD.n395 1084.97
R11144 VDD.n553 VDD.n394 1084.97
R11145 VDD.n556 VDD.n383 1084.97
R11146 VDD.n556 VDD.n384 1084.97
R11147 VDD.n563 VDD.n384 1084.97
R11148 VDD.n563 VDD.n383 1084.97
R11149 VDD.n566 VDD.n370 1084.97
R11150 VDD.n566 VDD.n371 1084.97
R11151 VDD.n573 VDD.n371 1084.97
R11152 VDD.n573 VDD.n370 1084.97
R11153 VDD.n576 VDD.n360 1084.97
R11154 VDD.n576 VDD.n361 1084.97
R11155 VDD.n583 VDD.n361 1084.97
R11156 VDD.n583 VDD.n360 1084.97
R11157 VDD.n586 VDD.n349 1084.97
R11158 VDD.n586 VDD.n350 1084.97
R11159 VDD.n593 VDD.n350 1084.97
R11160 VDD.n593 VDD.n349 1084.97
R11161 VDD.n482 VDD.n481 1084.97
R11162 VDD.n481 VDD.n475 1084.97
R11163 VDD.n475 VDD.n465 1084.97
R11164 VDD.n482 VDD.n465 1084.97
R11165 VDD.n492 VDD.n491 1084.97
R11166 VDD.n491 VDD.n462 1084.97
R11167 VDD.n462 VDD.n455 1084.97
R11168 VDD.n492 VDD.n455 1084.97
R11169 VDD.n502 VDD.n501 1084.97
R11170 VDD.n501 VDD.n452 1084.97
R11171 VDD.n452 VDD.n444 1084.97
R11172 VDD.n502 VDD.n444 1084.97
R11173 VDD.n512 VDD.n511 1084.97
R11174 VDD.n511 VDD.n441 1084.97
R11175 VDD.n441 VDD.n431 1084.97
R11176 VDD.n512 VDD.n431 1084.97
R11177 VDD.n522 VDD.n521 1084.97
R11178 VDD.n521 VDD.n428 1084.97
R11179 VDD.n428 VDD.n419 1084.97
R11180 VDD.n522 VDD.n419 1084.97
R11181 VDD.n529 VDD.n416 1084.97
R11182 VDD.n529 VDD.n417 1084.97
R11183 VDD.n533 VDD.n417 1084.97
R11184 VDD.n533 VDD.n416 1084.97
R11185 VDD.n539 VDD.n538 1084.97
R11186 VDD.n538 VDD.n413 1084.97
R11187 VDD.n413 VDD.n403 1084.97
R11188 VDD.n539 VDD.n403 1084.97
R11189 VDD.n549 VDD.n548 1084.97
R11190 VDD.n548 VDD.n400 1084.97
R11191 VDD.n400 VDD.n393 1084.97
R11192 VDD.n549 VDD.n393 1084.97
R11193 VDD.n559 VDD.n558 1084.97
R11194 VDD.n558 VDD.n390 1084.97
R11195 VDD.n390 VDD.n382 1084.97
R11196 VDD.n559 VDD.n382 1084.97
R11197 VDD.n569 VDD.n568 1084.97
R11198 VDD.n568 VDD.n379 1084.97
R11199 VDD.n379 VDD.n369 1084.97
R11200 VDD.n569 VDD.n369 1084.97
R11201 VDD.n579 VDD.n578 1084.97
R11202 VDD.n578 VDD.n366 1084.97
R11203 VDD.n366 VDD.n359 1084.97
R11204 VDD.n579 VDD.n359 1084.97
R11205 VDD.n589 VDD.n588 1084.97
R11206 VDD.n588 VDD.n356 1084.97
R11207 VDD.n356 VDD.n348 1084.97
R11208 VDD.n589 VDD.n348 1084.97
R11209 VDD.n346 VDD.n345 1084.97
R11210 VDD.n596 VDD.n345 1084.97
R11211 VDD.n596 VDD.n343 1084.97
R11212 VDD.n148 VDD.n143 1084.97
R11213 VDD.n152 VDD.n144 1084.97
R11214 VDD.n152 VDD.n143 1084.97
R11215 VDD.n155 VDD.n138 1084.97
R11216 VDD.n141 VDD.n140 1084.97
R11217 VDD.n155 VDD.n140 1084.97
R11218 VDD.n162 VDD.n130 1084.97
R11219 VDD.n166 VDD.n131 1084.97
R11220 VDD.n166 VDD.n130 1084.97
R11221 VDD.n169 VDD.n127 1084.97
R11222 VDD.n169 VDD.n128 1084.97
R11223 VDD.n173 VDD.n128 1084.97
R11224 VDD.n173 VDD.n127 1084.97
R11225 VDD.n176 VDD.n122 1084.97
R11226 VDD.n125 VDD.n124 1084.97
R11227 VDD.n176 VDD.n124 1084.97
R11228 VDD.n183 VDD.n118 1084.97
R11229 VDD.n187 VDD.n119 1084.97
R11230 VDD.n187 VDD.n118 1084.97
R11231 VDD.n190 VDD.n113 1084.97
R11232 VDD.n116 VDD.n115 1084.97
R11233 VDD.n190 VDD.n115 1084.97
R11234 VDD.n197 VDD.n105 1084.97
R11235 VDD.n201 VDD.n106 1084.97
R11236 VDD.n201 VDD.n105 1084.97
R11237 VDD.n204 VDD.n102 1084.97
R11238 VDD.n204 VDD.n103 1084.97
R11239 VDD.n208 VDD.n103 1084.97
R11240 VDD.n208 VDD.n102 1084.97
R11241 VDD.n211 VDD.n97 1084.97
R11242 VDD.n100 VDD.n99 1084.97
R11243 VDD.n211 VDD.n99 1084.97
R11244 VDD.n218 VDD.n93 1084.97
R11245 VDD.n222 VDD.n94 1084.97
R11246 VDD.n222 VDD.n93 1084.97
R11247 VDD.n225 VDD.n88 1084.97
R11248 VDD.n91 VDD.n90 1084.97
R11249 VDD.n225 VDD.n90 1084.97
R11250 VDD.n232 VDD.n80 1084.97
R11251 VDD.n236 VDD.n81 1084.97
R11252 VDD.n236 VDD.n80 1084.97
R11253 VDD.n239 VDD.n77 1084.97
R11254 VDD.n239 VDD.n78 1084.97
R11255 VDD.n243 VDD.n78 1084.97
R11256 VDD.n243 VDD.n77 1084.97
R11257 VDD.n246 VDD.n72 1084.97
R11258 VDD.n75 VDD.n74 1084.97
R11259 VDD.n246 VDD.n74 1084.97
R11260 VDD.n253 VDD.n68 1084.97
R11261 VDD.n257 VDD.n69 1084.97
R11262 VDD.n257 VDD.n68 1084.97
R11263 VDD.n260 VDD.n63 1084.97
R11264 VDD.n66 VDD.n65 1084.97
R11265 VDD.n260 VDD.n65 1084.97
R11266 VDD.n267 VDD.n55 1084.97
R11267 VDD.n271 VDD.n56 1084.97
R11268 VDD.n271 VDD.n55 1084.97
R11269 VDD.n274 VDD.n52 1084.97
R11270 VDD.n274 VDD.n53 1084.97
R11271 VDD.n278 VDD.n53 1084.97
R11272 VDD.n278 VDD.n52 1084.97
R11273 VDD.n281 VDD.n47 1084.97
R11274 VDD.n50 VDD.n49 1084.97
R11275 VDD.n281 VDD.n49 1084.97
R11276 VDD.n7395 VDD.n7382 1084.97
R11277 VDD.n7395 VDD.n7383 1084.97
R11278 VDD.n7402 VDD.n7383 1084.97
R11279 VDD.n7402 VDD.n7382 1084.97
R11280 VDD.n7405 VDD.n7372 1084.97
R11281 VDD.n7405 VDD.n7373 1084.97
R11282 VDD.n7412 VDD.n7373 1084.97
R11283 VDD.n7412 VDD.n7372 1084.97
R11284 VDD.n7415 VDD.n7361 1084.97
R11285 VDD.n7415 VDD.n7362 1084.97
R11286 VDD.n7422 VDD.n7362 1084.97
R11287 VDD.n7422 VDD.n7361 1084.97
R11288 VDD.n7425 VDD.n7348 1084.97
R11289 VDD.n7425 VDD.n7349 1084.97
R11290 VDD.n7432 VDD.n7349 1084.97
R11291 VDD.n7432 VDD.n7348 1084.97
R11292 VDD.n7435 VDD.n7336 1084.97
R11293 VDD.n7435 VDD.n7337 1084.97
R11294 VDD.n7442 VDD.n7337 1084.97
R11295 VDD.n7442 VDD.n7336 1084.97
R11296 VDD.n7452 VDD.n7320 1084.97
R11297 VDD.n7452 VDD.n7321 1084.97
R11298 VDD.n7459 VDD.n7321 1084.97
R11299 VDD.n7459 VDD.n7320 1084.97
R11300 VDD.n7462 VDD.n7310 1084.97
R11301 VDD.n7462 VDD.n7311 1084.97
R11302 VDD.n7469 VDD.n7311 1084.97
R11303 VDD.n7469 VDD.n7310 1084.97
R11304 VDD.n7472 VDD.n7299 1084.97
R11305 VDD.n7472 VDD.n7300 1084.97
R11306 VDD.n7479 VDD.n7300 1084.97
R11307 VDD.n7479 VDD.n7299 1084.97
R11308 VDD.n7482 VDD.n7286 1084.97
R11309 VDD.n7482 VDD.n7287 1084.97
R11310 VDD.n7489 VDD.n7287 1084.97
R11311 VDD.n7489 VDD.n7286 1084.97
R11312 VDD.n7492 VDD.n7276 1084.97
R11313 VDD.n7492 VDD.n7277 1084.97
R11314 VDD.n7499 VDD.n7277 1084.97
R11315 VDD.n7499 VDD.n7276 1084.97
R11316 VDD.n7502 VDD.n7265 1084.97
R11317 VDD.n7502 VDD.n7266 1084.97
R11318 VDD.n7509 VDD.n7266 1084.97
R11319 VDD.n7509 VDD.n7265 1084.97
R11320 VDD.n7398 VDD.n7397 1084.97
R11321 VDD.n7397 VDD.n7391 1084.97
R11322 VDD.n7391 VDD.n7381 1084.97
R11323 VDD.n7398 VDD.n7381 1084.97
R11324 VDD.n7408 VDD.n7407 1084.97
R11325 VDD.n7407 VDD.n7378 1084.97
R11326 VDD.n7378 VDD.n7371 1084.97
R11327 VDD.n7408 VDD.n7371 1084.97
R11328 VDD.n7418 VDD.n7417 1084.97
R11329 VDD.n7417 VDD.n7368 1084.97
R11330 VDD.n7368 VDD.n7360 1084.97
R11331 VDD.n7418 VDD.n7360 1084.97
R11332 VDD.n7428 VDD.n7427 1084.97
R11333 VDD.n7427 VDD.n7357 1084.97
R11334 VDD.n7357 VDD.n7347 1084.97
R11335 VDD.n7428 VDD.n7347 1084.97
R11336 VDD.n7438 VDD.n7437 1084.97
R11337 VDD.n7437 VDD.n7344 1084.97
R11338 VDD.n7344 VDD.n7335 1084.97
R11339 VDD.n7438 VDD.n7335 1084.97
R11340 VDD.n7445 VDD.n7332 1084.97
R11341 VDD.n7445 VDD.n7333 1084.97
R11342 VDD.n7449 VDD.n7333 1084.97
R11343 VDD.n7449 VDD.n7332 1084.97
R11344 VDD.n7455 VDD.n7454 1084.97
R11345 VDD.n7454 VDD.n7329 1084.97
R11346 VDD.n7329 VDD.n7319 1084.97
R11347 VDD.n7455 VDD.n7319 1084.97
R11348 VDD.n7465 VDD.n7464 1084.97
R11349 VDD.n7464 VDD.n7316 1084.97
R11350 VDD.n7316 VDD.n7309 1084.97
R11351 VDD.n7465 VDD.n7309 1084.97
R11352 VDD.n7475 VDD.n7474 1084.97
R11353 VDD.n7474 VDD.n7306 1084.97
R11354 VDD.n7306 VDD.n7298 1084.97
R11355 VDD.n7475 VDD.n7298 1084.97
R11356 VDD.n7485 VDD.n7484 1084.97
R11357 VDD.n7484 VDD.n7295 1084.97
R11358 VDD.n7295 VDD.n7285 1084.97
R11359 VDD.n7485 VDD.n7285 1084.97
R11360 VDD.n7495 VDD.n7494 1084.97
R11361 VDD.n7494 VDD.n7282 1084.97
R11362 VDD.n7282 VDD.n7275 1084.97
R11363 VDD.n7495 VDD.n7275 1084.97
R11364 VDD.n7505 VDD.n7504 1084.97
R11365 VDD.n7504 VDD.n7272 1084.97
R11366 VDD.n7272 VDD.n7264 1084.97
R11367 VDD.n7505 VDD.n7264 1084.97
R11368 VDD.n7262 VDD.n7261 1084.97
R11369 VDD.n7512 VDD.n7261 1084.97
R11370 VDD.n7512 VDD.n7259 1084.97
R11371 VDD.n7138 VDD.n2031 1084.97
R11372 VDD.n7138 VDD.n2032 1084.97
R11373 VDD.n7145 VDD.n2032 1084.97
R11374 VDD.n7145 VDD.n2031 1084.97
R11375 VDD.n7148 VDD.n2021 1084.97
R11376 VDD.n7148 VDD.n2022 1084.97
R11377 VDD.n7155 VDD.n2022 1084.97
R11378 VDD.n7155 VDD.n2021 1084.97
R11379 VDD.n7158 VDD.n2010 1084.97
R11380 VDD.n7158 VDD.n2011 1084.97
R11381 VDD.n7165 VDD.n2011 1084.97
R11382 VDD.n7165 VDD.n2010 1084.97
R11383 VDD.n7168 VDD.n1997 1084.97
R11384 VDD.n7168 VDD.n1998 1084.97
R11385 VDD.n7175 VDD.n1998 1084.97
R11386 VDD.n7175 VDD.n1997 1084.97
R11387 VDD.n7178 VDD.n1985 1084.97
R11388 VDD.n7178 VDD.n1986 1084.97
R11389 VDD.n7185 VDD.n1986 1084.97
R11390 VDD.n7185 VDD.n1985 1084.97
R11391 VDD.n7200 VDD.n7196 1084.97
R11392 VDD.n7196 VDD.n1965 1084.97
R11393 VDD.n7195 VDD.n1965 1084.97
R11394 VDD.n7200 VDD.n7195 1084.97
R11395 VDD.n7212 VDD.n1943 1084.97
R11396 VDD.n7212 VDD.n1944 1084.97
R11397 VDD.n7219 VDD.n1944 1084.97
R11398 VDD.n7219 VDD.n1943 1084.97
R11399 VDD.n7222 VDD.n1930 1084.97
R11400 VDD.n7222 VDD.n1931 1084.97
R11401 VDD.n7229 VDD.n1931 1084.97
R11402 VDD.n7229 VDD.n1930 1084.97
R11403 VDD.n7232 VDD.n1920 1084.97
R11404 VDD.n7232 VDD.n1921 1084.97
R11405 VDD.n7239 VDD.n1921 1084.97
R11406 VDD.n7239 VDD.n1920 1084.97
R11407 VDD.n7242 VDD.n1909 1084.97
R11408 VDD.n7242 VDD.n1910 1084.97
R11409 VDD.n7249 VDD.n1910 1084.97
R11410 VDD.n7249 VDD.n1909 1084.97
R11411 VDD.n7252 VDD.n1905 1084.97
R11412 VDD.n7252 VDD.n1903 1084.97
R11413 VDD.n1906 VDD.n1905 1084.97
R11414 VDD.n7141 VDD.n7140 1084.97
R11415 VDD.n7140 VDD.n7134 1084.97
R11416 VDD.n7134 VDD.n2030 1084.97
R11417 VDD.n7141 VDD.n2030 1084.97
R11418 VDD.n7151 VDD.n7150 1084.97
R11419 VDD.n7150 VDD.n2027 1084.97
R11420 VDD.n2027 VDD.n2020 1084.97
R11421 VDD.n7151 VDD.n2020 1084.97
R11422 VDD.n7161 VDD.n7160 1084.97
R11423 VDD.n7160 VDD.n2017 1084.97
R11424 VDD.n2017 VDD.n2009 1084.97
R11425 VDD.n7161 VDD.n2009 1084.97
R11426 VDD.n7171 VDD.n7170 1084.97
R11427 VDD.n7170 VDD.n2006 1084.97
R11428 VDD.n2006 VDD.n1996 1084.97
R11429 VDD.n7171 VDD.n1996 1084.97
R11430 VDD.n7181 VDD.n7180 1084.97
R11431 VDD.n7180 VDD.n1993 1084.97
R11432 VDD.n1993 VDD.n1984 1084.97
R11433 VDD.n7181 VDD.n1984 1084.97
R11434 VDD.n7188 VDD.n1981 1084.97
R11435 VDD.n7188 VDD.n1982 1084.97
R11436 VDD.n7192 VDD.n1982 1084.97
R11437 VDD.n7192 VDD.n1981 1084.97
R11438 VDD.n7201 VDD.n1968 1084.97
R11439 VDD.n1980 VDD.n1968 1084.97
R11440 VDD.n1980 VDD.n1967 1084.97
R11441 VDD.n7201 VDD.n1967 1084.97
R11442 VDD.n1960 VDD.n1954 1084.97
R11443 VDD.n1972 VDD.n1960 1084.97
R11444 VDD.n1972 VDD.n1969 1084.97
R11445 VDD.n1969 VDD.n1954 1084.97
R11446 VDD.n7215 VDD.n7214 1084.97
R11447 VDD.n7214 VDD.n1951 1084.97
R11448 VDD.n1951 VDD.n1942 1084.97
R11449 VDD.n7215 VDD.n1942 1084.97
R11450 VDD.n7225 VDD.n7224 1084.97
R11451 VDD.n7224 VDD.n1939 1084.97
R11452 VDD.n1939 VDD.n1929 1084.97
R11453 VDD.n7225 VDD.n1929 1084.97
R11454 VDD.n7235 VDD.n7234 1084.97
R11455 VDD.n7234 VDD.n1926 1084.97
R11456 VDD.n1926 VDD.n1919 1084.97
R11457 VDD.n7235 VDD.n1919 1084.97
R11458 VDD.n7245 VDD.n7244 1084.97
R11459 VDD.n7244 VDD.n1916 1084.97
R11460 VDD.n1916 VDD.n1908 1084.97
R11461 VDD.n7245 VDD.n1908 1084.97
R11462 VDD.n7209 VDD.n1955 1084.97
R11463 VDD.n1974 VDD.n1955 1084.97
R11464 VDD.n7209 VDD.n1956 1084.97
R11465 VDD.n1974 VDD.n1956 1084.97
R11466 VDD.n7116 VDD.n6907 1084.97
R11467 VDD.n7120 VDD.n6908 1084.97
R11468 VDD.n7120 VDD.n6907 1084.97
R11469 VDD.n7125 VDD.n6894 1084.97
R11470 VDD.n7124 VDD.n6894 1084.97
R11471 VDD.n7124 VDD.n6893 1084.97
R11472 VDD.n7125 VDD.n6893 1084.97
R11473 VDD.n6997 VDD.n6992 1084.97
R11474 VDD.n7001 VDD.n6993 1084.97
R11475 VDD.n7001 VDD.n6992 1084.97
R11476 VDD.n7004 VDD.n6987 1084.97
R11477 VDD.n6990 VDD.n6989 1084.97
R11478 VDD.n7004 VDD.n6989 1084.97
R11479 VDD.n7011 VDD.n6979 1084.97
R11480 VDD.n7015 VDD.n6980 1084.97
R11481 VDD.n7015 VDD.n6979 1084.97
R11482 VDD.n7018 VDD.n6976 1084.97
R11483 VDD.n7018 VDD.n6977 1084.97
R11484 VDD.n7022 VDD.n6977 1084.97
R11485 VDD.n7022 VDD.n6976 1084.97
R11486 VDD.n7025 VDD.n6971 1084.97
R11487 VDD.n6974 VDD.n6973 1084.97
R11488 VDD.n7025 VDD.n6973 1084.97
R11489 VDD.n7032 VDD.n6967 1084.97
R11490 VDD.n7036 VDD.n6968 1084.97
R11491 VDD.n7036 VDD.n6967 1084.97
R11492 VDD.n7039 VDD.n6962 1084.97
R11493 VDD.n6965 VDD.n6964 1084.97
R11494 VDD.n7039 VDD.n6964 1084.97
R11495 VDD.n7046 VDD.n6954 1084.97
R11496 VDD.n7050 VDD.n6955 1084.97
R11497 VDD.n7050 VDD.n6954 1084.97
R11498 VDD.n7053 VDD.n6951 1084.97
R11499 VDD.n7053 VDD.n6952 1084.97
R11500 VDD.n7057 VDD.n6952 1084.97
R11501 VDD.n7057 VDD.n6951 1084.97
R11502 VDD.n7060 VDD.n6946 1084.97
R11503 VDD.n6949 VDD.n6948 1084.97
R11504 VDD.n7060 VDD.n6948 1084.97
R11505 VDD.n7067 VDD.n6942 1084.97
R11506 VDD.n7071 VDD.n6943 1084.97
R11507 VDD.n7071 VDD.n6942 1084.97
R11508 VDD.n7074 VDD.n6937 1084.97
R11509 VDD.n6940 VDD.n6939 1084.97
R11510 VDD.n7074 VDD.n6939 1084.97
R11511 VDD.n7081 VDD.n6929 1084.97
R11512 VDD.n7085 VDD.n6930 1084.97
R11513 VDD.n7085 VDD.n6929 1084.97
R11514 VDD.n7088 VDD.n6926 1084.97
R11515 VDD.n7088 VDD.n6927 1084.97
R11516 VDD.n7092 VDD.n6927 1084.97
R11517 VDD.n7092 VDD.n6926 1084.97
R11518 VDD.n7095 VDD.n6921 1084.97
R11519 VDD.n6924 VDD.n6923 1084.97
R11520 VDD.n7095 VDD.n6923 1084.97
R11521 VDD.n7102 VDD.n6917 1084.97
R11522 VDD.n7106 VDD.n6918 1084.97
R11523 VDD.n7106 VDD.n6917 1084.97
R11524 VDD.n7109 VDD.n6912 1084.97
R11525 VDD.n6915 VDD.n6914 1084.97
R11526 VDD.n7109 VDD.n6914 1084.97
R11527 VDD.n6904 VDD.n6895 1084.97
R11528 VDD.n6900 VDD.n6896 1084.97
R11529 VDD.n6904 VDD.n6896 1084.97
R11530 VDD.n6023 VDD.n6019 1084.97
R11531 VDD.n6030 VDD.n6020 1084.97
R11532 VDD.n6030 VDD.n6019 1084.97
R11533 VDD.n6033 VDD.n6010 1084.97
R11534 VDD.n6033 VDD.n6011 1084.97
R11535 VDD.n6040 VDD.n6011 1084.97
R11536 VDD.n6040 VDD.n6010 1084.97
R11537 VDD.n6043 VDD.n5997 1084.97
R11538 VDD.n6043 VDD.n5998 1084.97
R11539 VDD.n6050 VDD.n5998 1084.97
R11540 VDD.n6050 VDD.n5997 1084.97
R11541 VDD.n6053 VDD.n5986 1084.97
R11542 VDD.n6053 VDD.n5987 1084.97
R11543 VDD.n6060 VDD.n5987 1084.97
R11544 VDD.n6060 VDD.n5986 1084.97
R11545 VDD.n6063 VDD.n5976 1084.97
R11546 VDD.n6063 VDD.n5977 1084.97
R11547 VDD.n6070 VDD.n5977 1084.97
R11548 VDD.n6070 VDD.n5976 1084.97
R11549 VDD.n6073 VDD.n5963 1084.97
R11550 VDD.n6073 VDD.n5964 1084.97
R11551 VDD.n6080 VDD.n5964 1084.97
R11552 VDD.n6080 VDD.n5963 1084.97
R11553 VDD.n6083 VDD.n5951 1084.97
R11554 VDD.n6083 VDD.n5952 1084.97
R11555 VDD.n6090 VDD.n5952 1084.97
R11556 VDD.n6090 VDD.n5951 1084.97
R11557 VDD.n6100 VDD.n5935 1084.97
R11558 VDD.n6100 VDD.n5936 1084.97
R11559 VDD.n6107 VDD.n5936 1084.97
R11560 VDD.n6107 VDD.n5935 1084.97
R11561 VDD.n6110 VDD.n5924 1084.97
R11562 VDD.n6110 VDD.n5925 1084.97
R11563 VDD.n6117 VDD.n5925 1084.97
R11564 VDD.n6117 VDD.n5924 1084.97
R11565 VDD.n6120 VDD.n5914 1084.97
R11566 VDD.n6120 VDD.n5915 1084.97
R11567 VDD.n6127 VDD.n5915 1084.97
R11568 VDD.n6127 VDD.n5914 1084.97
R11569 VDD.n6130 VDD.n5904 1084.97
R11570 VDD.n6130 VDD.n5905 1084.97
R11571 VDD.n6137 VDD.n5905 1084.97
R11572 VDD.n6137 VDD.n5904 1084.97
R11573 VDD.n6036 VDD.n6035 1084.97
R11574 VDD.n6035 VDD.n6016 1084.97
R11575 VDD.n6016 VDD.n6009 1084.97
R11576 VDD.n6036 VDD.n6009 1084.97
R11577 VDD.n6046 VDD.n6045 1084.97
R11578 VDD.n6045 VDD.n6006 1084.97
R11579 VDD.n6006 VDD.n5996 1084.97
R11580 VDD.n6046 VDD.n5996 1084.97
R11581 VDD.n6056 VDD.n6055 1084.97
R11582 VDD.n6055 VDD.n5993 1084.97
R11583 VDD.n5993 VDD.n5985 1084.97
R11584 VDD.n6056 VDD.n5985 1084.97
R11585 VDD.n6066 VDD.n6065 1084.97
R11586 VDD.n6065 VDD.n5982 1084.97
R11587 VDD.n5982 VDD.n5975 1084.97
R11588 VDD.n6066 VDD.n5975 1084.97
R11589 VDD.n6076 VDD.n6075 1084.97
R11590 VDD.n6075 VDD.n5972 1084.97
R11591 VDD.n5972 VDD.n5962 1084.97
R11592 VDD.n6076 VDD.n5962 1084.97
R11593 VDD.n6086 VDD.n6085 1084.97
R11594 VDD.n6085 VDD.n5959 1084.97
R11595 VDD.n5959 VDD.n5950 1084.97
R11596 VDD.n6086 VDD.n5950 1084.97
R11597 VDD.n6093 VDD.n5947 1084.97
R11598 VDD.n6093 VDD.n5948 1084.97
R11599 VDD.n6097 VDD.n5948 1084.97
R11600 VDD.n6097 VDD.n5947 1084.97
R11601 VDD.n6103 VDD.n6102 1084.97
R11602 VDD.n6102 VDD.n5944 1084.97
R11603 VDD.n5944 VDD.n5934 1084.97
R11604 VDD.n6103 VDD.n5934 1084.97
R11605 VDD.n6113 VDD.n6112 1084.97
R11606 VDD.n6112 VDD.n5931 1084.97
R11607 VDD.n5931 VDD.n5923 1084.97
R11608 VDD.n6113 VDD.n5923 1084.97
R11609 VDD.n6123 VDD.n6122 1084.97
R11610 VDD.n6122 VDD.n5920 1084.97
R11611 VDD.n5920 VDD.n5913 1084.97
R11612 VDD.n6123 VDD.n5913 1084.97
R11613 VDD.n6133 VDD.n6132 1084.97
R11614 VDD.n6132 VDD.n5910 1084.97
R11615 VDD.n5910 VDD.n5903 1084.97
R11616 VDD.n6133 VDD.n5903 1084.97
R11617 VDD.n6146 VDD.n5896 1084.97
R11618 VDD.n6146 VDD.n5897 1084.97
R11619 VDD.n5902 VDD.n5897 1084.97
R11620 VDD.n5902 VDD.n5896 1084.97
R11621 VDD.n6145 VDD.n6140 1084.97
R11622 VDD.n6145 VDD.n6141 1084.97
R11623 VDD.n6140 VDD.n5894 1084.97
R11624 VDD.n6141 VDD.n5894 1084.97
R11625 VDD.n5887 VDD.n5883 1084.97
R11626 VDD.n6153 VDD.n5884 1084.97
R11627 VDD.n6153 VDD.n5883 1084.97
R11628 VDD.n6156 VDD.n5874 1084.97
R11629 VDD.n6156 VDD.n5875 1084.97
R11630 VDD.n6163 VDD.n5875 1084.97
R11631 VDD.n6163 VDD.n5874 1084.97
R11632 VDD.n6166 VDD.n5861 1084.97
R11633 VDD.n6166 VDD.n5862 1084.97
R11634 VDD.n6173 VDD.n5862 1084.97
R11635 VDD.n6173 VDD.n5861 1084.97
R11636 VDD.n6176 VDD.n5850 1084.97
R11637 VDD.n6176 VDD.n5851 1084.97
R11638 VDD.n6183 VDD.n5851 1084.97
R11639 VDD.n6183 VDD.n5850 1084.97
R11640 VDD.n6186 VDD.n5840 1084.97
R11641 VDD.n6186 VDD.n5841 1084.97
R11642 VDD.n6193 VDD.n5841 1084.97
R11643 VDD.n6193 VDD.n5840 1084.97
R11644 VDD.n6196 VDD.n5827 1084.97
R11645 VDD.n6196 VDD.n5828 1084.97
R11646 VDD.n6203 VDD.n5828 1084.97
R11647 VDD.n6203 VDD.n5827 1084.97
R11648 VDD.n6206 VDD.n5815 1084.97
R11649 VDD.n6206 VDD.n5816 1084.97
R11650 VDD.n6213 VDD.n5816 1084.97
R11651 VDD.n6213 VDD.n5815 1084.97
R11652 VDD.n6223 VDD.n5799 1084.97
R11653 VDD.n6223 VDD.n5800 1084.97
R11654 VDD.n6230 VDD.n5800 1084.97
R11655 VDD.n6230 VDD.n5799 1084.97
R11656 VDD.n6233 VDD.n5788 1084.97
R11657 VDD.n6233 VDD.n5789 1084.97
R11658 VDD.n6240 VDD.n5789 1084.97
R11659 VDD.n6240 VDD.n5788 1084.97
R11660 VDD.n6243 VDD.n5778 1084.97
R11661 VDD.n6243 VDD.n5779 1084.97
R11662 VDD.n6250 VDD.n5779 1084.97
R11663 VDD.n6250 VDD.n5778 1084.97
R11664 VDD.n6253 VDD.n5768 1084.97
R11665 VDD.n6253 VDD.n5769 1084.97
R11666 VDD.n6260 VDD.n5769 1084.97
R11667 VDD.n6260 VDD.n5768 1084.97
R11668 VDD.n6159 VDD.n6158 1084.97
R11669 VDD.n6158 VDD.n5880 1084.97
R11670 VDD.n5880 VDD.n5873 1084.97
R11671 VDD.n6159 VDD.n5873 1084.97
R11672 VDD.n6169 VDD.n6168 1084.97
R11673 VDD.n6168 VDD.n5870 1084.97
R11674 VDD.n5870 VDD.n5860 1084.97
R11675 VDD.n6169 VDD.n5860 1084.97
R11676 VDD.n6179 VDD.n6178 1084.97
R11677 VDD.n6178 VDD.n5857 1084.97
R11678 VDD.n5857 VDD.n5849 1084.97
R11679 VDD.n6179 VDD.n5849 1084.97
R11680 VDD.n6189 VDD.n6188 1084.97
R11681 VDD.n6188 VDD.n5846 1084.97
R11682 VDD.n5846 VDD.n5839 1084.97
R11683 VDD.n6189 VDD.n5839 1084.97
R11684 VDD.n6199 VDD.n6198 1084.97
R11685 VDD.n6198 VDD.n5836 1084.97
R11686 VDD.n5836 VDD.n5826 1084.97
R11687 VDD.n6199 VDD.n5826 1084.97
R11688 VDD.n6209 VDD.n6208 1084.97
R11689 VDD.n6208 VDD.n5823 1084.97
R11690 VDD.n5823 VDD.n5814 1084.97
R11691 VDD.n6209 VDD.n5814 1084.97
R11692 VDD.n6216 VDD.n5811 1084.97
R11693 VDD.n6216 VDD.n5812 1084.97
R11694 VDD.n6220 VDD.n5812 1084.97
R11695 VDD.n6220 VDD.n5811 1084.97
R11696 VDD.n6226 VDD.n6225 1084.97
R11697 VDD.n6225 VDD.n5808 1084.97
R11698 VDD.n5808 VDD.n5798 1084.97
R11699 VDD.n6226 VDD.n5798 1084.97
R11700 VDD.n6236 VDD.n6235 1084.97
R11701 VDD.n6235 VDD.n5795 1084.97
R11702 VDD.n5795 VDD.n5787 1084.97
R11703 VDD.n6236 VDD.n5787 1084.97
R11704 VDD.n6246 VDD.n6245 1084.97
R11705 VDD.n6245 VDD.n5784 1084.97
R11706 VDD.n5784 VDD.n5777 1084.97
R11707 VDD.n6246 VDD.n5777 1084.97
R11708 VDD.n6256 VDD.n6255 1084.97
R11709 VDD.n6255 VDD.n5774 1084.97
R11710 VDD.n5774 VDD.n5767 1084.97
R11711 VDD.n6256 VDD.n5767 1084.97
R11712 VDD.n6269 VDD.n5760 1084.97
R11713 VDD.n6269 VDD.n5761 1084.97
R11714 VDD.n5766 VDD.n5761 1084.97
R11715 VDD.n5766 VDD.n5760 1084.97
R11716 VDD.n6268 VDD.n6263 1084.97
R11717 VDD.n6268 VDD.n6264 1084.97
R11718 VDD.n6263 VDD.n5758 1084.97
R11719 VDD.n6264 VDD.n5758 1084.97
R11720 VDD.n5751 VDD.n5747 1084.97
R11721 VDD.n6276 VDD.n5748 1084.97
R11722 VDD.n6276 VDD.n5747 1084.97
R11723 VDD.n6279 VDD.n5738 1084.97
R11724 VDD.n6279 VDD.n5739 1084.97
R11725 VDD.n6286 VDD.n5739 1084.97
R11726 VDD.n6286 VDD.n5738 1084.97
R11727 VDD.n6289 VDD.n5725 1084.97
R11728 VDD.n6289 VDD.n5726 1084.97
R11729 VDD.n6296 VDD.n5726 1084.97
R11730 VDD.n6296 VDD.n5725 1084.97
R11731 VDD.n6299 VDD.n5714 1084.97
R11732 VDD.n6299 VDD.n5715 1084.97
R11733 VDD.n6306 VDD.n5715 1084.97
R11734 VDD.n6306 VDD.n5714 1084.97
R11735 VDD.n6309 VDD.n5704 1084.97
R11736 VDD.n6309 VDD.n5705 1084.97
R11737 VDD.n6316 VDD.n5705 1084.97
R11738 VDD.n6316 VDD.n5704 1084.97
R11739 VDD.n6319 VDD.n5691 1084.97
R11740 VDD.n6319 VDD.n5692 1084.97
R11741 VDD.n6326 VDD.n5692 1084.97
R11742 VDD.n6326 VDD.n5691 1084.97
R11743 VDD.n6329 VDD.n5679 1084.97
R11744 VDD.n6329 VDD.n5680 1084.97
R11745 VDD.n6336 VDD.n5680 1084.97
R11746 VDD.n6336 VDD.n5679 1084.97
R11747 VDD.n6346 VDD.n5663 1084.97
R11748 VDD.n6346 VDD.n5664 1084.97
R11749 VDD.n6353 VDD.n5664 1084.97
R11750 VDD.n6353 VDD.n5663 1084.97
R11751 VDD.n6356 VDD.n5652 1084.97
R11752 VDD.n6356 VDD.n5653 1084.97
R11753 VDD.n6363 VDD.n5653 1084.97
R11754 VDD.n6363 VDD.n5652 1084.97
R11755 VDD.n6366 VDD.n5642 1084.97
R11756 VDD.n6366 VDD.n5643 1084.97
R11757 VDD.n6373 VDD.n5643 1084.97
R11758 VDD.n6373 VDD.n5642 1084.97
R11759 VDD.n6376 VDD.n5632 1084.97
R11760 VDD.n6376 VDD.n5633 1084.97
R11761 VDD.n6383 VDD.n5633 1084.97
R11762 VDD.n6383 VDD.n5632 1084.97
R11763 VDD.n6282 VDD.n6281 1084.97
R11764 VDD.n6281 VDD.n5744 1084.97
R11765 VDD.n5744 VDD.n5737 1084.97
R11766 VDD.n6282 VDD.n5737 1084.97
R11767 VDD.n6292 VDD.n6291 1084.97
R11768 VDD.n6291 VDD.n5734 1084.97
R11769 VDD.n5734 VDD.n5724 1084.97
R11770 VDD.n6292 VDD.n5724 1084.97
R11771 VDD.n6302 VDD.n6301 1084.97
R11772 VDD.n6301 VDD.n5721 1084.97
R11773 VDD.n5721 VDD.n5713 1084.97
R11774 VDD.n6302 VDD.n5713 1084.97
R11775 VDD.n6312 VDD.n6311 1084.97
R11776 VDD.n6311 VDD.n5710 1084.97
R11777 VDD.n5710 VDD.n5703 1084.97
R11778 VDD.n6312 VDD.n5703 1084.97
R11779 VDD.n6322 VDD.n6321 1084.97
R11780 VDD.n6321 VDD.n5700 1084.97
R11781 VDD.n5700 VDD.n5690 1084.97
R11782 VDD.n6322 VDD.n5690 1084.97
R11783 VDD.n6332 VDD.n6331 1084.97
R11784 VDD.n6331 VDD.n5687 1084.97
R11785 VDD.n5687 VDD.n5678 1084.97
R11786 VDD.n6332 VDD.n5678 1084.97
R11787 VDD.n6339 VDD.n5675 1084.97
R11788 VDD.n6339 VDD.n5676 1084.97
R11789 VDD.n6343 VDD.n5676 1084.97
R11790 VDD.n6343 VDD.n5675 1084.97
R11791 VDD.n6349 VDD.n6348 1084.97
R11792 VDD.n6348 VDD.n5672 1084.97
R11793 VDD.n5672 VDD.n5662 1084.97
R11794 VDD.n6349 VDD.n5662 1084.97
R11795 VDD.n6359 VDD.n6358 1084.97
R11796 VDD.n6358 VDD.n5659 1084.97
R11797 VDD.n5659 VDD.n5651 1084.97
R11798 VDD.n6359 VDD.n5651 1084.97
R11799 VDD.n6369 VDD.n6368 1084.97
R11800 VDD.n6368 VDD.n5648 1084.97
R11801 VDD.n5648 VDD.n5641 1084.97
R11802 VDD.n6369 VDD.n5641 1084.97
R11803 VDD.n6379 VDD.n6378 1084.97
R11804 VDD.n6378 VDD.n5638 1084.97
R11805 VDD.n5638 VDD.n5631 1084.97
R11806 VDD.n6379 VDD.n5631 1084.97
R11807 VDD.n6392 VDD.n5624 1084.97
R11808 VDD.n6392 VDD.n5625 1084.97
R11809 VDD.n5630 VDD.n5625 1084.97
R11810 VDD.n5630 VDD.n5624 1084.97
R11811 VDD.n6391 VDD.n6386 1084.97
R11812 VDD.n6391 VDD.n6387 1084.97
R11813 VDD.n6386 VDD.n5622 1084.97
R11814 VDD.n6387 VDD.n5622 1084.97
R11815 VDD.n5615 VDD.n5611 1084.97
R11816 VDD.n6399 VDD.n5612 1084.97
R11817 VDD.n6399 VDD.n5611 1084.97
R11818 VDD.n6402 VDD.n5602 1084.97
R11819 VDD.n6402 VDD.n5603 1084.97
R11820 VDD.n6409 VDD.n5603 1084.97
R11821 VDD.n6409 VDD.n5602 1084.97
R11822 VDD.n6412 VDD.n5589 1084.97
R11823 VDD.n6412 VDD.n5590 1084.97
R11824 VDD.n6419 VDD.n5590 1084.97
R11825 VDD.n6419 VDD.n5589 1084.97
R11826 VDD.n6422 VDD.n5578 1084.97
R11827 VDD.n6422 VDD.n5579 1084.97
R11828 VDD.n6429 VDD.n5579 1084.97
R11829 VDD.n6429 VDD.n5578 1084.97
R11830 VDD.n6432 VDD.n5568 1084.97
R11831 VDD.n6432 VDD.n5569 1084.97
R11832 VDD.n6439 VDD.n5569 1084.97
R11833 VDD.n6439 VDD.n5568 1084.97
R11834 VDD.n6442 VDD.n5555 1084.97
R11835 VDD.n6442 VDD.n5556 1084.97
R11836 VDD.n6449 VDD.n5556 1084.97
R11837 VDD.n6449 VDD.n5555 1084.97
R11838 VDD.n6452 VDD.n5543 1084.97
R11839 VDD.n6452 VDD.n5544 1084.97
R11840 VDD.n6459 VDD.n5544 1084.97
R11841 VDD.n6459 VDD.n5543 1084.97
R11842 VDD.n6469 VDD.n5527 1084.97
R11843 VDD.n6469 VDD.n5528 1084.97
R11844 VDD.n6476 VDD.n5528 1084.97
R11845 VDD.n6476 VDD.n5527 1084.97
R11846 VDD.n6479 VDD.n5516 1084.97
R11847 VDD.n6479 VDD.n5517 1084.97
R11848 VDD.n6486 VDD.n5517 1084.97
R11849 VDD.n6486 VDD.n5516 1084.97
R11850 VDD.n6489 VDD.n5506 1084.97
R11851 VDD.n6489 VDD.n5507 1084.97
R11852 VDD.n6496 VDD.n5507 1084.97
R11853 VDD.n6496 VDD.n5506 1084.97
R11854 VDD.n6499 VDD.n5496 1084.97
R11855 VDD.n6499 VDD.n5497 1084.97
R11856 VDD.n6506 VDD.n5497 1084.97
R11857 VDD.n6506 VDD.n5496 1084.97
R11858 VDD.n6405 VDD.n6404 1084.97
R11859 VDD.n6404 VDD.n5608 1084.97
R11860 VDD.n5608 VDD.n5601 1084.97
R11861 VDD.n6405 VDD.n5601 1084.97
R11862 VDD.n6415 VDD.n6414 1084.97
R11863 VDD.n6414 VDD.n5598 1084.97
R11864 VDD.n5598 VDD.n5588 1084.97
R11865 VDD.n6415 VDD.n5588 1084.97
R11866 VDD.n6425 VDD.n6424 1084.97
R11867 VDD.n6424 VDD.n5585 1084.97
R11868 VDD.n5585 VDD.n5577 1084.97
R11869 VDD.n6425 VDD.n5577 1084.97
R11870 VDD.n6435 VDD.n6434 1084.97
R11871 VDD.n6434 VDD.n5574 1084.97
R11872 VDD.n5574 VDD.n5567 1084.97
R11873 VDD.n6435 VDD.n5567 1084.97
R11874 VDD.n6445 VDD.n6444 1084.97
R11875 VDD.n6444 VDD.n5564 1084.97
R11876 VDD.n5564 VDD.n5554 1084.97
R11877 VDD.n6445 VDD.n5554 1084.97
R11878 VDD.n6455 VDD.n6454 1084.97
R11879 VDD.n6454 VDD.n5551 1084.97
R11880 VDD.n5551 VDD.n5542 1084.97
R11881 VDD.n6455 VDD.n5542 1084.97
R11882 VDD.n6462 VDD.n5539 1084.97
R11883 VDD.n6462 VDD.n5540 1084.97
R11884 VDD.n6466 VDD.n5540 1084.97
R11885 VDD.n6466 VDD.n5539 1084.97
R11886 VDD.n6472 VDD.n6471 1084.97
R11887 VDD.n6471 VDD.n5536 1084.97
R11888 VDD.n5536 VDD.n5526 1084.97
R11889 VDD.n6472 VDD.n5526 1084.97
R11890 VDD.n6482 VDD.n6481 1084.97
R11891 VDD.n6481 VDD.n5523 1084.97
R11892 VDD.n5523 VDD.n5515 1084.97
R11893 VDD.n6482 VDD.n5515 1084.97
R11894 VDD.n6492 VDD.n6491 1084.97
R11895 VDD.n6491 VDD.n5512 1084.97
R11896 VDD.n5512 VDD.n5505 1084.97
R11897 VDD.n6492 VDD.n5505 1084.97
R11898 VDD.n6502 VDD.n6501 1084.97
R11899 VDD.n6501 VDD.n5502 1084.97
R11900 VDD.n5502 VDD.n5495 1084.97
R11901 VDD.n6502 VDD.n5495 1084.97
R11902 VDD.n6515 VDD.n5488 1084.97
R11903 VDD.n6515 VDD.n5489 1084.97
R11904 VDD.n5494 VDD.n5489 1084.97
R11905 VDD.n5494 VDD.n5488 1084.97
R11906 VDD.n6514 VDD.n6509 1084.97
R11907 VDD.n6514 VDD.n6510 1084.97
R11908 VDD.n6509 VDD.n5486 1084.97
R11909 VDD.n6510 VDD.n5486 1084.97
R11910 VDD.n5479 VDD.n5475 1084.97
R11911 VDD.n6522 VDD.n5476 1084.97
R11912 VDD.n6522 VDD.n5475 1084.97
R11913 VDD.n6525 VDD.n5466 1084.97
R11914 VDD.n6525 VDD.n5467 1084.97
R11915 VDD.n6532 VDD.n5467 1084.97
R11916 VDD.n6532 VDD.n5466 1084.97
R11917 VDD.n6535 VDD.n5453 1084.97
R11918 VDD.n6535 VDD.n5454 1084.97
R11919 VDD.n6542 VDD.n5454 1084.97
R11920 VDD.n6542 VDD.n5453 1084.97
R11921 VDD.n6545 VDD.n5442 1084.97
R11922 VDD.n6545 VDD.n5443 1084.97
R11923 VDD.n6552 VDD.n5443 1084.97
R11924 VDD.n6552 VDD.n5442 1084.97
R11925 VDD.n6555 VDD.n5432 1084.97
R11926 VDD.n6555 VDD.n5433 1084.97
R11927 VDD.n6562 VDD.n5433 1084.97
R11928 VDD.n6562 VDD.n5432 1084.97
R11929 VDD.n6565 VDD.n5419 1084.97
R11930 VDD.n6565 VDD.n5420 1084.97
R11931 VDD.n6572 VDD.n5420 1084.97
R11932 VDD.n6572 VDD.n5419 1084.97
R11933 VDD.n6575 VDD.n5407 1084.97
R11934 VDD.n6575 VDD.n5408 1084.97
R11935 VDD.n6582 VDD.n5408 1084.97
R11936 VDD.n6582 VDD.n5407 1084.97
R11937 VDD.n6592 VDD.n5391 1084.97
R11938 VDD.n6592 VDD.n5392 1084.97
R11939 VDD.n6599 VDD.n5392 1084.97
R11940 VDD.n6599 VDD.n5391 1084.97
R11941 VDD.n6602 VDD.n5380 1084.97
R11942 VDD.n6602 VDD.n5381 1084.97
R11943 VDD.n6609 VDD.n5381 1084.97
R11944 VDD.n6609 VDD.n5380 1084.97
R11945 VDD.n6612 VDD.n5370 1084.97
R11946 VDD.n6612 VDD.n5371 1084.97
R11947 VDD.n6619 VDD.n5371 1084.97
R11948 VDD.n6619 VDD.n5370 1084.97
R11949 VDD.n6622 VDD.n5360 1084.97
R11950 VDD.n6622 VDD.n5361 1084.97
R11951 VDD.n6629 VDD.n5361 1084.97
R11952 VDD.n6629 VDD.n5360 1084.97
R11953 VDD.n6528 VDD.n6527 1084.97
R11954 VDD.n6527 VDD.n5472 1084.97
R11955 VDD.n5472 VDD.n5465 1084.97
R11956 VDD.n6528 VDD.n5465 1084.97
R11957 VDD.n6538 VDD.n6537 1084.97
R11958 VDD.n6537 VDD.n5462 1084.97
R11959 VDD.n5462 VDD.n5452 1084.97
R11960 VDD.n6538 VDD.n5452 1084.97
R11961 VDD.n6548 VDD.n6547 1084.97
R11962 VDD.n6547 VDD.n5449 1084.97
R11963 VDD.n5449 VDD.n5441 1084.97
R11964 VDD.n6548 VDD.n5441 1084.97
R11965 VDD.n6558 VDD.n6557 1084.97
R11966 VDD.n6557 VDD.n5438 1084.97
R11967 VDD.n5438 VDD.n5431 1084.97
R11968 VDD.n6558 VDD.n5431 1084.97
R11969 VDD.n6568 VDD.n6567 1084.97
R11970 VDD.n6567 VDD.n5428 1084.97
R11971 VDD.n5428 VDD.n5418 1084.97
R11972 VDD.n6568 VDD.n5418 1084.97
R11973 VDD.n6578 VDD.n6577 1084.97
R11974 VDD.n6577 VDD.n5415 1084.97
R11975 VDD.n5415 VDD.n5406 1084.97
R11976 VDD.n6578 VDD.n5406 1084.97
R11977 VDD.n6585 VDD.n5403 1084.97
R11978 VDD.n6585 VDD.n5404 1084.97
R11979 VDD.n6589 VDD.n5404 1084.97
R11980 VDD.n6589 VDD.n5403 1084.97
R11981 VDD.n6595 VDD.n6594 1084.97
R11982 VDD.n6594 VDD.n5400 1084.97
R11983 VDD.n5400 VDD.n5390 1084.97
R11984 VDD.n6595 VDD.n5390 1084.97
R11985 VDD.n6605 VDD.n6604 1084.97
R11986 VDD.n6604 VDD.n5387 1084.97
R11987 VDD.n5387 VDD.n5379 1084.97
R11988 VDD.n6605 VDD.n5379 1084.97
R11989 VDD.n6615 VDD.n6614 1084.97
R11990 VDD.n6614 VDD.n5376 1084.97
R11991 VDD.n5376 VDD.n5369 1084.97
R11992 VDD.n6615 VDD.n5369 1084.97
R11993 VDD.n6625 VDD.n6624 1084.97
R11994 VDD.n6624 VDD.n5366 1084.97
R11995 VDD.n5366 VDD.n5359 1084.97
R11996 VDD.n6625 VDD.n5359 1084.97
R11997 VDD.n6638 VDD.n5352 1084.97
R11998 VDD.n6638 VDD.n5353 1084.97
R11999 VDD.n5358 VDD.n5353 1084.97
R12000 VDD.n5358 VDD.n5352 1084.97
R12001 VDD.n6637 VDD.n6632 1084.97
R12002 VDD.n6637 VDD.n6633 1084.97
R12003 VDD.n6632 VDD.n5350 1084.97
R12004 VDD.n6633 VDD.n5350 1084.97
R12005 VDD.n5343 VDD.n5339 1084.97
R12006 VDD.n6645 VDD.n5340 1084.97
R12007 VDD.n6645 VDD.n5339 1084.97
R12008 VDD.n6648 VDD.n5330 1084.97
R12009 VDD.n6648 VDD.n5331 1084.97
R12010 VDD.n6655 VDD.n5331 1084.97
R12011 VDD.n6655 VDD.n5330 1084.97
R12012 VDD.n6658 VDD.n5317 1084.97
R12013 VDD.n6658 VDD.n5318 1084.97
R12014 VDD.n6665 VDD.n5318 1084.97
R12015 VDD.n6665 VDD.n5317 1084.97
R12016 VDD.n6668 VDD.n5306 1084.97
R12017 VDD.n6668 VDD.n5307 1084.97
R12018 VDD.n6675 VDD.n5307 1084.97
R12019 VDD.n6675 VDD.n5306 1084.97
R12020 VDD.n6678 VDD.n5296 1084.97
R12021 VDD.n6678 VDD.n5297 1084.97
R12022 VDD.n6685 VDD.n5297 1084.97
R12023 VDD.n6685 VDD.n5296 1084.97
R12024 VDD.n6688 VDD.n5283 1084.97
R12025 VDD.n6688 VDD.n5284 1084.97
R12026 VDD.n6695 VDD.n5284 1084.97
R12027 VDD.n6695 VDD.n5283 1084.97
R12028 VDD.n6698 VDD.n5271 1084.97
R12029 VDD.n6698 VDD.n5272 1084.97
R12030 VDD.n6705 VDD.n5272 1084.97
R12031 VDD.n6705 VDD.n5271 1084.97
R12032 VDD.n6715 VDD.n5255 1084.97
R12033 VDD.n6715 VDD.n5256 1084.97
R12034 VDD.n6722 VDD.n5256 1084.97
R12035 VDD.n6722 VDD.n5255 1084.97
R12036 VDD.n6725 VDD.n5244 1084.97
R12037 VDD.n6725 VDD.n5245 1084.97
R12038 VDD.n6732 VDD.n5245 1084.97
R12039 VDD.n6732 VDD.n5244 1084.97
R12040 VDD.n6735 VDD.n5234 1084.97
R12041 VDD.n6735 VDD.n5235 1084.97
R12042 VDD.n6742 VDD.n5235 1084.97
R12043 VDD.n6742 VDD.n5234 1084.97
R12044 VDD.n6745 VDD.n5224 1084.97
R12045 VDD.n6745 VDD.n5225 1084.97
R12046 VDD.n6752 VDD.n5225 1084.97
R12047 VDD.n6752 VDD.n5224 1084.97
R12048 VDD.n6651 VDD.n6650 1084.97
R12049 VDD.n6650 VDD.n5336 1084.97
R12050 VDD.n5336 VDD.n5329 1084.97
R12051 VDD.n6651 VDD.n5329 1084.97
R12052 VDD.n6661 VDD.n6660 1084.97
R12053 VDD.n6660 VDD.n5326 1084.97
R12054 VDD.n5326 VDD.n5316 1084.97
R12055 VDD.n6661 VDD.n5316 1084.97
R12056 VDD.n6671 VDD.n6670 1084.97
R12057 VDD.n6670 VDD.n5313 1084.97
R12058 VDD.n5313 VDD.n5305 1084.97
R12059 VDD.n6671 VDD.n5305 1084.97
R12060 VDD.n6681 VDD.n6680 1084.97
R12061 VDD.n6680 VDD.n5302 1084.97
R12062 VDD.n5302 VDD.n5295 1084.97
R12063 VDD.n6681 VDD.n5295 1084.97
R12064 VDD.n6691 VDD.n6690 1084.97
R12065 VDD.n6690 VDD.n5292 1084.97
R12066 VDD.n5292 VDD.n5282 1084.97
R12067 VDD.n6691 VDD.n5282 1084.97
R12068 VDD.n6701 VDD.n6700 1084.97
R12069 VDD.n6700 VDD.n5279 1084.97
R12070 VDD.n5279 VDD.n5270 1084.97
R12071 VDD.n6701 VDD.n5270 1084.97
R12072 VDD.n6708 VDD.n5267 1084.97
R12073 VDD.n6708 VDD.n5268 1084.97
R12074 VDD.n6712 VDD.n5268 1084.97
R12075 VDD.n6712 VDD.n5267 1084.97
R12076 VDD.n6718 VDD.n6717 1084.97
R12077 VDD.n6717 VDD.n5264 1084.97
R12078 VDD.n5264 VDD.n5254 1084.97
R12079 VDD.n6718 VDD.n5254 1084.97
R12080 VDD.n6728 VDD.n6727 1084.97
R12081 VDD.n6727 VDD.n5251 1084.97
R12082 VDD.n5251 VDD.n5243 1084.97
R12083 VDD.n6728 VDD.n5243 1084.97
R12084 VDD.n6738 VDD.n6737 1084.97
R12085 VDD.n6737 VDD.n5240 1084.97
R12086 VDD.n5240 VDD.n5233 1084.97
R12087 VDD.n6738 VDD.n5233 1084.97
R12088 VDD.n6748 VDD.n6747 1084.97
R12089 VDD.n6747 VDD.n5230 1084.97
R12090 VDD.n5230 VDD.n5223 1084.97
R12091 VDD.n6748 VDD.n5223 1084.97
R12092 VDD.n6761 VDD.n5216 1084.97
R12093 VDD.n6761 VDD.n5217 1084.97
R12094 VDD.n5222 VDD.n5217 1084.97
R12095 VDD.n5222 VDD.n5216 1084.97
R12096 VDD.n6760 VDD.n6755 1084.97
R12097 VDD.n6760 VDD.n6756 1084.97
R12098 VDD.n6755 VDD.n5214 1084.97
R12099 VDD.n6756 VDD.n5214 1084.97
R12100 VDD.n5207 VDD.n5203 1084.97
R12101 VDD.n6768 VDD.n5204 1084.97
R12102 VDD.n6768 VDD.n5203 1084.97
R12103 VDD.n6771 VDD.n5194 1084.97
R12104 VDD.n6771 VDD.n5195 1084.97
R12105 VDD.n6778 VDD.n5195 1084.97
R12106 VDD.n6778 VDD.n5194 1084.97
R12107 VDD.n6781 VDD.n5181 1084.97
R12108 VDD.n6781 VDD.n5182 1084.97
R12109 VDD.n6788 VDD.n5182 1084.97
R12110 VDD.n6788 VDD.n5181 1084.97
R12111 VDD.n6791 VDD.n5170 1084.97
R12112 VDD.n6791 VDD.n5171 1084.97
R12113 VDD.n6798 VDD.n5171 1084.97
R12114 VDD.n6798 VDD.n5170 1084.97
R12115 VDD.n6801 VDD.n5160 1084.97
R12116 VDD.n6801 VDD.n5161 1084.97
R12117 VDD.n6808 VDD.n5161 1084.97
R12118 VDD.n6808 VDD.n5160 1084.97
R12119 VDD.n6811 VDD.n5147 1084.97
R12120 VDD.n6811 VDD.n5148 1084.97
R12121 VDD.n6818 VDD.n5148 1084.97
R12122 VDD.n6818 VDD.n5147 1084.97
R12123 VDD.n6821 VDD.n5135 1084.97
R12124 VDD.n6821 VDD.n5136 1084.97
R12125 VDD.n6828 VDD.n5136 1084.97
R12126 VDD.n6828 VDD.n5135 1084.97
R12127 VDD.n6838 VDD.n5119 1084.97
R12128 VDD.n6838 VDD.n5120 1084.97
R12129 VDD.n6845 VDD.n5120 1084.97
R12130 VDD.n6845 VDD.n5119 1084.97
R12131 VDD.n6848 VDD.n5108 1084.97
R12132 VDD.n6848 VDD.n5109 1084.97
R12133 VDD.n6855 VDD.n5109 1084.97
R12134 VDD.n6855 VDD.n5108 1084.97
R12135 VDD.n6858 VDD.n5098 1084.97
R12136 VDD.n6858 VDD.n5099 1084.97
R12137 VDD.n6865 VDD.n5099 1084.97
R12138 VDD.n6865 VDD.n5098 1084.97
R12139 VDD.n6868 VDD.n5088 1084.97
R12140 VDD.n6868 VDD.n5089 1084.97
R12141 VDD.n6875 VDD.n5089 1084.97
R12142 VDD.n6875 VDD.n5088 1084.97
R12143 VDD.n6774 VDD.n6773 1084.97
R12144 VDD.n6773 VDD.n5200 1084.97
R12145 VDD.n5200 VDD.n5193 1084.97
R12146 VDD.n6774 VDD.n5193 1084.97
R12147 VDD.n6784 VDD.n6783 1084.97
R12148 VDD.n6783 VDD.n5190 1084.97
R12149 VDD.n5190 VDD.n5180 1084.97
R12150 VDD.n6784 VDD.n5180 1084.97
R12151 VDD.n6794 VDD.n6793 1084.97
R12152 VDD.n6793 VDD.n5177 1084.97
R12153 VDD.n5177 VDD.n5169 1084.97
R12154 VDD.n6794 VDD.n5169 1084.97
R12155 VDD.n6804 VDD.n6803 1084.97
R12156 VDD.n6803 VDD.n5166 1084.97
R12157 VDD.n5166 VDD.n5159 1084.97
R12158 VDD.n6804 VDD.n5159 1084.97
R12159 VDD.n6814 VDD.n6813 1084.97
R12160 VDD.n6813 VDD.n5156 1084.97
R12161 VDD.n5156 VDD.n5146 1084.97
R12162 VDD.n6814 VDD.n5146 1084.97
R12163 VDD.n6824 VDD.n6823 1084.97
R12164 VDD.n6823 VDD.n5143 1084.97
R12165 VDD.n5143 VDD.n5134 1084.97
R12166 VDD.n6824 VDD.n5134 1084.97
R12167 VDD.n6831 VDD.n5131 1084.97
R12168 VDD.n6831 VDD.n5132 1084.97
R12169 VDD.n6835 VDD.n5132 1084.97
R12170 VDD.n6835 VDD.n5131 1084.97
R12171 VDD.n6841 VDD.n6840 1084.97
R12172 VDD.n6840 VDD.n5128 1084.97
R12173 VDD.n5128 VDD.n5118 1084.97
R12174 VDD.n6841 VDD.n5118 1084.97
R12175 VDD.n6851 VDD.n6850 1084.97
R12176 VDD.n6850 VDD.n5115 1084.97
R12177 VDD.n5115 VDD.n5107 1084.97
R12178 VDD.n6851 VDD.n5107 1084.97
R12179 VDD.n6861 VDD.n6860 1084.97
R12180 VDD.n6860 VDD.n5104 1084.97
R12181 VDD.n5104 VDD.n5097 1084.97
R12182 VDD.n6861 VDD.n5097 1084.97
R12183 VDD.n6871 VDD.n6870 1084.97
R12184 VDD.n6870 VDD.n5094 1084.97
R12185 VDD.n5094 VDD.n5087 1084.97
R12186 VDD.n6871 VDD.n5087 1084.97
R12187 VDD.n6884 VDD.n5080 1084.97
R12188 VDD.n6884 VDD.n5081 1084.97
R12189 VDD.n5086 VDD.n5081 1084.97
R12190 VDD.n5086 VDD.n5080 1084.97
R12191 VDD.n6883 VDD.n6878 1084.97
R12192 VDD.n6883 VDD.n6879 1084.97
R12193 VDD.n6878 VDD.n5078 1084.97
R12194 VDD.n6879 VDD.n5078 1084.97
R12195 VDD.n5069 VDD.n4819 1084.97
R12196 VDD.n5066 VDD.n4817 1084.97
R12197 VDD.n5066 VDD.n4819 1084.97
R12198 VDD.n5064 VDD.n4821 1084.97
R12199 VDD.n5064 VDD.n4822 1084.97
R12200 VDD.n5057 VDD.n4822 1084.97
R12201 VDD.n5057 VDD.n4821 1084.97
R12202 VDD.n5054 VDD.n4832 1084.97
R12203 VDD.n5054 VDD.n4833 1084.97
R12204 VDD.n5047 VDD.n4833 1084.97
R12205 VDD.n5047 VDD.n4832 1084.97
R12206 VDD.n5044 VDD.n4842 1084.97
R12207 VDD.n5044 VDD.n4843 1084.97
R12208 VDD.n5037 VDD.n4843 1084.97
R12209 VDD.n5037 VDD.n4842 1084.97
R12210 VDD.n5034 VDD.n4855 1084.97
R12211 VDD.n5034 VDD.n4856 1084.97
R12212 VDD.n5027 VDD.n4856 1084.97
R12213 VDD.n5027 VDD.n4855 1084.97
R12214 VDD.n5024 VDD.n4866 1084.97
R12215 VDD.n5024 VDD.n4867 1084.97
R12216 VDD.n5017 VDD.n4867 1084.97
R12217 VDD.n5017 VDD.n4866 1084.97
R12218 VDD.n5014 VDD.n4876 1084.97
R12219 VDD.n5014 VDD.n4877 1084.97
R12220 VDD.n5007 VDD.n4877 1084.97
R12221 VDD.n5007 VDD.n4876 1084.97
R12222 VDD.n4997 VDD.n4892 1084.97
R12223 VDD.n4997 VDD.n4893 1084.97
R12224 VDD.n4990 VDD.n4893 1084.97
R12225 VDD.n4990 VDD.n4892 1084.97
R12226 VDD.n4987 VDD.n4904 1084.97
R12227 VDD.n4987 VDD.n4905 1084.97
R12228 VDD.n4980 VDD.n4905 1084.97
R12229 VDD.n4980 VDD.n4904 1084.97
R12230 VDD.n4977 VDD.n4917 1084.97
R12231 VDD.n4977 VDD.n4918 1084.97
R12232 VDD.n4970 VDD.n4918 1084.97
R12233 VDD.n4970 VDD.n4917 1084.97
R12234 VDD.n4967 VDD.n4928 1084.97
R12235 VDD.n4967 VDD.n4929 1084.97
R12236 VDD.n4960 VDD.n4929 1084.97
R12237 VDD.n4960 VDD.n4928 1084.97
R12238 VDD.n5060 VDD.n4820 1084.97
R12239 VDD.n4828 VDD.n4820 1084.97
R12240 VDD.n5059 VDD.n4828 1084.97
R12241 VDD.n5060 VDD.n5059 1084.97
R12242 VDD.n5050 VDD.n4831 1084.97
R12243 VDD.n4838 VDD.n4831 1084.97
R12244 VDD.n5049 VDD.n4838 1084.97
R12245 VDD.n5050 VDD.n5049 1084.97
R12246 VDD.n5040 VDD.n4841 1084.97
R12247 VDD.n4851 VDD.n4841 1084.97
R12248 VDD.n5039 VDD.n4851 1084.97
R12249 VDD.n5040 VDD.n5039 1084.97
R12250 VDD.n5030 VDD.n4854 1084.97
R12251 VDD.n4862 VDD.n4854 1084.97
R12252 VDD.n5029 VDD.n4862 1084.97
R12253 VDD.n5030 VDD.n5029 1084.97
R12254 VDD.n5020 VDD.n4865 1084.97
R12255 VDD.n4872 VDD.n4865 1084.97
R12256 VDD.n5019 VDD.n4872 1084.97
R12257 VDD.n5020 VDD.n5019 1084.97
R12258 VDD.n5010 VDD.n4875 1084.97
R12259 VDD.n4885 VDD.n4875 1084.97
R12260 VDD.n5009 VDD.n4885 1084.97
R12261 VDD.n5010 VDD.n5009 1084.97
R12262 VDD.n5004 VDD.n4888 1084.97
R12263 VDD.n5004 VDD.n4889 1084.97
R12264 VDD.n5000 VDD.n4889 1084.97
R12265 VDD.n5000 VDD.n4888 1084.97
R12266 VDD.n4993 VDD.n4891 1084.97
R12267 VDD.n4900 VDD.n4891 1084.97
R12268 VDD.n4992 VDD.n4900 1084.97
R12269 VDD.n4993 VDD.n4992 1084.97
R12270 VDD.n4983 VDD.n4903 1084.97
R12271 VDD.n4913 VDD.n4903 1084.97
R12272 VDD.n4982 VDD.n4913 1084.97
R12273 VDD.n4983 VDD.n4982 1084.97
R12274 VDD.n4973 VDD.n4916 1084.97
R12275 VDD.n4924 VDD.n4916 1084.97
R12276 VDD.n4972 VDD.n4924 1084.97
R12277 VDD.n4973 VDD.n4972 1084.97
R12278 VDD.n4963 VDD.n4927 1084.97
R12279 VDD.n4934 VDD.n4927 1084.97
R12280 VDD.n4962 VDD.n4934 1084.97
R12281 VDD.n4963 VDD.n4962 1084.97
R12282 VDD.n4950 VDD.n4949 1084.97
R12283 VDD.n4950 VDD.n4937 1084.97
R12284 VDD.n4943 VDD.n4937 1084.97
R12285 VDD.n4949 VDD.n4943 1084.97
R12286 VDD.n4947 VDD.n4938 1084.97
R12287 VDD.n4957 VDD.n4938 1084.97
R12288 VDD.n4947 VDD.n4939 1084.97
R12289 VDD.n4957 VDD.n4939 1084.97
R12290 VDD.n4697 VDD.n2167 1084.97
R12291 VDD.n4697 VDD.n2168 1084.97
R12292 VDD.n4704 VDD.n2168 1084.97
R12293 VDD.n4704 VDD.n2167 1084.97
R12294 VDD.n4707 VDD.n2157 1084.97
R12295 VDD.n4707 VDD.n2158 1084.97
R12296 VDD.n4714 VDD.n2158 1084.97
R12297 VDD.n4714 VDD.n2157 1084.97
R12298 VDD.n4717 VDD.n2146 1084.97
R12299 VDD.n4717 VDD.n2147 1084.97
R12300 VDD.n4724 VDD.n2147 1084.97
R12301 VDD.n4724 VDD.n2146 1084.97
R12302 VDD.n4727 VDD.n2133 1084.97
R12303 VDD.n4727 VDD.n2134 1084.97
R12304 VDD.n4734 VDD.n2134 1084.97
R12305 VDD.n4734 VDD.n2133 1084.97
R12306 VDD.n4737 VDD.n2121 1084.97
R12307 VDD.n4737 VDD.n2122 1084.97
R12308 VDD.n4744 VDD.n2122 1084.97
R12309 VDD.n4744 VDD.n2121 1084.97
R12310 VDD.n4759 VDD.n4755 1084.97
R12311 VDD.n4755 VDD.n2101 1084.97
R12312 VDD.n4754 VDD.n2101 1084.97
R12313 VDD.n4759 VDD.n4754 1084.97
R12314 VDD.n4771 VDD.n2079 1084.97
R12315 VDD.n4771 VDD.n2080 1084.97
R12316 VDD.n4778 VDD.n2080 1084.97
R12317 VDD.n4778 VDD.n2079 1084.97
R12318 VDD.n4781 VDD.n2066 1084.97
R12319 VDD.n4781 VDD.n2067 1084.97
R12320 VDD.n4788 VDD.n2067 1084.97
R12321 VDD.n4788 VDD.n2066 1084.97
R12322 VDD.n4791 VDD.n2056 1084.97
R12323 VDD.n4791 VDD.n2057 1084.97
R12324 VDD.n4798 VDD.n2057 1084.97
R12325 VDD.n4798 VDD.n2056 1084.97
R12326 VDD.n4801 VDD.n2045 1084.97
R12327 VDD.n4801 VDD.n2046 1084.97
R12328 VDD.n4808 VDD.n2046 1084.97
R12329 VDD.n4808 VDD.n2045 1084.97
R12330 VDD.n4811 VDD.n2041 1084.97
R12331 VDD.n4811 VDD.n2039 1084.97
R12332 VDD.n2042 VDD.n2041 1084.97
R12333 VDD.n4700 VDD.n4699 1084.97
R12334 VDD.n4699 VDD.n4693 1084.97
R12335 VDD.n4693 VDD.n2166 1084.97
R12336 VDD.n4700 VDD.n2166 1084.97
R12337 VDD.n4710 VDD.n4709 1084.97
R12338 VDD.n4709 VDD.n2163 1084.97
R12339 VDD.n2163 VDD.n2156 1084.97
R12340 VDD.n4710 VDD.n2156 1084.97
R12341 VDD.n4720 VDD.n4719 1084.97
R12342 VDD.n4719 VDD.n2153 1084.97
R12343 VDD.n2153 VDD.n2145 1084.97
R12344 VDD.n4720 VDD.n2145 1084.97
R12345 VDD.n4730 VDD.n4729 1084.97
R12346 VDD.n4729 VDD.n2142 1084.97
R12347 VDD.n2142 VDD.n2132 1084.97
R12348 VDD.n4730 VDD.n2132 1084.97
R12349 VDD.n4740 VDD.n4739 1084.97
R12350 VDD.n4739 VDD.n2129 1084.97
R12351 VDD.n2129 VDD.n2120 1084.97
R12352 VDD.n4740 VDD.n2120 1084.97
R12353 VDD.n4747 VDD.n2117 1084.97
R12354 VDD.n4747 VDD.n2118 1084.97
R12355 VDD.n4751 VDD.n2118 1084.97
R12356 VDD.n4751 VDD.n2117 1084.97
R12357 VDD.n4760 VDD.n2104 1084.97
R12358 VDD.n2116 VDD.n2104 1084.97
R12359 VDD.n2116 VDD.n2103 1084.97
R12360 VDD.n4760 VDD.n2103 1084.97
R12361 VDD.n2096 VDD.n2090 1084.97
R12362 VDD.n2108 VDD.n2096 1084.97
R12363 VDD.n2108 VDD.n2105 1084.97
R12364 VDD.n2105 VDD.n2090 1084.97
R12365 VDD.n4774 VDD.n4773 1084.97
R12366 VDD.n4773 VDD.n2087 1084.97
R12367 VDD.n2087 VDD.n2078 1084.97
R12368 VDD.n4774 VDD.n2078 1084.97
R12369 VDD.n4784 VDD.n4783 1084.97
R12370 VDD.n4783 VDD.n2075 1084.97
R12371 VDD.n2075 VDD.n2065 1084.97
R12372 VDD.n4784 VDD.n2065 1084.97
R12373 VDD.n4794 VDD.n4793 1084.97
R12374 VDD.n4793 VDD.n2062 1084.97
R12375 VDD.n2062 VDD.n2055 1084.97
R12376 VDD.n4794 VDD.n2055 1084.97
R12377 VDD.n4804 VDD.n4803 1084.97
R12378 VDD.n4803 VDD.n2052 1084.97
R12379 VDD.n2052 VDD.n2044 1084.97
R12380 VDD.n4804 VDD.n2044 1084.97
R12381 VDD.n4768 VDD.n2091 1084.97
R12382 VDD.n2110 VDD.n2091 1084.97
R12383 VDD.n4768 VDD.n2092 1084.97
R12384 VDD.n2110 VDD.n2092 1084.97
R12385 VDD.n4572 VDD.n2303 1084.97
R12386 VDD.n4572 VDD.n2304 1084.97
R12387 VDD.n4579 VDD.n2304 1084.97
R12388 VDD.n4579 VDD.n2303 1084.97
R12389 VDD.n4582 VDD.n2293 1084.97
R12390 VDD.n4582 VDD.n2294 1084.97
R12391 VDD.n4589 VDD.n2294 1084.97
R12392 VDD.n4589 VDD.n2293 1084.97
R12393 VDD.n4592 VDD.n2282 1084.97
R12394 VDD.n4592 VDD.n2283 1084.97
R12395 VDD.n4599 VDD.n2283 1084.97
R12396 VDD.n4599 VDD.n2282 1084.97
R12397 VDD.n4602 VDD.n2269 1084.97
R12398 VDD.n4602 VDD.n2270 1084.97
R12399 VDD.n4609 VDD.n2270 1084.97
R12400 VDD.n4609 VDD.n2269 1084.97
R12401 VDD.n4612 VDD.n2257 1084.97
R12402 VDD.n4612 VDD.n2258 1084.97
R12403 VDD.n4619 VDD.n2258 1084.97
R12404 VDD.n4619 VDD.n2257 1084.97
R12405 VDD.n4634 VDD.n4630 1084.97
R12406 VDD.n4630 VDD.n2237 1084.97
R12407 VDD.n4629 VDD.n2237 1084.97
R12408 VDD.n4634 VDD.n4629 1084.97
R12409 VDD.n4646 VDD.n2215 1084.97
R12410 VDD.n4646 VDD.n2216 1084.97
R12411 VDD.n4653 VDD.n2216 1084.97
R12412 VDD.n4653 VDD.n2215 1084.97
R12413 VDD.n4656 VDD.n2202 1084.97
R12414 VDD.n4656 VDD.n2203 1084.97
R12415 VDD.n4663 VDD.n2203 1084.97
R12416 VDD.n4663 VDD.n2202 1084.97
R12417 VDD.n4666 VDD.n2192 1084.97
R12418 VDD.n4666 VDD.n2193 1084.97
R12419 VDD.n4673 VDD.n2193 1084.97
R12420 VDD.n4673 VDD.n2192 1084.97
R12421 VDD.n4676 VDD.n2181 1084.97
R12422 VDD.n4676 VDD.n2182 1084.97
R12423 VDD.n4683 VDD.n2182 1084.97
R12424 VDD.n4683 VDD.n2181 1084.97
R12425 VDD.n4686 VDD.n2177 1084.97
R12426 VDD.n4686 VDD.n2175 1084.97
R12427 VDD.n2178 VDD.n2177 1084.97
R12428 VDD.n4575 VDD.n4574 1084.97
R12429 VDD.n4574 VDD.n4568 1084.97
R12430 VDD.n4568 VDD.n2302 1084.97
R12431 VDD.n4575 VDD.n2302 1084.97
R12432 VDD.n4585 VDD.n4584 1084.97
R12433 VDD.n4584 VDD.n2299 1084.97
R12434 VDD.n2299 VDD.n2292 1084.97
R12435 VDD.n4585 VDD.n2292 1084.97
R12436 VDD.n4595 VDD.n4594 1084.97
R12437 VDD.n4594 VDD.n2289 1084.97
R12438 VDD.n2289 VDD.n2281 1084.97
R12439 VDD.n4595 VDD.n2281 1084.97
R12440 VDD.n4605 VDD.n4604 1084.97
R12441 VDD.n4604 VDD.n2278 1084.97
R12442 VDD.n2278 VDD.n2268 1084.97
R12443 VDD.n4605 VDD.n2268 1084.97
R12444 VDD.n4615 VDD.n4614 1084.97
R12445 VDD.n4614 VDD.n2265 1084.97
R12446 VDD.n2265 VDD.n2256 1084.97
R12447 VDD.n4615 VDD.n2256 1084.97
R12448 VDD.n4622 VDD.n2253 1084.97
R12449 VDD.n4622 VDD.n2254 1084.97
R12450 VDD.n4626 VDD.n2254 1084.97
R12451 VDD.n4626 VDD.n2253 1084.97
R12452 VDD.n4635 VDD.n2240 1084.97
R12453 VDD.n2252 VDD.n2240 1084.97
R12454 VDD.n2252 VDD.n2239 1084.97
R12455 VDD.n4635 VDD.n2239 1084.97
R12456 VDD.n2232 VDD.n2226 1084.97
R12457 VDD.n2244 VDD.n2232 1084.97
R12458 VDD.n2244 VDD.n2241 1084.97
R12459 VDD.n2241 VDD.n2226 1084.97
R12460 VDD.n4649 VDD.n4648 1084.97
R12461 VDD.n4648 VDD.n2223 1084.97
R12462 VDD.n2223 VDD.n2214 1084.97
R12463 VDD.n4649 VDD.n2214 1084.97
R12464 VDD.n4659 VDD.n4658 1084.97
R12465 VDD.n4658 VDD.n2211 1084.97
R12466 VDD.n2211 VDD.n2201 1084.97
R12467 VDD.n4659 VDD.n2201 1084.97
R12468 VDD.n4669 VDD.n4668 1084.97
R12469 VDD.n4668 VDD.n2198 1084.97
R12470 VDD.n2198 VDD.n2191 1084.97
R12471 VDD.n4669 VDD.n2191 1084.97
R12472 VDD.n4679 VDD.n4678 1084.97
R12473 VDD.n4678 VDD.n2188 1084.97
R12474 VDD.n2188 VDD.n2180 1084.97
R12475 VDD.n4679 VDD.n2180 1084.97
R12476 VDD.n4643 VDD.n2227 1084.97
R12477 VDD.n2246 VDD.n2227 1084.97
R12478 VDD.n4643 VDD.n2228 1084.97
R12479 VDD.n2246 VDD.n2228 1084.97
R12480 VDD.n4447 VDD.n2439 1084.97
R12481 VDD.n4447 VDD.n2440 1084.97
R12482 VDD.n4454 VDD.n2440 1084.97
R12483 VDD.n4454 VDD.n2439 1084.97
R12484 VDD.n4457 VDD.n2429 1084.97
R12485 VDD.n4457 VDD.n2430 1084.97
R12486 VDD.n4464 VDD.n2430 1084.97
R12487 VDD.n4464 VDD.n2429 1084.97
R12488 VDD.n4467 VDD.n2418 1084.97
R12489 VDD.n4467 VDD.n2419 1084.97
R12490 VDD.n4474 VDD.n2419 1084.97
R12491 VDD.n4474 VDD.n2418 1084.97
R12492 VDD.n4477 VDD.n2405 1084.97
R12493 VDD.n4477 VDD.n2406 1084.97
R12494 VDD.n4484 VDD.n2406 1084.97
R12495 VDD.n4484 VDD.n2405 1084.97
R12496 VDD.n4487 VDD.n2393 1084.97
R12497 VDD.n4487 VDD.n2394 1084.97
R12498 VDD.n4494 VDD.n2394 1084.97
R12499 VDD.n4494 VDD.n2393 1084.97
R12500 VDD.n4509 VDD.n4505 1084.97
R12501 VDD.n4505 VDD.n2373 1084.97
R12502 VDD.n4504 VDD.n2373 1084.97
R12503 VDD.n4509 VDD.n4504 1084.97
R12504 VDD.n4521 VDD.n2351 1084.97
R12505 VDD.n4521 VDD.n2352 1084.97
R12506 VDD.n4528 VDD.n2352 1084.97
R12507 VDD.n4528 VDD.n2351 1084.97
R12508 VDD.n4531 VDD.n2338 1084.97
R12509 VDD.n4531 VDD.n2339 1084.97
R12510 VDD.n4538 VDD.n2339 1084.97
R12511 VDD.n4538 VDD.n2338 1084.97
R12512 VDD.n4541 VDD.n2328 1084.97
R12513 VDD.n4541 VDD.n2329 1084.97
R12514 VDD.n4548 VDD.n2329 1084.97
R12515 VDD.n4548 VDD.n2328 1084.97
R12516 VDD.n4551 VDD.n2317 1084.97
R12517 VDD.n4551 VDD.n2318 1084.97
R12518 VDD.n4558 VDD.n2318 1084.97
R12519 VDD.n4558 VDD.n2317 1084.97
R12520 VDD.n4561 VDD.n2313 1084.97
R12521 VDD.n4561 VDD.n2311 1084.97
R12522 VDD.n2314 VDD.n2313 1084.97
R12523 VDD.n4450 VDD.n4449 1084.97
R12524 VDD.n4449 VDD.n4443 1084.97
R12525 VDD.n4443 VDD.n2438 1084.97
R12526 VDD.n4450 VDD.n2438 1084.97
R12527 VDD.n4460 VDD.n4459 1084.97
R12528 VDD.n4459 VDD.n2435 1084.97
R12529 VDD.n2435 VDD.n2428 1084.97
R12530 VDD.n4460 VDD.n2428 1084.97
R12531 VDD.n4470 VDD.n4469 1084.97
R12532 VDD.n4469 VDD.n2425 1084.97
R12533 VDD.n2425 VDD.n2417 1084.97
R12534 VDD.n4470 VDD.n2417 1084.97
R12535 VDD.n4480 VDD.n4479 1084.97
R12536 VDD.n4479 VDD.n2414 1084.97
R12537 VDD.n2414 VDD.n2404 1084.97
R12538 VDD.n4480 VDD.n2404 1084.97
R12539 VDD.n4490 VDD.n4489 1084.97
R12540 VDD.n4489 VDD.n2401 1084.97
R12541 VDD.n2401 VDD.n2392 1084.97
R12542 VDD.n4490 VDD.n2392 1084.97
R12543 VDD.n4497 VDD.n2389 1084.97
R12544 VDD.n4497 VDD.n2390 1084.97
R12545 VDD.n4501 VDD.n2390 1084.97
R12546 VDD.n4501 VDD.n2389 1084.97
R12547 VDD.n4510 VDD.n2376 1084.97
R12548 VDD.n2388 VDD.n2376 1084.97
R12549 VDD.n2388 VDD.n2375 1084.97
R12550 VDD.n4510 VDD.n2375 1084.97
R12551 VDD.n2368 VDD.n2362 1084.97
R12552 VDD.n2380 VDD.n2368 1084.97
R12553 VDD.n2380 VDD.n2377 1084.97
R12554 VDD.n2377 VDD.n2362 1084.97
R12555 VDD.n4524 VDD.n4523 1084.97
R12556 VDD.n4523 VDD.n2359 1084.97
R12557 VDD.n2359 VDD.n2350 1084.97
R12558 VDD.n4524 VDD.n2350 1084.97
R12559 VDD.n4534 VDD.n4533 1084.97
R12560 VDD.n4533 VDD.n2347 1084.97
R12561 VDD.n2347 VDD.n2337 1084.97
R12562 VDD.n4534 VDD.n2337 1084.97
R12563 VDD.n4544 VDD.n4543 1084.97
R12564 VDD.n4543 VDD.n2334 1084.97
R12565 VDD.n2334 VDD.n2327 1084.97
R12566 VDD.n4544 VDD.n2327 1084.97
R12567 VDD.n4554 VDD.n4553 1084.97
R12568 VDD.n4553 VDD.n2324 1084.97
R12569 VDD.n2324 VDD.n2316 1084.97
R12570 VDD.n4554 VDD.n2316 1084.97
R12571 VDD.n4518 VDD.n2363 1084.97
R12572 VDD.n2382 VDD.n2363 1084.97
R12573 VDD.n4518 VDD.n2364 1084.97
R12574 VDD.n2382 VDD.n2364 1084.97
R12575 VDD.n4322 VDD.n2575 1084.97
R12576 VDD.n4322 VDD.n2576 1084.97
R12577 VDD.n4329 VDD.n2576 1084.97
R12578 VDD.n4329 VDD.n2575 1084.97
R12579 VDD.n4332 VDD.n2565 1084.97
R12580 VDD.n4332 VDD.n2566 1084.97
R12581 VDD.n4339 VDD.n2566 1084.97
R12582 VDD.n4339 VDD.n2565 1084.97
R12583 VDD.n4342 VDD.n2554 1084.97
R12584 VDD.n4342 VDD.n2555 1084.97
R12585 VDD.n4349 VDD.n2555 1084.97
R12586 VDD.n4349 VDD.n2554 1084.97
R12587 VDD.n4352 VDD.n2541 1084.97
R12588 VDD.n4352 VDD.n2542 1084.97
R12589 VDD.n4359 VDD.n2542 1084.97
R12590 VDD.n4359 VDD.n2541 1084.97
R12591 VDD.n4362 VDD.n2529 1084.97
R12592 VDD.n4362 VDD.n2530 1084.97
R12593 VDD.n4369 VDD.n2530 1084.97
R12594 VDD.n4369 VDD.n2529 1084.97
R12595 VDD.n4384 VDD.n4380 1084.97
R12596 VDD.n4380 VDD.n2509 1084.97
R12597 VDD.n4379 VDD.n2509 1084.97
R12598 VDD.n4384 VDD.n4379 1084.97
R12599 VDD.n4396 VDD.n2487 1084.97
R12600 VDD.n4396 VDD.n2488 1084.97
R12601 VDD.n4403 VDD.n2488 1084.97
R12602 VDD.n4403 VDD.n2487 1084.97
R12603 VDD.n4406 VDD.n2474 1084.97
R12604 VDD.n4406 VDD.n2475 1084.97
R12605 VDD.n4413 VDD.n2475 1084.97
R12606 VDD.n4413 VDD.n2474 1084.97
R12607 VDD.n4416 VDD.n2464 1084.97
R12608 VDD.n4416 VDD.n2465 1084.97
R12609 VDD.n4423 VDD.n2465 1084.97
R12610 VDD.n4423 VDD.n2464 1084.97
R12611 VDD.n4426 VDD.n2453 1084.97
R12612 VDD.n4426 VDD.n2454 1084.97
R12613 VDD.n4433 VDD.n2454 1084.97
R12614 VDD.n4433 VDD.n2453 1084.97
R12615 VDD.n4436 VDD.n2449 1084.97
R12616 VDD.n4436 VDD.n2447 1084.97
R12617 VDD.n2450 VDD.n2449 1084.97
R12618 VDD.n4325 VDD.n4324 1084.97
R12619 VDD.n4324 VDD.n4318 1084.97
R12620 VDD.n4318 VDD.n2574 1084.97
R12621 VDD.n4325 VDD.n2574 1084.97
R12622 VDD.n4335 VDD.n4334 1084.97
R12623 VDD.n4334 VDD.n2571 1084.97
R12624 VDD.n2571 VDD.n2564 1084.97
R12625 VDD.n4335 VDD.n2564 1084.97
R12626 VDD.n4345 VDD.n4344 1084.97
R12627 VDD.n4344 VDD.n2561 1084.97
R12628 VDD.n2561 VDD.n2553 1084.97
R12629 VDD.n4345 VDD.n2553 1084.97
R12630 VDD.n4355 VDD.n4354 1084.97
R12631 VDD.n4354 VDD.n2550 1084.97
R12632 VDD.n2550 VDD.n2540 1084.97
R12633 VDD.n4355 VDD.n2540 1084.97
R12634 VDD.n4365 VDD.n4364 1084.97
R12635 VDD.n4364 VDD.n2537 1084.97
R12636 VDD.n2537 VDD.n2528 1084.97
R12637 VDD.n4365 VDD.n2528 1084.97
R12638 VDD.n4372 VDD.n2525 1084.97
R12639 VDD.n4372 VDD.n2526 1084.97
R12640 VDD.n4376 VDD.n2526 1084.97
R12641 VDD.n4376 VDD.n2525 1084.97
R12642 VDD.n4385 VDD.n2512 1084.97
R12643 VDD.n2524 VDD.n2512 1084.97
R12644 VDD.n2524 VDD.n2511 1084.97
R12645 VDD.n4385 VDD.n2511 1084.97
R12646 VDD.n2504 VDD.n2498 1084.97
R12647 VDD.n2516 VDD.n2504 1084.97
R12648 VDD.n2516 VDD.n2513 1084.97
R12649 VDD.n2513 VDD.n2498 1084.97
R12650 VDD.n4399 VDD.n4398 1084.97
R12651 VDD.n4398 VDD.n2495 1084.97
R12652 VDD.n2495 VDD.n2486 1084.97
R12653 VDD.n4399 VDD.n2486 1084.97
R12654 VDD.n4409 VDD.n4408 1084.97
R12655 VDD.n4408 VDD.n2483 1084.97
R12656 VDD.n2483 VDD.n2473 1084.97
R12657 VDD.n4409 VDD.n2473 1084.97
R12658 VDD.n4419 VDD.n4418 1084.97
R12659 VDD.n4418 VDD.n2470 1084.97
R12660 VDD.n2470 VDD.n2463 1084.97
R12661 VDD.n4419 VDD.n2463 1084.97
R12662 VDD.n4429 VDD.n4428 1084.97
R12663 VDD.n4428 VDD.n2460 1084.97
R12664 VDD.n2460 VDD.n2452 1084.97
R12665 VDD.n4429 VDD.n2452 1084.97
R12666 VDD.n4393 VDD.n2499 1084.97
R12667 VDD.n2518 VDD.n2499 1084.97
R12668 VDD.n4393 VDD.n2500 1084.97
R12669 VDD.n2518 VDD.n2500 1084.97
R12670 VDD.n4197 VDD.n2711 1084.97
R12671 VDD.n4197 VDD.n2712 1084.97
R12672 VDD.n4204 VDD.n2712 1084.97
R12673 VDD.n4204 VDD.n2711 1084.97
R12674 VDD.n4207 VDD.n2701 1084.97
R12675 VDD.n4207 VDD.n2702 1084.97
R12676 VDD.n4214 VDD.n2702 1084.97
R12677 VDD.n4214 VDD.n2701 1084.97
R12678 VDD.n4217 VDD.n2690 1084.97
R12679 VDD.n4217 VDD.n2691 1084.97
R12680 VDD.n4224 VDD.n2691 1084.97
R12681 VDD.n4224 VDD.n2690 1084.97
R12682 VDD.n4227 VDD.n2677 1084.97
R12683 VDD.n4227 VDD.n2678 1084.97
R12684 VDD.n4234 VDD.n2678 1084.97
R12685 VDD.n4234 VDD.n2677 1084.97
R12686 VDD.n4237 VDD.n2665 1084.97
R12687 VDD.n4237 VDD.n2666 1084.97
R12688 VDD.n4244 VDD.n2666 1084.97
R12689 VDD.n4244 VDD.n2665 1084.97
R12690 VDD.n4259 VDD.n4255 1084.97
R12691 VDD.n4255 VDD.n2645 1084.97
R12692 VDD.n4254 VDD.n2645 1084.97
R12693 VDD.n4259 VDD.n4254 1084.97
R12694 VDD.n4271 VDD.n2623 1084.97
R12695 VDD.n4271 VDD.n2624 1084.97
R12696 VDD.n4278 VDD.n2624 1084.97
R12697 VDD.n4278 VDD.n2623 1084.97
R12698 VDD.n4281 VDD.n2610 1084.97
R12699 VDD.n4281 VDD.n2611 1084.97
R12700 VDD.n4288 VDD.n2611 1084.97
R12701 VDD.n4288 VDD.n2610 1084.97
R12702 VDD.n4291 VDD.n2600 1084.97
R12703 VDD.n4291 VDD.n2601 1084.97
R12704 VDD.n4298 VDD.n2601 1084.97
R12705 VDD.n4298 VDD.n2600 1084.97
R12706 VDD.n4301 VDD.n2589 1084.97
R12707 VDD.n4301 VDD.n2590 1084.97
R12708 VDD.n4308 VDD.n2590 1084.97
R12709 VDD.n4308 VDD.n2589 1084.97
R12710 VDD.n4311 VDD.n2585 1084.97
R12711 VDD.n4311 VDD.n2583 1084.97
R12712 VDD.n2586 VDD.n2585 1084.97
R12713 VDD.n4200 VDD.n4199 1084.97
R12714 VDD.n4199 VDD.n4193 1084.97
R12715 VDD.n4193 VDD.n2710 1084.97
R12716 VDD.n4200 VDD.n2710 1084.97
R12717 VDD.n4210 VDD.n4209 1084.97
R12718 VDD.n4209 VDD.n2707 1084.97
R12719 VDD.n2707 VDD.n2700 1084.97
R12720 VDD.n4210 VDD.n2700 1084.97
R12721 VDD.n4220 VDD.n4219 1084.97
R12722 VDD.n4219 VDD.n2697 1084.97
R12723 VDD.n2697 VDD.n2689 1084.97
R12724 VDD.n4220 VDD.n2689 1084.97
R12725 VDD.n4230 VDD.n4229 1084.97
R12726 VDD.n4229 VDD.n2686 1084.97
R12727 VDD.n2686 VDD.n2676 1084.97
R12728 VDD.n4230 VDD.n2676 1084.97
R12729 VDD.n4240 VDD.n4239 1084.97
R12730 VDD.n4239 VDD.n2673 1084.97
R12731 VDD.n2673 VDD.n2664 1084.97
R12732 VDD.n4240 VDD.n2664 1084.97
R12733 VDD.n4247 VDD.n2661 1084.97
R12734 VDD.n4247 VDD.n2662 1084.97
R12735 VDD.n4251 VDD.n2662 1084.97
R12736 VDD.n4251 VDD.n2661 1084.97
R12737 VDD.n4260 VDD.n2648 1084.97
R12738 VDD.n2660 VDD.n2648 1084.97
R12739 VDD.n2660 VDD.n2647 1084.97
R12740 VDD.n4260 VDD.n2647 1084.97
R12741 VDD.n2640 VDD.n2634 1084.97
R12742 VDD.n2652 VDD.n2640 1084.97
R12743 VDD.n2652 VDD.n2649 1084.97
R12744 VDD.n2649 VDD.n2634 1084.97
R12745 VDD.n4274 VDD.n4273 1084.97
R12746 VDD.n4273 VDD.n2631 1084.97
R12747 VDD.n2631 VDD.n2622 1084.97
R12748 VDD.n4274 VDD.n2622 1084.97
R12749 VDD.n4284 VDD.n4283 1084.97
R12750 VDD.n4283 VDD.n2619 1084.97
R12751 VDD.n2619 VDD.n2609 1084.97
R12752 VDD.n4284 VDD.n2609 1084.97
R12753 VDD.n4294 VDD.n4293 1084.97
R12754 VDD.n4293 VDD.n2606 1084.97
R12755 VDD.n2606 VDD.n2599 1084.97
R12756 VDD.n4294 VDD.n2599 1084.97
R12757 VDD.n4304 VDD.n4303 1084.97
R12758 VDD.n4303 VDD.n2596 1084.97
R12759 VDD.n2596 VDD.n2588 1084.97
R12760 VDD.n4304 VDD.n2588 1084.97
R12761 VDD.n4268 VDD.n2635 1084.97
R12762 VDD.n2654 VDD.n2635 1084.97
R12763 VDD.n4268 VDD.n2636 1084.97
R12764 VDD.n2654 VDD.n2636 1084.97
R12765 VDD.n4072 VDD.n2847 1084.97
R12766 VDD.n4072 VDD.n2848 1084.97
R12767 VDD.n4079 VDD.n2848 1084.97
R12768 VDD.n4079 VDD.n2847 1084.97
R12769 VDD.n4082 VDD.n2837 1084.97
R12770 VDD.n4082 VDD.n2838 1084.97
R12771 VDD.n4089 VDD.n2838 1084.97
R12772 VDD.n4089 VDD.n2837 1084.97
R12773 VDD.n4092 VDD.n2826 1084.97
R12774 VDD.n4092 VDD.n2827 1084.97
R12775 VDD.n4099 VDD.n2827 1084.97
R12776 VDD.n4099 VDD.n2826 1084.97
R12777 VDD.n4102 VDD.n2813 1084.97
R12778 VDD.n4102 VDD.n2814 1084.97
R12779 VDD.n4109 VDD.n2814 1084.97
R12780 VDD.n4109 VDD.n2813 1084.97
R12781 VDD.n4112 VDD.n2801 1084.97
R12782 VDD.n4112 VDD.n2802 1084.97
R12783 VDD.n4119 VDD.n2802 1084.97
R12784 VDD.n4119 VDD.n2801 1084.97
R12785 VDD.n4134 VDD.n4130 1084.97
R12786 VDD.n4130 VDD.n2781 1084.97
R12787 VDD.n4129 VDD.n2781 1084.97
R12788 VDD.n4134 VDD.n4129 1084.97
R12789 VDD.n4146 VDD.n2759 1084.97
R12790 VDD.n4146 VDD.n2760 1084.97
R12791 VDD.n4153 VDD.n2760 1084.97
R12792 VDD.n4153 VDD.n2759 1084.97
R12793 VDD.n4156 VDD.n2746 1084.97
R12794 VDD.n4156 VDD.n2747 1084.97
R12795 VDD.n4163 VDD.n2747 1084.97
R12796 VDD.n4163 VDD.n2746 1084.97
R12797 VDD.n4166 VDD.n2736 1084.97
R12798 VDD.n4166 VDD.n2737 1084.97
R12799 VDD.n4173 VDD.n2737 1084.97
R12800 VDD.n4173 VDD.n2736 1084.97
R12801 VDD.n4176 VDD.n2725 1084.97
R12802 VDD.n4176 VDD.n2726 1084.97
R12803 VDD.n4183 VDD.n2726 1084.97
R12804 VDD.n4183 VDD.n2725 1084.97
R12805 VDD.n4186 VDD.n2721 1084.97
R12806 VDD.n4186 VDD.n2719 1084.97
R12807 VDD.n2722 VDD.n2721 1084.97
R12808 VDD.n4075 VDD.n4074 1084.97
R12809 VDD.n4074 VDD.n4068 1084.97
R12810 VDD.n4068 VDD.n2846 1084.97
R12811 VDD.n4075 VDD.n2846 1084.97
R12812 VDD.n4085 VDD.n4084 1084.97
R12813 VDD.n4084 VDD.n2843 1084.97
R12814 VDD.n2843 VDD.n2836 1084.97
R12815 VDD.n4085 VDD.n2836 1084.97
R12816 VDD.n4095 VDD.n4094 1084.97
R12817 VDD.n4094 VDD.n2833 1084.97
R12818 VDD.n2833 VDD.n2825 1084.97
R12819 VDD.n4095 VDD.n2825 1084.97
R12820 VDD.n4105 VDD.n4104 1084.97
R12821 VDD.n4104 VDD.n2822 1084.97
R12822 VDD.n2822 VDD.n2812 1084.97
R12823 VDD.n4105 VDD.n2812 1084.97
R12824 VDD.n4115 VDD.n4114 1084.97
R12825 VDD.n4114 VDD.n2809 1084.97
R12826 VDD.n2809 VDD.n2800 1084.97
R12827 VDD.n4115 VDD.n2800 1084.97
R12828 VDD.n4122 VDD.n2797 1084.97
R12829 VDD.n4122 VDD.n2798 1084.97
R12830 VDD.n4126 VDD.n2798 1084.97
R12831 VDD.n4126 VDD.n2797 1084.97
R12832 VDD.n4135 VDD.n2784 1084.97
R12833 VDD.n2796 VDD.n2784 1084.97
R12834 VDD.n2796 VDD.n2783 1084.97
R12835 VDD.n4135 VDD.n2783 1084.97
R12836 VDD.n2776 VDD.n2770 1084.97
R12837 VDD.n2788 VDD.n2776 1084.97
R12838 VDD.n2788 VDD.n2785 1084.97
R12839 VDD.n2785 VDD.n2770 1084.97
R12840 VDD.n4149 VDD.n4148 1084.97
R12841 VDD.n4148 VDD.n2767 1084.97
R12842 VDD.n2767 VDD.n2758 1084.97
R12843 VDD.n4149 VDD.n2758 1084.97
R12844 VDD.n4159 VDD.n4158 1084.97
R12845 VDD.n4158 VDD.n2755 1084.97
R12846 VDD.n2755 VDD.n2745 1084.97
R12847 VDD.n4159 VDD.n2745 1084.97
R12848 VDD.n4169 VDD.n4168 1084.97
R12849 VDD.n4168 VDD.n2742 1084.97
R12850 VDD.n2742 VDD.n2735 1084.97
R12851 VDD.n4169 VDD.n2735 1084.97
R12852 VDD.n4179 VDD.n4178 1084.97
R12853 VDD.n4178 VDD.n2732 1084.97
R12854 VDD.n2732 VDD.n2724 1084.97
R12855 VDD.n4179 VDD.n2724 1084.97
R12856 VDD.n4143 VDD.n2771 1084.97
R12857 VDD.n2790 VDD.n2771 1084.97
R12858 VDD.n4143 VDD.n2772 1084.97
R12859 VDD.n2790 VDD.n2772 1084.97
R12860 VDD.n3947 VDD.n2983 1084.97
R12861 VDD.n3947 VDD.n2984 1084.97
R12862 VDD.n3954 VDD.n2984 1084.97
R12863 VDD.n3954 VDD.n2983 1084.97
R12864 VDD.n3957 VDD.n2973 1084.97
R12865 VDD.n3957 VDD.n2974 1084.97
R12866 VDD.n3964 VDD.n2974 1084.97
R12867 VDD.n3964 VDD.n2973 1084.97
R12868 VDD.n3967 VDD.n2962 1084.97
R12869 VDD.n3967 VDD.n2963 1084.97
R12870 VDD.n3974 VDD.n2963 1084.97
R12871 VDD.n3974 VDD.n2962 1084.97
R12872 VDD.n3977 VDD.n2949 1084.97
R12873 VDD.n3977 VDD.n2950 1084.97
R12874 VDD.n3984 VDD.n2950 1084.97
R12875 VDD.n3984 VDD.n2949 1084.97
R12876 VDD.n3987 VDD.n2937 1084.97
R12877 VDD.n3987 VDD.n2938 1084.97
R12878 VDD.n3994 VDD.n2938 1084.97
R12879 VDD.n3994 VDD.n2937 1084.97
R12880 VDD.n4009 VDD.n4005 1084.97
R12881 VDD.n4005 VDD.n2917 1084.97
R12882 VDD.n4004 VDD.n2917 1084.97
R12883 VDD.n4009 VDD.n4004 1084.97
R12884 VDD.n4021 VDD.n2895 1084.97
R12885 VDD.n4021 VDD.n2896 1084.97
R12886 VDD.n4028 VDD.n2896 1084.97
R12887 VDD.n4028 VDD.n2895 1084.97
R12888 VDD.n4031 VDD.n2882 1084.97
R12889 VDD.n4031 VDD.n2883 1084.97
R12890 VDD.n4038 VDD.n2883 1084.97
R12891 VDD.n4038 VDD.n2882 1084.97
R12892 VDD.n4041 VDD.n2872 1084.97
R12893 VDD.n4041 VDD.n2873 1084.97
R12894 VDD.n4048 VDD.n2873 1084.97
R12895 VDD.n4048 VDD.n2872 1084.97
R12896 VDD.n4051 VDD.n2861 1084.97
R12897 VDD.n4051 VDD.n2862 1084.97
R12898 VDD.n4058 VDD.n2862 1084.97
R12899 VDD.n4058 VDD.n2861 1084.97
R12900 VDD.n4061 VDD.n2857 1084.97
R12901 VDD.n4061 VDD.n2855 1084.97
R12902 VDD.n2858 VDD.n2857 1084.97
R12903 VDD.n3950 VDD.n3949 1084.97
R12904 VDD.n3949 VDD.n3943 1084.97
R12905 VDD.n3943 VDD.n2982 1084.97
R12906 VDD.n3950 VDD.n2982 1084.97
R12907 VDD.n3960 VDD.n3959 1084.97
R12908 VDD.n3959 VDD.n2979 1084.97
R12909 VDD.n2979 VDD.n2972 1084.97
R12910 VDD.n3960 VDD.n2972 1084.97
R12911 VDD.n3970 VDD.n3969 1084.97
R12912 VDD.n3969 VDD.n2969 1084.97
R12913 VDD.n2969 VDD.n2961 1084.97
R12914 VDD.n3970 VDD.n2961 1084.97
R12915 VDD.n3980 VDD.n3979 1084.97
R12916 VDD.n3979 VDD.n2958 1084.97
R12917 VDD.n2958 VDD.n2948 1084.97
R12918 VDD.n3980 VDD.n2948 1084.97
R12919 VDD.n3990 VDD.n3989 1084.97
R12920 VDD.n3989 VDD.n2945 1084.97
R12921 VDD.n2945 VDD.n2936 1084.97
R12922 VDD.n3990 VDD.n2936 1084.97
R12923 VDD.n3997 VDD.n2933 1084.97
R12924 VDD.n3997 VDD.n2934 1084.97
R12925 VDD.n4001 VDD.n2934 1084.97
R12926 VDD.n4001 VDD.n2933 1084.97
R12927 VDD.n4010 VDD.n2920 1084.97
R12928 VDD.n2932 VDD.n2920 1084.97
R12929 VDD.n2932 VDD.n2919 1084.97
R12930 VDD.n4010 VDD.n2919 1084.97
R12931 VDD.n2912 VDD.n2906 1084.97
R12932 VDD.n2924 VDD.n2912 1084.97
R12933 VDD.n2924 VDD.n2921 1084.97
R12934 VDD.n2921 VDD.n2906 1084.97
R12935 VDD.n4024 VDD.n4023 1084.97
R12936 VDD.n4023 VDD.n2903 1084.97
R12937 VDD.n2903 VDD.n2894 1084.97
R12938 VDD.n4024 VDD.n2894 1084.97
R12939 VDD.n4034 VDD.n4033 1084.97
R12940 VDD.n4033 VDD.n2891 1084.97
R12941 VDD.n2891 VDD.n2881 1084.97
R12942 VDD.n4034 VDD.n2881 1084.97
R12943 VDD.n4044 VDD.n4043 1084.97
R12944 VDD.n4043 VDD.n2878 1084.97
R12945 VDD.n2878 VDD.n2871 1084.97
R12946 VDD.n4044 VDD.n2871 1084.97
R12947 VDD.n4054 VDD.n4053 1084.97
R12948 VDD.n4053 VDD.n2868 1084.97
R12949 VDD.n2868 VDD.n2860 1084.97
R12950 VDD.n4054 VDD.n2860 1084.97
R12951 VDD.n4018 VDD.n2907 1084.97
R12952 VDD.n2926 VDD.n2907 1084.97
R12953 VDD.n4018 VDD.n2908 1084.97
R12954 VDD.n2926 VDD.n2908 1084.97
R12955 VDD.n3599 VDD.n3277 1084.97
R12956 VDD.n3599 VDD.n3278 1084.97
R12957 VDD.n3606 VDD.n3278 1084.97
R12958 VDD.n3606 VDD.n3277 1084.97
R12959 VDD.n3614 VDD.n3610 1084.97
R12960 VDD.n3610 VDD.n3267 1084.97
R12961 VDD.n3609 VDD.n3267 1084.97
R12962 VDD.n3614 VDD.n3609 1084.97
R12963 VDD.n3299 VDD.n3286 1084.97
R12964 VDD.n3299 VDD.n3298 1084.97
R12965 VDD.n3298 VDD.n3292 1084.97
R12966 VDD.n3292 VDD.n3286 1084.97
R12967 VDD.n3602 VDD.n3601 1084.97
R12968 VDD.n3601 VDD.n3283 1084.97
R12969 VDD.n3283 VDD.n3276 1084.97
R12970 VDD.n3602 VDD.n3276 1084.97
R12971 VDD.n3615 VDD.n3270 1084.97
R12972 VDD.n3275 VDD.n3270 1084.97
R12973 VDD.n3275 VDD.n3269 1084.97
R12974 VDD.n3615 VDD.n3269 1084.97
R12975 VDD.n3596 VDD.n3287 1084.97
R12976 VDD.n3296 VDD.n3287 1084.97
R12977 VDD.n3596 VDD.n3288 1084.97
R12978 VDD.n3296 VDD.n3288 1084.97
R12979 VDD.n3446 VDD.n3346 1084.97
R12980 VDD.n3443 VDD.n3344 1084.97
R12981 VDD.n3443 VDD.n3346 1084.97
R12982 VDD.n3441 VDD.n3347 1084.97
R12983 VDD.n3441 VDD.n3348 1084.97
R12984 VDD.n3429 VDD.n3348 1084.97
R12985 VDD.n3429 VDD.n3347 1084.97
R12986 VDD.n3427 VDD.n3426 1084.97
R12987 VDD.n3432 VDD.n3426 1084.97
R12988 VDD.n3432 VDD.n3424 1084.97
R12989 VDD.n3483 VDD.n3455 1084.97
R12990 VDD.n3480 VDD.n3453 1084.97
R12991 VDD.n3480 VDD.n3455 1084.97
R12992 VDD.n3478 VDD.n3456 1084.97
R12993 VDD.n3478 VDD.n3457 1084.97
R12994 VDD.n3467 VDD.n3457 1084.97
R12995 VDD.n3467 VDD.n3456 1084.97
R12996 VDD.n3465 VDD.n3464 1084.97
R12997 VDD.n3470 VDD.n3464 1084.97
R12998 VDD.n3470 VDD.n3462 1084.97
R12999 VDD.n3335 VDD.n3329 1084.97
R13000 VDD.n3332 VDD.n3327 1084.97
R13001 VDD.n3332 VDD.n3329 1084.97
R13002 VDD.n3330 VDD.n3322 1084.97
R13003 VDD.n3330 VDD.n3323 1084.97
R13004 VDD.n3507 VDD.n3323 1084.97
R13005 VDD.n3507 VDD.n3322 1084.97
R13006 VDD.n3320 VDD.n3319 1084.97
R13007 VDD.n3510 VDD.n3319 1084.97
R13008 VDD.n3510 VDD.n3317 1084.97
R13009 VDD.n3541 VDD.n3309 1084.97
R13010 VDD.n3538 VDD.n3307 1084.97
R13011 VDD.n3538 VDD.n3309 1084.97
R13012 VDD.n3536 VDD.n3310 1084.97
R13013 VDD.n3536 VDD.n3311 1084.97
R13014 VDD.n3524 VDD.n3311 1084.97
R13015 VDD.n3524 VDD.n3310 1084.97
R13016 VDD.n3522 VDD.n3521 1084.97
R13017 VDD.n3527 VDD.n3521 1084.97
R13018 VDD.n3527 VDD.n3519 1084.97
R13019 VDD.n3577 VDD.n3549 1084.97
R13020 VDD.n3574 VDD.n3547 1084.97
R13021 VDD.n3574 VDD.n3549 1084.97
R13022 VDD.n3572 VDD.n3550 1084.97
R13023 VDD.n3572 VDD.n3551 1084.97
R13024 VDD.n3561 VDD.n3551 1084.97
R13025 VDD.n3561 VDD.n3550 1084.97
R13026 VDD.n3559 VDD.n3558 1084.97
R13027 VDD.n3564 VDD.n3558 1084.97
R13028 VDD.n3564 VDD.n3556 1084.97
R13029 VDD.n3391 VDD.n3385 1084.97
R13030 VDD.n3388 VDD.n3383 1084.97
R13031 VDD.n3388 VDD.n3385 1084.97
R13032 VDD.n3386 VDD.n3378 1084.97
R13033 VDD.n3386 VDD.n3379 1084.97
R13034 VDD.n3412 VDD.n3379 1084.97
R13035 VDD.n3412 VDD.n3378 1084.97
R13036 VDD.n3376 VDD.n3375 1084.97
R13037 VDD.n3415 VDD.n3375 1084.97
R13038 VDD.n3415 VDD.n3373 1084.97
R13039 VDD.n3822 VDD.n3809 1084.97
R13040 VDD.n3822 VDD.n3810 1084.97
R13041 VDD.n3829 VDD.n3810 1084.97
R13042 VDD.n3829 VDD.n3809 1084.97
R13043 VDD.n3832 VDD.n3799 1084.97
R13044 VDD.n3832 VDD.n3800 1084.97
R13045 VDD.n3839 VDD.n3800 1084.97
R13046 VDD.n3839 VDD.n3799 1084.97
R13047 VDD.n3842 VDD.n3788 1084.97
R13048 VDD.n3842 VDD.n3789 1084.97
R13049 VDD.n3849 VDD.n3789 1084.97
R13050 VDD.n3849 VDD.n3788 1084.97
R13051 VDD.n3852 VDD.n3775 1084.97
R13052 VDD.n3852 VDD.n3776 1084.97
R13053 VDD.n3859 VDD.n3776 1084.97
R13054 VDD.n3859 VDD.n3775 1084.97
R13055 VDD.n3862 VDD.n3763 1084.97
R13056 VDD.n3862 VDD.n3764 1084.97
R13057 VDD.n3869 VDD.n3764 1084.97
R13058 VDD.n3869 VDD.n3763 1084.97
R13059 VDD.n3884 VDD.n3880 1084.97
R13060 VDD.n3880 VDD.n3743 1084.97
R13061 VDD.n3879 VDD.n3743 1084.97
R13062 VDD.n3884 VDD.n3879 1084.97
R13063 VDD.n3896 VDD.n3031 1084.97
R13064 VDD.n3896 VDD.n3032 1084.97
R13065 VDD.n3903 VDD.n3032 1084.97
R13066 VDD.n3903 VDD.n3031 1084.97
R13067 VDD.n3906 VDD.n3018 1084.97
R13068 VDD.n3906 VDD.n3019 1084.97
R13069 VDD.n3913 VDD.n3019 1084.97
R13070 VDD.n3913 VDD.n3018 1084.97
R13071 VDD.n3916 VDD.n3008 1084.97
R13072 VDD.n3916 VDD.n3009 1084.97
R13073 VDD.n3923 VDD.n3009 1084.97
R13074 VDD.n3923 VDD.n3008 1084.97
R13075 VDD.n3926 VDD.n2997 1084.97
R13076 VDD.n3926 VDD.n2998 1084.97
R13077 VDD.n3933 VDD.n2998 1084.97
R13078 VDD.n3933 VDD.n2997 1084.97
R13079 VDD.n3936 VDD.n2993 1084.97
R13080 VDD.n3936 VDD.n2991 1084.97
R13081 VDD.n2994 VDD.n2993 1084.97
R13082 VDD.n3825 VDD.n3824 1084.97
R13083 VDD.n3824 VDD.n3818 1084.97
R13084 VDD.n3818 VDD.n3808 1084.97
R13085 VDD.n3825 VDD.n3808 1084.97
R13086 VDD.n3835 VDD.n3834 1084.97
R13087 VDD.n3834 VDD.n3805 1084.97
R13088 VDD.n3805 VDD.n3798 1084.97
R13089 VDD.n3835 VDD.n3798 1084.97
R13090 VDD.n3845 VDD.n3844 1084.97
R13091 VDD.n3844 VDD.n3795 1084.97
R13092 VDD.n3795 VDD.n3787 1084.97
R13093 VDD.n3845 VDD.n3787 1084.97
R13094 VDD.n3855 VDD.n3854 1084.97
R13095 VDD.n3854 VDD.n3784 1084.97
R13096 VDD.n3784 VDD.n3774 1084.97
R13097 VDD.n3855 VDD.n3774 1084.97
R13098 VDD.n3865 VDD.n3864 1084.97
R13099 VDD.n3864 VDD.n3771 1084.97
R13100 VDD.n3771 VDD.n3762 1084.97
R13101 VDD.n3865 VDD.n3762 1084.97
R13102 VDD.n3872 VDD.n3759 1084.97
R13103 VDD.n3872 VDD.n3760 1084.97
R13104 VDD.n3876 VDD.n3760 1084.97
R13105 VDD.n3876 VDD.n3759 1084.97
R13106 VDD.n3885 VDD.n3746 1084.97
R13107 VDD.n3758 VDD.n3746 1084.97
R13108 VDD.n3758 VDD.n3745 1084.97
R13109 VDD.n3885 VDD.n3745 1084.97
R13110 VDD.n3738 VDD.n3732 1084.97
R13111 VDD.n3750 VDD.n3738 1084.97
R13112 VDD.n3750 VDD.n3747 1084.97
R13113 VDD.n3747 VDD.n3732 1084.97
R13114 VDD.n3899 VDD.n3898 1084.97
R13115 VDD.n3898 VDD.n3729 1084.97
R13116 VDD.n3729 VDD.n3030 1084.97
R13117 VDD.n3899 VDD.n3030 1084.97
R13118 VDD.n3909 VDD.n3908 1084.97
R13119 VDD.n3908 VDD.n3027 1084.97
R13120 VDD.n3027 VDD.n3017 1084.97
R13121 VDD.n3909 VDD.n3017 1084.97
R13122 VDD.n3919 VDD.n3918 1084.97
R13123 VDD.n3918 VDD.n3014 1084.97
R13124 VDD.n3014 VDD.n3007 1084.97
R13125 VDD.n3919 VDD.n3007 1084.97
R13126 VDD.n3929 VDD.n3928 1084.97
R13127 VDD.n3928 VDD.n3004 1084.97
R13128 VDD.n3004 VDD.n2996 1084.97
R13129 VDD.n3929 VDD.n2996 1084.97
R13130 VDD.n3893 VDD.n3733 1084.97
R13131 VDD.n3752 VDD.n3733 1084.97
R13132 VDD.n3893 VDD.n3734 1084.97
R13133 VDD.n3752 VDD.n3734 1084.97
R13134 VDD.n328 VDD.n303 516.932
R13135 VDD.n303 VDD.n294 516.932
R13136 VDD.n330 VDD.n300 516.932
R13137 VDD.n300 VDD.n295 516.932
R13138 VDD.n175 VDD.n174 295.125
R13139 VDD.n210 VDD.n209 295.125
R13140 VDD.n245 VDD.n244 295.125
R13141 VDD.n280 VDD.n279 295.125
R13142 VDD.n7024 VDD.n7023 295.125
R13143 VDD.n7059 VDD.n7058 295.125
R13144 VDD.n7094 VDD.n7093 295.125
R13145 VDD.n6906 VDD.n6905 295.125
R13146 VDD.n154 VDD.t370 253.119
R13147 VDD.n153 VDD.t213 253.119
R13148 VDD.n175 VDD.t846 253.119
R13149 VDD.n174 VDD.t1072 253.119
R13150 VDD.n168 VDD.t1072 253.119
R13151 VDD.n167 VDD.t654 253.119
R13152 VDD.n189 VDD.t128 253.119
R13153 VDD.n188 VDD.t619 253.119
R13154 VDD.n210 VDD.t170 253.119
R13155 VDD.n209 VDD.t1026 253.119
R13156 VDD.n203 VDD.t1026 253.119
R13157 VDD.n202 VDD.t976 253.119
R13158 VDD.n224 VDD.t921 253.119
R13159 VDD.n223 VDD.t838 253.119
R13160 VDD.n245 VDD.t878 253.119
R13161 VDD.n244 VDD.t1065 253.119
R13162 VDD.n238 VDD.t1065 253.119
R13163 VDD.n237 VDD.t957 253.119
R13164 VDD.n259 VDD.t646 253.119
R13165 VDD.n258 VDD.t351 253.119
R13166 VDD.n280 VDD.t629 253.119
R13167 VDD.n279 VDD.t1089 253.119
R13168 VDD.n273 VDD.t1089 253.119
R13169 VDD.n272 VDD.t77 253.119
R13170 VDD.n7003 VDD.t968 253.119
R13171 VDD.n7002 VDD.t939 253.119
R13172 VDD.n7024 VDD.t931 253.119
R13173 VDD.n7023 VDD.t954 253.119
R13174 VDD.n7017 VDD.t954 253.119
R13175 VDD.n7016 VDD.t1036 253.119
R13176 VDD.n7038 VDD.t71 253.119
R13177 VDD.n7037 VDD.t126 253.119
R13178 VDD.n7059 VDD.t189 253.119
R13179 VDD.n7058 VDD.t420 253.119
R13180 VDD.n7052 VDD.t420 253.119
R13181 VDD.n7051 VDD.t1012 253.119
R13182 VDD.n7073 VDD.t791 253.119
R13183 VDD.n7072 VDD.t798 253.119
R13184 VDD.n7094 VDD.t583 253.119
R13185 VDD.n7093 VDD.t399 253.119
R13186 VDD.n7087 VDD.t399 253.119
R13187 VDD.n7086 VDD.t1040 253.119
R13188 VDD.n7108 VDD.t276 253.119
R13189 VDD.n7107 VDD.t773 253.119
R13190 VDD.n6905 VDD.t301 253.119
R13191 VDD.t950 VDD.n6906 253.119
R13192 VDD.t950 VDD.n7122 253.119
R13193 VDD.n7121 VDD.t1008 253.119
R13194 VDD.n3431 VDD.t854 253.119
R13195 VDD.n3430 VDD.t176 253.119
R13196 VDD.n3442 VDD.t176 253.119
R13197 VDD.t985 VDD.n3444 253.119
R13198 VDD.n3469 VDD.t810 253.119
R13199 VDD.n3468 VDD.t812 253.119
R13200 VDD.n3479 VDD.t812 253.119
R13201 VDD.t131 VDD.n3481 253.119
R13202 VDD.n3509 VDD.t271 253.119
R13203 VDD.n3508 VDD.t256 253.119
R13204 VDD.n3331 VDD.t256 253.119
R13205 VDD.t884 VDD.n3333 253.119
R13206 VDD.n3526 VDD.t996 253.119
R13207 VDD.n3525 VDD.t998 253.119
R13208 VDD.n3537 VDD.t998 253.119
R13209 VDD.t122 VDD.n3539 253.119
R13210 VDD.n3563 VDD.t408 253.119
R13211 VDD.n3562 VDD.t410 253.119
R13212 VDD.n3573 VDD.t410 253.119
R13213 VDD.t137 VDD.n3575 253.119
R13214 VDD.n3414 VDD.t782 253.119
R13215 VDD.n3413 VDD.t784 253.119
R13216 VDD.n3387 VDD.t784 253.119
R13217 VDD.t206 VDD.n3389 253.119
R13218 VDD.n148 VDD.n147 214.357
R13219 VDD.n142 VDD.n141 214.357
R13220 VDD.n162 VDD.n161 214.357
R13221 VDD.n126 VDD.n125 214.357
R13222 VDD.n183 VDD.n182 214.357
R13223 VDD.n117 VDD.n116 214.357
R13224 VDD.n197 VDD.n196 214.357
R13225 VDD.n101 VDD.n100 214.357
R13226 VDD.n218 VDD.n217 214.357
R13227 VDD.n92 VDD.n91 214.357
R13228 VDD.n232 VDD.n231 214.357
R13229 VDD.n76 VDD.n75 214.357
R13230 VDD.n253 VDD.n252 214.357
R13231 VDD.n67 VDD.n66 214.357
R13232 VDD.n267 VDD.n266 214.357
R13233 VDD.n51 VDD.n50 214.357
R13234 VDD.n7116 VDD.n7115 214.357
R13235 VDD.n6997 VDD.n6996 214.357
R13236 VDD.n6991 VDD.n6990 214.357
R13237 VDD.n7011 VDD.n7010 214.357
R13238 VDD.n6975 VDD.n6974 214.357
R13239 VDD.n7032 VDD.n7031 214.357
R13240 VDD.n6966 VDD.n6965 214.357
R13241 VDD.n7046 VDD.n7045 214.357
R13242 VDD.n6950 VDD.n6949 214.357
R13243 VDD.n7067 VDD.n7066 214.357
R13244 VDD.n6941 VDD.n6940 214.357
R13245 VDD.n7081 VDD.n7080 214.357
R13246 VDD.n6925 VDD.n6924 214.357
R13247 VDD.n7102 VDD.n7101 214.357
R13248 VDD.n6916 VDD.n6915 214.357
R13249 VDD.n6900 VDD.n6899 214.357
R13250 VDD.n3446 VDD.n3445 214.357
R13251 VDD.n3428 VDD.n3427 214.357
R13252 VDD.n3483 VDD.n3482 214.357
R13253 VDD.n3466 VDD.n3465 214.357
R13254 VDD.n3335 VDD.n3334 214.357
R13255 VDD.n3321 VDD.n3320 214.357
R13256 VDD.n3541 VDD.n3540 214.357
R13257 VDD.n3523 VDD.n3522 214.357
R13258 VDD.n3577 VDD.n3576 214.357
R13259 VDD.n3560 VDD.n3559 214.357
R13260 VDD.n3391 VDD.n3390 214.357
R13261 VDD.n3377 VDD.n3376 214.357
R13262 VDD.n7644 VDD.n7643 212.329
R13263 VDD.n7643 VDD.n7636 212.329
R13264 VDD.n7645 VDD.n7635 212.329
R13265 VDD.n7652 VDD.n7635 212.329
R13266 VDD.n7631 VDD.n7630 212.329
R13267 VDD.n7630 VDD.n7626 212.329
R13268 VDD.n7655 VDD.n7625 212.329
R13269 VDD.n7662 VDD.n7625 212.329
R13270 VDD.n7621 VDD.n7620 212.329
R13271 VDD.n7620 VDD.n7615 212.329
R13272 VDD.n7665 VDD.n7614 212.329
R13273 VDD.n7672 VDD.n7614 212.329
R13274 VDD.n7610 VDD.n7609 212.329
R13275 VDD.n7609 VDD.n7602 212.329
R13276 VDD.n7675 VDD.n7601 212.329
R13277 VDD.n7682 VDD.n7601 212.329
R13278 VDD.n7597 VDD.n7596 212.329
R13279 VDD.n7596 VDD.n7590 212.329
R13280 VDD.n7685 VDD.n7589 212.329
R13281 VDD.n7692 VDD.n7589 212.329
R13282 VDD.n7698 VDD.n7697 212.329
R13283 VDD.n7699 VDD.n7698 212.329
R13284 VDD.n7582 VDD.n7581 212.329
R13285 VDD.n7581 VDD.n7574 212.329
R13286 VDD.n7702 VDD.n7573 212.329
R13287 VDD.n7709 VDD.n7573 212.329
R13288 VDD.n7569 VDD.n7568 212.329
R13289 VDD.n7568 VDD.n7565 212.329
R13290 VDD.n7712 VDD.n7564 212.329
R13291 VDD.n7719 VDD.n7564 212.329
R13292 VDD.n7559 VDD.n7558 212.329
R13293 VDD.n7559 VDD.n7557 212.329
R13294 VDD.n7727 VDD.n7726 212.329
R13295 VDD.n7727 VDD.n7725 212.329
R13296 VDD.n14 VDD.n11 212.329
R13297 VDD.n15 VDD.n14 212.329
R13298 VDD.n7553 VDD.n10 212.329
R13299 VDD.n7546 VDD.n10 212.329
R13300 VDD.n27 VDD.n20 212.329
R13301 VDD.n28 VDD.n27 212.329
R13302 VDD.n7543 VDD.n19 212.329
R13303 VDD.n7536 VDD.n19 212.329
R13304 VDD.n37 VDD.n33 212.329
R13305 VDD.n38 VDD.n37 212.329
R13306 VDD.n7533 VDD.n32 212.329
R13307 VDD.n7526 VDD.n32 212.329
R13308 VDD.n7523 VDD.n41 212.329
R13309 VDD.n44 VDD.n41 212.329
R13310 VDD.n1777 VDD.n1776 212.329
R13311 VDD.n1776 VDD.n1769 212.329
R13312 VDD.n1778 VDD.n1768 212.329
R13313 VDD.n1785 VDD.n1768 212.329
R13314 VDD.n1764 VDD.n1763 212.329
R13315 VDD.n1763 VDD.n1759 212.329
R13316 VDD.n1788 VDD.n1758 212.329
R13317 VDD.n1795 VDD.n1758 212.329
R13318 VDD.n1754 VDD.n1753 212.329
R13319 VDD.n1753 VDD.n1748 212.329
R13320 VDD.n1798 VDD.n1747 212.329
R13321 VDD.n1805 VDD.n1747 212.329
R13322 VDD.n1743 VDD.n1742 212.329
R13323 VDD.n1742 VDD.n1735 212.329
R13324 VDD.n1808 VDD.n1734 212.329
R13325 VDD.n1815 VDD.n1734 212.329
R13326 VDD.n1730 VDD.n1729 212.329
R13327 VDD.n1729 VDD.n1723 212.329
R13328 VDD.n1818 VDD.n1722 212.329
R13329 VDD.n1825 VDD.n1722 212.329
R13330 VDD.n1831 VDD.n1830 212.329
R13331 VDD.n1832 VDD.n1831 212.329
R13332 VDD.n1715 VDD.n1714 212.329
R13333 VDD.n1714 VDD.n1707 212.329
R13334 VDD.n1835 VDD.n1706 212.329
R13335 VDD.n1842 VDD.n1706 212.329
R13336 VDD.n1702 VDD.n1701 212.329
R13337 VDD.n1701 VDD.n1697 212.329
R13338 VDD.n1845 VDD.n1696 212.329
R13339 VDD.n1852 VDD.n1696 212.329
R13340 VDD.n1692 VDD.n1691 212.329
R13341 VDD.n1691 VDD.n1686 212.329
R13342 VDD.n1855 VDD.n1685 212.329
R13343 VDD.n1862 VDD.n1685 212.329
R13344 VDD.n1681 VDD.n1680 212.329
R13345 VDD.n1680 VDD.n1673 212.329
R13346 VDD.n1865 VDD.n1672 212.329
R13347 VDD.n1872 VDD.n1672 212.329
R13348 VDD.n1668 VDD.n1667 212.329
R13349 VDD.n1667 VDD.n1663 212.329
R13350 VDD.n1875 VDD.n1662 212.329
R13351 VDD.n1882 VDD.n1662 212.329
R13352 VDD.n1658 VDD.n1657 212.329
R13353 VDD.n1657 VDD.n1652 212.329
R13354 VDD.n1885 VDD.n1651 212.329
R13355 VDD.n1892 VDD.n1651 212.329
R13356 VDD.n1897 VDD.n1644 212.329
R13357 VDD.n1644 VDD.n1642 212.329
R13358 VDD.n1517 VDD.n1516 212.329
R13359 VDD.n1516 VDD.n1509 212.329
R13360 VDD.n1518 VDD.n1508 212.329
R13361 VDD.n1525 VDD.n1508 212.329
R13362 VDD.n1504 VDD.n1503 212.329
R13363 VDD.n1503 VDD.n1499 212.329
R13364 VDD.n1528 VDD.n1498 212.329
R13365 VDD.n1535 VDD.n1498 212.329
R13366 VDD.n1494 VDD.n1493 212.329
R13367 VDD.n1493 VDD.n1488 212.329
R13368 VDD.n1538 VDD.n1487 212.329
R13369 VDD.n1545 VDD.n1487 212.329
R13370 VDD.n1483 VDD.n1482 212.329
R13371 VDD.n1482 VDD.n1475 212.329
R13372 VDD.n1548 VDD.n1474 212.329
R13373 VDD.n1555 VDD.n1474 212.329
R13374 VDD.n1470 VDD.n1469 212.329
R13375 VDD.n1469 VDD.n1463 212.329
R13376 VDD.n1558 VDD.n1462 212.329
R13377 VDD.n1565 VDD.n1462 212.329
R13378 VDD.n1571 VDD.n1570 212.329
R13379 VDD.n1572 VDD.n1571 212.329
R13380 VDD.n1455 VDD.n1454 212.329
R13381 VDD.n1454 VDD.n1447 212.329
R13382 VDD.n1575 VDD.n1446 212.329
R13383 VDD.n1582 VDD.n1446 212.329
R13384 VDD.n1442 VDD.n1441 212.329
R13385 VDD.n1441 VDD.n1437 212.329
R13386 VDD.n1585 VDD.n1436 212.329
R13387 VDD.n1592 VDD.n1436 212.329
R13388 VDD.n1432 VDD.n1431 212.329
R13389 VDD.n1431 VDD.n1426 212.329
R13390 VDD.n1595 VDD.n1425 212.329
R13391 VDD.n1602 VDD.n1425 212.329
R13392 VDD.n1421 VDD.n1420 212.329
R13393 VDD.n1420 VDD.n1413 212.329
R13394 VDD.n1605 VDD.n1412 212.329
R13395 VDD.n1612 VDD.n1412 212.329
R13396 VDD.n1408 VDD.n1407 212.329
R13397 VDD.n1407 VDD.n1403 212.329
R13398 VDD.n1615 VDD.n1402 212.329
R13399 VDD.n1622 VDD.n1402 212.329
R13400 VDD.n1398 VDD.n1397 212.329
R13401 VDD.n1397 VDD.n1392 212.329
R13402 VDD.n1625 VDD.n1391 212.329
R13403 VDD.n1632 VDD.n1391 212.329
R13404 VDD.n1637 VDD.n1384 212.329
R13405 VDD.n1384 VDD.n1382 212.329
R13406 VDD.n1257 VDD.n1256 212.329
R13407 VDD.n1256 VDD.n1249 212.329
R13408 VDD.n1258 VDD.n1248 212.329
R13409 VDD.n1265 VDD.n1248 212.329
R13410 VDD.n1244 VDD.n1243 212.329
R13411 VDD.n1243 VDD.n1239 212.329
R13412 VDD.n1268 VDD.n1238 212.329
R13413 VDD.n1275 VDD.n1238 212.329
R13414 VDD.n1234 VDD.n1233 212.329
R13415 VDD.n1233 VDD.n1228 212.329
R13416 VDD.n1278 VDD.n1227 212.329
R13417 VDD.n1285 VDD.n1227 212.329
R13418 VDD.n1223 VDD.n1222 212.329
R13419 VDD.n1222 VDD.n1215 212.329
R13420 VDD.n1288 VDD.n1214 212.329
R13421 VDD.n1295 VDD.n1214 212.329
R13422 VDD.n1210 VDD.n1209 212.329
R13423 VDD.n1209 VDD.n1203 212.329
R13424 VDD.n1298 VDD.n1202 212.329
R13425 VDD.n1305 VDD.n1202 212.329
R13426 VDD.n1311 VDD.n1310 212.329
R13427 VDD.n1312 VDD.n1311 212.329
R13428 VDD.n1195 VDD.n1194 212.329
R13429 VDD.n1194 VDD.n1187 212.329
R13430 VDD.n1315 VDD.n1186 212.329
R13431 VDD.n1322 VDD.n1186 212.329
R13432 VDD.n1182 VDD.n1181 212.329
R13433 VDD.n1181 VDD.n1177 212.329
R13434 VDD.n1325 VDD.n1176 212.329
R13435 VDD.n1332 VDD.n1176 212.329
R13436 VDD.n1172 VDD.n1171 212.329
R13437 VDD.n1171 VDD.n1166 212.329
R13438 VDD.n1335 VDD.n1165 212.329
R13439 VDD.n1342 VDD.n1165 212.329
R13440 VDD.n1161 VDD.n1160 212.329
R13441 VDD.n1160 VDD.n1153 212.329
R13442 VDD.n1345 VDD.n1152 212.329
R13443 VDD.n1352 VDD.n1152 212.329
R13444 VDD.n1148 VDD.n1147 212.329
R13445 VDD.n1147 VDD.n1143 212.329
R13446 VDD.n1355 VDD.n1142 212.329
R13447 VDD.n1362 VDD.n1142 212.329
R13448 VDD.n1138 VDD.n1137 212.329
R13449 VDD.n1137 VDD.n1132 212.329
R13450 VDD.n1365 VDD.n1131 212.329
R13451 VDD.n1372 VDD.n1131 212.329
R13452 VDD.n1377 VDD.n1124 212.329
R13453 VDD.n1124 VDD.n1122 212.329
R13454 VDD.n997 VDD.n996 212.329
R13455 VDD.n996 VDD.n989 212.329
R13456 VDD.n998 VDD.n988 212.329
R13457 VDD.n1005 VDD.n988 212.329
R13458 VDD.n984 VDD.n983 212.329
R13459 VDD.n983 VDD.n979 212.329
R13460 VDD.n1008 VDD.n978 212.329
R13461 VDD.n1015 VDD.n978 212.329
R13462 VDD.n974 VDD.n973 212.329
R13463 VDD.n973 VDD.n968 212.329
R13464 VDD.n1018 VDD.n967 212.329
R13465 VDD.n1025 VDD.n967 212.329
R13466 VDD.n963 VDD.n962 212.329
R13467 VDD.n962 VDD.n955 212.329
R13468 VDD.n1028 VDD.n954 212.329
R13469 VDD.n1035 VDD.n954 212.329
R13470 VDD.n950 VDD.n949 212.329
R13471 VDD.n949 VDD.n943 212.329
R13472 VDD.n1038 VDD.n942 212.329
R13473 VDD.n1045 VDD.n942 212.329
R13474 VDD.n1051 VDD.n1050 212.329
R13475 VDD.n1052 VDD.n1051 212.329
R13476 VDD.n935 VDD.n934 212.329
R13477 VDD.n934 VDD.n927 212.329
R13478 VDD.n1055 VDD.n926 212.329
R13479 VDD.n1062 VDD.n926 212.329
R13480 VDD.n922 VDD.n921 212.329
R13481 VDD.n921 VDD.n917 212.329
R13482 VDD.n1065 VDD.n916 212.329
R13483 VDD.n1072 VDD.n916 212.329
R13484 VDD.n912 VDD.n911 212.329
R13485 VDD.n911 VDD.n906 212.329
R13486 VDD.n1075 VDD.n905 212.329
R13487 VDD.n1082 VDD.n905 212.329
R13488 VDD.n901 VDD.n900 212.329
R13489 VDD.n900 VDD.n893 212.329
R13490 VDD.n1085 VDD.n892 212.329
R13491 VDD.n1092 VDD.n892 212.329
R13492 VDD.n888 VDD.n887 212.329
R13493 VDD.n887 VDD.n883 212.329
R13494 VDD.n1095 VDD.n882 212.329
R13495 VDD.n1102 VDD.n882 212.329
R13496 VDD.n878 VDD.n877 212.329
R13497 VDD.n877 VDD.n872 212.329
R13498 VDD.n1105 VDD.n871 212.329
R13499 VDD.n1112 VDD.n871 212.329
R13500 VDD.n1117 VDD.n864 212.329
R13501 VDD.n864 VDD.n862 212.329
R13502 VDD.n737 VDD.n736 212.329
R13503 VDD.n736 VDD.n729 212.329
R13504 VDD.n738 VDD.n728 212.329
R13505 VDD.n745 VDD.n728 212.329
R13506 VDD.n724 VDD.n723 212.329
R13507 VDD.n723 VDD.n719 212.329
R13508 VDD.n748 VDD.n718 212.329
R13509 VDD.n755 VDD.n718 212.329
R13510 VDD.n714 VDD.n713 212.329
R13511 VDD.n713 VDD.n708 212.329
R13512 VDD.n758 VDD.n707 212.329
R13513 VDD.n765 VDD.n707 212.329
R13514 VDD.n703 VDD.n702 212.329
R13515 VDD.n702 VDD.n695 212.329
R13516 VDD.n768 VDD.n694 212.329
R13517 VDD.n775 VDD.n694 212.329
R13518 VDD.n690 VDD.n689 212.329
R13519 VDD.n689 VDD.n683 212.329
R13520 VDD.n778 VDD.n682 212.329
R13521 VDD.n785 VDD.n682 212.329
R13522 VDD.n791 VDD.n790 212.329
R13523 VDD.n792 VDD.n791 212.329
R13524 VDD.n675 VDD.n674 212.329
R13525 VDD.n674 VDD.n667 212.329
R13526 VDD.n795 VDD.n666 212.329
R13527 VDD.n802 VDD.n666 212.329
R13528 VDD.n662 VDD.n661 212.329
R13529 VDD.n661 VDD.n657 212.329
R13530 VDD.n805 VDD.n656 212.329
R13531 VDD.n812 VDD.n656 212.329
R13532 VDD.n652 VDD.n651 212.329
R13533 VDD.n651 VDD.n646 212.329
R13534 VDD.n815 VDD.n645 212.329
R13535 VDD.n822 VDD.n645 212.329
R13536 VDD.n641 VDD.n640 212.329
R13537 VDD.n640 VDD.n633 212.329
R13538 VDD.n825 VDD.n632 212.329
R13539 VDD.n832 VDD.n632 212.329
R13540 VDD.n628 VDD.n627 212.329
R13541 VDD.n627 VDD.n623 212.329
R13542 VDD.n835 VDD.n622 212.329
R13543 VDD.n842 VDD.n622 212.329
R13544 VDD.n618 VDD.n617 212.329
R13545 VDD.n617 VDD.n612 212.329
R13546 VDD.n845 VDD.n611 212.329
R13547 VDD.n852 VDD.n611 212.329
R13548 VDD.n857 VDD.n604 212.329
R13549 VDD.n604 VDD.n602 212.329
R13550 VDD.n477 VDD.n476 212.329
R13551 VDD.n476 VDD.n469 212.329
R13552 VDD.n478 VDD.n468 212.329
R13553 VDD.n485 VDD.n468 212.329
R13554 VDD.n464 VDD.n463 212.329
R13555 VDD.n463 VDD.n459 212.329
R13556 VDD.n488 VDD.n458 212.329
R13557 VDD.n495 VDD.n458 212.329
R13558 VDD.n454 VDD.n453 212.329
R13559 VDD.n453 VDD.n448 212.329
R13560 VDD.n498 VDD.n447 212.329
R13561 VDD.n505 VDD.n447 212.329
R13562 VDD.n443 VDD.n442 212.329
R13563 VDD.n442 VDD.n435 212.329
R13564 VDD.n508 VDD.n434 212.329
R13565 VDD.n515 VDD.n434 212.329
R13566 VDD.n430 VDD.n429 212.329
R13567 VDD.n429 VDD.n423 212.329
R13568 VDD.n518 VDD.n422 212.329
R13569 VDD.n525 VDD.n422 212.329
R13570 VDD.n531 VDD.n530 212.329
R13571 VDD.n532 VDD.n531 212.329
R13572 VDD.n415 VDD.n414 212.329
R13573 VDD.n414 VDD.n407 212.329
R13574 VDD.n535 VDD.n406 212.329
R13575 VDD.n542 VDD.n406 212.329
R13576 VDD.n402 VDD.n401 212.329
R13577 VDD.n401 VDD.n397 212.329
R13578 VDD.n545 VDD.n396 212.329
R13579 VDD.n552 VDD.n396 212.329
R13580 VDD.n392 VDD.n391 212.329
R13581 VDD.n391 VDD.n386 212.329
R13582 VDD.n555 VDD.n385 212.329
R13583 VDD.n562 VDD.n385 212.329
R13584 VDD.n381 VDD.n380 212.329
R13585 VDD.n380 VDD.n373 212.329
R13586 VDD.n565 VDD.n372 212.329
R13587 VDD.n572 VDD.n372 212.329
R13588 VDD.n368 VDD.n367 212.329
R13589 VDD.n367 VDD.n363 212.329
R13590 VDD.n575 VDD.n362 212.329
R13591 VDD.n582 VDD.n362 212.329
R13592 VDD.n358 VDD.n357 212.329
R13593 VDD.n357 VDD.n352 212.329
R13594 VDD.n585 VDD.n351 212.329
R13595 VDD.n592 VDD.n351 212.329
R13596 VDD.n597 VDD.n344 212.329
R13597 VDD.n344 VDD.n342 212.329
R13598 VDD.n150 VDD.n149 212.329
R13599 VDD.n151 VDD.n150 212.329
R13600 VDD.n156 VDD.n139 212.329
R13601 VDD.n139 VDD.n137 212.329
R13602 VDD.n164 VDD.n163 212.329
R13603 VDD.n165 VDD.n164 212.329
R13604 VDD.n171 VDD.n170 212.329
R13605 VDD.n172 VDD.n171 212.329
R13606 VDD.n177 VDD.n123 212.329
R13607 VDD.n123 VDD.n121 212.329
R13608 VDD.n185 VDD.n184 212.329
R13609 VDD.n186 VDD.n185 212.329
R13610 VDD.n191 VDD.n114 212.329
R13611 VDD.n114 VDD.n112 212.329
R13612 VDD.n199 VDD.n198 212.329
R13613 VDD.n200 VDD.n199 212.329
R13614 VDD.n206 VDD.n205 212.329
R13615 VDD.n207 VDD.n206 212.329
R13616 VDD.n212 VDD.n98 212.329
R13617 VDD.n98 VDD.n96 212.329
R13618 VDD.n220 VDD.n219 212.329
R13619 VDD.n221 VDD.n220 212.329
R13620 VDD.n226 VDD.n89 212.329
R13621 VDD.n89 VDD.n87 212.329
R13622 VDD.n234 VDD.n233 212.329
R13623 VDD.n235 VDD.n234 212.329
R13624 VDD.n241 VDD.n240 212.329
R13625 VDD.n242 VDD.n241 212.329
R13626 VDD.n247 VDD.n73 212.329
R13627 VDD.n73 VDD.n71 212.329
R13628 VDD.n255 VDD.n254 212.329
R13629 VDD.n256 VDD.n255 212.329
R13630 VDD.n261 VDD.n64 212.329
R13631 VDD.n64 VDD.n62 212.329
R13632 VDD.n269 VDD.n268 212.329
R13633 VDD.n270 VDD.n269 212.329
R13634 VDD.n276 VDD.n275 212.329
R13635 VDD.n277 VDD.n276 212.329
R13636 VDD.n282 VDD.n48 212.329
R13637 VDD.n48 VDD.n46 212.329
R13638 VDD.n7393 VDD.n7392 212.329
R13639 VDD.n7392 VDD.n7385 212.329
R13640 VDD.n7394 VDD.n7384 212.329
R13641 VDD.n7401 VDD.n7384 212.329
R13642 VDD.n7380 VDD.n7379 212.329
R13643 VDD.n7379 VDD.n7375 212.329
R13644 VDD.n7404 VDD.n7374 212.329
R13645 VDD.n7411 VDD.n7374 212.329
R13646 VDD.n7370 VDD.n7369 212.329
R13647 VDD.n7369 VDD.n7364 212.329
R13648 VDD.n7414 VDD.n7363 212.329
R13649 VDD.n7421 VDD.n7363 212.329
R13650 VDD.n7359 VDD.n7358 212.329
R13651 VDD.n7358 VDD.n7351 212.329
R13652 VDD.n7424 VDD.n7350 212.329
R13653 VDD.n7431 VDD.n7350 212.329
R13654 VDD.n7346 VDD.n7345 212.329
R13655 VDD.n7345 VDD.n7339 212.329
R13656 VDD.n7434 VDD.n7338 212.329
R13657 VDD.n7441 VDD.n7338 212.329
R13658 VDD.n7447 VDD.n7446 212.329
R13659 VDD.n7448 VDD.n7447 212.329
R13660 VDD.n7331 VDD.n7330 212.329
R13661 VDD.n7330 VDD.n7323 212.329
R13662 VDD.n7451 VDD.n7322 212.329
R13663 VDD.n7458 VDD.n7322 212.329
R13664 VDD.n7318 VDD.n7317 212.329
R13665 VDD.n7317 VDD.n7313 212.329
R13666 VDD.n7461 VDD.n7312 212.329
R13667 VDD.n7468 VDD.n7312 212.329
R13668 VDD.n7308 VDD.n7307 212.329
R13669 VDD.n7307 VDD.n7302 212.329
R13670 VDD.n7471 VDD.n7301 212.329
R13671 VDD.n7478 VDD.n7301 212.329
R13672 VDD.n7297 VDD.n7296 212.329
R13673 VDD.n7296 VDD.n7289 212.329
R13674 VDD.n7481 VDD.n7288 212.329
R13675 VDD.n7488 VDD.n7288 212.329
R13676 VDD.n7284 VDD.n7283 212.329
R13677 VDD.n7283 VDD.n7279 212.329
R13678 VDD.n7491 VDD.n7278 212.329
R13679 VDD.n7498 VDD.n7278 212.329
R13680 VDD.n7274 VDD.n7273 212.329
R13681 VDD.n7273 VDD.n7268 212.329
R13682 VDD.n7501 VDD.n7267 212.329
R13683 VDD.n7508 VDD.n7267 212.329
R13684 VDD.n7513 VDD.n7260 212.329
R13685 VDD.n7260 VDD.n7258 212.329
R13686 VDD.n7253 VDD.n1904 212.329
R13687 VDD.n1904 VDD.n1902 212.329
R13688 VDD.n7136 VDD.n7135 212.329
R13689 VDD.n7135 VDD.n2034 212.329
R13690 VDD.n7137 VDD.n2033 212.329
R13691 VDD.n7144 VDD.n2033 212.329
R13692 VDD.n2029 VDD.n2028 212.329
R13693 VDD.n2028 VDD.n2024 212.329
R13694 VDD.n7147 VDD.n2023 212.329
R13695 VDD.n7154 VDD.n2023 212.329
R13696 VDD.n2019 VDD.n2018 212.329
R13697 VDD.n2018 VDD.n2013 212.329
R13698 VDD.n7157 VDD.n2012 212.329
R13699 VDD.n7164 VDD.n2012 212.329
R13700 VDD.n2008 VDD.n2007 212.329
R13701 VDD.n2007 VDD.n2000 212.329
R13702 VDD.n7167 VDD.n1999 212.329
R13703 VDD.n7174 VDD.n1999 212.329
R13704 VDD.n1995 VDD.n1994 212.329
R13705 VDD.n1994 VDD.n1988 212.329
R13706 VDD.n7177 VDD.n1987 212.329
R13707 VDD.n7184 VDD.n1987 212.329
R13708 VDD.n7190 VDD.n7189 212.329
R13709 VDD.n7191 VDD.n7190 212.329
R13710 VDD.n1979 VDD.n1978 212.329
R13711 VDD.n1979 VDD.n1977 212.329
R13712 VDD.n7199 VDD.n7198 212.329
R13713 VDD.n7199 VDD.n7197 212.329
R13714 VDD.n1971 VDD.n1970 212.329
R13715 VDD.n1970 VDD.n1958 212.329
R13716 VDD.n1953 VDD.n1952 212.329
R13717 VDD.n1952 VDD.n1946 212.329
R13718 VDD.n7211 VDD.n1945 212.329
R13719 VDD.n7218 VDD.n1945 212.329
R13720 VDD.n1941 VDD.n1940 212.329
R13721 VDD.n1940 VDD.n1933 212.329
R13722 VDD.n7221 VDD.n1932 212.329
R13723 VDD.n7228 VDD.n1932 212.329
R13724 VDD.n1928 VDD.n1927 212.329
R13725 VDD.n1927 VDD.n1923 212.329
R13726 VDD.n7231 VDD.n1922 212.329
R13727 VDD.n7238 VDD.n1922 212.329
R13728 VDD.n1918 VDD.n1917 212.329
R13729 VDD.n1917 VDD.n1912 212.329
R13730 VDD.n7241 VDD.n1911 212.329
R13731 VDD.n7248 VDD.n1911 212.329
R13732 VDD.n1973 VDD.n1957 212.329
R13733 VDD.n7208 VDD.n1957 212.329
R13734 VDD.n6999 VDD.n6998 212.329
R13735 VDD.n7000 VDD.n6999 212.329
R13736 VDD.n7005 VDD.n6988 212.329
R13737 VDD.n6988 VDD.n6986 212.329
R13738 VDD.n7013 VDD.n7012 212.329
R13739 VDD.n7014 VDD.n7013 212.329
R13740 VDD.n7020 VDD.n7019 212.329
R13741 VDD.n7021 VDD.n7020 212.329
R13742 VDD.n7026 VDD.n6972 212.329
R13743 VDD.n6972 VDD.n6970 212.329
R13744 VDD.n7034 VDD.n7033 212.329
R13745 VDD.n7035 VDD.n7034 212.329
R13746 VDD.n7040 VDD.n6963 212.329
R13747 VDD.n6963 VDD.n6961 212.329
R13748 VDD.n7048 VDD.n7047 212.329
R13749 VDD.n7049 VDD.n7048 212.329
R13750 VDD.n7055 VDD.n7054 212.329
R13751 VDD.n7056 VDD.n7055 212.329
R13752 VDD.n7061 VDD.n6947 212.329
R13753 VDD.n6947 VDD.n6945 212.329
R13754 VDD.n7069 VDD.n7068 212.329
R13755 VDD.n7070 VDD.n7069 212.329
R13756 VDD.n7075 VDD.n6938 212.329
R13757 VDD.n6938 VDD.n6936 212.329
R13758 VDD.n7083 VDD.n7082 212.329
R13759 VDD.n7084 VDD.n7083 212.329
R13760 VDD.n7090 VDD.n7089 212.329
R13761 VDD.n7091 VDD.n7090 212.329
R13762 VDD.n7096 VDD.n6922 212.329
R13763 VDD.n6922 VDD.n6920 212.329
R13764 VDD.n7104 VDD.n7103 212.329
R13765 VDD.n7105 VDD.n7104 212.329
R13766 VDD.n7110 VDD.n6913 212.329
R13767 VDD.n6913 VDD.n6911 212.329
R13768 VDD.n7118 VDD.n7117 212.329
R13769 VDD.n7119 VDD.n7118 212.329
R13770 VDD.n7123 VDD.n6892 212.329
R13771 VDD.n7123 VDD.n6891 212.329
R13772 VDD.n6903 VDD.n6902 212.329
R13773 VDD.n6902 VDD.n6901 212.329
R13774 VDD.n6024 VDD.n6021 212.329
R13775 VDD.n6029 VDD.n6021 212.329
R13776 VDD.n6018 VDD.n6017 212.329
R13777 VDD.n6017 VDD.n6013 212.329
R13778 VDD.n6032 VDD.n6012 212.329
R13779 VDD.n6039 VDD.n6012 212.329
R13780 VDD.n6008 VDD.n6007 212.329
R13781 VDD.n6007 VDD.n6000 212.329
R13782 VDD.n6042 VDD.n5999 212.329
R13783 VDD.n6049 VDD.n5999 212.329
R13784 VDD.n5995 VDD.n5994 212.329
R13785 VDD.n5994 VDD.n5989 212.329
R13786 VDD.n6052 VDD.n5988 212.329
R13787 VDD.n6059 VDD.n5988 212.329
R13788 VDD.n5984 VDD.n5983 212.329
R13789 VDD.n5983 VDD.n5979 212.329
R13790 VDD.n6062 VDD.n5978 212.329
R13791 VDD.n6069 VDD.n5978 212.329
R13792 VDD.n5974 VDD.n5973 212.329
R13793 VDD.n5973 VDD.n5966 212.329
R13794 VDD.n6072 VDD.n5965 212.329
R13795 VDD.n6079 VDD.n5965 212.329
R13796 VDD.n5961 VDD.n5960 212.329
R13797 VDD.n5960 VDD.n5954 212.329
R13798 VDD.n6082 VDD.n5953 212.329
R13799 VDD.n6089 VDD.n5953 212.329
R13800 VDD.n6095 VDD.n6094 212.329
R13801 VDD.n6096 VDD.n6095 212.329
R13802 VDD.n5946 VDD.n5945 212.329
R13803 VDD.n5945 VDD.n5938 212.329
R13804 VDD.n6099 VDD.n5937 212.329
R13805 VDD.n6106 VDD.n5937 212.329
R13806 VDD.n5933 VDD.n5932 212.329
R13807 VDD.n5932 VDD.n5927 212.329
R13808 VDD.n6109 VDD.n5926 212.329
R13809 VDD.n6116 VDD.n5926 212.329
R13810 VDD.n5922 VDD.n5921 212.329
R13811 VDD.n5921 VDD.n5917 212.329
R13812 VDD.n6119 VDD.n5916 212.329
R13813 VDD.n6126 VDD.n5916 212.329
R13814 VDD.n5912 VDD.n5911 212.329
R13815 VDD.n5911 VDD.n5907 212.329
R13816 VDD.n6129 VDD.n5906 212.329
R13817 VDD.n6136 VDD.n5906 212.329
R13818 VDD.n5901 VDD.n5900 212.329
R13819 VDD.n5901 VDD.n5899 212.329
R13820 VDD.n6144 VDD.n6143 212.329
R13821 VDD.n6144 VDD.n6142 212.329
R13822 VDD.n5888 VDD.n5885 212.329
R13823 VDD.n6152 VDD.n5885 212.329
R13824 VDD.n5882 VDD.n5881 212.329
R13825 VDD.n5881 VDD.n5877 212.329
R13826 VDD.n6155 VDD.n5876 212.329
R13827 VDD.n6162 VDD.n5876 212.329
R13828 VDD.n5872 VDD.n5871 212.329
R13829 VDD.n5871 VDD.n5864 212.329
R13830 VDD.n6165 VDD.n5863 212.329
R13831 VDD.n6172 VDD.n5863 212.329
R13832 VDD.n5859 VDD.n5858 212.329
R13833 VDD.n5858 VDD.n5853 212.329
R13834 VDD.n6175 VDD.n5852 212.329
R13835 VDD.n6182 VDD.n5852 212.329
R13836 VDD.n5848 VDD.n5847 212.329
R13837 VDD.n5847 VDD.n5843 212.329
R13838 VDD.n6185 VDD.n5842 212.329
R13839 VDD.n6192 VDD.n5842 212.329
R13840 VDD.n5838 VDD.n5837 212.329
R13841 VDD.n5837 VDD.n5830 212.329
R13842 VDD.n6195 VDD.n5829 212.329
R13843 VDD.n6202 VDD.n5829 212.329
R13844 VDD.n5825 VDD.n5824 212.329
R13845 VDD.n5824 VDD.n5818 212.329
R13846 VDD.n6205 VDD.n5817 212.329
R13847 VDD.n6212 VDD.n5817 212.329
R13848 VDD.n6218 VDD.n6217 212.329
R13849 VDD.n6219 VDD.n6218 212.329
R13850 VDD.n5810 VDD.n5809 212.329
R13851 VDD.n5809 VDD.n5802 212.329
R13852 VDD.n6222 VDD.n5801 212.329
R13853 VDD.n6229 VDD.n5801 212.329
R13854 VDD.n5797 VDD.n5796 212.329
R13855 VDD.n5796 VDD.n5791 212.329
R13856 VDD.n6232 VDD.n5790 212.329
R13857 VDD.n6239 VDD.n5790 212.329
R13858 VDD.n5786 VDD.n5785 212.329
R13859 VDD.n5785 VDD.n5781 212.329
R13860 VDD.n6242 VDD.n5780 212.329
R13861 VDD.n6249 VDD.n5780 212.329
R13862 VDD.n5776 VDD.n5775 212.329
R13863 VDD.n5775 VDD.n5771 212.329
R13864 VDD.n6252 VDD.n5770 212.329
R13865 VDD.n6259 VDD.n5770 212.329
R13866 VDD.n5765 VDD.n5764 212.329
R13867 VDD.n5765 VDD.n5763 212.329
R13868 VDD.n6267 VDD.n6266 212.329
R13869 VDD.n6267 VDD.n6265 212.329
R13870 VDD.n5752 VDD.n5749 212.329
R13871 VDD.n6275 VDD.n5749 212.329
R13872 VDD.n5746 VDD.n5745 212.329
R13873 VDD.n5745 VDD.n5741 212.329
R13874 VDD.n6278 VDD.n5740 212.329
R13875 VDD.n6285 VDD.n5740 212.329
R13876 VDD.n5736 VDD.n5735 212.329
R13877 VDD.n5735 VDD.n5728 212.329
R13878 VDD.n6288 VDD.n5727 212.329
R13879 VDD.n6295 VDD.n5727 212.329
R13880 VDD.n5723 VDD.n5722 212.329
R13881 VDD.n5722 VDD.n5717 212.329
R13882 VDD.n6298 VDD.n5716 212.329
R13883 VDD.n6305 VDD.n5716 212.329
R13884 VDD.n5712 VDD.n5711 212.329
R13885 VDD.n5711 VDD.n5707 212.329
R13886 VDD.n6308 VDD.n5706 212.329
R13887 VDD.n6315 VDD.n5706 212.329
R13888 VDD.n5702 VDD.n5701 212.329
R13889 VDD.n5701 VDD.n5694 212.329
R13890 VDD.n6318 VDD.n5693 212.329
R13891 VDD.n6325 VDD.n5693 212.329
R13892 VDD.n5689 VDD.n5688 212.329
R13893 VDD.n5688 VDD.n5682 212.329
R13894 VDD.n6328 VDD.n5681 212.329
R13895 VDD.n6335 VDD.n5681 212.329
R13896 VDD.n6341 VDD.n6340 212.329
R13897 VDD.n6342 VDD.n6341 212.329
R13898 VDD.n5674 VDD.n5673 212.329
R13899 VDD.n5673 VDD.n5666 212.329
R13900 VDD.n6345 VDD.n5665 212.329
R13901 VDD.n6352 VDD.n5665 212.329
R13902 VDD.n5661 VDD.n5660 212.329
R13903 VDD.n5660 VDD.n5655 212.329
R13904 VDD.n6355 VDD.n5654 212.329
R13905 VDD.n6362 VDD.n5654 212.329
R13906 VDD.n5650 VDD.n5649 212.329
R13907 VDD.n5649 VDD.n5645 212.329
R13908 VDD.n6365 VDD.n5644 212.329
R13909 VDD.n6372 VDD.n5644 212.329
R13910 VDD.n5640 VDD.n5639 212.329
R13911 VDD.n5639 VDD.n5635 212.329
R13912 VDD.n6375 VDD.n5634 212.329
R13913 VDD.n6382 VDD.n5634 212.329
R13914 VDD.n5629 VDD.n5628 212.329
R13915 VDD.n5629 VDD.n5627 212.329
R13916 VDD.n6390 VDD.n6389 212.329
R13917 VDD.n6390 VDD.n6388 212.329
R13918 VDD.n5616 VDD.n5613 212.329
R13919 VDD.n6398 VDD.n5613 212.329
R13920 VDD.n5610 VDD.n5609 212.329
R13921 VDD.n5609 VDD.n5605 212.329
R13922 VDD.n6401 VDD.n5604 212.329
R13923 VDD.n6408 VDD.n5604 212.329
R13924 VDD.n5600 VDD.n5599 212.329
R13925 VDD.n5599 VDD.n5592 212.329
R13926 VDD.n6411 VDD.n5591 212.329
R13927 VDD.n6418 VDD.n5591 212.329
R13928 VDD.n5587 VDD.n5586 212.329
R13929 VDD.n5586 VDD.n5581 212.329
R13930 VDD.n6421 VDD.n5580 212.329
R13931 VDD.n6428 VDD.n5580 212.329
R13932 VDD.n5576 VDD.n5575 212.329
R13933 VDD.n5575 VDD.n5571 212.329
R13934 VDD.n6431 VDD.n5570 212.329
R13935 VDD.n6438 VDD.n5570 212.329
R13936 VDD.n5566 VDD.n5565 212.329
R13937 VDD.n5565 VDD.n5558 212.329
R13938 VDD.n6441 VDD.n5557 212.329
R13939 VDD.n6448 VDD.n5557 212.329
R13940 VDD.n5553 VDD.n5552 212.329
R13941 VDD.n5552 VDD.n5546 212.329
R13942 VDD.n6451 VDD.n5545 212.329
R13943 VDD.n6458 VDD.n5545 212.329
R13944 VDD.n6464 VDD.n6463 212.329
R13945 VDD.n6465 VDD.n6464 212.329
R13946 VDD.n5538 VDD.n5537 212.329
R13947 VDD.n5537 VDD.n5530 212.329
R13948 VDD.n6468 VDD.n5529 212.329
R13949 VDD.n6475 VDD.n5529 212.329
R13950 VDD.n5525 VDD.n5524 212.329
R13951 VDD.n5524 VDD.n5519 212.329
R13952 VDD.n6478 VDD.n5518 212.329
R13953 VDD.n6485 VDD.n5518 212.329
R13954 VDD.n5514 VDD.n5513 212.329
R13955 VDD.n5513 VDD.n5509 212.329
R13956 VDD.n6488 VDD.n5508 212.329
R13957 VDD.n6495 VDD.n5508 212.329
R13958 VDD.n5504 VDD.n5503 212.329
R13959 VDD.n5503 VDD.n5499 212.329
R13960 VDD.n6498 VDD.n5498 212.329
R13961 VDD.n6505 VDD.n5498 212.329
R13962 VDD.n5493 VDD.n5492 212.329
R13963 VDD.n5493 VDD.n5491 212.329
R13964 VDD.n6513 VDD.n6512 212.329
R13965 VDD.n6513 VDD.n6511 212.329
R13966 VDD.n5480 VDD.n5477 212.329
R13967 VDD.n6521 VDD.n5477 212.329
R13968 VDD.n5474 VDD.n5473 212.329
R13969 VDD.n5473 VDD.n5469 212.329
R13970 VDD.n6524 VDD.n5468 212.329
R13971 VDD.n6531 VDD.n5468 212.329
R13972 VDD.n5464 VDD.n5463 212.329
R13973 VDD.n5463 VDD.n5456 212.329
R13974 VDD.n6534 VDD.n5455 212.329
R13975 VDD.n6541 VDD.n5455 212.329
R13976 VDD.n5451 VDD.n5450 212.329
R13977 VDD.n5450 VDD.n5445 212.329
R13978 VDD.n6544 VDD.n5444 212.329
R13979 VDD.n6551 VDD.n5444 212.329
R13980 VDD.n5440 VDD.n5439 212.329
R13981 VDD.n5439 VDD.n5435 212.329
R13982 VDD.n6554 VDD.n5434 212.329
R13983 VDD.n6561 VDD.n5434 212.329
R13984 VDD.n5430 VDD.n5429 212.329
R13985 VDD.n5429 VDD.n5422 212.329
R13986 VDD.n6564 VDD.n5421 212.329
R13987 VDD.n6571 VDD.n5421 212.329
R13988 VDD.n5417 VDD.n5416 212.329
R13989 VDD.n5416 VDD.n5410 212.329
R13990 VDD.n6574 VDD.n5409 212.329
R13991 VDD.n6581 VDD.n5409 212.329
R13992 VDD.n6587 VDD.n6586 212.329
R13993 VDD.n6588 VDD.n6587 212.329
R13994 VDD.n5402 VDD.n5401 212.329
R13995 VDD.n5401 VDD.n5394 212.329
R13996 VDD.n6591 VDD.n5393 212.329
R13997 VDD.n6598 VDD.n5393 212.329
R13998 VDD.n5389 VDD.n5388 212.329
R13999 VDD.n5388 VDD.n5383 212.329
R14000 VDD.n6601 VDD.n5382 212.329
R14001 VDD.n6608 VDD.n5382 212.329
R14002 VDD.n5378 VDD.n5377 212.329
R14003 VDD.n5377 VDD.n5373 212.329
R14004 VDD.n6611 VDD.n5372 212.329
R14005 VDD.n6618 VDD.n5372 212.329
R14006 VDD.n5368 VDD.n5367 212.329
R14007 VDD.n5367 VDD.n5363 212.329
R14008 VDD.n6621 VDD.n5362 212.329
R14009 VDD.n6628 VDD.n5362 212.329
R14010 VDD.n5357 VDD.n5356 212.329
R14011 VDD.n5357 VDD.n5355 212.329
R14012 VDD.n6636 VDD.n6635 212.329
R14013 VDD.n6636 VDD.n6634 212.329
R14014 VDD.n5344 VDD.n5341 212.329
R14015 VDD.n6644 VDD.n5341 212.329
R14016 VDD.n5338 VDD.n5337 212.329
R14017 VDD.n5337 VDD.n5333 212.329
R14018 VDD.n6647 VDD.n5332 212.329
R14019 VDD.n6654 VDD.n5332 212.329
R14020 VDD.n5328 VDD.n5327 212.329
R14021 VDD.n5327 VDD.n5320 212.329
R14022 VDD.n6657 VDD.n5319 212.329
R14023 VDD.n6664 VDD.n5319 212.329
R14024 VDD.n5315 VDD.n5314 212.329
R14025 VDD.n5314 VDD.n5309 212.329
R14026 VDD.n6667 VDD.n5308 212.329
R14027 VDD.n6674 VDD.n5308 212.329
R14028 VDD.n5304 VDD.n5303 212.329
R14029 VDD.n5303 VDD.n5299 212.329
R14030 VDD.n6677 VDD.n5298 212.329
R14031 VDD.n6684 VDD.n5298 212.329
R14032 VDD.n5294 VDD.n5293 212.329
R14033 VDD.n5293 VDD.n5286 212.329
R14034 VDD.n6687 VDD.n5285 212.329
R14035 VDD.n6694 VDD.n5285 212.329
R14036 VDD.n5281 VDD.n5280 212.329
R14037 VDD.n5280 VDD.n5274 212.329
R14038 VDD.n6697 VDD.n5273 212.329
R14039 VDD.n6704 VDD.n5273 212.329
R14040 VDD.n6710 VDD.n6709 212.329
R14041 VDD.n6711 VDD.n6710 212.329
R14042 VDD.n5266 VDD.n5265 212.329
R14043 VDD.n5265 VDD.n5258 212.329
R14044 VDD.n6714 VDD.n5257 212.329
R14045 VDD.n6721 VDD.n5257 212.329
R14046 VDD.n5253 VDD.n5252 212.329
R14047 VDD.n5252 VDD.n5247 212.329
R14048 VDD.n6724 VDD.n5246 212.329
R14049 VDD.n6731 VDD.n5246 212.329
R14050 VDD.n5242 VDD.n5241 212.329
R14051 VDD.n5241 VDD.n5237 212.329
R14052 VDD.n6734 VDD.n5236 212.329
R14053 VDD.n6741 VDD.n5236 212.329
R14054 VDD.n5232 VDD.n5231 212.329
R14055 VDD.n5231 VDD.n5227 212.329
R14056 VDD.n6744 VDD.n5226 212.329
R14057 VDD.n6751 VDD.n5226 212.329
R14058 VDD.n5221 VDD.n5220 212.329
R14059 VDD.n5221 VDD.n5219 212.329
R14060 VDD.n6759 VDD.n6758 212.329
R14061 VDD.n6759 VDD.n6757 212.329
R14062 VDD.n5208 VDD.n5205 212.329
R14063 VDD.n6767 VDD.n5205 212.329
R14064 VDD.n5202 VDD.n5201 212.329
R14065 VDD.n5201 VDD.n5197 212.329
R14066 VDD.n6770 VDD.n5196 212.329
R14067 VDD.n6777 VDD.n5196 212.329
R14068 VDD.n5192 VDD.n5191 212.329
R14069 VDD.n5191 VDD.n5184 212.329
R14070 VDD.n6780 VDD.n5183 212.329
R14071 VDD.n6787 VDD.n5183 212.329
R14072 VDD.n5179 VDD.n5178 212.329
R14073 VDD.n5178 VDD.n5173 212.329
R14074 VDD.n6790 VDD.n5172 212.329
R14075 VDD.n6797 VDD.n5172 212.329
R14076 VDD.n5168 VDD.n5167 212.329
R14077 VDD.n5167 VDD.n5163 212.329
R14078 VDD.n6800 VDD.n5162 212.329
R14079 VDD.n6807 VDD.n5162 212.329
R14080 VDD.n5158 VDD.n5157 212.329
R14081 VDD.n5157 VDD.n5150 212.329
R14082 VDD.n6810 VDD.n5149 212.329
R14083 VDD.n6817 VDD.n5149 212.329
R14084 VDD.n5145 VDD.n5144 212.329
R14085 VDD.n5144 VDD.n5138 212.329
R14086 VDD.n6820 VDD.n5137 212.329
R14087 VDD.n6827 VDD.n5137 212.329
R14088 VDD.n6833 VDD.n6832 212.329
R14089 VDD.n6834 VDD.n6833 212.329
R14090 VDD.n5130 VDD.n5129 212.329
R14091 VDD.n5129 VDD.n5122 212.329
R14092 VDD.n6837 VDD.n5121 212.329
R14093 VDD.n6844 VDD.n5121 212.329
R14094 VDD.n5117 VDD.n5116 212.329
R14095 VDD.n5116 VDD.n5111 212.329
R14096 VDD.n6847 VDD.n5110 212.329
R14097 VDD.n6854 VDD.n5110 212.329
R14098 VDD.n5106 VDD.n5105 212.329
R14099 VDD.n5105 VDD.n5101 212.329
R14100 VDD.n6857 VDD.n5100 212.329
R14101 VDD.n6864 VDD.n5100 212.329
R14102 VDD.n5096 VDD.n5095 212.329
R14103 VDD.n5095 VDD.n5091 212.329
R14104 VDD.n6867 VDD.n5090 212.329
R14105 VDD.n6874 VDD.n5090 212.329
R14106 VDD.n5085 VDD.n5084 212.329
R14107 VDD.n5085 VDD.n5083 212.329
R14108 VDD.n6882 VDD.n6881 212.329
R14109 VDD.n6882 VDD.n6880 212.329
R14110 VDD.n5070 VDD.n4818 212.329
R14111 VDD.n4818 VDD.n4816 212.329
R14112 VDD.n4829 VDD.n4824 212.329
R14113 VDD.n4830 VDD.n4829 212.329
R14114 VDD.n5063 VDD.n4823 212.329
R14115 VDD.n5056 VDD.n4823 212.329
R14116 VDD.n4839 VDD.n4835 212.329
R14117 VDD.n4840 VDD.n4839 212.329
R14118 VDD.n5053 VDD.n4834 212.329
R14119 VDD.n5046 VDD.n4834 212.329
R14120 VDD.n4852 VDD.n4845 212.329
R14121 VDD.n4853 VDD.n4852 212.329
R14122 VDD.n5043 VDD.n4844 212.329
R14123 VDD.n5036 VDD.n4844 212.329
R14124 VDD.n4863 VDD.n4858 212.329
R14125 VDD.n4864 VDD.n4863 212.329
R14126 VDD.n5033 VDD.n4857 212.329
R14127 VDD.n5026 VDD.n4857 212.329
R14128 VDD.n4873 VDD.n4869 212.329
R14129 VDD.n4874 VDD.n4873 212.329
R14130 VDD.n5023 VDD.n4868 212.329
R14131 VDD.n5016 VDD.n4868 212.329
R14132 VDD.n4886 VDD.n4879 212.329
R14133 VDD.n4887 VDD.n4886 212.329
R14134 VDD.n5013 VDD.n4878 212.329
R14135 VDD.n5006 VDD.n4878 212.329
R14136 VDD.n5003 VDD.n5002 212.329
R14137 VDD.n5002 VDD.n5001 212.329
R14138 VDD.n4901 VDD.n4895 212.329
R14139 VDD.n4902 VDD.n4901 212.329
R14140 VDD.n4996 VDD.n4894 212.329
R14141 VDD.n4989 VDD.n4894 212.329
R14142 VDD.n4914 VDD.n4907 212.329
R14143 VDD.n4915 VDD.n4914 212.329
R14144 VDD.n4986 VDD.n4906 212.329
R14145 VDD.n4979 VDD.n4906 212.329
R14146 VDD.n4925 VDD.n4920 212.329
R14147 VDD.n4926 VDD.n4925 212.329
R14148 VDD.n4976 VDD.n4919 212.329
R14149 VDD.n4969 VDD.n4919 212.329
R14150 VDD.n4935 VDD.n4931 212.329
R14151 VDD.n4936 VDD.n4935 212.329
R14152 VDD.n4966 VDD.n4930 212.329
R14153 VDD.n4959 VDD.n4930 212.329
R14154 VDD.n4944 VDD.n4941 212.329
R14155 VDD.n4945 VDD.n4944 212.329
R14156 VDD.n4956 VDD.n4940 212.329
R14157 VDD.n4946 VDD.n4940 212.329
R14158 VDD.n4812 VDD.n2040 212.329
R14159 VDD.n2040 VDD.n2038 212.329
R14160 VDD.n4695 VDD.n4694 212.329
R14161 VDD.n4694 VDD.n2170 212.329
R14162 VDD.n4696 VDD.n2169 212.329
R14163 VDD.n4703 VDD.n2169 212.329
R14164 VDD.n2165 VDD.n2164 212.329
R14165 VDD.n2164 VDD.n2160 212.329
R14166 VDD.n4706 VDD.n2159 212.329
R14167 VDD.n4713 VDD.n2159 212.329
R14168 VDD.n2155 VDD.n2154 212.329
R14169 VDD.n2154 VDD.n2149 212.329
R14170 VDD.n4716 VDD.n2148 212.329
R14171 VDD.n4723 VDD.n2148 212.329
R14172 VDD.n2144 VDD.n2143 212.329
R14173 VDD.n2143 VDD.n2136 212.329
R14174 VDD.n4726 VDD.n2135 212.329
R14175 VDD.n4733 VDD.n2135 212.329
R14176 VDD.n2131 VDD.n2130 212.329
R14177 VDD.n2130 VDD.n2124 212.329
R14178 VDD.n4736 VDD.n2123 212.329
R14179 VDD.n4743 VDD.n2123 212.329
R14180 VDD.n4749 VDD.n4748 212.329
R14181 VDD.n4750 VDD.n4749 212.329
R14182 VDD.n2115 VDD.n2114 212.329
R14183 VDD.n2115 VDD.n2113 212.329
R14184 VDD.n4758 VDD.n4757 212.329
R14185 VDD.n4758 VDD.n4756 212.329
R14186 VDD.n2107 VDD.n2106 212.329
R14187 VDD.n2106 VDD.n2094 212.329
R14188 VDD.n2089 VDD.n2088 212.329
R14189 VDD.n2088 VDD.n2082 212.329
R14190 VDD.n4770 VDD.n2081 212.329
R14191 VDD.n4777 VDD.n2081 212.329
R14192 VDD.n2077 VDD.n2076 212.329
R14193 VDD.n2076 VDD.n2069 212.329
R14194 VDD.n4780 VDD.n2068 212.329
R14195 VDD.n4787 VDD.n2068 212.329
R14196 VDD.n2064 VDD.n2063 212.329
R14197 VDD.n2063 VDD.n2059 212.329
R14198 VDD.n4790 VDD.n2058 212.329
R14199 VDD.n4797 VDD.n2058 212.329
R14200 VDD.n2054 VDD.n2053 212.329
R14201 VDD.n2053 VDD.n2048 212.329
R14202 VDD.n4800 VDD.n2047 212.329
R14203 VDD.n4807 VDD.n2047 212.329
R14204 VDD.n2109 VDD.n2093 212.329
R14205 VDD.n4767 VDD.n2093 212.329
R14206 VDD.n4687 VDD.n2176 212.329
R14207 VDD.n2176 VDD.n2174 212.329
R14208 VDD.n4570 VDD.n4569 212.329
R14209 VDD.n4569 VDD.n2306 212.329
R14210 VDD.n4571 VDD.n2305 212.329
R14211 VDD.n4578 VDD.n2305 212.329
R14212 VDD.n2301 VDD.n2300 212.329
R14213 VDD.n2300 VDD.n2296 212.329
R14214 VDD.n4581 VDD.n2295 212.329
R14215 VDD.n4588 VDD.n2295 212.329
R14216 VDD.n2291 VDD.n2290 212.329
R14217 VDD.n2290 VDD.n2285 212.329
R14218 VDD.n4591 VDD.n2284 212.329
R14219 VDD.n4598 VDD.n2284 212.329
R14220 VDD.n2280 VDD.n2279 212.329
R14221 VDD.n2279 VDD.n2272 212.329
R14222 VDD.n4601 VDD.n2271 212.329
R14223 VDD.n4608 VDD.n2271 212.329
R14224 VDD.n2267 VDD.n2266 212.329
R14225 VDD.n2266 VDD.n2260 212.329
R14226 VDD.n4611 VDD.n2259 212.329
R14227 VDD.n4618 VDD.n2259 212.329
R14228 VDD.n4624 VDD.n4623 212.329
R14229 VDD.n4625 VDD.n4624 212.329
R14230 VDD.n2251 VDD.n2250 212.329
R14231 VDD.n2251 VDD.n2249 212.329
R14232 VDD.n4633 VDD.n4632 212.329
R14233 VDD.n4633 VDD.n4631 212.329
R14234 VDD.n2243 VDD.n2242 212.329
R14235 VDD.n2242 VDD.n2230 212.329
R14236 VDD.n2225 VDD.n2224 212.329
R14237 VDD.n2224 VDD.n2218 212.329
R14238 VDD.n4645 VDD.n2217 212.329
R14239 VDD.n4652 VDD.n2217 212.329
R14240 VDD.n2213 VDD.n2212 212.329
R14241 VDD.n2212 VDD.n2205 212.329
R14242 VDD.n4655 VDD.n2204 212.329
R14243 VDD.n4662 VDD.n2204 212.329
R14244 VDD.n2200 VDD.n2199 212.329
R14245 VDD.n2199 VDD.n2195 212.329
R14246 VDD.n4665 VDD.n2194 212.329
R14247 VDD.n4672 VDD.n2194 212.329
R14248 VDD.n2190 VDD.n2189 212.329
R14249 VDD.n2189 VDD.n2184 212.329
R14250 VDD.n4675 VDD.n2183 212.329
R14251 VDD.n4682 VDD.n2183 212.329
R14252 VDD.n2245 VDD.n2229 212.329
R14253 VDD.n4642 VDD.n2229 212.329
R14254 VDD.n4562 VDD.n2312 212.329
R14255 VDD.n2312 VDD.n2310 212.329
R14256 VDD.n4445 VDD.n4444 212.329
R14257 VDD.n4444 VDD.n2442 212.329
R14258 VDD.n4446 VDD.n2441 212.329
R14259 VDD.n4453 VDD.n2441 212.329
R14260 VDD.n2437 VDD.n2436 212.329
R14261 VDD.n2436 VDD.n2432 212.329
R14262 VDD.n4456 VDD.n2431 212.329
R14263 VDD.n4463 VDD.n2431 212.329
R14264 VDD.n2427 VDD.n2426 212.329
R14265 VDD.n2426 VDD.n2421 212.329
R14266 VDD.n4466 VDD.n2420 212.329
R14267 VDD.n4473 VDD.n2420 212.329
R14268 VDD.n2416 VDD.n2415 212.329
R14269 VDD.n2415 VDD.n2408 212.329
R14270 VDD.n4476 VDD.n2407 212.329
R14271 VDD.n4483 VDD.n2407 212.329
R14272 VDD.n2403 VDD.n2402 212.329
R14273 VDD.n2402 VDD.n2396 212.329
R14274 VDD.n4486 VDD.n2395 212.329
R14275 VDD.n4493 VDD.n2395 212.329
R14276 VDD.n4499 VDD.n4498 212.329
R14277 VDD.n4500 VDD.n4499 212.329
R14278 VDD.n2387 VDD.n2386 212.329
R14279 VDD.n2387 VDD.n2385 212.329
R14280 VDD.n4508 VDD.n4507 212.329
R14281 VDD.n4508 VDD.n4506 212.329
R14282 VDD.n2379 VDD.n2378 212.329
R14283 VDD.n2378 VDD.n2366 212.329
R14284 VDD.n2361 VDD.n2360 212.329
R14285 VDD.n2360 VDD.n2354 212.329
R14286 VDD.n4520 VDD.n2353 212.329
R14287 VDD.n4527 VDD.n2353 212.329
R14288 VDD.n2349 VDD.n2348 212.329
R14289 VDD.n2348 VDD.n2341 212.329
R14290 VDD.n4530 VDD.n2340 212.329
R14291 VDD.n4537 VDD.n2340 212.329
R14292 VDD.n2336 VDD.n2335 212.329
R14293 VDD.n2335 VDD.n2331 212.329
R14294 VDD.n4540 VDD.n2330 212.329
R14295 VDD.n4547 VDD.n2330 212.329
R14296 VDD.n2326 VDD.n2325 212.329
R14297 VDD.n2325 VDD.n2320 212.329
R14298 VDD.n4550 VDD.n2319 212.329
R14299 VDD.n4557 VDD.n2319 212.329
R14300 VDD.n2381 VDD.n2365 212.329
R14301 VDD.n4517 VDD.n2365 212.329
R14302 VDD.n4437 VDD.n2448 212.329
R14303 VDD.n2448 VDD.n2446 212.329
R14304 VDD.n4320 VDD.n4319 212.329
R14305 VDD.n4319 VDD.n2578 212.329
R14306 VDD.n4321 VDD.n2577 212.329
R14307 VDD.n4328 VDD.n2577 212.329
R14308 VDD.n2573 VDD.n2572 212.329
R14309 VDD.n2572 VDD.n2568 212.329
R14310 VDD.n4331 VDD.n2567 212.329
R14311 VDD.n4338 VDD.n2567 212.329
R14312 VDD.n2563 VDD.n2562 212.329
R14313 VDD.n2562 VDD.n2557 212.329
R14314 VDD.n4341 VDD.n2556 212.329
R14315 VDD.n4348 VDD.n2556 212.329
R14316 VDD.n2552 VDD.n2551 212.329
R14317 VDD.n2551 VDD.n2544 212.329
R14318 VDD.n4351 VDD.n2543 212.329
R14319 VDD.n4358 VDD.n2543 212.329
R14320 VDD.n2539 VDD.n2538 212.329
R14321 VDD.n2538 VDD.n2532 212.329
R14322 VDD.n4361 VDD.n2531 212.329
R14323 VDD.n4368 VDD.n2531 212.329
R14324 VDD.n4374 VDD.n4373 212.329
R14325 VDD.n4375 VDD.n4374 212.329
R14326 VDD.n2523 VDD.n2522 212.329
R14327 VDD.n2523 VDD.n2521 212.329
R14328 VDD.n4383 VDD.n4382 212.329
R14329 VDD.n4383 VDD.n4381 212.329
R14330 VDD.n2515 VDD.n2514 212.329
R14331 VDD.n2514 VDD.n2502 212.329
R14332 VDD.n2497 VDD.n2496 212.329
R14333 VDD.n2496 VDD.n2490 212.329
R14334 VDD.n4395 VDD.n2489 212.329
R14335 VDD.n4402 VDD.n2489 212.329
R14336 VDD.n2485 VDD.n2484 212.329
R14337 VDD.n2484 VDD.n2477 212.329
R14338 VDD.n4405 VDD.n2476 212.329
R14339 VDD.n4412 VDD.n2476 212.329
R14340 VDD.n2472 VDD.n2471 212.329
R14341 VDD.n2471 VDD.n2467 212.329
R14342 VDD.n4415 VDD.n2466 212.329
R14343 VDD.n4422 VDD.n2466 212.329
R14344 VDD.n2462 VDD.n2461 212.329
R14345 VDD.n2461 VDD.n2456 212.329
R14346 VDD.n4425 VDD.n2455 212.329
R14347 VDD.n4432 VDD.n2455 212.329
R14348 VDD.n2517 VDD.n2501 212.329
R14349 VDD.n4392 VDD.n2501 212.329
R14350 VDD.n4312 VDD.n2584 212.329
R14351 VDD.n2584 VDD.n2582 212.329
R14352 VDD.n4195 VDD.n4194 212.329
R14353 VDD.n4194 VDD.n2714 212.329
R14354 VDD.n4196 VDD.n2713 212.329
R14355 VDD.n4203 VDD.n2713 212.329
R14356 VDD.n2709 VDD.n2708 212.329
R14357 VDD.n2708 VDD.n2704 212.329
R14358 VDD.n4206 VDD.n2703 212.329
R14359 VDD.n4213 VDD.n2703 212.329
R14360 VDD.n2699 VDD.n2698 212.329
R14361 VDD.n2698 VDD.n2693 212.329
R14362 VDD.n4216 VDD.n2692 212.329
R14363 VDD.n4223 VDD.n2692 212.329
R14364 VDD.n2688 VDD.n2687 212.329
R14365 VDD.n2687 VDD.n2680 212.329
R14366 VDD.n4226 VDD.n2679 212.329
R14367 VDD.n4233 VDD.n2679 212.329
R14368 VDD.n2675 VDD.n2674 212.329
R14369 VDD.n2674 VDD.n2668 212.329
R14370 VDD.n4236 VDD.n2667 212.329
R14371 VDD.n4243 VDD.n2667 212.329
R14372 VDD.n4249 VDD.n4248 212.329
R14373 VDD.n4250 VDD.n4249 212.329
R14374 VDD.n2659 VDD.n2658 212.329
R14375 VDD.n2659 VDD.n2657 212.329
R14376 VDD.n4258 VDD.n4257 212.329
R14377 VDD.n4258 VDD.n4256 212.329
R14378 VDD.n2651 VDD.n2650 212.329
R14379 VDD.n2650 VDD.n2638 212.329
R14380 VDD.n2633 VDD.n2632 212.329
R14381 VDD.n2632 VDD.n2626 212.329
R14382 VDD.n4270 VDD.n2625 212.329
R14383 VDD.n4277 VDD.n2625 212.329
R14384 VDD.n2621 VDD.n2620 212.329
R14385 VDD.n2620 VDD.n2613 212.329
R14386 VDD.n4280 VDD.n2612 212.329
R14387 VDD.n4287 VDD.n2612 212.329
R14388 VDD.n2608 VDD.n2607 212.329
R14389 VDD.n2607 VDD.n2603 212.329
R14390 VDD.n4290 VDD.n2602 212.329
R14391 VDD.n4297 VDD.n2602 212.329
R14392 VDD.n2598 VDD.n2597 212.329
R14393 VDD.n2597 VDD.n2592 212.329
R14394 VDD.n4300 VDD.n2591 212.329
R14395 VDD.n4307 VDD.n2591 212.329
R14396 VDD.n2653 VDD.n2637 212.329
R14397 VDD.n4267 VDD.n2637 212.329
R14398 VDD.n4187 VDD.n2720 212.329
R14399 VDD.n2720 VDD.n2718 212.329
R14400 VDD.n4070 VDD.n4069 212.329
R14401 VDD.n4069 VDD.n2850 212.329
R14402 VDD.n4071 VDD.n2849 212.329
R14403 VDD.n4078 VDD.n2849 212.329
R14404 VDD.n2845 VDD.n2844 212.329
R14405 VDD.n2844 VDD.n2840 212.329
R14406 VDD.n4081 VDD.n2839 212.329
R14407 VDD.n4088 VDD.n2839 212.329
R14408 VDD.n2835 VDD.n2834 212.329
R14409 VDD.n2834 VDD.n2829 212.329
R14410 VDD.n4091 VDD.n2828 212.329
R14411 VDD.n4098 VDD.n2828 212.329
R14412 VDD.n2824 VDD.n2823 212.329
R14413 VDD.n2823 VDD.n2816 212.329
R14414 VDD.n4101 VDD.n2815 212.329
R14415 VDD.n4108 VDD.n2815 212.329
R14416 VDD.n2811 VDD.n2810 212.329
R14417 VDD.n2810 VDD.n2804 212.329
R14418 VDD.n4111 VDD.n2803 212.329
R14419 VDD.n4118 VDD.n2803 212.329
R14420 VDD.n4124 VDD.n4123 212.329
R14421 VDD.n4125 VDD.n4124 212.329
R14422 VDD.n2795 VDD.n2794 212.329
R14423 VDD.n2795 VDD.n2793 212.329
R14424 VDD.n4133 VDD.n4132 212.329
R14425 VDD.n4133 VDD.n4131 212.329
R14426 VDD.n2787 VDD.n2786 212.329
R14427 VDD.n2786 VDD.n2774 212.329
R14428 VDD.n2769 VDD.n2768 212.329
R14429 VDD.n2768 VDD.n2762 212.329
R14430 VDD.n4145 VDD.n2761 212.329
R14431 VDD.n4152 VDD.n2761 212.329
R14432 VDD.n2757 VDD.n2756 212.329
R14433 VDD.n2756 VDD.n2749 212.329
R14434 VDD.n4155 VDD.n2748 212.329
R14435 VDD.n4162 VDD.n2748 212.329
R14436 VDD.n2744 VDD.n2743 212.329
R14437 VDD.n2743 VDD.n2739 212.329
R14438 VDD.n4165 VDD.n2738 212.329
R14439 VDD.n4172 VDD.n2738 212.329
R14440 VDD.n2734 VDD.n2733 212.329
R14441 VDD.n2733 VDD.n2728 212.329
R14442 VDD.n4175 VDD.n2727 212.329
R14443 VDD.n4182 VDD.n2727 212.329
R14444 VDD.n2789 VDD.n2773 212.329
R14445 VDD.n4142 VDD.n2773 212.329
R14446 VDD.n4062 VDD.n2856 212.329
R14447 VDD.n2856 VDD.n2854 212.329
R14448 VDD.n3945 VDD.n3944 212.329
R14449 VDD.n3944 VDD.n2986 212.329
R14450 VDD.n3946 VDD.n2985 212.329
R14451 VDD.n3953 VDD.n2985 212.329
R14452 VDD.n2981 VDD.n2980 212.329
R14453 VDD.n2980 VDD.n2976 212.329
R14454 VDD.n3956 VDD.n2975 212.329
R14455 VDD.n3963 VDD.n2975 212.329
R14456 VDD.n2971 VDD.n2970 212.329
R14457 VDD.n2970 VDD.n2965 212.329
R14458 VDD.n3966 VDD.n2964 212.329
R14459 VDD.n3973 VDD.n2964 212.329
R14460 VDD.n2960 VDD.n2959 212.329
R14461 VDD.n2959 VDD.n2952 212.329
R14462 VDD.n3976 VDD.n2951 212.329
R14463 VDD.n3983 VDD.n2951 212.329
R14464 VDD.n2947 VDD.n2946 212.329
R14465 VDD.n2946 VDD.n2940 212.329
R14466 VDD.n3986 VDD.n2939 212.329
R14467 VDD.n3993 VDD.n2939 212.329
R14468 VDD.n3999 VDD.n3998 212.329
R14469 VDD.n4000 VDD.n3999 212.329
R14470 VDD.n2931 VDD.n2930 212.329
R14471 VDD.n2931 VDD.n2929 212.329
R14472 VDD.n4008 VDD.n4007 212.329
R14473 VDD.n4008 VDD.n4006 212.329
R14474 VDD.n2923 VDD.n2922 212.329
R14475 VDD.n2922 VDD.n2910 212.329
R14476 VDD.n2905 VDD.n2904 212.329
R14477 VDD.n2904 VDD.n2898 212.329
R14478 VDD.n4020 VDD.n2897 212.329
R14479 VDD.n4027 VDD.n2897 212.329
R14480 VDD.n2893 VDD.n2892 212.329
R14481 VDD.n2892 VDD.n2885 212.329
R14482 VDD.n4030 VDD.n2884 212.329
R14483 VDD.n4037 VDD.n2884 212.329
R14484 VDD.n2880 VDD.n2879 212.329
R14485 VDD.n2879 VDD.n2875 212.329
R14486 VDD.n4040 VDD.n2874 212.329
R14487 VDD.n4047 VDD.n2874 212.329
R14488 VDD.n2870 VDD.n2869 212.329
R14489 VDD.n2869 VDD.n2864 212.329
R14490 VDD.n4050 VDD.n2863 212.329
R14491 VDD.n4057 VDD.n2863 212.329
R14492 VDD.n2925 VDD.n2909 212.329
R14493 VDD.n4017 VDD.n2909 212.329
R14494 VDD.n3294 VDD.n3293 212.329
R14495 VDD.n3293 VDD.n3290 212.329
R14496 VDD.n3285 VDD.n3284 212.329
R14497 VDD.n3284 VDD.n3280 212.329
R14498 VDD.n3598 VDD.n3279 212.329
R14499 VDD.n3605 VDD.n3279 212.329
R14500 VDD.n3274 VDD.n3273 212.329
R14501 VDD.n3274 VDD.n3272 212.329
R14502 VDD.n3613 VDD.n3612 212.329
R14503 VDD.n3613 VDD.n3611 212.329
R14504 VDD.n3295 VDD.n3289 212.329
R14505 VDD.n3595 VDD.n3289 212.329
R14506 VDD.n3447 VDD.n3345 212.329
R14507 VDD.n3345 VDD.n3343 212.329
R14508 VDD.n3440 VDD.n3349 212.329
R14509 VDD.n3350 VDD.n3349 212.329
R14510 VDD.n3433 VDD.n3425 212.329
R14511 VDD.n3425 VDD.n3423 212.329
R14512 VDD.n3484 VDD.n3454 212.329
R14513 VDD.n3454 VDD.n3452 212.329
R14514 VDD.n3477 VDD.n3458 212.329
R14515 VDD.n3459 VDD.n3458 212.329
R14516 VDD.n3471 VDD.n3463 212.329
R14517 VDD.n3463 VDD.n3461 212.329
R14518 VDD.n3336 VDD.n3328 212.329
R14519 VDD.n3328 VDD.n3326 212.329
R14520 VDD.n3325 VDD.n3324 212.329
R14521 VDD.n3506 VDD.n3324 212.329
R14522 VDD.n3511 VDD.n3318 212.329
R14523 VDD.n3318 VDD.n3316 212.329
R14524 VDD.n3542 VDD.n3308 212.329
R14525 VDD.n3308 VDD.n3306 212.329
R14526 VDD.n3535 VDD.n3312 212.329
R14527 VDD.n3313 VDD.n3312 212.329
R14528 VDD.n3528 VDD.n3520 212.329
R14529 VDD.n3520 VDD.n3518 212.329
R14530 VDD.n3578 VDD.n3548 212.329
R14531 VDD.n3548 VDD.n3546 212.329
R14532 VDD.n3571 VDD.n3552 212.329
R14533 VDD.n3553 VDD.n3552 212.329
R14534 VDD.n3565 VDD.n3557 212.329
R14535 VDD.n3557 VDD.n3555 212.329
R14536 VDD.n3392 VDD.n3384 212.329
R14537 VDD.n3384 VDD.n3382 212.329
R14538 VDD.n3381 VDD.n3380 212.329
R14539 VDD.n3411 VDD.n3380 212.329
R14540 VDD.n3416 VDD.n3374 212.329
R14541 VDD.n3374 VDD.n3372 212.329
R14542 VDD.n3937 VDD.n2992 212.329
R14543 VDD.n2992 VDD.n2990 212.329
R14544 VDD.n3820 VDD.n3819 212.329
R14545 VDD.n3819 VDD.n3812 212.329
R14546 VDD.n3821 VDD.n3811 212.329
R14547 VDD.n3828 VDD.n3811 212.329
R14548 VDD.n3807 VDD.n3806 212.329
R14549 VDD.n3806 VDD.n3802 212.329
R14550 VDD.n3831 VDD.n3801 212.329
R14551 VDD.n3838 VDD.n3801 212.329
R14552 VDD.n3797 VDD.n3796 212.329
R14553 VDD.n3796 VDD.n3791 212.329
R14554 VDD.n3841 VDD.n3790 212.329
R14555 VDD.n3848 VDD.n3790 212.329
R14556 VDD.n3786 VDD.n3785 212.329
R14557 VDD.n3785 VDD.n3778 212.329
R14558 VDD.n3851 VDD.n3777 212.329
R14559 VDD.n3858 VDD.n3777 212.329
R14560 VDD.n3773 VDD.n3772 212.329
R14561 VDD.n3772 VDD.n3766 212.329
R14562 VDD.n3861 VDD.n3765 212.329
R14563 VDD.n3868 VDD.n3765 212.329
R14564 VDD.n3874 VDD.n3873 212.329
R14565 VDD.n3875 VDD.n3874 212.329
R14566 VDD.n3757 VDD.n3756 212.329
R14567 VDD.n3757 VDD.n3755 212.329
R14568 VDD.n3883 VDD.n3882 212.329
R14569 VDD.n3883 VDD.n3881 212.329
R14570 VDD.n3749 VDD.n3748 212.329
R14571 VDD.n3748 VDD.n3736 212.329
R14572 VDD.n3731 VDD.n3730 212.329
R14573 VDD.n3730 VDD.n3034 212.329
R14574 VDD.n3895 VDD.n3033 212.329
R14575 VDD.n3902 VDD.n3033 212.329
R14576 VDD.n3029 VDD.n3028 212.329
R14577 VDD.n3028 VDD.n3021 212.329
R14578 VDD.n3905 VDD.n3020 212.329
R14579 VDD.n3912 VDD.n3020 212.329
R14580 VDD.n3016 VDD.n3015 212.329
R14581 VDD.n3015 VDD.n3011 212.329
R14582 VDD.n3915 VDD.n3010 212.329
R14583 VDD.n3922 VDD.n3010 212.329
R14584 VDD.n3006 VDD.n3005 212.329
R14585 VDD.n3005 VDD.n3000 212.329
R14586 VDD.n3925 VDD.n2999 212.329
R14587 VDD.n3932 VDD.n2999 212.329
R14588 VDD.n3751 VDD.n3735 212.329
R14589 VDD.n3892 VDD.n3735 212.329
R14590 VDD.n3397 VDD.t207 176.65
R14591 VDD.n3402 VDD.t986 176.65
R14592 VDD.n3339 VDD.t132 176.65
R14593 VDD.n3492 VDD.t885 176.65
R14594 VDD.n3497 VDD.t123 176.65
R14595 VDD.n3302 VDD.t138 176.65
R14596 VDD.n3586 VDD.t569 176.65
R14597 VDD.n3589 VDD.t22 176.65
R14598 VDD.n1900 VDD.t864 169.018
R14599 VDD.n1653 VDD.t793 169.018
R14600 VDD.n1653 VDD.t244 169.018
R14601 VDD.n1687 VDD.t359 169.018
R14602 VDD.n1687 VDD.t790 169.018
R14603 VDD.n1749 VDD.t383 169.018
R14604 VDD.n1749 VDD.t28 169.018
R14605 VDD.n1724 VDD.t926 169.018
R14606 VDD.n1640 VDD.t610 169.018
R14607 VDD.n1393 VDD.t419 169.018
R14608 VDD.n1393 VDD.t641 169.018
R14609 VDD.n1427 VDD.t16 169.018
R14610 VDD.n1427 VDD.t417 169.018
R14611 VDD.n1489 VDD.t645 169.018
R14612 VDD.n1489 VDD.t895 169.018
R14613 VDD.n1464 VDD.t7 169.018
R14614 VDD.n1380 VDD.t962 169.018
R14615 VDD.n1133 VDD.t883 169.018
R14616 VDD.n1133 VDD.t481 169.018
R14617 VDD.n1167 VDD.t539 169.018
R14618 VDD.n1167 VDD.t880 169.018
R14619 VDD.n1229 VDD.t477 169.018
R14620 VDD.n1229 VDD.t212 169.018
R14621 VDD.n1204 VDD.t104 169.018
R14622 VDD.n1120 VDD.t866 169.018
R14623 VDD.n873 VDD.t624 169.018
R14624 VDD.n873 VDD.t248 169.018
R14625 VDD.n907 VDD.t643 169.018
R14626 VDD.n907 VDD.t873 169.018
R14627 VDD.n969 VDD.t10 169.018
R14628 VDD.n969 VDD.t625 169.018
R14629 VDD.n944 VDD.t660 169.018
R14630 VDD.n860 VDD.t606 169.018
R14631 VDD.n613 VDD.t843 169.018
R14632 VDD.n613 VDD.t354 169.018
R14633 VDD.n647 VDD.t385 169.018
R14634 VDD.n647 VDD.t842 169.018
R14635 VDD.n709 VDD.t357 169.018
R14636 VDD.n709 VDD.t844 169.018
R14637 VDD.n684 VDD.t44 169.018
R14638 VDD.n600 VDD.t964 169.018
R14639 VDD.n353 VDD.t79 169.018
R14640 VDD.n353 VDD.t12 169.018
R14641 VDD.n387 VDD.t250 169.018
R14642 VDD.n387 VDD.t577 169.018
R14643 VDD.n449 VDD.t340 169.018
R14644 VDD.n449 VDD.t959 169.018
R14645 VDD.n424 VDD.t59 169.018
R14646 VDD.n120 VDD.t847 169.018
R14647 VDD.n95 VDD.t171 169.018
R14648 VDD.n70 VDD.t879 169.018
R14649 VDD.n45 VDD.t630 169.018
R14650 VDD.n7516 VDD.t608 169.018
R14651 VDD.n7269 VDD.t156 169.018
R14652 VDD.n7269 VDD.t355 169.018
R14653 VDD.n7303 VDD.t14 169.018
R14654 VDD.n7303 VDD.t561 169.018
R14655 VDD.n7365 VDD.t640 169.018
R14656 VDD.n7365 VDD.t970 169.018
R14657 VDD.n7340 VDD.t914 169.018
R14658 VDD.n6969 VDD.t932 169.018
R14659 VDD.n6944 VDD.t190 169.018
R14660 VDD.n6919 VDD.t584 169.018
R14661 VDD.n6897 VDD.t302 169.018
R14662 VDD.n5112 VDD.t707 169.018
R14663 VDD.n5112 VDD.t434 169.018
R14664 VDD.n5174 VDD.t675 169.018
R14665 VDD.n5174 VDD.t511 169.018
R14666 VDD.n5209 VDD.t458 169.018
R14667 VDD.n5209 VDD.t753 169.018
R14668 VDD.n6764 VDD.t920 169.018
R14669 VDD.n5248 VDD.t757 169.018
R14670 VDD.n5248 VDD.t483 169.018
R14671 VDD.n5310 VDD.t681 169.018
R14672 VDD.n5310 VDD.t521 169.018
R14673 VDD.n5345 VDD.t466 169.018
R14674 VDD.n5345 VDD.t759 169.018
R14675 VDD.n6641 VDD.t841 169.018
R14676 VDD.n5384 VDD.t663 169.018
R14677 VDD.n5384 VDD.t493 169.018
R14678 VDD.n5446 VDD.t745 169.018
R14679 VDD.n5446 VDD.t476 169.018
R14680 VDD.n5481 VDD.t479 169.018
R14681 VDD.n5481 VDD.t673 169.018
R14682 VDD.n6518 VDD.t24 169.018
R14683 VDD.n5520 VDD.t735 169.018
R14684 VDD.n5520 VDD.t460 169.018
R14685 VDD.n5582 VDD.t763 169.018
R14686 VDD.n5582 VDD.t491 169.018
R14687 VDD.n5617 VDD.t444 169.018
R14688 VDD.n5617 VDD.t737 169.018
R14689 VDD.n6395 VDD.t622 169.018
R14690 VDD.n5656 VDD.t679 169.018
R14691 VDD.n5656 VDD.t507 169.018
R14692 VDD.n5718 VDD.t721 169.018
R14693 VDD.n5718 VDD.t454 169.018
R14694 VDD.n5753 VDD.t464 169.018
R14695 VDD.n5753 VDD.t755 169.018
R14696 VDD.n6272 VDD.t917 169.018
R14697 VDD.n5792 VDD.t705 169.018
R14698 VDD.n5792 VDD.t436 169.018
R14699 VDD.n5854 VDD.t741 169.018
R14700 VDD.n5854 VDD.t472 169.018
R14701 VDD.n5889 VDD.t517 169.018
R14702 VDD.n5889 VDD.t709 169.018
R14703 VDD.n6149 VDD.t882 169.018
R14704 VDD.n5928 VDD.t531 169.018
R14705 VDD.n5928 VDD.t727 169.018
R14706 VDD.n5990 VDD.t535 169.018
R14707 VDD.n5990 VDD.t729 169.018
R14708 VDD.n6025 VDD.t667 169.018
R14709 VDD.n6025 VDD.t495 169.018
R14710 VDD.n6026 VDD.t889 169.018
R14711 VDD.n5956 VDD.t1025 169.018
R14712 VDD.n5820 VDD.t1080 169.018
R14713 VDD.n5684 VDD.t1055 169.018
R14714 VDD.n5548 VDD.t1097 169.018
R14715 VDD.n5412 VDD.t1085 169.018
R14716 VDD.n5276 VDD.t1059 169.018
R14717 VDD.n5140 VDD.t1077 169.018
R14718 VDD.n4922 VDD.t677 169.018
R14719 VDD.n4922 VDD.t513 169.018
R14720 VDD.n4860 VDD.t761 169.018
R14721 VDD.n4860 VDD.t487 169.018
R14722 VDD.n4826 VDD.t497 169.018
R14723 VDD.n4826 VDD.t693 169.018
R14724 VDD.n5073 VDD.t575 169.018
R14725 VDD.n4897 VDD.t1053 169.018
R14726 VDD.n3792 VDD.t719 169.018
R14727 VDD.n3792 VDD.t446 169.018
R14728 VDD.n3767 VDD.t1092 169.018
R14729 VDD.n2966 VDD.t725 169.018
R14730 VDD.n2966 VDD.t448 169.018
R14731 VDD.n3940 VDD.t942 169.018
R14732 VDD.n3001 VDD.t529 169.018
R14733 VDD.n3001 VDD.t713 169.018
R14734 VDD.n3035 VDD.t665 169.018
R14735 VDD.n3035 VDD.t485 169.018
R14736 VDD.n2941 VDD.t1035 169.018
R14737 VDD.n2830 VDD.t699 169.018
R14738 VDD.n2830 VDD.t525 169.018
R14739 VDD.n4065 VDD.t154 169.018
R14740 VDD.n2865 VDD.t503 169.018
R14741 VDD.n2865 VDD.t687 169.018
R14742 VDD.n2899 VDD.t711 169.018
R14743 VDD.n2899 VDD.t438 169.018
R14744 VDD.n2805 VDD.t1007 169.018
R14745 VDD.n2694 VDD.t747 169.018
R14746 VDD.n2694 VDD.t470 169.018
R14747 VDD.n4190 VDD.t125 169.018
R14748 VDD.n2729 VDD.t456 169.018
R14749 VDD.n2729 VDD.t739 169.018
R14750 VDD.n2763 VDD.t683 169.018
R14751 VDD.n2763 VDD.t515 169.018
R14752 VDD.n2669 VDD.t1063 169.018
R14753 VDD.n2558 VDD.t731 169.018
R14754 VDD.n2558 VDD.t452 169.018
R14755 VDD.n4315 VDD.t765 169.018
R14756 VDD.n2593 VDD.t537 169.018
R14757 VDD.n2593 VDD.t717 169.018
R14758 VDD.n2627 VDD.t669 169.018
R14759 VDD.n2627 VDD.t489 169.018
R14760 VDD.n2533 VDD.t1039 169.018
R14761 VDD.n2422 VDD.t703 169.018
R14762 VDD.n2422 VDD.t533 169.018
R14763 VDD.n4440 VDD.t797 169.018
R14764 VDD.n2457 VDD.t505 169.018
R14765 VDD.n2457 VDD.t691 169.018
R14766 VDD.n2491 VDD.t715 169.018
R14767 VDD.n2491 VDD.t442 169.018
R14768 VDD.n2397 VDD.t1011 169.018
R14769 VDD.n2286 VDD.t751 169.018
R14770 VDD.n2286 VDD.t474 169.018
R14771 VDD.n4565 VDD.t26 169.018
R14772 VDD.n2321 VDD.t509 169.018
R14773 VDD.n2321 VDD.t697 169.018
R14774 VDD.n2355 VDD.t689 169.018
R14775 VDD.n2355 VDD.t519 169.018
R14776 VDD.n2261 VDD.t1083 169.018
R14777 VDD.n2150 VDD.t743 169.018
R14778 VDD.n2150 VDD.t468 169.018
R14779 VDD.n4690 VDD.t66 169.018
R14780 VDD.n2185 VDD.t499 169.018
R14781 VDD.n2185 VDD.t685 169.018
R14782 VDD.n2219 VDD.t723 169.018
R14783 VDD.n2219 VDD.t450 169.018
R14784 VDD.n2125 VDD.t1069 169.018
R14785 VDD.n4815 VDD.t304 169.018
R14786 VDD.n2049 VDD.t462 169.018
R14787 VDD.n2049 VDD.t749 169.018
R14788 VDD.n2083 VDD.t701 169.018
R14789 VDD.n2083 VDD.t527 169.018
R14790 VDD.n2014 VDD.t695 169.018
R14791 VDD.n2014 VDD.t523 169.018
R14792 VDD.n1989 VDD.t1075 169.018
R14793 VDD.n7256 VDD.t650 169.018
R14794 VDD.n1913 VDD.t440 169.018
R14795 VDD.n1913 VDD.t733 169.018
R14796 VDD.n1947 VDD.t671 169.018
R14797 VDD.n1947 VDD.t501 169.018
R14798 VDD.n7519 VDD.t868 169.018
R14799 VDD.n7520 VDD.t242 169.018
R14800 VDD.n7520 VDD.t251 169.018
R14801 VDD.n7732 VDD.t343 169.018
R14802 VDD.n7732 VDD.t240 169.018
R14803 VDD.n7616 VDD.t210 169.018
R14804 VDD.n7616 VDD.t74 169.018
R14805 VDD.n7591 VDD.t833 169.018
R14806 VDD.n3436 VDD.t855 169.012
R14807 VDD.n3474 VDD.t811 169.012
R14808 VDD.n3315 VDD.t272 169.012
R14809 VDD.n3531 VDD.t997 169.012
R14810 VDD.n3568 VDD.t409 169.012
R14811 VDD.n3371 VDD.t783 169.012
R14812 VDD.n3265 VDD.t87 169.012
R14813 VDD.n3265 VDD.t903 169.012
R14814 VDD.n1675 VDD.t927 168.635
R14815 VDD.n1675 VDD.t875 168.635
R14816 VDD.n1674 VDD.t600 168.635
R14817 VDD.n1674 VDD.t924 168.635
R14818 VDD.n1709 VDD.t598 168.635
R14819 VDD.n1709 VDD.t979 168.635
R14820 VDD.n1708 VDD.t568 168.635
R14821 VDD.n1708 VDD.t991 168.635
R14822 VDD.n1737 VDD.t159 168.635
R14823 VDD.n1737 VDD.t992 168.635
R14824 VDD.n1736 VDD.t596 168.635
R14825 VDD.n1736 VDD.t158 168.635
R14826 VDD.n1771 VDD.t55 168.635
R14827 VDD.n1771 VDD.t936 168.635
R14828 VDD.n1770 VDD.t423 168.635
R14829 VDD.n1770 VDD.t265 168.635
R14830 VDD.n1415 VDD.t8 168.635
R14831 VDD.n1415 VDD.t982 168.635
R14832 VDD.n1414 VDD.t807 168.635
R14833 VDD.n1414 VDD.t5 168.635
R14834 VDD.n1449 VDD.t929 168.635
R14835 VDD.n1449 VDD.t94 168.635
R14836 VDD.n1448 VDD.t392 168.635
R14837 VDD.n1448 VDD.t770 168.635
R14838 VDD.n1477 VDD.t816 168.635
R14839 VDD.n1477 VDD.t772 168.635
R14840 VDD.n1476 VDD.t928 168.635
R14841 VDD.n1476 VDD.t817 168.635
R14842 VDD.n1511 VDD.t995 168.635
R14843 VDD.n1511 VDD.t826 168.635
R14844 VDD.n1510 VDD.t299 168.635
R14845 VDD.n1510 VDD.t1107 168.635
R14846 VDD.n1155 VDD.t275 168.635
R14847 VDD.n1155 VDD.t638 168.635
R14848 VDD.n1154 VDD.t394 168.635
R14849 VDD.n1154 VDD.t102 168.635
R14850 VDD.n1189 VDD.t966 168.635
R14851 VDD.n1189 VDD.t550 168.635
R14852 VDD.n1188 VDD.t413 168.635
R14853 VDD.n1188 VDD.t779 168.635
R14854 VDD.n1217 VDD.t179 168.635
R14855 VDD.n1217 VDD.t777 168.635
R14856 VDD.n1216 VDD.t192 168.635
R14857 VDD.n1216 VDD.t180 168.635
R14858 VDD.n1251 VDD.t269 168.635
R14859 VDD.n1251 VDD.t361 168.635
R14860 VDD.n1250 VDD.t615 168.635
R14861 VDD.n1250 VDD.t115 168.635
R14862 VDD.n895 VDD.t766 168.635
R14863 VDD.n895 VDD.t631 168.635
R14864 VDD.n894 VDD.t602 168.635
R14865 VDD.n894 VDD.t658 168.635
R14866 VDD.n929 VDD.t175 168.635
R14867 VDD.n929 VDD.t430 168.635
R14868 VDD.n928 VDD.t824 168.635
R14869 VDD.n928 VDD.t910 168.635
R14870 VDD.n957 VDD.t348 168.635
R14871 VDD.n957 VDD.t909 168.635
R14872 VDD.n956 VDD.t173 168.635
R14873 VDD.n956 VDD.t347 168.635
R14874 VDD.n991 VDD.t809 168.635
R14875 VDD.n991 VDD.t319 168.635
R14876 VDD.n990 VDD.t540 168.635
R14877 VDD.n990 VDD.t825 168.635
R14878 VDD.n635 VDD.t45 168.635
R14879 VDD.n635 VDD.t121 168.635
R14880 VDD.n634 VDD.t965 168.635
R14881 VDD.n634 VDD.t42 168.635
R14882 VDD.n669 VDD.t167 168.635
R14883 VDD.n669 VDD.t853 168.635
R14884 VDD.n668 VDD.t221 168.635
R14885 VDD.n668 VDD.t613 168.635
R14886 VDD.n697 VDD.t61 168.635
R14887 VDD.n697 VDD.t614 168.635
R14888 VDD.n696 VDD.t165 168.635
R14889 VDD.n696 VDD.t62 168.635
R14890 VDD.n731 VDD.t279 168.635
R14891 VDD.n731 VDD.t294 168.635
R14892 VDD.n730 VDD.t64 168.635
R14893 VDD.n730 VDD.t560 168.635
R14894 VDD.n375 VDD.t556 168.635
R14895 VDD.n375 VDD.t334 168.635
R14896 VDD.n374 VDD.t395 168.635
R14897 VDD.n374 VDD.t557 168.635
R14898 VDD.n409 VDD.t234 168.635
R14899 VDD.n409 VDD.t108 168.635
R14900 VDD.n408 VDD.t76 168.635
R14901 VDD.n408 VDD.t975 168.635
R14902 VDD.n437 VDD.t989 168.635
R14903 VDD.n437 VDD.t273 168.635
R14904 VDD.n436 VDD.t205 168.635
R14905 VDD.n436 VDD.t990 168.635
R14906 VDD.n471 VDD.t785 168.635
R14907 VDD.n471 VDD.t336 168.635
R14908 VDD.n470 VDD.t398 168.635
R14909 VDD.n470 VDD.t363 168.635
R14910 VDD.n135 VDD.t214 168.635
R14911 VDD.n135 VDD.t371 168.635
R14912 VDD.n132 VDD.t655 168.635
R14913 VDD.n132 VDD.t1073 168.635
R14914 VDD.n110 VDD.t620 168.635
R14915 VDD.n110 VDD.t129 168.635
R14916 VDD.n107 VDD.t977 168.635
R14917 VDD.n107 VDD.t1027 168.635
R14918 VDD.n85 VDD.t839 168.635
R14919 VDD.n85 VDD.t922 168.635
R14920 VDD.n82 VDD.t958 168.635
R14921 VDD.n82 VDD.t1066 168.635
R14922 VDD.n60 VDD.t352 168.635
R14923 VDD.n60 VDD.t647 168.635
R14924 VDD.n57 VDD.t78 168.635
R14925 VDD.n57 VDD.t1090 168.635
R14926 VDD.n7291 VDD.t915 168.635
R14927 VDD.n7291 VDD.t981 168.635
R14928 VDD.n7290 VDD.t338 168.635
R14929 VDD.n7290 VDD.t912 168.635
R14930 VDD.n7325 VDD.t972 168.635
R14931 VDD.n7325 VDD.t113 168.635
R14932 VDD.n7324 VDD.t288 168.635
R14933 VDD.n7324 VDD.t949 168.635
R14934 VDD.n7353 VDD.t49 168.635
R14935 VDD.n7353 VDD.t223 168.635
R14936 VDD.n7352 VDD.t971 168.635
R14937 VDD.n7352 VDD.t50 168.635
R14938 VDD.n7387 VDD.t545 168.635
R14939 VDD.n7387 VDD.t803 168.635
R14940 VDD.n7386 VDD.t653 168.635
R14941 VDD.n7386 VDD.t874 168.635
R14942 VDD.n6984 VDD.t940 168.635
R14943 VDD.n6984 VDD.t969 168.635
R14944 VDD.n6981 VDD.t1037 168.635
R14945 VDD.n6981 VDD.t955 168.635
R14946 VDD.n6959 VDD.t127 168.635
R14947 VDD.n6959 VDD.t72 168.635
R14948 VDD.n6956 VDD.t1013 168.635
R14949 VDD.n6956 VDD.t421 168.635
R14950 VDD.n6934 VDD.t799 168.635
R14951 VDD.n6934 VDD.t792 168.635
R14952 VDD.n6931 VDD.t1041 168.635
R14953 VDD.n6931 VDD.t400 168.635
R14954 VDD.n6909 VDD.t774 168.635
R14955 VDD.n6909 VDD.t277 168.635
R14956 VDD.n6889 VDD.t1009 168.635
R14957 VDD.n6889 VDD.t951 168.635
R14958 VDD.n5075 VDD.t850 168.635
R14959 VDD.n5075 VDD.t350 168.635
R14960 VDD.n5074 VDD.t930 168.635
R14961 VDD.n5074 VDD.t432 168.635
R14962 VDD.n5124 VDD.t286 168.635
R14963 VDD.n5124 VDD.t851 168.635
R14964 VDD.n5123 VDD.t331 168.635
R14965 VDD.n5123 VDD.t229 168.635
R14966 VDD.n5152 VDD.t612 168.635
R14967 VDD.n5152 VDD.t227 168.635
R14968 VDD.n5151 VDD.t287 168.635
R14969 VDD.n5151 VDD.t163 168.635
R14970 VDD.n5186 VDD.t391 168.635
R14971 VDD.n5186 VDD.t1031 168.635
R14972 VDD.n5185 VDD.t1095 168.635
R14973 VDD.n5185 VDD.t780 168.635
R14974 VDD.n5211 VDD.t321 168.635
R14975 VDD.n5211 VDD.t918 168.635
R14976 VDD.n5210 VDD.t306 168.635
R14977 VDD.n5210 VDD.t587 168.635
R14978 VDD.n5260 VDD.t317 168.635
R14979 VDD.n5260 VDD.t543 168.635
R14980 VDD.n5259 VDD.t379 168.635
R14981 VDD.n5259 VDD.t376 168.635
R14982 VDD.n5288 VDD.t367 168.635
R14983 VDD.n5288 VDD.t377 168.635
R14984 VDD.n5287 VDD.t315 168.635
R14985 VDD.n5287 VDD.t661 168.635
R14986 VDD.n5322 VDD.t904 168.635
R14987 VDD.n5322 VDD.t1078 168.635
R14988 VDD.n5321 VDD.t1033 168.635
R14989 VDD.n5321 VDD.t836 168.635
R14990 VDD.n5347 VDD.t195 168.635
R14991 VDD.n5347 VDD.t837 168.635
R14992 VDD.n5346 VDD.t313 168.635
R14993 VDD.n5346 VDD.t34 168.635
R14994 VDD.n5396 VDD.t209 168.635
R14995 VDD.n5396 VDD.t551 168.635
R14996 VDD.n5395 VDD.t140 168.635
R14997 VDD.n5395 VDD.t282 168.635
R14998 VDD.n5424 VDD.t18 168.635
R14999 VDD.n5424 VDD.t281 168.635
R15000 VDD.n5423 VDD.t585 168.635
R15001 VDD.n5423 VDD.t274 168.635
R15002 VDD.n5458 VDD.t426 168.635
R15003 VDD.n5458 VDD.t1093 168.635
R15004 VDD.n5457 VDD.t1061 168.635
R15005 VDD.n5457 VDD.t804 168.635
R15006 VDD.n5483 VDD.t656 168.635
R15007 VDD.n5483 VDD.t130 168.635
R15008 VDD.n5482 VDD.t47 168.635
R15009 VDD.n5482 VDD.t254 168.635
R15010 VDD.n5532 VDD.t258 168.635
R15011 VDD.n5532 VDD.t960 168.635
R15012 VDD.n5531 VDD.t238 168.635
R15013 VDD.n5531 VDD.t891 168.635
R15014 VDD.n5560 VDD.t795 168.635
R15015 VDD.n5560 VDD.t908 168.635
R15016 VDD.n5559 VDD.t136 168.635
R15017 VDD.n5559 VDD.t983 168.635
R15018 VDD.n5594 VDD.t886 168.635
R15019 VDD.n5594 VDD.t1047 168.635
R15020 VDD.n5593 VDD.t1003 168.635
R15021 VDD.n5593 VDD.t872 168.635
R15022 VDD.n5619 VDD.t110 168.635
R15023 VDD.n5619 VDD.t623 168.635
R15024 VDD.n5618 VDD.t365 168.635
R15025 VDD.n5618 VDD.t252 168.635
R15026 VDD.n5668 VDD.t146 168.635
R15027 VDD.n5668 VDD.t554 168.635
R15028 VDD.n5667 VDD.t553 168.635
R15029 VDD.n5667 VDD.t268 168.635
R15030 VDD.n5696 VDD.t869 168.635
R15031 VDD.n5696 VDD.t820 168.635
R15032 VDD.n5695 VDD.t148 168.635
R15033 VDD.n5695 VDD.t117 168.635
R15034 VDD.n5730 VDD.t980 168.635
R15035 VDD.n5730 VDD.t1070 168.635
R15036 VDD.n5729 VDD.t1029 168.635
R15037 VDD.n5729 VDD.t369 168.635
R15038 VDD.n5755 VDD.t264 168.635
R15039 VDD.n5755 VDD.t372 168.635
R15040 VDD.n5754 VDD.t142 168.635
R15041 VDD.n5754 VDD.t424 168.635
R15042 VDD.n5804 VDD.t945 168.635
R15043 VDD.n5804 VDD.t828 168.635
R15044 VDD.n5803 VDD.t829 168.635
R15045 VDD.n5803 VDD.t987 168.635
R15046 VDD.n5832 VDD.t978 168.635
R15047 VDD.n5832 VDD.t633 168.635
R15048 VDD.n5831 VDD.t946 168.635
R15049 VDD.n5831 VDD.t188 168.635
R15050 VDD.n5866 VDD.t414 168.635
R15051 VDD.n5866 VDD.t1088 168.635
R15052 VDD.n5865 VDD.t1057 168.635
R15053 VDD.n5865 VDD.t342 168.635
R15054 VDD.n5891 VDD.t411 168.635
R15055 VDD.n5891 VDD.t246 168.635
R15056 VDD.n5890 VDD.t819 168.635
R15057 VDD.n5890 VDD.t38 168.635
R15058 VDD.n5940 VDD.t323 168.635
R15059 VDD.n5940 VDD.t57 168.635
R15060 VDD.n5939 VDD.t295 168.635
R15061 VDD.n5939 VDD.t973 168.635
R15062 VDD.n5968 VDD.t860 168.635
R15063 VDD.n5968 VDD.t974 168.635
R15064 VDD.n5967 VDD.t325 168.635
R15065 VDD.n5967 VDD.t203 168.635
R15066 VDD.n6002 VDD.t186 168.635
R15067 VDD.n6002 VDD.t1044 168.635
R15068 VDD.n6001 VDD.t1001 168.635
R15069 VDD.n6001 VDD.t887 168.635
R15070 VDD.n4952 VDD.t332 168.635
R15071 VDD.n4952 VDD.t648 168.635
R15072 VDD.n4951 VDD.t184 168.635
R15073 VDD.n4951 VDD.t182 168.635
R15074 VDD.n4910 VDD.t291 168.635
R15075 VDD.n4910 VDD.t382 168.635
R15076 VDD.n4909 VDD.t381 168.635
R15077 VDD.n4909 VDD.t119 168.635
R15078 VDD.n4882 VDD.t898 168.635
R15079 VDD.n4882 VDD.t85 168.635
R15080 VDD.n4881 VDD.t947 168.635
R15081 VDD.n4881 VDD.t260 168.635
R15082 VDD.n4848 VDD.t290 168.635
R15083 VDD.n4848 VDD.t1005 168.635
R15084 VDD.n4847 VDD.t1081 168.635
R15085 VDD.n4847 VDD.t576 168.635
R15086 VDD.n3741 VDD.t232 168.635
R15087 VDD.n3741 VDD.t111 168.635
R15088 VDD.n3740 VDD.t52 168.635
R15089 VDD.n3740 VDD.t283 168.635
R15090 VDD.n3780 VDD.t967 168.635
R15091 VDD.n3780 VDD.t285 168.635
R15092 VDD.n3779 VDD.t570 168.635
R15093 VDD.n3779 VDD.t559 168.635
R15094 VDD.n3814 VDD.t890 168.635
R15095 VDD.n3814 VDD.t862 168.635
R15096 VDD.n3813 VDD.t428 168.635
R15097 VDD.n3813 VDD.t236 168.635
R15098 VDD.n2915 VDD.t1104 168.635
R15099 VDD.n2915 VDD.t822 168.635
R15100 VDD.n2914 VDD.t956 168.635
R15101 VDD.n2914 VDD.t311 168.635
R15102 VDD.n2954 VDD.t197 168.635
R15103 VDD.n2954 VDD.t309 168.635
R15104 VDD.n2953 VDD.t1105 168.635
R15105 VDD.n2953 VDD.t198 168.635
R15106 VDD.n2988 VDD.t943 168.635
R15107 VDD.n2988 VDD.t327 168.635
R15108 VDD.n2987 VDD.t297 168.635
R15109 VDD.n2987 VDD.t627 168.635
R15110 VDD.n3023 VDD.t1064 168.635
R15111 VDD.n3023 VDD.t152 168.635
R15112 VDD.n3022 VDD.t938 168.635
R15113 VDD.n3022 VDD.t1015 168.635
R15114 VDD.n2779 VDD.t81 168.635
R15115 VDD.n2779 VDD.t611 168.635
R15116 VDD.n2778 VDD.t374 168.635
R15117 VDD.n2778 VDD.t201 168.635
R15118 VDD.n2818 VDD.t326 168.635
R15119 VDD.n2818 VDD.t588 168.635
R15120 VDD.n2817 VDD.t83 168.635
R15121 VDD.n2817 VDD.t169 168.635
R15122 VDD.n2852 VDD.t953 168.635
R15123 VDD.n2852 VDD.t100 168.635
R15124 VDD.n2851 VDD.t861 168.635
R15125 VDD.n2851 VDD.t293 168.635
R15126 VDD.n2887 VDD.t1046 168.635
R15127 VDD.n2887 VDD.t935 168.635
R15128 VDD.n2886 VDD.t952 168.635
R15129 VDD.n2886 VDD.t1099 168.635
R15130 VDD.n2643 VDD.t387 168.635
R15131 VDD.n2643 VDD.t894 168.635
R15132 VDD.n2642 VDD.t32 168.635
R15133 VDD.n2642 VDD.t617 168.635
R15134 VDD.n2682 VDD.t1103 168.635
R15135 VDD.n2682 VDD.t618 168.635
R15136 VDD.n2681 VDD.t389 168.635
R15137 VDD.n2681 VDD.t345 168.635
R15138 VDD.n2716 VDD.t3 168.635
R15139 VDD.n2716 VDD.t893 168.635
R15140 VDD.n2715 VDD.t1101 168.635
R15141 VDD.n2715 VDD.t900 168.635
R15142 VDD.n2751 VDD.t1019 168.635
R15143 VDD.n2751 VDD.t230 168.635
R15144 VDD.n2750 VDD.t1 168.635
R15145 VDD.n2750 VDD.t1087 168.635
R15146 VDD.n2507 VDD.t592 168.635
R15147 VDD.n2507 VDD.t1102 168.635
R15148 VDD.n2506 VDD.t329 168.635
R15149 VDD.n2506 VDD.t20 168.635
R15150 VDD.n2546 VDD.t200 168.635
R15151 VDD.n2546 VDD.t905 168.635
R15152 VDD.n2545 VDD.t594 168.635
R15153 VDD.n2545 VDD.t767 168.635
R15154 VDD.n2580 VDD.t70 168.635
R15155 VDD.n2580 VDD.t40 168.635
R15156 VDD.n2579 VDD.t628 168.635
R15157 VDD.n2579 VDD.t375 168.635
R15158 VDD.n2615 VDD.t1071 168.635
R15159 VDD.n2615 VDD.t586 168.635
R15160 VDD.n2614 VDD.t68 168.635
R15161 VDD.n2614 VDD.t1023 168.635
R15162 VDD.n2371 VDD.t216 168.635
R15163 VDD.n2371 VDD.t267 168.635
R15164 VDD.n2370 VDD.t582 168.635
R15165 VDD.n2370 VDD.t219 168.635
R15166 VDD.n2410 VDD.t616 168.635
R15167 VDD.n2410 VDD.t589 168.635
R15168 VDD.n2409 VDD.t218 168.635
R15169 VDD.n2409 VDD.t92 168.635
R15170 VDD.n2444 VDD.t802 168.635
R15171 VDD.n2444 VDD.t899 168.635
R15172 VDD.n2443 VDD.t161 168.635
R15173 VDD.n2443 VDD.t591 168.635
R15174 VDD.n2479 VDD.t1049 168.635
R15175 VDD.n2479 VDD.t876 168.635
R15176 VDD.n2478 VDD.t801 168.635
R15177 VDD.n2478 VDD.t1100 168.635
R15178 VDD.n2235 VDD.t96 168.635
R15179 VDD.n2235 VDD.t134 168.635
R15180 VDD.n2234 VDD.t300 168.635
R15181 VDD.n2234 VDD.t255 168.635
R15182 VDD.n2274 VDD.t933 168.635
R15183 VDD.n2274 VDD.t776 168.635
R15184 VDD.n2273 VDD.t98 168.635
R15185 VDD.n2273 VDD.t144 168.635
R15186 VDD.n2308 VDD.t789 168.635
R15187 VDD.n2308 VDD.t870 168.635
R15188 VDD.n2307 VDD.t542 168.635
R15189 VDD.n2307 VDD.t897 168.635
R15190 VDD.n2343 VDD.t1094 168.635
R15191 VDD.n2343 VDD.t859 168.635
R15192 VDD.n2342 VDD.t937 168.635
R15193 VDD.n2342 VDD.t1051 168.635
R15194 VDD.n2099 VDD.t906 168.635
R15195 VDD.n2099 VDD.t262 168.635
R15196 VDD.n2098 VDD.t877 168.635
R15197 VDD.n2098 VDD.t563 168.635
R15198 VDD.n2138 VDD.t1106 168.635
R15199 VDD.n2138 VDD.t565 168.635
R15200 VDD.n2137 VDD.t907 168.635
R15201 VDD.n2137 VDD.t849 168.635
R15202 VDD.n2172 VDD.t775 168.635
R15203 VDD.n2172 VDD.t635 168.635
R15204 VDD.n2171 VDD.t818 168.635
R15205 VDD.n2171 VDD.t549 168.635
R15206 VDD.n2207 VDD.t1043 168.635
R15207 VDD.n2207 VDD.t397 168.635
R15208 VDD.n2206 VDD.t814 168.635
R15209 VDD.n2206 VDD.t1098 168.635
R15210 VDD.n2071 VDD.t1017 168.635
R15211 VDD.n2071 VDD.t984 168.635
R15212 VDD.n2070 VDD.t416 168.635
R15213 VDD.n2070 VDD.t1086 168.635
R15214 VDD.n1963 VDD.t105 168.635
R15215 VDD.n1963 VDD.t150 168.635
R15216 VDD.n1962 VDD.t571 168.635
R15217 VDD.n1962 VDD.t36 168.635
R15218 VDD.n2002 VDD.t999 168.635
R15219 VDD.n2002 VDD.t107 168.635
R15220 VDD.n2001 VDD.t768 168.635
R15221 VDD.n2001 VDD.t30 168.635
R15222 VDD.n2036 VDD.t896 168.635
R15223 VDD.n2036 VDD.t194 168.635
R15224 VDD.n2035 VDD.t307 168.635
R15225 VDD.n2035 VDD.t547 168.635
R15226 VDD.n1935 VDD.t1067 168.635
R15227 VDD.n1935 VDD.t573 168.635
R15228 VDD.n1934 VDD.t651 168.635
R15229 VDD.n1934 VDD.t1021 168.635
R15230 VDD.n23 VDD.t834 168.635
R15231 VDD.n23 VDD.t852 168.635
R15232 VDD.n22 VDD.t604 168.635
R15233 VDD.n22 VDD.t831 168.635
R15234 VDD.n7576 VDD.t637 168.635
R15235 VDD.n7576 VDD.t225 168.635
R15236 VDD.n7575 VDD.t823 168.635
R15237 VDD.n7575 VDD.t579 168.635
R15238 VDD.n7604 VDD.t407 168.635
R15239 VDD.n7604 VDD.t581 168.635
R15240 VDD.n7603 VDD.t636 168.635
R15241 VDD.n7603 VDD.t406 168.635
R15242 VDD.n7638 VDD.t901 168.635
R15243 VDD.n7638 VDD.t404 168.635
R15244 VDD.n7637 VDD.t845 168.635
R15245 VDD.n7637 VDD.t857 168.635
R15246 VDD.n7697 VDD.n7585 166.238
R15247 VDD.n7699 VDD.n7585 166.238
R15248 VDD.n7523 VDD.n7522 166.238
R15249 VDD.n7522 VDD.n44 166.238
R15250 VDD.n1830 VDD.n1718 166.238
R15251 VDD.n1832 VDD.n1718 166.238
R15252 VDD.n1898 VDD.n1897 166.238
R15253 VDD.n1898 VDD.n1642 166.238
R15254 VDD.n1570 VDD.n1458 166.238
R15255 VDD.n1572 VDD.n1458 166.238
R15256 VDD.n1638 VDD.n1637 166.238
R15257 VDD.n1638 VDD.n1382 166.238
R15258 VDD.n1310 VDD.n1198 166.238
R15259 VDD.n1312 VDD.n1198 166.238
R15260 VDD.n1378 VDD.n1377 166.238
R15261 VDD.n1378 VDD.n1122 166.238
R15262 VDD.n1050 VDD.n938 166.238
R15263 VDD.n1052 VDD.n938 166.238
R15264 VDD.n1118 VDD.n1117 166.238
R15265 VDD.n1118 VDD.n862 166.238
R15266 VDD.n790 VDD.n678 166.238
R15267 VDD.n792 VDD.n678 166.238
R15268 VDD.n858 VDD.n857 166.238
R15269 VDD.n858 VDD.n602 166.238
R15270 VDD.n530 VDD.n418 166.238
R15271 VDD.n532 VDD.n418 166.238
R15272 VDD.n598 VDD.n597 166.238
R15273 VDD.n598 VDD.n342 166.238
R15274 VDD.n149 VDD.n146 166.238
R15275 VDD.n151 VDD.n146 166.238
R15276 VDD.n157 VDD.n156 166.238
R15277 VDD.n157 VDD.n137 166.238
R15278 VDD.n163 VDD.n160 166.238
R15279 VDD.n165 VDD.n160 166.238
R15280 VDD.n170 VDD.n129 166.238
R15281 VDD.n172 VDD.n129 166.238
R15282 VDD.n178 VDD.n177 166.238
R15283 VDD.n178 VDD.n121 166.238
R15284 VDD.n184 VDD.n181 166.238
R15285 VDD.n186 VDD.n181 166.238
R15286 VDD.n192 VDD.n191 166.238
R15287 VDD.n192 VDD.n112 166.238
R15288 VDD.n198 VDD.n195 166.238
R15289 VDD.n200 VDD.n195 166.238
R15290 VDD.n205 VDD.n104 166.238
R15291 VDD.n207 VDD.n104 166.238
R15292 VDD.n213 VDD.n212 166.238
R15293 VDD.n213 VDD.n96 166.238
R15294 VDD.n219 VDD.n216 166.238
R15295 VDD.n221 VDD.n216 166.238
R15296 VDD.n227 VDD.n226 166.238
R15297 VDD.n227 VDD.n87 166.238
R15298 VDD.n233 VDD.n230 166.238
R15299 VDD.n235 VDD.n230 166.238
R15300 VDD.n240 VDD.n79 166.238
R15301 VDD.n242 VDD.n79 166.238
R15302 VDD.n248 VDD.n247 166.238
R15303 VDD.n248 VDD.n71 166.238
R15304 VDD.n254 VDD.n251 166.238
R15305 VDD.n256 VDD.n251 166.238
R15306 VDD.n262 VDD.n261 166.238
R15307 VDD.n262 VDD.n62 166.238
R15308 VDD.n268 VDD.n265 166.238
R15309 VDD.n270 VDD.n265 166.238
R15310 VDD.n275 VDD.n54 166.238
R15311 VDD.n277 VDD.n54 166.238
R15312 VDD.n283 VDD.n282 166.238
R15313 VDD.n283 VDD.n46 166.238
R15314 VDD.n7446 VDD.n7334 166.238
R15315 VDD.n7448 VDD.n7334 166.238
R15316 VDD.n7514 VDD.n7513 166.238
R15317 VDD.n7514 VDD.n7258 166.238
R15318 VDD.n7254 VDD.n7253 166.238
R15319 VDD.n7254 VDD.n1902 166.238
R15320 VDD.n7189 VDD.n1983 166.238
R15321 VDD.n7191 VDD.n1983 166.238
R15322 VDD.n6998 VDD.n6995 166.238
R15323 VDD.n7000 VDD.n6995 166.238
R15324 VDD.n7006 VDD.n7005 166.238
R15325 VDD.n7006 VDD.n6986 166.238
R15326 VDD.n7012 VDD.n7009 166.238
R15327 VDD.n7014 VDD.n7009 166.238
R15328 VDD.n7019 VDD.n6978 166.238
R15329 VDD.n7021 VDD.n6978 166.238
R15330 VDD.n7027 VDD.n7026 166.238
R15331 VDD.n7027 VDD.n6970 166.238
R15332 VDD.n7033 VDD.n7030 166.238
R15333 VDD.n7035 VDD.n7030 166.238
R15334 VDD.n7041 VDD.n7040 166.238
R15335 VDD.n7041 VDD.n6961 166.238
R15336 VDD.n7047 VDD.n7044 166.238
R15337 VDD.n7049 VDD.n7044 166.238
R15338 VDD.n7054 VDD.n6953 166.238
R15339 VDD.n7056 VDD.n6953 166.238
R15340 VDD.n7062 VDD.n7061 166.238
R15341 VDD.n7062 VDD.n6945 166.238
R15342 VDD.n7068 VDD.n7065 166.238
R15343 VDD.n7070 VDD.n7065 166.238
R15344 VDD.n7076 VDD.n7075 166.238
R15345 VDD.n7076 VDD.n6936 166.238
R15346 VDD.n7082 VDD.n7079 166.238
R15347 VDD.n7084 VDD.n7079 166.238
R15348 VDD.n7089 VDD.n6928 166.238
R15349 VDD.n7091 VDD.n6928 166.238
R15350 VDD.n7097 VDD.n7096 166.238
R15351 VDD.n7097 VDD.n6920 166.238
R15352 VDD.n7103 VDD.n7100 166.238
R15353 VDD.n7105 VDD.n7100 166.238
R15354 VDD.n7111 VDD.n7110 166.238
R15355 VDD.n7111 VDD.n6911 166.238
R15356 VDD.n7117 VDD.n7114 166.238
R15357 VDD.n7119 VDD.n7114 166.238
R15358 VDD.n7126 VDD.n6892 166.238
R15359 VDD.n7126 VDD.n6891 166.238
R15360 VDD.n6903 VDD.n6898 166.238
R15361 VDD.n6901 VDD.n6898 166.238
R15362 VDD.n6028 VDD.n6024 166.238
R15363 VDD.n6029 VDD.n6028 166.238
R15364 VDD.n6094 VDD.n5949 166.238
R15365 VDD.n6096 VDD.n5949 166.238
R15366 VDD.n6151 VDD.n5888 166.238
R15367 VDD.n6152 VDD.n6151 166.238
R15368 VDD.n6217 VDD.n5813 166.238
R15369 VDD.n6219 VDD.n5813 166.238
R15370 VDD.n6274 VDD.n5752 166.238
R15371 VDD.n6275 VDD.n6274 166.238
R15372 VDD.n6340 VDD.n5677 166.238
R15373 VDD.n6342 VDD.n5677 166.238
R15374 VDD.n6397 VDD.n5616 166.238
R15375 VDD.n6398 VDD.n6397 166.238
R15376 VDD.n6463 VDD.n5541 166.238
R15377 VDD.n6465 VDD.n5541 166.238
R15378 VDD.n6520 VDD.n5480 166.238
R15379 VDD.n6521 VDD.n6520 166.238
R15380 VDD.n6586 VDD.n5405 166.238
R15381 VDD.n6588 VDD.n5405 166.238
R15382 VDD.n6643 VDD.n5344 166.238
R15383 VDD.n6644 VDD.n6643 166.238
R15384 VDD.n6709 VDD.n5269 166.238
R15385 VDD.n6711 VDD.n5269 166.238
R15386 VDD.n6766 VDD.n5208 166.238
R15387 VDD.n6767 VDD.n6766 166.238
R15388 VDD.n6832 VDD.n5133 166.238
R15389 VDD.n6834 VDD.n5133 166.238
R15390 VDD.n5071 VDD.n5070 166.238
R15391 VDD.n5071 VDD.n4816 166.238
R15392 VDD.n5003 VDD.n4890 166.238
R15393 VDD.n5001 VDD.n4890 166.238
R15394 VDD.n4813 VDD.n4812 166.238
R15395 VDD.n4813 VDD.n2038 166.238
R15396 VDD.n4748 VDD.n2119 166.238
R15397 VDD.n4750 VDD.n2119 166.238
R15398 VDD.n4688 VDD.n4687 166.238
R15399 VDD.n4688 VDD.n2174 166.238
R15400 VDD.n4623 VDD.n2255 166.238
R15401 VDD.n4625 VDD.n2255 166.238
R15402 VDD.n4563 VDD.n4562 166.238
R15403 VDD.n4563 VDD.n2310 166.238
R15404 VDD.n4498 VDD.n2391 166.238
R15405 VDD.n4500 VDD.n2391 166.238
R15406 VDD.n4438 VDD.n4437 166.238
R15407 VDD.n4438 VDD.n2446 166.238
R15408 VDD.n4373 VDD.n2527 166.238
R15409 VDD.n4375 VDD.n2527 166.238
R15410 VDD.n4313 VDD.n4312 166.238
R15411 VDD.n4313 VDD.n2582 166.238
R15412 VDD.n4248 VDD.n2663 166.238
R15413 VDD.n4250 VDD.n2663 166.238
R15414 VDD.n4188 VDD.n4187 166.238
R15415 VDD.n4188 VDD.n2718 166.238
R15416 VDD.n4123 VDD.n2799 166.238
R15417 VDD.n4125 VDD.n2799 166.238
R15418 VDD.n4063 VDD.n4062 166.238
R15419 VDD.n4063 VDD.n2854 166.238
R15420 VDD.n3998 VDD.n2935 166.238
R15421 VDD.n4000 VDD.n2935 166.238
R15422 VDD.n3448 VDD.n3447 166.238
R15423 VDD.n3448 VDD.n3343 166.238
R15424 VDD.n3440 VDD.n3439 166.238
R15425 VDD.n3439 VDD.n3350 166.238
R15426 VDD.n3434 VDD.n3433 166.238
R15427 VDD.n3434 VDD.n3423 166.238
R15428 VDD.n3485 VDD.n3484 166.238
R15429 VDD.n3485 VDD.n3452 166.238
R15430 VDD.n3477 VDD.n3476 166.238
R15431 VDD.n3476 VDD.n3459 166.238
R15432 VDD.n3472 VDD.n3471 166.238
R15433 VDD.n3472 VDD.n3461 166.238
R15434 VDD.n3337 VDD.n3336 166.238
R15435 VDD.n3337 VDD.n3326 166.238
R15436 VDD.n3505 VDD.n3325 166.238
R15437 VDD.n3506 VDD.n3505 166.238
R15438 VDD.n3512 VDD.n3511 166.238
R15439 VDD.n3512 VDD.n3316 166.238
R15440 VDD.n3543 VDD.n3542 166.238
R15441 VDD.n3543 VDD.n3306 166.238
R15442 VDD.n3535 VDD.n3534 166.238
R15443 VDD.n3534 VDD.n3313 166.238
R15444 VDD.n3529 VDD.n3528 166.238
R15445 VDD.n3529 VDD.n3518 166.238
R15446 VDD.n3579 VDD.n3578 166.238
R15447 VDD.n3579 VDD.n3546 166.238
R15448 VDD.n3571 VDD.n3570 166.238
R15449 VDD.n3570 VDD.n3553 166.238
R15450 VDD.n3566 VDD.n3565 166.238
R15451 VDD.n3566 VDD.n3555 166.238
R15452 VDD.n3393 VDD.n3392 166.238
R15453 VDD.n3393 VDD.n3382 166.238
R15454 VDD.n3410 VDD.n3381 166.238
R15455 VDD.n3411 VDD.n3410 166.238
R15456 VDD.n3417 VDD.n3416 166.238
R15457 VDD.n3417 VDD.n3372 166.238
R15458 VDD.n3938 VDD.n3937 166.238
R15459 VDD.n3938 VDD.n2990 166.238
R15460 VDD.n3873 VDD.n3761 166.238
R15461 VDD.n3875 VDD.n3761 166.238
R15462 VDD.n3145 VDD.t752 158.988
R15463 VDD.n3161 VDD.t748 158.988
R15464 VDD.n3209 VDD.t758 158.988
R15465 VDD.n3225 VDD.t684 158.988
R15466 VDD.n3106 VDD.t672 158.988
R15467 VDD.n3249 VDD.t696 158.988
R15468 VDD.n3360 VDD.t736 158.988
R15469 VDD.n3626 VDD.t690 158.988
R15470 VDD.n3067 VDD.t754 158.988
R15471 VDD.n3083 VDD.t716 158.988
R15472 VDD.n3654 VDD.t708 158.988
R15473 VDD.n3670 VDD.t738 158.988
R15474 VDD.n3693 VDD.t686 158.988
R15475 VDD.n3125 VDD.t692 158.988
R15476 VDD.n3180 VDD.t732 158.988
R15477 VDD.n3714 VDD.t712 158.988
R15478 VDD VDD.t666 158.581
R15479 VDD.n3173 VDD.t700 158.379
R15480 VDD.n3237 VDD.t722 158.379
R15481 VDD.n3261 VDD.t688 158.379
R15482 VDD.n3638 VDD.t714 158.379
R15483 VDD.n3095 VDD.t668 158.379
R15484 VDD.n3682 VDD.t682 158.379
R15485 VDD.n3705 VDD.t710 158.379
R15486 VDD.n3192 VDD.t670 158.379
R15487 VDD.n3726 VDD.t664 158.379
R15488 VDD.n154 VDD.n153 155.102
R15489 VDD.n168 VDD.n167 155.102
R15490 VDD.n189 VDD.n188 155.102
R15491 VDD.n203 VDD.n202 155.102
R15492 VDD.n224 VDD.n223 155.102
R15493 VDD.n238 VDD.n237 155.102
R15494 VDD.n259 VDD.n258 155.102
R15495 VDD.n273 VDD.n272 155.102
R15496 VDD.n7003 VDD.n7002 155.102
R15497 VDD.n7017 VDD.n7016 155.102
R15498 VDD.n7038 VDD.n7037 155.102
R15499 VDD.n7052 VDD.n7051 155.102
R15500 VDD.n7073 VDD.n7072 155.102
R15501 VDD.n7087 VDD.n7086 155.102
R15502 VDD.n7108 VDD.n7107 155.102
R15503 VDD.n7122 VDD.n7121 155.102
R15504 VDD.n3431 VDD.n3430 155.102
R15505 VDD.n3444 VDD.n3442 155.102
R15506 VDD.n3469 VDD.n3468 155.102
R15507 VDD.n3481 VDD.n3479 155.102
R15508 VDD.n3509 VDD.n3508 155.102
R15509 VDD.n3333 VDD.n3331 155.102
R15510 VDD.n3526 VDD.n3525 155.102
R15511 VDD.n3539 VDD.n3537 155.102
R15512 VDD.n3563 VDD.n3562 155.102
R15513 VDD.n3575 VDD.n3573 155.102
R15514 VDD.n3414 VDD.n3413 155.102
R15515 VDD.n3389 VDD.n3387 155.102
R15516 VDD.n7644 VDD.n7641 153.601
R15517 VDD.n7651 VDD.n7636 153.601
R15518 VDD.n7645 VDD.n7641 153.601
R15519 VDD.n7652 VDD.n7651 153.601
R15520 VDD.n7631 VDD.n7628 153.601
R15521 VDD.n7661 VDD.n7626 153.601
R15522 VDD.n7655 VDD.n7628 153.601
R15523 VDD.n7662 VDD.n7661 153.601
R15524 VDD.n7621 VDD.n7618 153.601
R15525 VDD.n7671 VDD.n7615 153.601
R15526 VDD.n7665 VDD.n7618 153.601
R15527 VDD.n7672 VDD.n7671 153.601
R15528 VDD.n7610 VDD.n7607 153.601
R15529 VDD.n7681 VDD.n7602 153.601
R15530 VDD.n7675 VDD.n7607 153.601
R15531 VDD.n7682 VDD.n7681 153.601
R15532 VDD.n7597 VDD.n7594 153.601
R15533 VDD.n7691 VDD.n7590 153.601
R15534 VDD.n7685 VDD.n7594 153.601
R15535 VDD.n7692 VDD.n7691 153.601
R15536 VDD.n7582 VDD.n7579 153.601
R15537 VDD.n7708 VDD.n7574 153.601
R15538 VDD.n7702 VDD.n7579 153.601
R15539 VDD.n7709 VDD.n7708 153.601
R15540 VDD.n7569 VDD.n7566 153.601
R15541 VDD.n7718 VDD.n7565 153.601
R15542 VDD.n7712 VDD.n7566 153.601
R15543 VDD.n7719 VDD.n7718 153.601
R15544 VDD.n7558 VDD.n4 153.601
R15545 VDD.n7557 VDD.n2 153.601
R15546 VDD.n7726 VDD.n4 153.601
R15547 VDD.n7725 VDD.n2 153.601
R15548 VDD.n7552 VDD.n11 153.601
R15549 VDD.n15 VDD.n12 153.601
R15550 VDD.n7553 VDD.n7552 153.601
R15551 VDD.n7546 VDD.n12 153.601
R15552 VDD.n7542 VDD.n20 153.601
R15553 VDD.n28 VDD.n21 153.601
R15554 VDD.n7543 VDD.n7542 153.601
R15555 VDD.n7536 VDD.n21 153.601
R15556 VDD.n7532 VDD.n33 153.601
R15557 VDD.n38 VDD.n34 153.601
R15558 VDD.n7533 VDD.n7532 153.601
R15559 VDD.n7526 VDD.n34 153.601
R15560 VDD.n1777 VDD.n1774 153.601
R15561 VDD.n1784 VDD.n1769 153.601
R15562 VDD.n1778 VDD.n1774 153.601
R15563 VDD.n1785 VDD.n1784 153.601
R15564 VDD.n1764 VDD.n1761 153.601
R15565 VDD.n1794 VDD.n1759 153.601
R15566 VDD.n1788 VDD.n1761 153.601
R15567 VDD.n1795 VDD.n1794 153.601
R15568 VDD.n1754 VDD.n1751 153.601
R15569 VDD.n1804 VDD.n1748 153.601
R15570 VDD.n1798 VDD.n1751 153.601
R15571 VDD.n1805 VDD.n1804 153.601
R15572 VDD.n1743 VDD.n1740 153.601
R15573 VDD.n1814 VDD.n1735 153.601
R15574 VDD.n1808 VDD.n1740 153.601
R15575 VDD.n1815 VDD.n1814 153.601
R15576 VDD.n1730 VDD.n1727 153.601
R15577 VDD.n1824 VDD.n1723 153.601
R15578 VDD.n1818 VDD.n1727 153.601
R15579 VDD.n1825 VDD.n1824 153.601
R15580 VDD.n1715 VDD.n1712 153.601
R15581 VDD.n1841 VDD.n1707 153.601
R15582 VDD.n1835 VDD.n1712 153.601
R15583 VDD.n1842 VDD.n1841 153.601
R15584 VDD.n1702 VDD.n1699 153.601
R15585 VDD.n1851 VDD.n1697 153.601
R15586 VDD.n1845 VDD.n1699 153.601
R15587 VDD.n1852 VDD.n1851 153.601
R15588 VDD.n1692 VDD.n1689 153.601
R15589 VDD.n1861 VDD.n1686 153.601
R15590 VDD.n1855 VDD.n1689 153.601
R15591 VDD.n1862 VDD.n1861 153.601
R15592 VDD.n1681 VDD.n1678 153.601
R15593 VDD.n1871 VDD.n1673 153.601
R15594 VDD.n1865 VDD.n1678 153.601
R15595 VDD.n1872 VDD.n1871 153.601
R15596 VDD.n1668 VDD.n1665 153.601
R15597 VDD.n1881 VDD.n1663 153.601
R15598 VDD.n1875 VDD.n1665 153.601
R15599 VDD.n1882 VDD.n1881 153.601
R15600 VDD.n1658 VDD.n1655 153.601
R15601 VDD.n1891 VDD.n1652 153.601
R15602 VDD.n1885 VDD.n1655 153.601
R15603 VDD.n1892 VDD.n1891 153.601
R15604 VDD.n1517 VDD.n1514 153.601
R15605 VDD.n1524 VDD.n1509 153.601
R15606 VDD.n1518 VDD.n1514 153.601
R15607 VDD.n1525 VDD.n1524 153.601
R15608 VDD.n1504 VDD.n1501 153.601
R15609 VDD.n1534 VDD.n1499 153.601
R15610 VDD.n1528 VDD.n1501 153.601
R15611 VDD.n1535 VDD.n1534 153.601
R15612 VDD.n1494 VDD.n1491 153.601
R15613 VDD.n1544 VDD.n1488 153.601
R15614 VDD.n1538 VDD.n1491 153.601
R15615 VDD.n1545 VDD.n1544 153.601
R15616 VDD.n1483 VDD.n1480 153.601
R15617 VDD.n1554 VDD.n1475 153.601
R15618 VDD.n1548 VDD.n1480 153.601
R15619 VDD.n1555 VDD.n1554 153.601
R15620 VDD.n1470 VDD.n1467 153.601
R15621 VDD.n1564 VDD.n1463 153.601
R15622 VDD.n1558 VDD.n1467 153.601
R15623 VDD.n1565 VDD.n1564 153.601
R15624 VDD.n1455 VDD.n1452 153.601
R15625 VDD.n1581 VDD.n1447 153.601
R15626 VDD.n1575 VDD.n1452 153.601
R15627 VDD.n1582 VDD.n1581 153.601
R15628 VDD.n1442 VDD.n1439 153.601
R15629 VDD.n1591 VDD.n1437 153.601
R15630 VDD.n1585 VDD.n1439 153.601
R15631 VDD.n1592 VDD.n1591 153.601
R15632 VDD.n1432 VDD.n1429 153.601
R15633 VDD.n1601 VDD.n1426 153.601
R15634 VDD.n1595 VDD.n1429 153.601
R15635 VDD.n1602 VDD.n1601 153.601
R15636 VDD.n1421 VDD.n1418 153.601
R15637 VDD.n1611 VDD.n1413 153.601
R15638 VDD.n1605 VDD.n1418 153.601
R15639 VDD.n1612 VDD.n1611 153.601
R15640 VDD.n1408 VDD.n1405 153.601
R15641 VDD.n1621 VDD.n1403 153.601
R15642 VDD.n1615 VDD.n1405 153.601
R15643 VDD.n1622 VDD.n1621 153.601
R15644 VDD.n1398 VDD.n1395 153.601
R15645 VDD.n1631 VDD.n1392 153.601
R15646 VDD.n1625 VDD.n1395 153.601
R15647 VDD.n1632 VDD.n1631 153.601
R15648 VDD.n1257 VDD.n1254 153.601
R15649 VDD.n1264 VDD.n1249 153.601
R15650 VDD.n1258 VDD.n1254 153.601
R15651 VDD.n1265 VDD.n1264 153.601
R15652 VDD.n1244 VDD.n1241 153.601
R15653 VDD.n1274 VDD.n1239 153.601
R15654 VDD.n1268 VDD.n1241 153.601
R15655 VDD.n1275 VDD.n1274 153.601
R15656 VDD.n1234 VDD.n1231 153.601
R15657 VDD.n1284 VDD.n1228 153.601
R15658 VDD.n1278 VDD.n1231 153.601
R15659 VDD.n1285 VDD.n1284 153.601
R15660 VDD.n1223 VDD.n1220 153.601
R15661 VDD.n1294 VDD.n1215 153.601
R15662 VDD.n1288 VDD.n1220 153.601
R15663 VDD.n1295 VDD.n1294 153.601
R15664 VDD.n1210 VDD.n1207 153.601
R15665 VDD.n1304 VDD.n1203 153.601
R15666 VDD.n1298 VDD.n1207 153.601
R15667 VDD.n1305 VDD.n1304 153.601
R15668 VDD.n1195 VDD.n1192 153.601
R15669 VDD.n1321 VDD.n1187 153.601
R15670 VDD.n1315 VDD.n1192 153.601
R15671 VDD.n1322 VDD.n1321 153.601
R15672 VDD.n1182 VDD.n1179 153.601
R15673 VDD.n1331 VDD.n1177 153.601
R15674 VDD.n1325 VDD.n1179 153.601
R15675 VDD.n1332 VDD.n1331 153.601
R15676 VDD.n1172 VDD.n1169 153.601
R15677 VDD.n1341 VDD.n1166 153.601
R15678 VDD.n1335 VDD.n1169 153.601
R15679 VDD.n1342 VDD.n1341 153.601
R15680 VDD.n1161 VDD.n1158 153.601
R15681 VDD.n1351 VDD.n1153 153.601
R15682 VDD.n1345 VDD.n1158 153.601
R15683 VDD.n1352 VDD.n1351 153.601
R15684 VDD.n1148 VDD.n1145 153.601
R15685 VDD.n1361 VDD.n1143 153.601
R15686 VDD.n1355 VDD.n1145 153.601
R15687 VDD.n1362 VDD.n1361 153.601
R15688 VDD.n1138 VDD.n1135 153.601
R15689 VDD.n1371 VDD.n1132 153.601
R15690 VDD.n1365 VDD.n1135 153.601
R15691 VDD.n1372 VDD.n1371 153.601
R15692 VDD.n997 VDD.n994 153.601
R15693 VDD.n1004 VDD.n989 153.601
R15694 VDD.n998 VDD.n994 153.601
R15695 VDD.n1005 VDD.n1004 153.601
R15696 VDD.n984 VDD.n981 153.601
R15697 VDD.n1014 VDD.n979 153.601
R15698 VDD.n1008 VDD.n981 153.601
R15699 VDD.n1015 VDD.n1014 153.601
R15700 VDD.n974 VDD.n971 153.601
R15701 VDD.n1024 VDD.n968 153.601
R15702 VDD.n1018 VDD.n971 153.601
R15703 VDD.n1025 VDD.n1024 153.601
R15704 VDD.n963 VDD.n960 153.601
R15705 VDD.n1034 VDD.n955 153.601
R15706 VDD.n1028 VDD.n960 153.601
R15707 VDD.n1035 VDD.n1034 153.601
R15708 VDD.n950 VDD.n947 153.601
R15709 VDD.n1044 VDD.n943 153.601
R15710 VDD.n1038 VDD.n947 153.601
R15711 VDD.n1045 VDD.n1044 153.601
R15712 VDD.n935 VDD.n932 153.601
R15713 VDD.n1061 VDD.n927 153.601
R15714 VDD.n1055 VDD.n932 153.601
R15715 VDD.n1062 VDD.n1061 153.601
R15716 VDD.n922 VDD.n919 153.601
R15717 VDD.n1071 VDD.n917 153.601
R15718 VDD.n1065 VDD.n919 153.601
R15719 VDD.n1072 VDD.n1071 153.601
R15720 VDD.n912 VDD.n909 153.601
R15721 VDD.n1081 VDD.n906 153.601
R15722 VDD.n1075 VDD.n909 153.601
R15723 VDD.n1082 VDD.n1081 153.601
R15724 VDD.n901 VDD.n898 153.601
R15725 VDD.n1091 VDD.n893 153.601
R15726 VDD.n1085 VDD.n898 153.601
R15727 VDD.n1092 VDD.n1091 153.601
R15728 VDD.n888 VDD.n885 153.601
R15729 VDD.n1101 VDD.n883 153.601
R15730 VDD.n1095 VDD.n885 153.601
R15731 VDD.n1102 VDD.n1101 153.601
R15732 VDD.n878 VDD.n875 153.601
R15733 VDD.n1111 VDD.n872 153.601
R15734 VDD.n1105 VDD.n875 153.601
R15735 VDD.n1112 VDD.n1111 153.601
R15736 VDD.n737 VDD.n734 153.601
R15737 VDD.n744 VDD.n729 153.601
R15738 VDD.n738 VDD.n734 153.601
R15739 VDD.n745 VDD.n744 153.601
R15740 VDD.n724 VDD.n721 153.601
R15741 VDD.n754 VDD.n719 153.601
R15742 VDD.n748 VDD.n721 153.601
R15743 VDD.n755 VDD.n754 153.601
R15744 VDD.n714 VDD.n711 153.601
R15745 VDD.n764 VDD.n708 153.601
R15746 VDD.n758 VDD.n711 153.601
R15747 VDD.n765 VDD.n764 153.601
R15748 VDD.n703 VDD.n700 153.601
R15749 VDD.n774 VDD.n695 153.601
R15750 VDD.n768 VDD.n700 153.601
R15751 VDD.n775 VDD.n774 153.601
R15752 VDD.n690 VDD.n687 153.601
R15753 VDD.n784 VDD.n683 153.601
R15754 VDD.n778 VDD.n687 153.601
R15755 VDD.n785 VDD.n784 153.601
R15756 VDD.n675 VDD.n672 153.601
R15757 VDD.n801 VDD.n667 153.601
R15758 VDD.n795 VDD.n672 153.601
R15759 VDD.n802 VDD.n801 153.601
R15760 VDD.n662 VDD.n659 153.601
R15761 VDD.n811 VDD.n657 153.601
R15762 VDD.n805 VDD.n659 153.601
R15763 VDD.n812 VDD.n811 153.601
R15764 VDD.n652 VDD.n649 153.601
R15765 VDD.n821 VDD.n646 153.601
R15766 VDD.n815 VDD.n649 153.601
R15767 VDD.n822 VDD.n821 153.601
R15768 VDD.n641 VDD.n638 153.601
R15769 VDD.n831 VDD.n633 153.601
R15770 VDD.n825 VDD.n638 153.601
R15771 VDD.n832 VDD.n831 153.601
R15772 VDD.n628 VDD.n625 153.601
R15773 VDD.n841 VDD.n623 153.601
R15774 VDD.n835 VDD.n625 153.601
R15775 VDD.n842 VDD.n841 153.601
R15776 VDD.n618 VDD.n615 153.601
R15777 VDD.n851 VDD.n612 153.601
R15778 VDD.n845 VDD.n615 153.601
R15779 VDD.n852 VDD.n851 153.601
R15780 VDD.n477 VDD.n474 153.601
R15781 VDD.n484 VDD.n469 153.601
R15782 VDD.n478 VDD.n474 153.601
R15783 VDD.n485 VDD.n484 153.601
R15784 VDD.n464 VDD.n461 153.601
R15785 VDD.n494 VDD.n459 153.601
R15786 VDD.n488 VDD.n461 153.601
R15787 VDD.n495 VDD.n494 153.601
R15788 VDD.n454 VDD.n451 153.601
R15789 VDD.n504 VDD.n448 153.601
R15790 VDD.n498 VDD.n451 153.601
R15791 VDD.n505 VDD.n504 153.601
R15792 VDD.n443 VDD.n440 153.601
R15793 VDD.n514 VDD.n435 153.601
R15794 VDD.n508 VDD.n440 153.601
R15795 VDD.n515 VDD.n514 153.601
R15796 VDD.n430 VDD.n427 153.601
R15797 VDD.n524 VDD.n423 153.601
R15798 VDD.n518 VDD.n427 153.601
R15799 VDD.n525 VDD.n524 153.601
R15800 VDD.n415 VDD.n412 153.601
R15801 VDD.n541 VDD.n407 153.601
R15802 VDD.n535 VDD.n412 153.601
R15803 VDD.n542 VDD.n541 153.601
R15804 VDD.n402 VDD.n399 153.601
R15805 VDD.n551 VDD.n397 153.601
R15806 VDD.n545 VDD.n399 153.601
R15807 VDD.n552 VDD.n551 153.601
R15808 VDD.n392 VDD.n389 153.601
R15809 VDD.n561 VDD.n386 153.601
R15810 VDD.n555 VDD.n389 153.601
R15811 VDD.n562 VDD.n561 153.601
R15812 VDD.n381 VDD.n378 153.601
R15813 VDD.n571 VDD.n373 153.601
R15814 VDD.n565 VDD.n378 153.601
R15815 VDD.n572 VDD.n571 153.601
R15816 VDD.n368 VDD.n365 153.601
R15817 VDD.n581 VDD.n363 153.601
R15818 VDD.n575 VDD.n365 153.601
R15819 VDD.n582 VDD.n581 153.601
R15820 VDD.n358 VDD.n355 153.601
R15821 VDD.n591 VDD.n352 153.601
R15822 VDD.n585 VDD.n355 153.601
R15823 VDD.n592 VDD.n591 153.601
R15824 VDD.n7393 VDD.n7390 153.601
R15825 VDD.n7400 VDD.n7385 153.601
R15826 VDD.n7394 VDD.n7390 153.601
R15827 VDD.n7401 VDD.n7400 153.601
R15828 VDD.n7380 VDD.n7377 153.601
R15829 VDD.n7410 VDD.n7375 153.601
R15830 VDD.n7404 VDD.n7377 153.601
R15831 VDD.n7411 VDD.n7410 153.601
R15832 VDD.n7370 VDD.n7367 153.601
R15833 VDD.n7420 VDD.n7364 153.601
R15834 VDD.n7414 VDD.n7367 153.601
R15835 VDD.n7421 VDD.n7420 153.601
R15836 VDD.n7359 VDD.n7356 153.601
R15837 VDD.n7430 VDD.n7351 153.601
R15838 VDD.n7424 VDD.n7356 153.601
R15839 VDD.n7431 VDD.n7430 153.601
R15840 VDD.n7346 VDD.n7343 153.601
R15841 VDD.n7440 VDD.n7339 153.601
R15842 VDD.n7434 VDD.n7343 153.601
R15843 VDD.n7441 VDD.n7440 153.601
R15844 VDD.n7331 VDD.n7328 153.601
R15845 VDD.n7457 VDD.n7323 153.601
R15846 VDD.n7451 VDD.n7328 153.601
R15847 VDD.n7458 VDD.n7457 153.601
R15848 VDD.n7318 VDD.n7315 153.601
R15849 VDD.n7467 VDD.n7313 153.601
R15850 VDD.n7461 VDD.n7315 153.601
R15851 VDD.n7468 VDD.n7467 153.601
R15852 VDD.n7308 VDD.n7305 153.601
R15853 VDD.n7477 VDD.n7302 153.601
R15854 VDD.n7471 VDD.n7305 153.601
R15855 VDD.n7478 VDD.n7477 153.601
R15856 VDD.n7297 VDD.n7294 153.601
R15857 VDD.n7487 VDD.n7289 153.601
R15858 VDD.n7481 VDD.n7294 153.601
R15859 VDD.n7488 VDD.n7487 153.601
R15860 VDD.n7284 VDD.n7281 153.601
R15861 VDD.n7497 VDD.n7279 153.601
R15862 VDD.n7491 VDD.n7281 153.601
R15863 VDD.n7498 VDD.n7497 153.601
R15864 VDD.n7274 VDD.n7271 153.601
R15865 VDD.n7507 VDD.n7268 153.601
R15866 VDD.n7501 VDD.n7271 153.601
R15867 VDD.n7508 VDD.n7507 153.601
R15868 VDD.n7136 VDD.n7133 153.601
R15869 VDD.n7143 VDD.n2034 153.601
R15870 VDD.n7137 VDD.n7133 153.601
R15871 VDD.n7144 VDD.n7143 153.601
R15872 VDD.n2029 VDD.n2026 153.601
R15873 VDD.n7153 VDD.n2024 153.601
R15874 VDD.n7147 VDD.n2026 153.601
R15875 VDD.n7154 VDD.n7153 153.601
R15876 VDD.n2019 VDD.n2016 153.601
R15877 VDD.n7163 VDD.n2013 153.601
R15878 VDD.n7157 VDD.n2016 153.601
R15879 VDD.n7164 VDD.n7163 153.601
R15880 VDD.n2008 VDD.n2005 153.601
R15881 VDD.n7173 VDD.n2000 153.601
R15882 VDD.n7167 VDD.n2005 153.601
R15883 VDD.n7174 VDD.n7173 153.601
R15884 VDD.n1995 VDD.n1992 153.601
R15885 VDD.n7183 VDD.n1988 153.601
R15886 VDD.n7177 VDD.n1992 153.601
R15887 VDD.n7184 VDD.n7183 153.601
R15888 VDD.n1978 VDD.n1966 153.601
R15889 VDD.n1977 VDD.n1964 153.601
R15890 VDD.n7198 VDD.n1966 153.601
R15891 VDD.n7197 VDD.n1964 153.601
R15892 VDD.n1971 VDD.n1959 153.601
R15893 VDD.n7207 VDD.n1958 153.601
R15894 VDD.n1953 VDD.n1950 153.601
R15895 VDD.n7217 VDD.n1946 153.601
R15896 VDD.n7211 VDD.n1950 153.601
R15897 VDD.n7218 VDD.n7217 153.601
R15898 VDD.n1941 VDD.n1938 153.601
R15899 VDD.n7227 VDD.n1933 153.601
R15900 VDD.n7221 VDD.n1938 153.601
R15901 VDD.n7228 VDD.n7227 153.601
R15902 VDD.n1928 VDD.n1925 153.601
R15903 VDD.n7237 VDD.n1923 153.601
R15904 VDD.n7231 VDD.n1925 153.601
R15905 VDD.n7238 VDD.n7237 153.601
R15906 VDD.n1918 VDD.n1915 153.601
R15907 VDD.n7247 VDD.n1912 153.601
R15908 VDD.n7241 VDD.n1915 153.601
R15909 VDD.n7248 VDD.n7247 153.601
R15910 VDD.n1973 VDD.n1959 153.601
R15911 VDD.n7208 VDD.n7207 153.601
R15912 VDD.n6018 VDD.n6015 153.601
R15913 VDD.n6038 VDD.n6013 153.601
R15914 VDD.n6032 VDD.n6015 153.601
R15915 VDD.n6039 VDD.n6038 153.601
R15916 VDD.n6008 VDD.n6005 153.601
R15917 VDD.n6048 VDD.n6000 153.601
R15918 VDD.n6042 VDD.n6005 153.601
R15919 VDD.n6049 VDD.n6048 153.601
R15920 VDD.n5995 VDD.n5992 153.601
R15921 VDD.n6058 VDD.n5989 153.601
R15922 VDD.n6052 VDD.n5992 153.601
R15923 VDD.n6059 VDD.n6058 153.601
R15924 VDD.n5984 VDD.n5981 153.601
R15925 VDD.n6068 VDD.n5979 153.601
R15926 VDD.n6062 VDD.n5981 153.601
R15927 VDD.n6069 VDD.n6068 153.601
R15928 VDD.n5974 VDD.n5971 153.601
R15929 VDD.n6078 VDD.n5966 153.601
R15930 VDD.n6072 VDD.n5971 153.601
R15931 VDD.n6079 VDD.n6078 153.601
R15932 VDD.n5961 VDD.n5958 153.601
R15933 VDD.n6088 VDD.n5954 153.601
R15934 VDD.n6082 VDD.n5958 153.601
R15935 VDD.n6089 VDD.n6088 153.601
R15936 VDD.n5946 VDD.n5943 153.601
R15937 VDD.n6105 VDD.n5938 153.601
R15938 VDD.n6099 VDD.n5943 153.601
R15939 VDD.n6106 VDD.n6105 153.601
R15940 VDD.n5933 VDD.n5930 153.601
R15941 VDD.n6115 VDD.n5927 153.601
R15942 VDD.n6109 VDD.n5930 153.601
R15943 VDD.n6116 VDD.n6115 153.601
R15944 VDD.n5922 VDD.n5919 153.601
R15945 VDD.n6125 VDD.n5917 153.601
R15946 VDD.n6119 VDD.n5919 153.601
R15947 VDD.n6126 VDD.n6125 153.601
R15948 VDD.n5912 VDD.n5909 153.601
R15949 VDD.n6135 VDD.n5907 153.601
R15950 VDD.n6129 VDD.n5909 153.601
R15951 VDD.n6136 VDD.n6135 153.601
R15952 VDD.n5900 VDD.n5895 153.601
R15953 VDD.n5899 VDD.n5893 153.601
R15954 VDD.n6143 VDD.n5895 153.601
R15955 VDD.n6142 VDD.n5893 153.601
R15956 VDD.n5882 VDD.n5879 153.601
R15957 VDD.n6161 VDD.n5877 153.601
R15958 VDD.n6155 VDD.n5879 153.601
R15959 VDD.n6162 VDD.n6161 153.601
R15960 VDD.n5872 VDD.n5869 153.601
R15961 VDD.n6171 VDD.n5864 153.601
R15962 VDD.n6165 VDD.n5869 153.601
R15963 VDD.n6172 VDD.n6171 153.601
R15964 VDD.n5859 VDD.n5856 153.601
R15965 VDD.n6181 VDD.n5853 153.601
R15966 VDD.n6175 VDD.n5856 153.601
R15967 VDD.n6182 VDD.n6181 153.601
R15968 VDD.n5848 VDD.n5845 153.601
R15969 VDD.n6191 VDD.n5843 153.601
R15970 VDD.n6185 VDD.n5845 153.601
R15971 VDD.n6192 VDD.n6191 153.601
R15972 VDD.n5838 VDD.n5835 153.601
R15973 VDD.n6201 VDD.n5830 153.601
R15974 VDD.n6195 VDD.n5835 153.601
R15975 VDD.n6202 VDD.n6201 153.601
R15976 VDD.n5825 VDD.n5822 153.601
R15977 VDD.n6211 VDD.n5818 153.601
R15978 VDD.n6205 VDD.n5822 153.601
R15979 VDD.n6212 VDD.n6211 153.601
R15980 VDD.n5810 VDD.n5807 153.601
R15981 VDD.n6228 VDD.n5802 153.601
R15982 VDD.n6222 VDD.n5807 153.601
R15983 VDD.n6229 VDD.n6228 153.601
R15984 VDD.n5797 VDD.n5794 153.601
R15985 VDD.n6238 VDD.n5791 153.601
R15986 VDD.n6232 VDD.n5794 153.601
R15987 VDD.n6239 VDD.n6238 153.601
R15988 VDD.n5786 VDD.n5783 153.601
R15989 VDD.n6248 VDD.n5781 153.601
R15990 VDD.n6242 VDD.n5783 153.601
R15991 VDD.n6249 VDD.n6248 153.601
R15992 VDD.n5776 VDD.n5773 153.601
R15993 VDD.n6258 VDD.n5771 153.601
R15994 VDD.n6252 VDD.n5773 153.601
R15995 VDD.n6259 VDD.n6258 153.601
R15996 VDD.n5764 VDD.n5759 153.601
R15997 VDD.n5763 VDD.n5757 153.601
R15998 VDD.n6266 VDD.n5759 153.601
R15999 VDD.n6265 VDD.n5757 153.601
R16000 VDD.n5746 VDD.n5743 153.601
R16001 VDD.n6284 VDD.n5741 153.601
R16002 VDD.n6278 VDD.n5743 153.601
R16003 VDD.n6285 VDD.n6284 153.601
R16004 VDD.n5736 VDD.n5733 153.601
R16005 VDD.n6294 VDD.n5728 153.601
R16006 VDD.n6288 VDD.n5733 153.601
R16007 VDD.n6295 VDD.n6294 153.601
R16008 VDD.n5723 VDD.n5720 153.601
R16009 VDD.n6304 VDD.n5717 153.601
R16010 VDD.n6298 VDD.n5720 153.601
R16011 VDD.n6305 VDD.n6304 153.601
R16012 VDD.n5712 VDD.n5709 153.601
R16013 VDD.n6314 VDD.n5707 153.601
R16014 VDD.n6308 VDD.n5709 153.601
R16015 VDD.n6315 VDD.n6314 153.601
R16016 VDD.n5702 VDD.n5699 153.601
R16017 VDD.n6324 VDD.n5694 153.601
R16018 VDD.n6318 VDD.n5699 153.601
R16019 VDD.n6325 VDD.n6324 153.601
R16020 VDD.n5689 VDD.n5686 153.601
R16021 VDD.n6334 VDD.n5682 153.601
R16022 VDD.n6328 VDD.n5686 153.601
R16023 VDD.n6335 VDD.n6334 153.601
R16024 VDD.n5674 VDD.n5671 153.601
R16025 VDD.n6351 VDD.n5666 153.601
R16026 VDD.n6345 VDD.n5671 153.601
R16027 VDD.n6352 VDD.n6351 153.601
R16028 VDD.n5661 VDD.n5658 153.601
R16029 VDD.n6361 VDD.n5655 153.601
R16030 VDD.n6355 VDD.n5658 153.601
R16031 VDD.n6362 VDD.n6361 153.601
R16032 VDD.n5650 VDD.n5647 153.601
R16033 VDD.n6371 VDD.n5645 153.601
R16034 VDD.n6365 VDD.n5647 153.601
R16035 VDD.n6372 VDD.n6371 153.601
R16036 VDD.n5640 VDD.n5637 153.601
R16037 VDD.n6381 VDD.n5635 153.601
R16038 VDD.n6375 VDD.n5637 153.601
R16039 VDD.n6382 VDD.n6381 153.601
R16040 VDD.n5628 VDD.n5623 153.601
R16041 VDD.n5627 VDD.n5621 153.601
R16042 VDD.n6389 VDD.n5623 153.601
R16043 VDD.n6388 VDD.n5621 153.601
R16044 VDD.n5610 VDD.n5607 153.601
R16045 VDD.n6407 VDD.n5605 153.601
R16046 VDD.n6401 VDD.n5607 153.601
R16047 VDD.n6408 VDD.n6407 153.601
R16048 VDD.n5600 VDD.n5597 153.601
R16049 VDD.n6417 VDD.n5592 153.601
R16050 VDD.n6411 VDD.n5597 153.601
R16051 VDD.n6418 VDD.n6417 153.601
R16052 VDD.n5587 VDD.n5584 153.601
R16053 VDD.n6427 VDD.n5581 153.601
R16054 VDD.n6421 VDD.n5584 153.601
R16055 VDD.n6428 VDD.n6427 153.601
R16056 VDD.n5576 VDD.n5573 153.601
R16057 VDD.n6437 VDD.n5571 153.601
R16058 VDD.n6431 VDD.n5573 153.601
R16059 VDD.n6438 VDD.n6437 153.601
R16060 VDD.n5566 VDD.n5563 153.601
R16061 VDD.n6447 VDD.n5558 153.601
R16062 VDD.n6441 VDD.n5563 153.601
R16063 VDD.n6448 VDD.n6447 153.601
R16064 VDD.n5553 VDD.n5550 153.601
R16065 VDD.n6457 VDD.n5546 153.601
R16066 VDD.n6451 VDD.n5550 153.601
R16067 VDD.n6458 VDD.n6457 153.601
R16068 VDD.n5538 VDD.n5535 153.601
R16069 VDD.n6474 VDD.n5530 153.601
R16070 VDD.n6468 VDD.n5535 153.601
R16071 VDD.n6475 VDD.n6474 153.601
R16072 VDD.n5525 VDD.n5522 153.601
R16073 VDD.n6484 VDD.n5519 153.601
R16074 VDD.n6478 VDD.n5522 153.601
R16075 VDD.n6485 VDD.n6484 153.601
R16076 VDD.n5514 VDD.n5511 153.601
R16077 VDD.n6494 VDD.n5509 153.601
R16078 VDD.n6488 VDD.n5511 153.601
R16079 VDD.n6495 VDD.n6494 153.601
R16080 VDD.n5504 VDD.n5501 153.601
R16081 VDD.n6504 VDD.n5499 153.601
R16082 VDD.n6498 VDD.n5501 153.601
R16083 VDD.n6505 VDD.n6504 153.601
R16084 VDD.n5492 VDD.n5487 153.601
R16085 VDD.n5491 VDD.n5485 153.601
R16086 VDD.n6512 VDD.n5487 153.601
R16087 VDD.n6511 VDD.n5485 153.601
R16088 VDD.n5474 VDD.n5471 153.601
R16089 VDD.n6530 VDD.n5469 153.601
R16090 VDD.n6524 VDD.n5471 153.601
R16091 VDD.n6531 VDD.n6530 153.601
R16092 VDD.n5464 VDD.n5461 153.601
R16093 VDD.n6540 VDD.n5456 153.601
R16094 VDD.n6534 VDD.n5461 153.601
R16095 VDD.n6541 VDD.n6540 153.601
R16096 VDD.n5451 VDD.n5448 153.601
R16097 VDD.n6550 VDD.n5445 153.601
R16098 VDD.n6544 VDD.n5448 153.601
R16099 VDD.n6551 VDD.n6550 153.601
R16100 VDD.n5440 VDD.n5437 153.601
R16101 VDD.n6560 VDD.n5435 153.601
R16102 VDD.n6554 VDD.n5437 153.601
R16103 VDD.n6561 VDD.n6560 153.601
R16104 VDD.n5430 VDD.n5427 153.601
R16105 VDD.n6570 VDD.n5422 153.601
R16106 VDD.n6564 VDD.n5427 153.601
R16107 VDD.n6571 VDD.n6570 153.601
R16108 VDD.n5417 VDD.n5414 153.601
R16109 VDD.n6580 VDD.n5410 153.601
R16110 VDD.n6574 VDD.n5414 153.601
R16111 VDD.n6581 VDD.n6580 153.601
R16112 VDD.n5402 VDD.n5399 153.601
R16113 VDD.n6597 VDD.n5394 153.601
R16114 VDD.n6591 VDD.n5399 153.601
R16115 VDD.n6598 VDD.n6597 153.601
R16116 VDD.n5389 VDD.n5386 153.601
R16117 VDD.n6607 VDD.n5383 153.601
R16118 VDD.n6601 VDD.n5386 153.601
R16119 VDD.n6608 VDD.n6607 153.601
R16120 VDD.n5378 VDD.n5375 153.601
R16121 VDD.n6617 VDD.n5373 153.601
R16122 VDD.n6611 VDD.n5375 153.601
R16123 VDD.n6618 VDD.n6617 153.601
R16124 VDD.n5368 VDD.n5365 153.601
R16125 VDD.n6627 VDD.n5363 153.601
R16126 VDD.n6621 VDD.n5365 153.601
R16127 VDD.n6628 VDD.n6627 153.601
R16128 VDD.n5356 VDD.n5351 153.601
R16129 VDD.n5355 VDD.n5349 153.601
R16130 VDD.n6635 VDD.n5351 153.601
R16131 VDD.n6634 VDD.n5349 153.601
R16132 VDD.n5338 VDD.n5335 153.601
R16133 VDD.n6653 VDD.n5333 153.601
R16134 VDD.n6647 VDD.n5335 153.601
R16135 VDD.n6654 VDD.n6653 153.601
R16136 VDD.n5328 VDD.n5325 153.601
R16137 VDD.n6663 VDD.n5320 153.601
R16138 VDD.n6657 VDD.n5325 153.601
R16139 VDD.n6664 VDD.n6663 153.601
R16140 VDD.n5315 VDD.n5312 153.601
R16141 VDD.n6673 VDD.n5309 153.601
R16142 VDD.n6667 VDD.n5312 153.601
R16143 VDD.n6674 VDD.n6673 153.601
R16144 VDD.n5304 VDD.n5301 153.601
R16145 VDD.n6683 VDD.n5299 153.601
R16146 VDD.n6677 VDD.n5301 153.601
R16147 VDD.n6684 VDD.n6683 153.601
R16148 VDD.n5294 VDD.n5291 153.601
R16149 VDD.n6693 VDD.n5286 153.601
R16150 VDD.n6687 VDD.n5291 153.601
R16151 VDD.n6694 VDD.n6693 153.601
R16152 VDD.n5281 VDD.n5278 153.601
R16153 VDD.n6703 VDD.n5274 153.601
R16154 VDD.n6697 VDD.n5278 153.601
R16155 VDD.n6704 VDD.n6703 153.601
R16156 VDD.n5266 VDD.n5263 153.601
R16157 VDD.n6720 VDD.n5258 153.601
R16158 VDD.n6714 VDD.n5263 153.601
R16159 VDD.n6721 VDD.n6720 153.601
R16160 VDD.n5253 VDD.n5250 153.601
R16161 VDD.n6730 VDD.n5247 153.601
R16162 VDD.n6724 VDD.n5250 153.601
R16163 VDD.n6731 VDD.n6730 153.601
R16164 VDD.n5242 VDD.n5239 153.601
R16165 VDD.n6740 VDD.n5237 153.601
R16166 VDD.n6734 VDD.n5239 153.601
R16167 VDD.n6741 VDD.n6740 153.601
R16168 VDD.n5232 VDD.n5229 153.601
R16169 VDD.n6750 VDD.n5227 153.601
R16170 VDD.n6744 VDD.n5229 153.601
R16171 VDD.n6751 VDD.n6750 153.601
R16172 VDD.n5220 VDD.n5215 153.601
R16173 VDD.n5219 VDD.n5213 153.601
R16174 VDD.n6758 VDD.n5215 153.601
R16175 VDD.n6757 VDD.n5213 153.601
R16176 VDD.n5202 VDD.n5199 153.601
R16177 VDD.n6776 VDD.n5197 153.601
R16178 VDD.n6770 VDD.n5199 153.601
R16179 VDD.n6777 VDD.n6776 153.601
R16180 VDD.n5192 VDD.n5189 153.601
R16181 VDD.n6786 VDD.n5184 153.601
R16182 VDD.n6780 VDD.n5189 153.601
R16183 VDD.n6787 VDD.n6786 153.601
R16184 VDD.n5179 VDD.n5176 153.601
R16185 VDD.n6796 VDD.n5173 153.601
R16186 VDD.n6790 VDD.n5176 153.601
R16187 VDD.n6797 VDD.n6796 153.601
R16188 VDD.n5168 VDD.n5165 153.601
R16189 VDD.n6806 VDD.n5163 153.601
R16190 VDD.n6800 VDD.n5165 153.601
R16191 VDD.n6807 VDD.n6806 153.601
R16192 VDD.n5158 VDD.n5155 153.601
R16193 VDD.n6816 VDD.n5150 153.601
R16194 VDD.n6810 VDD.n5155 153.601
R16195 VDD.n6817 VDD.n6816 153.601
R16196 VDD.n5145 VDD.n5142 153.601
R16197 VDD.n6826 VDD.n5138 153.601
R16198 VDD.n6820 VDD.n5142 153.601
R16199 VDD.n6827 VDD.n6826 153.601
R16200 VDD.n5130 VDD.n5127 153.601
R16201 VDD.n6843 VDD.n5122 153.601
R16202 VDD.n6837 VDD.n5127 153.601
R16203 VDD.n6844 VDD.n6843 153.601
R16204 VDD.n5117 VDD.n5114 153.601
R16205 VDD.n6853 VDD.n5111 153.601
R16206 VDD.n6847 VDD.n5114 153.601
R16207 VDD.n6854 VDD.n6853 153.601
R16208 VDD.n5106 VDD.n5103 153.601
R16209 VDD.n6863 VDD.n5101 153.601
R16210 VDD.n6857 VDD.n5103 153.601
R16211 VDD.n6864 VDD.n6863 153.601
R16212 VDD.n5096 VDD.n5093 153.601
R16213 VDD.n6873 VDD.n5091 153.601
R16214 VDD.n6867 VDD.n5093 153.601
R16215 VDD.n6874 VDD.n6873 153.601
R16216 VDD.n5084 VDD.n5079 153.601
R16217 VDD.n5083 VDD.n5077 153.601
R16218 VDD.n6881 VDD.n5079 153.601
R16219 VDD.n6880 VDD.n5077 153.601
R16220 VDD.n5062 VDD.n4824 153.601
R16221 VDD.n4830 VDD.n4825 153.601
R16222 VDD.n5063 VDD.n5062 153.601
R16223 VDD.n5056 VDD.n4825 153.601
R16224 VDD.n5052 VDD.n4835 153.601
R16225 VDD.n4840 VDD.n4836 153.601
R16226 VDD.n5053 VDD.n5052 153.601
R16227 VDD.n5046 VDD.n4836 153.601
R16228 VDD.n5042 VDD.n4845 153.601
R16229 VDD.n4853 VDD.n4846 153.601
R16230 VDD.n5043 VDD.n5042 153.601
R16231 VDD.n5036 VDD.n4846 153.601
R16232 VDD.n5032 VDD.n4858 153.601
R16233 VDD.n4864 VDD.n4859 153.601
R16234 VDD.n5033 VDD.n5032 153.601
R16235 VDD.n5026 VDD.n4859 153.601
R16236 VDD.n5022 VDD.n4869 153.601
R16237 VDD.n4874 VDD.n4870 153.601
R16238 VDD.n5023 VDD.n5022 153.601
R16239 VDD.n5016 VDD.n4870 153.601
R16240 VDD.n5012 VDD.n4879 153.601
R16241 VDD.n4887 VDD.n4880 153.601
R16242 VDD.n5013 VDD.n5012 153.601
R16243 VDD.n5006 VDD.n4880 153.601
R16244 VDD.n4995 VDD.n4895 153.601
R16245 VDD.n4902 VDD.n4896 153.601
R16246 VDD.n4996 VDD.n4995 153.601
R16247 VDD.n4989 VDD.n4896 153.601
R16248 VDD.n4985 VDD.n4907 153.601
R16249 VDD.n4915 VDD.n4908 153.601
R16250 VDD.n4986 VDD.n4985 153.601
R16251 VDD.n4979 VDD.n4908 153.601
R16252 VDD.n4975 VDD.n4920 153.601
R16253 VDD.n4926 VDD.n4921 153.601
R16254 VDD.n4976 VDD.n4975 153.601
R16255 VDD.n4969 VDD.n4921 153.601
R16256 VDD.n4965 VDD.n4931 153.601
R16257 VDD.n4936 VDD.n4932 153.601
R16258 VDD.n4966 VDD.n4965 153.601
R16259 VDD.n4959 VDD.n4932 153.601
R16260 VDD.n4955 VDD.n4941 153.601
R16261 VDD.n4945 VDD.n4942 153.601
R16262 VDD.n4956 VDD.n4955 153.601
R16263 VDD.n4946 VDD.n4942 153.601
R16264 VDD.n4695 VDD.n4692 153.601
R16265 VDD.n4702 VDD.n2170 153.601
R16266 VDD.n4696 VDD.n4692 153.601
R16267 VDD.n4703 VDD.n4702 153.601
R16268 VDD.n2165 VDD.n2162 153.601
R16269 VDD.n4712 VDD.n2160 153.601
R16270 VDD.n4706 VDD.n2162 153.601
R16271 VDD.n4713 VDD.n4712 153.601
R16272 VDD.n2155 VDD.n2152 153.601
R16273 VDD.n4722 VDD.n2149 153.601
R16274 VDD.n4716 VDD.n2152 153.601
R16275 VDD.n4723 VDD.n4722 153.601
R16276 VDD.n2144 VDD.n2141 153.601
R16277 VDD.n4732 VDD.n2136 153.601
R16278 VDD.n4726 VDD.n2141 153.601
R16279 VDD.n4733 VDD.n4732 153.601
R16280 VDD.n2131 VDD.n2128 153.601
R16281 VDD.n4742 VDD.n2124 153.601
R16282 VDD.n4736 VDD.n2128 153.601
R16283 VDD.n4743 VDD.n4742 153.601
R16284 VDD.n2114 VDD.n2102 153.601
R16285 VDD.n2113 VDD.n2100 153.601
R16286 VDD.n4757 VDD.n2102 153.601
R16287 VDD.n4756 VDD.n2100 153.601
R16288 VDD.n2107 VDD.n2095 153.601
R16289 VDD.n4766 VDD.n2094 153.601
R16290 VDD.n2089 VDD.n2086 153.601
R16291 VDD.n4776 VDD.n2082 153.601
R16292 VDD.n4770 VDD.n2086 153.601
R16293 VDD.n4777 VDD.n4776 153.601
R16294 VDD.n2077 VDD.n2074 153.601
R16295 VDD.n4786 VDD.n2069 153.601
R16296 VDD.n4780 VDD.n2074 153.601
R16297 VDD.n4787 VDD.n4786 153.601
R16298 VDD.n2064 VDD.n2061 153.601
R16299 VDD.n4796 VDD.n2059 153.601
R16300 VDD.n4790 VDD.n2061 153.601
R16301 VDD.n4797 VDD.n4796 153.601
R16302 VDD.n2054 VDD.n2051 153.601
R16303 VDD.n4806 VDD.n2048 153.601
R16304 VDD.n4800 VDD.n2051 153.601
R16305 VDD.n4807 VDD.n4806 153.601
R16306 VDD.n2109 VDD.n2095 153.601
R16307 VDD.n4767 VDD.n4766 153.601
R16308 VDD.n4570 VDD.n4567 153.601
R16309 VDD.n4577 VDD.n2306 153.601
R16310 VDD.n4571 VDD.n4567 153.601
R16311 VDD.n4578 VDD.n4577 153.601
R16312 VDD.n2301 VDD.n2298 153.601
R16313 VDD.n4587 VDD.n2296 153.601
R16314 VDD.n4581 VDD.n2298 153.601
R16315 VDD.n4588 VDD.n4587 153.601
R16316 VDD.n2291 VDD.n2288 153.601
R16317 VDD.n4597 VDD.n2285 153.601
R16318 VDD.n4591 VDD.n2288 153.601
R16319 VDD.n4598 VDD.n4597 153.601
R16320 VDD.n2280 VDD.n2277 153.601
R16321 VDD.n4607 VDD.n2272 153.601
R16322 VDD.n4601 VDD.n2277 153.601
R16323 VDD.n4608 VDD.n4607 153.601
R16324 VDD.n2267 VDD.n2264 153.601
R16325 VDD.n4617 VDD.n2260 153.601
R16326 VDD.n4611 VDD.n2264 153.601
R16327 VDD.n4618 VDD.n4617 153.601
R16328 VDD.n2250 VDD.n2238 153.601
R16329 VDD.n2249 VDD.n2236 153.601
R16330 VDD.n4632 VDD.n2238 153.601
R16331 VDD.n4631 VDD.n2236 153.601
R16332 VDD.n2243 VDD.n2231 153.601
R16333 VDD.n4641 VDD.n2230 153.601
R16334 VDD.n2225 VDD.n2222 153.601
R16335 VDD.n4651 VDD.n2218 153.601
R16336 VDD.n4645 VDD.n2222 153.601
R16337 VDD.n4652 VDD.n4651 153.601
R16338 VDD.n2213 VDD.n2210 153.601
R16339 VDD.n4661 VDD.n2205 153.601
R16340 VDD.n4655 VDD.n2210 153.601
R16341 VDD.n4662 VDD.n4661 153.601
R16342 VDD.n2200 VDD.n2197 153.601
R16343 VDD.n4671 VDD.n2195 153.601
R16344 VDD.n4665 VDD.n2197 153.601
R16345 VDD.n4672 VDD.n4671 153.601
R16346 VDD.n2190 VDD.n2187 153.601
R16347 VDD.n4681 VDD.n2184 153.601
R16348 VDD.n4675 VDD.n2187 153.601
R16349 VDD.n4682 VDD.n4681 153.601
R16350 VDD.n2245 VDD.n2231 153.601
R16351 VDD.n4642 VDD.n4641 153.601
R16352 VDD.n4445 VDD.n4442 153.601
R16353 VDD.n4452 VDD.n2442 153.601
R16354 VDD.n4446 VDD.n4442 153.601
R16355 VDD.n4453 VDD.n4452 153.601
R16356 VDD.n2437 VDD.n2434 153.601
R16357 VDD.n4462 VDD.n2432 153.601
R16358 VDD.n4456 VDD.n2434 153.601
R16359 VDD.n4463 VDD.n4462 153.601
R16360 VDD.n2427 VDD.n2424 153.601
R16361 VDD.n4472 VDD.n2421 153.601
R16362 VDD.n4466 VDD.n2424 153.601
R16363 VDD.n4473 VDD.n4472 153.601
R16364 VDD.n2416 VDD.n2413 153.601
R16365 VDD.n4482 VDD.n2408 153.601
R16366 VDD.n4476 VDD.n2413 153.601
R16367 VDD.n4483 VDD.n4482 153.601
R16368 VDD.n2403 VDD.n2400 153.601
R16369 VDD.n4492 VDD.n2396 153.601
R16370 VDD.n4486 VDD.n2400 153.601
R16371 VDD.n4493 VDD.n4492 153.601
R16372 VDD.n2386 VDD.n2374 153.601
R16373 VDD.n2385 VDD.n2372 153.601
R16374 VDD.n4507 VDD.n2374 153.601
R16375 VDD.n4506 VDD.n2372 153.601
R16376 VDD.n2379 VDD.n2367 153.601
R16377 VDD.n4516 VDD.n2366 153.601
R16378 VDD.n2361 VDD.n2358 153.601
R16379 VDD.n4526 VDD.n2354 153.601
R16380 VDD.n4520 VDD.n2358 153.601
R16381 VDD.n4527 VDD.n4526 153.601
R16382 VDD.n2349 VDD.n2346 153.601
R16383 VDD.n4536 VDD.n2341 153.601
R16384 VDD.n4530 VDD.n2346 153.601
R16385 VDD.n4537 VDD.n4536 153.601
R16386 VDD.n2336 VDD.n2333 153.601
R16387 VDD.n4546 VDD.n2331 153.601
R16388 VDD.n4540 VDD.n2333 153.601
R16389 VDD.n4547 VDD.n4546 153.601
R16390 VDD.n2326 VDD.n2323 153.601
R16391 VDD.n4556 VDD.n2320 153.601
R16392 VDD.n4550 VDD.n2323 153.601
R16393 VDD.n4557 VDD.n4556 153.601
R16394 VDD.n2381 VDD.n2367 153.601
R16395 VDD.n4517 VDD.n4516 153.601
R16396 VDD.n4320 VDD.n4317 153.601
R16397 VDD.n4327 VDD.n2578 153.601
R16398 VDD.n4321 VDD.n4317 153.601
R16399 VDD.n4328 VDD.n4327 153.601
R16400 VDD.n2573 VDD.n2570 153.601
R16401 VDD.n4337 VDD.n2568 153.601
R16402 VDD.n4331 VDD.n2570 153.601
R16403 VDD.n4338 VDD.n4337 153.601
R16404 VDD.n2563 VDD.n2560 153.601
R16405 VDD.n4347 VDD.n2557 153.601
R16406 VDD.n4341 VDD.n2560 153.601
R16407 VDD.n4348 VDD.n4347 153.601
R16408 VDD.n2552 VDD.n2549 153.601
R16409 VDD.n4357 VDD.n2544 153.601
R16410 VDD.n4351 VDD.n2549 153.601
R16411 VDD.n4358 VDD.n4357 153.601
R16412 VDD.n2539 VDD.n2536 153.601
R16413 VDD.n4367 VDD.n2532 153.601
R16414 VDD.n4361 VDD.n2536 153.601
R16415 VDD.n4368 VDD.n4367 153.601
R16416 VDD.n2522 VDD.n2510 153.601
R16417 VDD.n2521 VDD.n2508 153.601
R16418 VDD.n4382 VDD.n2510 153.601
R16419 VDD.n4381 VDD.n2508 153.601
R16420 VDD.n2515 VDD.n2503 153.601
R16421 VDD.n4391 VDD.n2502 153.601
R16422 VDD.n2497 VDD.n2494 153.601
R16423 VDD.n4401 VDD.n2490 153.601
R16424 VDD.n4395 VDD.n2494 153.601
R16425 VDD.n4402 VDD.n4401 153.601
R16426 VDD.n2485 VDD.n2482 153.601
R16427 VDD.n4411 VDD.n2477 153.601
R16428 VDD.n4405 VDD.n2482 153.601
R16429 VDD.n4412 VDD.n4411 153.601
R16430 VDD.n2472 VDD.n2469 153.601
R16431 VDD.n4421 VDD.n2467 153.601
R16432 VDD.n4415 VDD.n2469 153.601
R16433 VDD.n4422 VDD.n4421 153.601
R16434 VDD.n2462 VDD.n2459 153.601
R16435 VDD.n4431 VDD.n2456 153.601
R16436 VDD.n4425 VDD.n2459 153.601
R16437 VDD.n4432 VDD.n4431 153.601
R16438 VDD.n2517 VDD.n2503 153.601
R16439 VDD.n4392 VDD.n4391 153.601
R16440 VDD.n4195 VDD.n4192 153.601
R16441 VDD.n4202 VDD.n2714 153.601
R16442 VDD.n4196 VDD.n4192 153.601
R16443 VDD.n4203 VDD.n4202 153.601
R16444 VDD.n2709 VDD.n2706 153.601
R16445 VDD.n4212 VDD.n2704 153.601
R16446 VDD.n4206 VDD.n2706 153.601
R16447 VDD.n4213 VDD.n4212 153.601
R16448 VDD.n2699 VDD.n2696 153.601
R16449 VDD.n4222 VDD.n2693 153.601
R16450 VDD.n4216 VDD.n2696 153.601
R16451 VDD.n4223 VDD.n4222 153.601
R16452 VDD.n2688 VDD.n2685 153.601
R16453 VDD.n4232 VDD.n2680 153.601
R16454 VDD.n4226 VDD.n2685 153.601
R16455 VDD.n4233 VDD.n4232 153.601
R16456 VDD.n2675 VDD.n2672 153.601
R16457 VDD.n4242 VDD.n2668 153.601
R16458 VDD.n4236 VDD.n2672 153.601
R16459 VDD.n4243 VDD.n4242 153.601
R16460 VDD.n2658 VDD.n2646 153.601
R16461 VDD.n2657 VDD.n2644 153.601
R16462 VDD.n4257 VDD.n2646 153.601
R16463 VDD.n4256 VDD.n2644 153.601
R16464 VDD.n2651 VDD.n2639 153.601
R16465 VDD.n4266 VDD.n2638 153.601
R16466 VDD.n2633 VDD.n2630 153.601
R16467 VDD.n4276 VDD.n2626 153.601
R16468 VDD.n4270 VDD.n2630 153.601
R16469 VDD.n4277 VDD.n4276 153.601
R16470 VDD.n2621 VDD.n2618 153.601
R16471 VDD.n4286 VDD.n2613 153.601
R16472 VDD.n4280 VDD.n2618 153.601
R16473 VDD.n4287 VDD.n4286 153.601
R16474 VDD.n2608 VDD.n2605 153.601
R16475 VDD.n4296 VDD.n2603 153.601
R16476 VDD.n4290 VDD.n2605 153.601
R16477 VDD.n4297 VDD.n4296 153.601
R16478 VDD.n2598 VDD.n2595 153.601
R16479 VDD.n4306 VDD.n2592 153.601
R16480 VDD.n4300 VDD.n2595 153.601
R16481 VDD.n4307 VDD.n4306 153.601
R16482 VDD.n2653 VDD.n2639 153.601
R16483 VDD.n4267 VDD.n4266 153.601
R16484 VDD.n4070 VDD.n4067 153.601
R16485 VDD.n4077 VDD.n2850 153.601
R16486 VDD.n4071 VDD.n4067 153.601
R16487 VDD.n4078 VDD.n4077 153.601
R16488 VDD.n2845 VDD.n2842 153.601
R16489 VDD.n4087 VDD.n2840 153.601
R16490 VDD.n4081 VDD.n2842 153.601
R16491 VDD.n4088 VDD.n4087 153.601
R16492 VDD.n2835 VDD.n2832 153.601
R16493 VDD.n4097 VDD.n2829 153.601
R16494 VDD.n4091 VDD.n2832 153.601
R16495 VDD.n4098 VDD.n4097 153.601
R16496 VDD.n2824 VDD.n2821 153.601
R16497 VDD.n4107 VDD.n2816 153.601
R16498 VDD.n4101 VDD.n2821 153.601
R16499 VDD.n4108 VDD.n4107 153.601
R16500 VDD.n2811 VDD.n2808 153.601
R16501 VDD.n4117 VDD.n2804 153.601
R16502 VDD.n4111 VDD.n2808 153.601
R16503 VDD.n4118 VDD.n4117 153.601
R16504 VDD.n2794 VDD.n2782 153.601
R16505 VDD.n2793 VDD.n2780 153.601
R16506 VDD.n4132 VDD.n2782 153.601
R16507 VDD.n4131 VDD.n2780 153.601
R16508 VDD.n2787 VDD.n2775 153.601
R16509 VDD.n4141 VDD.n2774 153.601
R16510 VDD.n2769 VDD.n2766 153.601
R16511 VDD.n4151 VDD.n2762 153.601
R16512 VDD.n4145 VDD.n2766 153.601
R16513 VDD.n4152 VDD.n4151 153.601
R16514 VDD.n2757 VDD.n2754 153.601
R16515 VDD.n4161 VDD.n2749 153.601
R16516 VDD.n4155 VDD.n2754 153.601
R16517 VDD.n4162 VDD.n4161 153.601
R16518 VDD.n2744 VDD.n2741 153.601
R16519 VDD.n4171 VDD.n2739 153.601
R16520 VDD.n4165 VDD.n2741 153.601
R16521 VDD.n4172 VDD.n4171 153.601
R16522 VDD.n2734 VDD.n2731 153.601
R16523 VDD.n4181 VDD.n2728 153.601
R16524 VDD.n4175 VDD.n2731 153.601
R16525 VDD.n4182 VDD.n4181 153.601
R16526 VDD.n2789 VDD.n2775 153.601
R16527 VDD.n4142 VDD.n4141 153.601
R16528 VDD.n3945 VDD.n3942 153.601
R16529 VDD.n3952 VDD.n2986 153.601
R16530 VDD.n3946 VDD.n3942 153.601
R16531 VDD.n3953 VDD.n3952 153.601
R16532 VDD.n2981 VDD.n2978 153.601
R16533 VDD.n3962 VDD.n2976 153.601
R16534 VDD.n3956 VDD.n2978 153.601
R16535 VDD.n3963 VDD.n3962 153.601
R16536 VDD.n2971 VDD.n2968 153.601
R16537 VDD.n3972 VDD.n2965 153.601
R16538 VDD.n3966 VDD.n2968 153.601
R16539 VDD.n3973 VDD.n3972 153.601
R16540 VDD.n2960 VDD.n2957 153.601
R16541 VDD.n3982 VDD.n2952 153.601
R16542 VDD.n3976 VDD.n2957 153.601
R16543 VDD.n3983 VDD.n3982 153.601
R16544 VDD.n2947 VDD.n2944 153.601
R16545 VDD.n3992 VDD.n2940 153.601
R16546 VDD.n3986 VDD.n2944 153.601
R16547 VDD.n3993 VDD.n3992 153.601
R16548 VDD.n2930 VDD.n2918 153.601
R16549 VDD.n2929 VDD.n2916 153.601
R16550 VDD.n4007 VDD.n2918 153.601
R16551 VDD.n4006 VDD.n2916 153.601
R16552 VDD.n2923 VDD.n2911 153.601
R16553 VDD.n4016 VDD.n2910 153.601
R16554 VDD.n2905 VDD.n2902 153.601
R16555 VDD.n4026 VDD.n2898 153.601
R16556 VDD.n4020 VDD.n2902 153.601
R16557 VDD.n4027 VDD.n4026 153.601
R16558 VDD.n2893 VDD.n2890 153.601
R16559 VDD.n4036 VDD.n2885 153.601
R16560 VDD.n4030 VDD.n2890 153.601
R16561 VDD.n4037 VDD.n4036 153.601
R16562 VDD.n2880 VDD.n2877 153.601
R16563 VDD.n4046 VDD.n2875 153.601
R16564 VDD.n4040 VDD.n2877 153.601
R16565 VDD.n4047 VDD.n4046 153.601
R16566 VDD.n2870 VDD.n2867 153.601
R16567 VDD.n4056 VDD.n2864 153.601
R16568 VDD.n4050 VDD.n2867 153.601
R16569 VDD.n4057 VDD.n4056 153.601
R16570 VDD.n2925 VDD.n2911 153.601
R16571 VDD.n4017 VDD.n4016 153.601
R16572 VDD.n3294 VDD.n3291 153.601
R16573 VDD.n3594 VDD.n3290 153.601
R16574 VDD.n3285 VDD.n3282 153.601
R16575 VDD.n3604 VDD.n3280 153.601
R16576 VDD.n3598 VDD.n3282 153.601
R16577 VDD.n3605 VDD.n3604 153.601
R16578 VDD.n3273 VDD.n3268 153.601
R16579 VDD.n3272 VDD.n3266 153.601
R16580 VDD.n3612 VDD.n3268 153.601
R16581 VDD.n3611 VDD.n3266 153.601
R16582 VDD.n3295 VDD.n3291 153.601
R16583 VDD.n3595 VDD.n3594 153.601
R16584 VDD.n3820 VDD.n3817 153.601
R16585 VDD.n3827 VDD.n3812 153.601
R16586 VDD.n3821 VDD.n3817 153.601
R16587 VDD.n3828 VDD.n3827 153.601
R16588 VDD.n3807 VDD.n3804 153.601
R16589 VDD.n3837 VDD.n3802 153.601
R16590 VDD.n3831 VDD.n3804 153.601
R16591 VDD.n3838 VDD.n3837 153.601
R16592 VDD.n3797 VDD.n3794 153.601
R16593 VDD.n3847 VDD.n3791 153.601
R16594 VDD.n3841 VDD.n3794 153.601
R16595 VDD.n3848 VDD.n3847 153.601
R16596 VDD.n3786 VDD.n3783 153.601
R16597 VDD.n3857 VDD.n3778 153.601
R16598 VDD.n3851 VDD.n3783 153.601
R16599 VDD.n3858 VDD.n3857 153.601
R16600 VDD.n3773 VDD.n3770 153.601
R16601 VDD.n3867 VDD.n3766 153.601
R16602 VDD.n3861 VDD.n3770 153.601
R16603 VDD.n3868 VDD.n3867 153.601
R16604 VDD.n3756 VDD.n3744 153.601
R16605 VDD.n3755 VDD.n3742 153.601
R16606 VDD.n3882 VDD.n3744 153.601
R16607 VDD.n3881 VDD.n3742 153.601
R16608 VDD.n3749 VDD.n3737 153.601
R16609 VDD.n3891 VDD.n3736 153.601
R16610 VDD.n3731 VDD.n3728 153.601
R16611 VDD.n3901 VDD.n3034 153.601
R16612 VDD.n3895 VDD.n3728 153.601
R16613 VDD.n3902 VDD.n3901 153.601
R16614 VDD.n3029 VDD.n3026 153.601
R16615 VDD.n3911 VDD.n3021 153.601
R16616 VDD.n3905 VDD.n3026 153.601
R16617 VDD.n3912 VDD.n3911 153.601
R16618 VDD.n3016 VDD.n3013 153.601
R16619 VDD.n3921 VDD.n3011 153.601
R16620 VDD.n3915 VDD.n3013 153.601
R16621 VDD.n3922 VDD.n3921 153.601
R16622 VDD.n3006 VDD.n3003 153.601
R16623 VDD.n3931 VDD.n3000 153.601
R16624 VDD.n3925 VDD.n3003 153.601
R16625 VDD.n3932 VDD.n3931 153.601
R16626 VDD.n3751 VDD.n3737 153.601
R16627 VDD.n3892 VDD.n3891 153.601
R16628 VDD.n3147 VDD.t674 150.293
R16629 VDD.n3136 VDD.t706 150.293
R16630 VDD.n3163 VDD.t742 150.293
R16631 VDD.t700 VDD.n3172 150.293
R16632 VDD.n3211 VDD.t680 150.293
R16633 VDD.n3200 VDD.t756 150.293
R16634 VDD.n3227 VDD.t750 150.293
R16635 VDD.t722 VDD.n3236 150.293
R16636 VDD.n3108 VDD.t744 150.293
R16637 VDD.n3097 VDD.t662 150.293
R16638 VDD.n3251 VDD.t702 150.293
R16639 VDD.t688 VDD.n3260 150.293
R16640 VDD.n3362 VDD.t762 150.293
R16641 VDD.n3351 VDD.t734 150.293
R16642 VDD.n3628 VDD.t730 150.293
R16643 VDD.t714 VDD.n3637 150.293
R16644 VDD.n3069 VDD.t720 150.293
R16645 VDD.n3058 VDD.t678 150.293
R16646 VDD.n3085 VDD.t746 150.293
R16647 VDD.t668 VDD.n3094 150.293
R16648 VDD.n3656 VDD.t740 150.293
R16649 VDD.n3645 VDD.t704 150.293
R16650 VDD.n3672 VDD.t698 150.293
R16651 VDD.t682 VDD.n3681 150.293
R16652 VDD.t666 VDD.n3046 150.293
R16653 VDD.n3695 VDD.t724 150.293
R16654 VDD.t710 VDD.n3704 150.293
R16655 VDD.n3127 VDD.t760 150.293
R16656 VDD.n3116 VDD.t676 150.293
R16657 VDD.n3182 VDD.t694 150.293
R16658 VDD.t670 VDD.n3191 150.293
R16659 VDD.n3716 VDD.t718 150.293
R16660 VDD.t664 VDD.n3725 150.293
R16661 VDD.t752 VDD.n3144 150.273
R16662 VDD.t748 VDD.n3160 150.273
R16663 VDD.t758 VDD.n3208 150.273
R16664 VDD.t684 VDD.n3224 150.273
R16665 VDD.t672 VDD.n3105 150.273
R16666 VDD.t696 VDD.n3248 150.273
R16667 VDD.t736 VDD.n3359 150.273
R16668 VDD.t690 VDD.n3625 150.273
R16669 VDD.t754 VDD.n3066 150.273
R16670 VDD.t716 VDD.n3082 150.273
R16671 VDD.t708 VDD.n3653 150.273
R16672 VDD.t738 VDD.n3669 150.273
R16673 VDD.n3051 VDD.t728 150.273
R16674 VDD.n3040 VDD.t726 150.273
R16675 VDD.t686 VDD.n3692 150.273
R16676 VDD.t692 VDD.n3124 150.273
R16677 VDD.t732 VDD.n3179 150.273
R16678 VDD.t712 VDD.n3713 150.273
R16679 VDD.n7528 VDD.n7525 143.812
R16680 VDD.n7556 VDD.n7555 143.812
R16681 VDD.n7704 VDD.n7701 143.812
R16682 VDD.n7695 VDD.n7694 143.812
R16683 VDD.n7677 VDD.n7674 143.812
R16684 VDD.n1895 VDD.n1894 143.812
R16685 VDD.n1867 VDD.n1864 143.812
R16686 VDD.n1837 VDD.n1834 143.812
R16687 VDD.n1828 VDD.n1827 143.812
R16688 VDD.n1810 VDD.n1807 143.812
R16689 VDD.n1635 VDD.n1634 143.812
R16690 VDD.n1607 VDD.n1604 143.812
R16691 VDD.n1577 VDD.n1574 143.812
R16692 VDD.n1568 VDD.n1567 143.812
R16693 VDD.n1550 VDD.n1547 143.812
R16694 VDD.n1375 VDD.n1374 143.812
R16695 VDD.n1347 VDD.n1344 143.812
R16696 VDD.n1317 VDD.n1314 143.812
R16697 VDD.n1308 VDD.n1307 143.812
R16698 VDD.n1290 VDD.n1287 143.812
R16699 VDD.n1115 VDD.n1114 143.812
R16700 VDD.n1087 VDD.n1084 143.812
R16701 VDD.n1057 VDD.n1054 143.812
R16702 VDD.n1048 VDD.n1047 143.812
R16703 VDD.n1030 VDD.n1027 143.812
R16704 VDD.n855 VDD.n854 143.812
R16705 VDD.n827 VDD.n824 143.812
R16706 VDD.n797 VDD.n794 143.812
R16707 VDD.n788 VDD.n787 143.812
R16708 VDD.n770 VDD.n767 143.812
R16709 VDD.n595 VDD.n594 143.812
R16710 VDD.n567 VDD.n564 143.812
R16711 VDD.n537 VDD.n534 143.812
R16712 VDD.n528 VDD.n527 143.812
R16713 VDD.n510 VDD.n507 143.812
R16714 VDD.n7511 VDD.n7510 143.812
R16715 VDD.n7483 VDD.n7480 143.812
R16716 VDD.n7453 VDD.n7450 143.812
R16717 VDD.n7444 VDD.n7443 143.812
R16718 VDD.n7426 VDD.n7423 143.812
R16719 VDD.n7251 VDD.n7250 143.812
R16720 VDD.n7223 VDD.n7220 143.812
R16721 VDD.n7194 VDD.n7193 143.812
R16722 VDD.n7187 VDD.n7186 143.812
R16723 VDD.n7169 VDD.n7166 143.812
R16724 VDD.n6121 VDD.n6118 143.812
R16725 VDD.n6101 VDD.n6098 143.812
R16726 VDD.n6092 VDD.n6091 143.812
R16727 VDD.n6064 VDD.n6061 143.812
R16728 VDD.n6034 VDD.n6031 143.812
R16729 VDD.n6244 VDD.n6241 143.812
R16730 VDD.n6224 VDD.n6221 143.812
R16731 VDD.n6215 VDD.n6214 143.812
R16732 VDD.n6187 VDD.n6184 143.812
R16733 VDD.n6157 VDD.n6154 143.812
R16734 VDD.n6367 VDD.n6364 143.812
R16735 VDD.n6347 VDD.n6344 143.812
R16736 VDD.n6338 VDD.n6337 143.812
R16737 VDD.n6310 VDD.n6307 143.812
R16738 VDD.n6280 VDD.n6277 143.812
R16739 VDD.n6490 VDD.n6487 143.812
R16740 VDD.n6470 VDD.n6467 143.812
R16741 VDD.n6461 VDD.n6460 143.812
R16742 VDD.n6433 VDD.n6430 143.812
R16743 VDD.n6403 VDD.n6400 143.812
R16744 VDD.n6613 VDD.n6610 143.812
R16745 VDD.n6593 VDD.n6590 143.812
R16746 VDD.n6584 VDD.n6583 143.812
R16747 VDD.n6556 VDD.n6553 143.812
R16748 VDD.n6526 VDD.n6523 143.812
R16749 VDD.n6736 VDD.n6733 143.812
R16750 VDD.n6716 VDD.n6713 143.812
R16751 VDD.n6707 VDD.n6706 143.812
R16752 VDD.n6679 VDD.n6676 143.812
R16753 VDD.n6649 VDD.n6646 143.812
R16754 VDD.n6859 VDD.n6856 143.812
R16755 VDD.n6839 VDD.n6836 143.812
R16756 VDD.n6830 VDD.n6829 143.812
R16757 VDD.n6802 VDD.n6799 143.812
R16758 VDD.n6772 VDD.n6769 143.812
R16759 VDD.n4981 VDD.n4978 143.812
R16760 VDD.n4999 VDD.n4998 143.812
R16761 VDD.n5008 VDD.n5005 143.812
R16762 VDD.n5038 VDD.n5035 143.812
R16763 VDD.n5067 VDD.n5065 143.812
R16764 VDD.n4810 VDD.n4809 143.812
R16765 VDD.n4782 VDD.n4779 143.812
R16766 VDD.n4753 VDD.n4752 143.812
R16767 VDD.n4746 VDD.n4745 143.812
R16768 VDD.n4728 VDD.n4725 143.812
R16769 VDD.n4685 VDD.n4684 143.812
R16770 VDD.n4657 VDD.n4654 143.812
R16771 VDD.n4628 VDD.n4627 143.812
R16772 VDD.n4621 VDD.n4620 143.812
R16773 VDD.n4603 VDD.n4600 143.812
R16774 VDD.n4560 VDD.n4559 143.812
R16775 VDD.n4532 VDD.n4529 143.812
R16776 VDD.n4503 VDD.n4502 143.812
R16777 VDD.n4496 VDD.n4495 143.812
R16778 VDD.n4478 VDD.n4475 143.812
R16779 VDD.n4435 VDD.n4434 143.812
R16780 VDD.n4407 VDD.n4404 143.812
R16781 VDD.n4378 VDD.n4377 143.812
R16782 VDD.n4371 VDD.n4370 143.812
R16783 VDD.n4353 VDD.n4350 143.812
R16784 VDD.n4310 VDD.n4309 143.812
R16785 VDD.n4282 VDD.n4279 143.812
R16786 VDD.n4253 VDD.n4252 143.812
R16787 VDD.n4246 VDD.n4245 143.812
R16788 VDD.n4228 VDD.n4225 143.812
R16789 VDD.n4185 VDD.n4184 143.812
R16790 VDD.n4157 VDD.n4154 143.812
R16791 VDD.n4128 VDD.n4127 143.812
R16792 VDD.n4121 VDD.n4120 143.812
R16793 VDD.n4103 VDD.n4100 143.812
R16794 VDD.n4060 VDD.n4059 143.812
R16795 VDD.n4032 VDD.n4029 143.812
R16796 VDD.n4003 VDD.n4002 143.812
R16797 VDD.n3996 VDD.n3995 143.812
R16798 VDD.n3978 VDD.n3975 143.812
R16799 VDD.n3935 VDD.n3934 143.812
R16800 VDD.n3907 VDD.n3904 143.812
R16801 VDD.n3878 VDD.n3877 143.812
R16802 VDD.n3871 VDD.n3870 143.812
R16803 VDD.n3853 VDD.n3850 143.812
R16804 VDD.n43 VDD.n42 125.284
R16805 VDD.n1647 VDD.n1646 125.284
R16806 VDD.n1387 VDD.n1386 125.284
R16807 VDD.n1127 VDD.n1126 125.284
R16808 VDD.n867 VDD.n866 125.284
R16809 VDD.n607 VDD.n606 125.284
R16810 VDD.n347 VDD.n346 125.284
R16811 VDD.n7263 VDD.n7262 125.284
R16812 VDD.n1907 VDD.n1906 125.284
R16813 VDD.n6023 VDD.n6022 125.284
R16814 VDD.n5887 VDD.n5886 125.284
R16815 VDD.n5751 VDD.n5750 125.284
R16816 VDD.n5615 VDD.n5614 125.284
R16817 VDD.n5479 VDD.n5478 125.284
R16818 VDD.n5343 VDD.n5342 125.284
R16819 VDD.n5207 VDD.n5206 125.284
R16820 VDD.n5069 VDD.n5068 125.284
R16821 VDD.n2043 VDD.n2042 125.284
R16822 VDD.n2179 VDD.n2178 125.284
R16823 VDD.n2315 VDD.n2314 125.284
R16824 VDD.n2451 VDD.n2450 125.284
R16825 VDD.n2587 VDD.n2586 125.284
R16826 VDD.n2723 VDD.n2722 125.284
R16827 VDD.n2859 VDD.n2858 125.284
R16828 VDD.n2995 VDD.n2994 125.284
R16829 VDD.n7525 VDD.t867 123.344
R16830 VDD.n7528 VDD.t241 123.344
R16831 VDD.n7535 VDD.t241 123.344
R16832 VDD.n7538 VDD.t603 123.344
R16833 VDD.n7545 VDD.t603 123.344
R16834 VDD.n7548 VDD.t830 123.344
R16835 VDD.n7555 VDD.t830 123.344
R16836 VDD.t239 VDD.n7556 123.344
R16837 VDD.t239 VDD.n7722 123.344
R16838 VDD.n7721 VDD.t224 123.344
R16839 VDD.n7714 VDD.t224 123.344
R16840 VDD.n7711 VDD.t578 123.344
R16841 VDD.n7704 VDD.t578 123.344
R16842 VDD.n7701 VDD.t832 123.344
R16843 VDD.n7695 VDD.t832 123.344
R16844 VDD.n7694 VDD.t580 123.344
R16845 VDD.n7687 VDD.t580 123.344
R16846 VDD.n7684 VDD.t405 123.344
R16847 VDD.n7677 VDD.t405 123.344
R16848 VDD.n7674 VDD.t73 123.344
R16849 VDD.n7667 VDD.t73 123.344
R16850 VDD.n7664 VDD.t403 123.344
R16851 VDD.n7657 VDD.t403 123.344
R16852 VDD.n7654 VDD.t856 123.344
R16853 VDD.n7647 VDD.t856 123.344
R16854 VDD.n1895 VDD.t863 123.344
R16855 VDD.n1894 VDD.t243 123.344
R16856 VDD.n1887 VDD.t243 123.344
R16857 VDD.n1884 VDD.t599 123.344
R16858 VDD.n1877 VDD.t599 123.344
R16859 VDD.n1874 VDD.t923 123.344
R16860 VDD.n1867 VDD.t923 123.344
R16861 VDD.n1864 VDD.t358 123.344
R16862 VDD.n1857 VDD.t358 123.344
R16863 VDD.n1854 VDD.t567 123.344
R16864 VDD.n1847 VDD.t567 123.344
R16865 VDD.n1844 VDD.t597 123.344
R16866 VDD.n1837 VDD.t597 123.344
R16867 VDD.n1834 VDD.t925 123.344
R16868 VDD.n1828 VDD.t925 123.344
R16869 VDD.n1827 VDD.t595 123.344
R16870 VDD.n1820 VDD.t595 123.344
R16871 VDD.n1817 VDD.t157 123.344
R16872 VDD.n1810 VDD.t157 123.344
R16873 VDD.n1807 VDD.t27 123.344
R16874 VDD.n1800 VDD.t27 123.344
R16875 VDD.n1797 VDD.t422 123.344
R16876 VDD.n1790 VDD.t422 123.344
R16877 VDD.n1787 VDD.t54 123.344
R16878 VDD.n1780 VDD.t54 123.344
R16879 VDD.n1635 VDD.t609 123.344
R16880 VDD.n1634 VDD.t418 123.344
R16881 VDD.n1627 VDD.t418 123.344
R16882 VDD.n1624 VDD.t806 123.344
R16883 VDD.n1617 VDD.t806 123.344
R16884 VDD.n1614 VDD.t4 123.344
R16885 VDD.n1607 VDD.t4 123.344
R16886 VDD.n1604 VDD.t15 123.344
R16887 VDD.n1597 VDD.t15 123.344
R16888 VDD.n1594 VDD.t93 123.344
R16889 VDD.n1587 VDD.t93 123.344
R16890 VDD.n1584 VDD.t769 123.344
R16891 VDD.n1577 VDD.t769 123.344
R16892 VDD.n1574 VDD.t6 123.344
R16893 VDD.n1568 VDD.t6 123.344
R16894 VDD.n1567 VDD.t771 123.344
R16895 VDD.n1560 VDD.t771 123.344
R16896 VDD.n1557 VDD.t815 123.344
R16897 VDD.n1550 VDD.t815 123.344
R16898 VDD.n1547 VDD.t644 123.344
R16899 VDD.n1540 VDD.t644 123.344
R16900 VDD.n1537 VDD.t298 123.344
R16901 VDD.n1530 VDD.t298 123.344
R16902 VDD.n1527 VDD.t994 123.344
R16903 VDD.n1520 VDD.t994 123.344
R16904 VDD.n1375 VDD.t961 123.344
R16905 VDD.n1374 VDD.t480 123.344
R16906 VDD.n1367 VDD.t480 123.344
R16907 VDD.n1364 VDD.t393 123.344
R16908 VDD.n1357 VDD.t393 123.344
R16909 VDD.n1354 VDD.t101 123.344
R16910 VDD.n1347 VDD.t101 123.344
R16911 VDD.n1344 VDD.t538 123.344
R16912 VDD.n1337 VDD.t538 123.344
R16913 VDD.n1334 VDD.t412 123.344
R16914 VDD.n1327 VDD.t412 123.344
R16915 VDD.n1324 VDD.t778 123.344
R16916 VDD.n1317 VDD.t778 123.344
R16917 VDD.n1314 VDD.t103 123.344
R16918 VDD.n1308 VDD.t103 123.344
R16919 VDD.n1307 VDD.t191 123.344
R16920 VDD.n1300 VDD.t191 123.344
R16921 VDD.n1297 VDD.t178 123.344
R16922 VDD.n1290 VDD.t178 123.344
R16923 VDD.n1287 VDD.t211 123.344
R16924 VDD.n1280 VDD.t211 123.344
R16925 VDD.n1277 VDD.t360 123.344
R16926 VDD.n1270 VDD.t360 123.344
R16927 VDD.n1267 VDD.t114 123.344
R16928 VDD.n1260 VDD.t114 123.344
R16929 VDD.n1115 VDD.t865 123.344
R16930 VDD.n1114 VDD.t247 123.344
R16931 VDD.n1107 VDD.t247 123.344
R16932 VDD.n1104 VDD.t601 123.344
R16933 VDD.n1097 VDD.t601 123.344
R16934 VDD.n1094 VDD.t657 123.344
R16935 VDD.n1087 VDD.t657 123.344
R16936 VDD.n1084 VDD.t642 123.344
R16937 VDD.n1077 VDD.t642 123.344
R16938 VDD.n1074 VDD.t429 123.344
R16939 VDD.n1067 VDD.t429 123.344
R16940 VDD.n1064 VDD.t174 123.344
R16941 VDD.n1057 VDD.t174 123.344
R16942 VDD.n1054 VDD.t659 123.344
R16943 VDD.n1048 VDD.t659 123.344
R16944 VDD.n1047 VDD.t172 123.344
R16945 VDD.n1040 VDD.t172 123.344
R16946 VDD.n1037 VDD.t346 123.344
R16947 VDD.n1030 VDD.t346 123.344
R16948 VDD.n1027 VDD.t9 123.344
R16949 VDD.n1020 VDD.t9 123.344
R16950 VDD.n1017 VDD.t318 123.344
R16951 VDD.n1010 VDD.t318 123.344
R16952 VDD.n1007 VDD.t808 123.344
R16953 VDD.n1000 VDD.t808 123.344
R16954 VDD.n855 VDD.t605 123.344
R16955 VDD.n854 VDD.t353 123.344
R16956 VDD.n847 VDD.t353 123.344
R16957 VDD.n844 VDD.t120 123.344
R16958 VDD.n837 VDD.t120 123.344
R16959 VDD.n834 VDD.t41 123.344
R16960 VDD.n827 VDD.t41 123.344
R16961 VDD.n824 VDD.t384 123.344
R16962 VDD.n817 VDD.t384 123.344
R16963 VDD.n814 VDD.t220 123.344
R16964 VDD.n807 VDD.t220 123.344
R16965 VDD.n804 VDD.t166 123.344
R16966 VDD.n797 VDD.t166 123.344
R16967 VDD.n794 VDD.t43 123.344
R16968 VDD.n788 VDD.t43 123.344
R16969 VDD.n787 VDD.t164 123.344
R16970 VDD.n780 VDD.t164 123.344
R16971 VDD.n777 VDD.t60 123.344
R16972 VDD.n770 VDD.t60 123.344
R16973 VDD.n767 VDD.t356 123.344
R16974 VDD.n760 VDD.t356 123.344
R16975 VDD.n757 VDD.t63 123.344
R16976 VDD.n750 VDD.t63 123.344
R16977 VDD.n747 VDD.t278 123.344
R16978 VDD.n740 VDD.t278 123.344
R16979 VDD.n595 VDD.t963 123.344
R16980 VDD.n594 VDD.t11 123.344
R16981 VDD.n587 VDD.t11 123.344
R16982 VDD.n584 VDD.t333 123.344
R16983 VDD.n577 VDD.t333 123.344
R16984 VDD.n574 VDD.t555 123.344
R16985 VDD.n567 VDD.t555 123.344
R16986 VDD.n564 VDD.t249 123.344
R16987 VDD.n557 VDD.t249 123.344
R16988 VDD.n554 VDD.t75 123.344
R16989 VDD.n547 VDD.t75 123.344
R16990 VDD.n544 VDD.t233 123.344
R16991 VDD.n537 VDD.t233 123.344
R16992 VDD.n534 VDD.t58 123.344
R16993 VDD.n528 VDD.t58 123.344
R16994 VDD.n527 VDD.t204 123.344
R16995 VDD.n520 VDD.t204 123.344
R16996 VDD.n517 VDD.t988 123.344
R16997 VDD.n510 VDD.t988 123.344
R16998 VDD.n507 VDD.t339 123.344
R16999 VDD.n500 VDD.t339 123.344
R17000 VDD.n497 VDD.t335 123.344
R17001 VDD.n490 VDD.t335 123.344
R17002 VDD.n487 VDD.t362 123.344
R17003 VDD.n480 VDD.t362 123.344
R17004 VDD.n7511 VDD.t607 123.344
R17005 VDD.n7510 VDD.t155 123.344
R17006 VDD.n7503 VDD.t155 123.344
R17007 VDD.n7500 VDD.t337 123.344
R17008 VDD.n7493 VDD.t337 123.344
R17009 VDD.n7490 VDD.t911 123.344
R17010 VDD.n7483 VDD.t911 123.344
R17011 VDD.n7480 VDD.t13 123.344
R17012 VDD.n7473 VDD.t13 123.344
R17013 VDD.n7470 VDD.t112 123.344
R17014 VDD.n7463 VDD.t112 123.344
R17015 VDD.n7460 VDD.t948 123.344
R17016 VDD.n7453 VDD.t948 123.344
R17017 VDD.n7450 VDD.t913 123.344
R17018 VDD.n7444 VDD.t913 123.344
R17019 VDD.n7443 VDD.t222 123.344
R17020 VDD.n7436 VDD.t222 123.344
R17021 VDD.n7433 VDD.t48 123.344
R17022 VDD.n7426 VDD.t48 123.344
R17023 VDD.n7423 VDD.t639 123.344
R17024 VDD.n7416 VDD.t639 123.344
R17025 VDD.n7413 VDD.t652 123.344
R17026 VDD.n7406 VDD.t652 123.344
R17027 VDD.n7403 VDD.t544 123.344
R17028 VDD.n7396 VDD.t544 123.344
R17029 VDD.n7251 VDD.t649 123.344
R17030 VDD.n7250 VDD.t439 123.344
R17031 VDD.n7243 VDD.t439 123.344
R17032 VDD.n7240 VDD.t572 123.344
R17033 VDD.n7233 VDD.t572 123.344
R17034 VDD.n7230 VDD.t1020 123.344
R17035 VDD.n7223 VDD.t1020 123.344
R17036 VDD.n7220 VDD.t500 123.344
R17037 VDD.n7213 VDD.t500 123.344
R17038 VDD.n7210 VDD.t149 123.344
R17039 VDD.n1975 VDD.t149 123.344
R17040 VDD.t35 VDD.n1976 123.344
R17041 VDD.t35 VDD.n7194 123.344
R17042 VDD.n7193 VDD.t1074 123.344
R17043 VDD.n7187 VDD.t1074 123.344
R17044 VDD.n7186 VDD.t106 123.344
R17045 VDD.n7179 VDD.t106 123.344
R17046 VDD.n7176 VDD.t29 123.344
R17047 VDD.n7169 VDD.t29 123.344
R17048 VDD.n7166 VDD.t522 123.344
R17049 VDD.n7159 VDD.t522 123.344
R17050 VDD.n7156 VDD.t193 123.344
R17051 VDD.n7149 VDD.t193 123.344
R17052 VDD.n7146 VDD.t546 123.344
R17053 VDD.n7139 VDD.t546 123.344
R17054 VDD.t245 VDD.n5898 123.344
R17055 VDD.t245 VDD.n6139 123.344
R17056 VDD.n6138 VDD.t37 123.344
R17057 VDD.n6131 VDD.t37 123.344
R17058 VDD.n6128 VDD.t530 123.344
R17059 VDD.n6121 VDD.t530 123.344
R17060 VDD.n6118 VDD.t56 123.344
R17061 VDD.n6111 VDD.t56 123.344
R17062 VDD.n6108 VDD.t322 123.344
R17063 VDD.n6101 VDD.t322 123.344
R17064 VDD.n6098 VDD.t1024 123.344
R17065 VDD.n6092 VDD.t1024 123.344
R17066 VDD.n6091 VDD.t324 123.344
R17067 VDD.n6084 VDD.t324 123.344
R17068 VDD.n6081 VDD.t202 123.344
R17069 VDD.n6074 VDD.t202 123.344
R17070 VDD.n6071 VDD.t534 123.344
R17071 VDD.n6064 VDD.t534 123.344
R17072 VDD.n6061 VDD.t1000 123.344
R17073 VDD.n6054 VDD.t1000 123.344
R17074 VDD.n6051 VDD.t185 123.344
R17075 VDD.n6044 VDD.t185 123.344
R17076 VDD.n6041 VDD.t494 123.344
R17077 VDD.n6034 VDD.t494 123.344
R17078 VDD.n6031 VDD.t888 123.344
R17079 VDD.t141 VDD.n5762 123.344
R17080 VDD.t141 VDD.n6262 123.344
R17081 VDD.n6261 VDD.t263 123.344
R17082 VDD.n6254 VDD.t263 123.344
R17083 VDD.n6251 VDD.t435 123.344
R17084 VDD.n6244 VDD.t435 123.344
R17085 VDD.n6241 VDD.t827 123.344
R17086 VDD.n6234 VDD.t827 123.344
R17087 VDD.n6231 VDD.t944 123.344
R17088 VDD.n6224 VDD.t944 123.344
R17089 VDD.n6221 VDD.t1079 123.344
R17090 VDD.n6215 VDD.t1079 123.344
R17091 VDD.n6214 VDD.t632 123.344
R17092 VDD.n6207 VDD.t632 123.344
R17093 VDD.n6204 VDD.t187 123.344
R17094 VDD.n6197 VDD.t187 123.344
R17095 VDD.n6194 VDD.t471 123.344
R17096 VDD.n6187 VDD.t471 123.344
R17097 VDD.n6184 VDD.t1056 123.344
R17098 VDD.n6177 VDD.t1056 123.344
R17099 VDD.n6174 VDD.t341 123.344
R17100 VDD.n6167 VDD.t341 123.344
R17101 VDD.n6164 VDD.t516 123.344
R17102 VDD.n6157 VDD.t516 123.344
R17103 VDD.n6154 VDD.t881 123.344
R17104 VDD.t364 VDD.n5626 123.344
R17105 VDD.t364 VDD.n6385 123.344
R17106 VDD.n6384 VDD.t109 123.344
R17107 VDD.n6377 VDD.t109 123.344
R17108 VDD.n6374 VDD.t506 123.344
R17109 VDD.n6367 VDD.t506 123.344
R17110 VDD.n6364 VDD.t552 123.344
R17111 VDD.n6357 VDD.t552 123.344
R17112 VDD.n6354 VDD.t145 123.344
R17113 VDD.n6347 VDD.t145 123.344
R17114 VDD.n6344 VDD.t1054 123.344
R17115 VDD.n6338 VDD.t1054 123.344
R17116 VDD.n6337 VDD.t147 123.344
R17117 VDD.n6330 VDD.t147 123.344
R17118 VDD.n6327 VDD.t116 123.344
R17119 VDD.n6320 VDD.t116 123.344
R17120 VDD.n6317 VDD.t453 123.344
R17121 VDD.n6310 VDD.t453 123.344
R17122 VDD.n6307 VDD.t1028 123.344
R17123 VDD.n6300 VDD.t1028 123.344
R17124 VDD.n6297 VDD.t368 123.344
R17125 VDD.n6290 VDD.t368 123.344
R17126 VDD.n6287 VDD.t463 123.344
R17127 VDD.n6280 VDD.t463 123.344
R17128 VDD.n6277 VDD.t916 123.344
R17129 VDD.t46 VDD.n5490 123.344
R17130 VDD.t46 VDD.n6508 123.344
R17131 VDD.n6507 VDD.t253 123.344
R17132 VDD.n6500 VDD.t253 123.344
R17133 VDD.n6497 VDD.t459 123.344
R17134 VDD.n6490 VDD.t459 123.344
R17135 VDD.n6487 VDD.t237 123.344
R17136 VDD.n6480 VDD.t237 123.344
R17137 VDD.n6477 VDD.t257 123.344
R17138 VDD.n6470 VDD.t257 123.344
R17139 VDD.n6467 VDD.t1096 123.344
R17140 VDD.n6461 VDD.t1096 123.344
R17141 VDD.n6460 VDD.t135 123.344
R17142 VDD.n6453 VDD.t135 123.344
R17143 VDD.n6450 VDD.t794 123.344
R17144 VDD.n6443 VDD.t794 123.344
R17145 VDD.n6440 VDD.t490 123.344
R17146 VDD.n6433 VDD.t490 123.344
R17147 VDD.n6430 VDD.t1002 123.344
R17148 VDD.n6423 VDD.t1002 123.344
R17149 VDD.n6420 VDD.t871 123.344
R17150 VDD.n6413 VDD.t871 123.344
R17151 VDD.n6410 VDD.t443 123.344
R17152 VDD.n6403 VDD.t443 123.344
R17153 VDD.n6400 VDD.t621 123.344
R17154 VDD.t312 VDD.n5354 123.344
R17155 VDD.t312 VDD.n6631 123.344
R17156 VDD.n6630 VDD.t33 123.344
R17157 VDD.n6623 VDD.t33 123.344
R17158 VDD.n6620 VDD.t492 123.344
R17159 VDD.n6613 VDD.t492 123.344
R17160 VDD.n6610 VDD.t139 123.344
R17161 VDD.n6603 VDD.t139 123.344
R17162 VDD.n6600 VDD.t208 123.344
R17163 VDD.n6593 VDD.t208 123.344
R17164 VDD.n6590 VDD.t1084 123.344
R17165 VDD.n6584 VDD.t1084 123.344
R17166 VDD.n6583 VDD.t280 123.344
R17167 VDD.n6576 VDD.t280 123.344
R17168 VDD.n6573 VDD.t17 123.344
R17169 VDD.n6566 VDD.t17 123.344
R17170 VDD.n6563 VDD.t475 123.344
R17171 VDD.n6556 VDD.t475 123.344
R17172 VDD.n6553 VDD.t1060 123.344
R17173 VDD.n6546 VDD.t1060 123.344
R17174 VDD.n6543 VDD.t425 123.344
R17175 VDD.n6536 VDD.t425 123.344
R17176 VDD.n6533 VDD.t478 123.344
R17177 VDD.n6526 VDD.t478 123.344
R17178 VDD.n6523 VDD.t23 123.344
R17179 VDD.t305 VDD.n5218 123.344
R17180 VDD.t305 VDD.n6754 123.344
R17181 VDD.n6753 VDD.t320 123.344
R17182 VDD.n6746 VDD.t320 123.344
R17183 VDD.n6743 VDD.t482 123.344
R17184 VDD.n6736 VDD.t482 123.344
R17185 VDD.n6733 VDD.t378 123.344
R17186 VDD.n6726 VDD.t378 123.344
R17187 VDD.n6723 VDD.t316 123.344
R17188 VDD.n6716 VDD.t316 123.344
R17189 VDD.n6713 VDD.t1058 123.344
R17190 VDD.n6707 VDD.t1058 123.344
R17191 VDD.n6706 VDD.t314 123.344
R17192 VDD.n6699 VDD.t314 123.344
R17193 VDD.n6696 VDD.t366 123.344
R17194 VDD.n6689 VDD.t366 123.344
R17195 VDD.n6686 VDD.t520 123.344
R17196 VDD.n6679 VDD.t520 123.344
R17197 VDD.n6676 VDD.t1032 123.344
R17198 VDD.n6669 VDD.t1032 123.344
R17199 VDD.n6666 VDD.t835 123.344
R17200 VDD.n6659 VDD.t835 123.344
R17201 VDD.n6656 VDD.t465 123.344
R17202 VDD.n6649 VDD.t465 123.344
R17203 VDD.n6646 VDD.t840 123.344
R17204 VDD.t349 VDD.n5082 123.344
R17205 VDD.t349 VDD.n6877 123.344
R17206 VDD.n6876 VDD.t431 123.344
R17207 VDD.n6869 VDD.t431 123.344
R17208 VDD.n6866 VDD.t433 123.344
R17209 VDD.n6859 VDD.t433 123.344
R17210 VDD.n6856 VDD.t330 123.344
R17211 VDD.n6849 VDD.t330 123.344
R17212 VDD.n6846 VDD.t228 123.344
R17213 VDD.n6839 VDD.t228 123.344
R17214 VDD.n6836 VDD.t1076 123.344
R17215 VDD.n6830 VDD.t1076 123.344
R17216 VDD.n6829 VDD.t226 123.344
R17217 VDD.n6822 VDD.t226 123.344
R17218 VDD.n6819 VDD.t162 123.344
R17219 VDD.n6812 VDD.t162 123.344
R17220 VDD.n6809 VDD.t510 123.344
R17221 VDD.n6802 VDD.t510 123.344
R17222 VDD.n6799 VDD.t1030 123.344
R17223 VDD.n6792 VDD.t1030 123.344
R17224 VDD.n6789 VDD.t390 123.344
R17225 VDD.n6782 VDD.t390 123.344
R17226 VDD.n6779 VDD.t457 123.344
R17227 VDD.n6772 VDD.t457 123.344
R17228 VDD.n6769 VDD.t919 123.344
R17229 VDD.n4948 VDD.t183 123.344
R17230 VDD.n4958 VDD.t183 123.344
R17231 VDD.n4961 VDD.t181 123.344
R17232 VDD.n4968 VDD.t181 123.344
R17233 VDD.n4971 VDD.t512 123.344
R17234 VDD.n4978 VDD.t512 123.344
R17235 VDD.n4981 VDD.t380 123.344
R17236 VDD.n4988 VDD.t380 123.344
R17237 VDD.n4991 VDD.t118 123.344
R17238 VDD.n4998 VDD.t118 123.344
R17239 VDD.n4999 VDD.t1052 123.344
R17240 VDD.n5005 VDD.t1052 123.344
R17241 VDD.n5008 VDD.t84 123.344
R17242 VDD.n5015 VDD.t84 123.344
R17243 VDD.n5018 VDD.t259 123.344
R17244 VDD.n5025 VDD.t259 123.344
R17245 VDD.n5028 VDD.t486 123.344
R17246 VDD.n5035 VDD.t486 123.344
R17247 VDD.n5038 VDD.t1004 123.344
R17248 VDD.n5045 VDD.t1004 123.344
R17249 VDD.n5048 VDD.t289 123.344
R17250 VDD.n5055 VDD.t289 123.344
R17251 VDD.n5058 VDD.t496 123.344
R17252 VDD.n5065 VDD.t496 123.344
R17253 VDD.t574 VDD.n5067 123.344
R17254 VDD.n4810 VDD.t303 123.344
R17255 VDD.n4809 VDD.t461 123.344
R17256 VDD.n4802 VDD.t461 123.344
R17257 VDD.n4799 VDD.t415 123.344
R17258 VDD.n4792 VDD.t415 123.344
R17259 VDD.n4789 VDD.t1016 123.344
R17260 VDD.n4782 VDD.t1016 123.344
R17261 VDD.n4779 VDD.t526 123.344
R17262 VDD.n4772 VDD.t526 123.344
R17263 VDD.n4769 VDD.t261 123.344
R17264 VDD.n2111 VDD.t261 123.344
R17265 VDD.t562 VDD.n2112 123.344
R17266 VDD.t562 VDD.n4753 123.344
R17267 VDD.n4752 VDD.t1068 123.344
R17268 VDD.n4746 VDD.t1068 123.344
R17269 VDD.n4745 VDD.t564 123.344
R17270 VDD.n4738 VDD.t564 123.344
R17271 VDD.n4735 VDD.t848 123.344
R17272 VDD.n4728 VDD.t848 123.344
R17273 VDD.n4725 VDD.t467 123.344
R17274 VDD.n4718 VDD.t467 123.344
R17275 VDD.n4715 VDD.t634 123.344
R17276 VDD.n4708 VDD.t634 123.344
R17277 VDD.n4705 VDD.t548 123.344
R17278 VDD.n4698 VDD.t548 123.344
R17279 VDD.n4685 VDD.t65 123.344
R17280 VDD.n4684 VDD.t498 123.344
R17281 VDD.n4677 VDD.t498 123.344
R17282 VDD.n4674 VDD.t396 123.344
R17283 VDD.n4667 VDD.t396 123.344
R17284 VDD.n4664 VDD.t1042 123.344
R17285 VDD.n4657 VDD.t1042 123.344
R17286 VDD.n4654 VDD.t449 123.344
R17287 VDD.n4647 VDD.t449 123.344
R17288 VDD.n4644 VDD.t133 123.344
R17289 VDD.n2247 VDD.t133 123.344
R17290 VDD.t95 VDD.n2248 123.344
R17291 VDD.t95 VDD.n4628 123.344
R17292 VDD.n4627 VDD.t1082 123.344
R17293 VDD.n4621 VDD.t1082 123.344
R17294 VDD.n4620 VDD.t97 123.344
R17295 VDD.n4613 VDD.t97 123.344
R17296 VDD.n4610 VDD.t143 123.344
R17297 VDD.n4603 VDD.t143 123.344
R17298 VDD.n4600 VDD.t473 123.344
R17299 VDD.n4593 VDD.t473 123.344
R17300 VDD.n4590 VDD.t541 123.344
R17301 VDD.n4583 VDD.t541 123.344
R17302 VDD.n4580 VDD.t788 123.344
R17303 VDD.n4573 VDD.t788 123.344
R17304 VDD.n4560 VDD.t25 123.344
R17305 VDD.n4559 VDD.t508 123.344
R17306 VDD.n4552 VDD.t508 123.344
R17307 VDD.n4549 VDD.t858 123.344
R17308 VDD.n4542 VDD.t858 123.344
R17309 VDD.n4539 VDD.t1050 123.344
R17310 VDD.n4532 VDD.t1050 123.344
R17311 VDD.n4529 VDD.t518 123.344
R17312 VDD.n4522 VDD.t518 123.344
R17313 VDD.n4519 VDD.t266 123.344
R17314 VDD.n2383 VDD.t266 123.344
R17315 VDD.t215 VDD.n2384 123.344
R17316 VDD.t215 VDD.n4503 123.344
R17317 VDD.n4502 VDD.t1010 123.344
R17318 VDD.n4496 VDD.t1010 123.344
R17319 VDD.n4495 VDD.t217 123.344
R17320 VDD.n4488 VDD.t217 123.344
R17321 VDD.n4485 VDD.t91 123.344
R17322 VDD.n4478 VDD.t91 123.344
R17323 VDD.n4475 VDD.t532 123.344
R17324 VDD.n4468 VDD.t532 123.344
R17325 VDD.n4465 VDD.t160 123.344
R17326 VDD.n4458 VDD.t160 123.344
R17327 VDD.n4455 VDD.t590 123.344
R17328 VDD.n4448 VDD.t590 123.344
R17329 VDD.n4435 VDD.t796 123.344
R17330 VDD.n4434 VDD.t504 123.344
R17331 VDD.n4427 VDD.t504 123.344
R17332 VDD.n4424 VDD.t800 123.344
R17333 VDD.n4417 VDD.t800 123.344
R17334 VDD.n4414 VDD.t1048 123.344
R17335 VDD.n4407 VDD.t1048 123.344
R17336 VDD.n4404 VDD.t441 123.344
R17337 VDD.n4397 VDD.t441 123.344
R17338 VDD.n4394 VDD.t328 123.344
R17339 VDD.n2519 VDD.t328 123.344
R17340 VDD.t19 VDD.n2520 123.344
R17341 VDD.t19 VDD.n4378 123.344
R17342 VDD.n4377 VDD.t1038 123.344
R17343 VDD.n4371 VDD.t1038 123.344
R17344 VDD.n4370 VDD.t593 123.344
R17345 VDD.n4363 VDD.t593 123.344
R17346 VDD.n4360 VDD.t199 123.344
R17347 VDD.n4353 VDD.t199 123.344
R17348 VDD.n4350 VDD.t451 123.344
R17349 VDD.n4343 VDD.t451 123.344
R17350 VDD.n4340 VDD.t39 123.344
R17351 VDD.n4333 VDD.t39 123.344
R17352 VDD.n4330 VDD.t69 123.344
R17353 VDD.n4323 VDD.t69 123.344
R17354 VDD.n4310 VDD.t764 123.344
R17355 VDD.n4309 VDD.t536 123.344
R17356 VDD.n4302 VDD.t536 123.344
R17357 VDD.n4299 VDD.t67 123.344
R17358 VDD.n4292 VDD.t67 123.344
R17359 VDD.n4289 VDD.t1022 123.344
R17360 VDD.n4282 VDD.t1022 123.344
R17361 VDD.n4279 VDD.t488 123.344
R17362 VDD.n4272 VDD.t488 123.344
R17363 VDD.n4269 VDD.t31 123.344
R17364 VDD.n2655 VDD.t31 123.344
R17365 VDD.t386 VDD.n2656 123.344
R17366 VDD.t386 VDD.n4253 123.344
R17367 VDD.n4252 VDD.t1062 123.344
R17368 VDD.n4246 VDD.t1062 123.344
R17369 VDD.n4245 VDD.t388 123.344
R17370 VDD.n4238 VDD.t388 123.344
R17371 VDD.n4235 VDD.t344 123.344
R17372 VDD.n4228 VDD.t344 123.344
R17373 VDD.n4225 VDD.t469 123.344
R17374 VDD.n4218 VDD.t469 123.344
R17375 VDD.n4215 VDD.t892 123.344
R17376 VDD.n4208 VDD.t892 123.344
R17377 VDD.n4205 VDD.t2 123.344
R17378 VDD.n4198 VDD.t2 123.344
R17379 VDD.n4185 VDD.t124 123.344
R17380 VDD.n4184 VDD.t455 123.344
R17381 VDD.n4177 VDD.t455 123.344
R17382 VDD.n4174 VDD.t0 123.344
R17383 VDD.n4167 VDD.t0 123.344
R17384 VDD.n4164 VDD.t1018 123.344
R17385 VDD.n4157 VDD.t1018 123.344
R17386 VDD.n4154 VDD.t514 123.344
R17387 VDD.n4147 VDD.t514 123.344
R17388 VDD.n4144 VDD.t373 123.344
R17389 VDD.n2791 VDD.t373 123.344
R17390 VDD.t80 VDD.n2792 123.344
R17391 VDD.t80 VDD.n4128 123.344
R17392 VDD.n4127 VDD.t1006 123.344
R17393 VDD.n4121 VDD.t1006 123.344
R17394 VDD.n4120 VDD.t82 123.344
R17395 VDD.n4113 VDD.t82 123.344
R17396 VDD.n4110 VDD.t168 123.344
R17397 VDD.n4103 VDD.t168 123.344
R17398 VDD.n4100 VDD.t524 123.344
R17399 VDD.n4093 VDD.t524 123.344
R17400 VDD.n4090 VDD.t99 123.344
R17401 VDD.n4083 VDD.t99 123.344
R17402 VDD.n4080 VDD.t292 123.344
R17403 VDD.n4073 VDD.t292 123.344
R17404 VDD.n4060 VDD.t153 123.344
R17405 VDD.n4059 VDD.t502 123.344
R17406 VDD.n4052 VDD.t502 123.344
R17407 VDD.n4049 VDD.t934 123.344
R17408 VDD.n4042 VDD.t934 123.344
R17409 VDD.n4039 VDD.t1045 123.344
R17410 VDD.n4032 VDD.t1045 123.344
R17411 VDD.n4029 VDD.t437 123.344
R17412 VDD.n4022 VDD.t437 123.344
R17413 VDD.n4019 VDD.t821 123.344
R17414 VDD.n2927 VDD.t821 123.344
R17415 VDD.t310 VDD.n2928 123.344
R17416 VDD.t310 VDD.n4003 123.344
R17417 VDD.n4002 VDD.t1034 123.344
R17418 VDD.n3996 VDD.t1034 123.344
R17419 VDD.n3995 VDD.t308 123.344
R17420 VDD.n3988 VDD.t308 123.344
R17421 VDD.n3985 VDD.t196 123.344
R17422 VDD.n3978 VDD.t196 123.344
R17423 VDD.n3975 VDD.t447 123.344
R17424 VDD.n3968 VDD.t447 123.344
R17425 VDD.n3965 VDD.t296 123.344
R17426 VDD.n3958 VDD.t296 123.344
R17427 VDD.n3955 VDD.t626 123.344
R17428 VDD.n3948 VDD.t626 123.344
R17429 VDD.t86 VDD.n3271 123.344
R17430 VDD.t86 VDD.n3608 123.344
R17431 VDD.n3607 VDD.t88 123.344
R17432 VDD.n3600 VDD.t88 123.344
R17433 VDD.n3597 VDD.t21 123.344
R17434 VDD.n3297 VDD.t21 123.344
R17435 VDD.n3935 VDD.t941 123.344
R17436 VDD.n3934 VDD.t528 123.344
R17437 VDD.n3927 VDD.t528 123.344
R17438 VDD.n3924 VDD.t151 123.344
R17439 VDD.n3917 VDD.t151 123.344
R17440 VDD.n3914 VDD.t1014 123.344
R17441 VDD.n3907 VDD.t1014 123.344
R17442 VDD.n3904 VDD.t484 123.344
R17443 VDD.n3897 VDD.t484 123.344
R17444 VDD.n3894 VDD.t51 123.344
R17445 VDD.n3753 VDD.t51 123.344
R17446 VDD.t231 VDD.n3754 123.344
R17447 VDD.t231 VDD.n3878 123.344
R17448 VDD.n3877 VDD.t1091 123.344
R17449 VDD.n3871 VDD.t1091 123.344
R17450 VDD.n3870 VDD.t284 123.344
R17451 VDD.n3863 VDD.t284 123.344
R17452 VDD.n3860 VDD.t558 123.344
R17453 VDD.n3853 VDD.t558 123.344
R17454 VDD.n3850 VDD.t445 123.344
R17455 VDD.n3843 VDD.t445 123.344
R17456 VDD.n3840 VDD.t427 123.344
R17457 VDD.n3833 VDD.t427 123.344
R17458 VDD.n3830 VDD.t235 123.344
R17459 VDD.n3823 VDD.t235 123.344
R17460 VDD.n332 VDD.n331 99.0123
R17461 VDD.n333 VDD.n332 99.0123
R17462 VDD.n7538 VDD.n7535 75.5806
R17463 VDD.n7548 VDD.n7545 75.5806
R17464 VDD.n7722 VDD.n7721 75.5806
R17465 VDD.n7714 VDD.n7711 75.5806
R17466 VDD.n7687 VDD.n7684 75.5806
R17467 VDD.n7667 VDD.n7664 75.5806
R17468 VDD.n7657 VDD.n7654 75.5806
R17469 VDD.n1887 VDD.n1884 75.5806
R17470 VDD.n1877 VDD.n1874 75.5806
R17471 VDD.n1857 VDD.n1854 75.5806
R17472 VDD.n1847 VDD.n1844 75.5806
R17473 VDD.n1820 VDD.n1817 75.5806
R17474 VDD.n1800 VDD.n1797 75.5806
R17475 VDD.n1790 VDD.n1787 75.5806
R17476 VDD.n1627 VDD.n1624 75.5806
R17477 VDD.n1617 VDD.n1614 75.5806
R17478 VDD.n1597 VDD.n1594 75.5806
R17479 VDD.n1587 VDD.n1584 75.5806
R17480 VDD.n1560 VDD.n1557 75.5806
R17481 VDD.n1540 VDD.n1537 75.5806
R17482 VDD.n1530 VDD.n1527 75.5806
R17483 VDD.n1367 VDD.n1364 75.5806
R17484 VDD.n1357 VDD.n1354 75.5806
R17485 VDD.n1337 VDD.n1334 75.5806
R17486 VDD.n1327 VDD.n1324 75.5806
R17487 VDD.n1300 VDD.n1297 75.5806
R17488 VDD.n1280 VDD.n1277 75.5806
R17489 VDD.n1270 VDD.n1267 75.5806
R17490 VDD.n1107 VDD.n1104 75.5806
R17491 VDD.n1097 VDD.n1094 75.5806
R17492 VDD.n1077 VDD.n1074 75.5806
R17493 VDD.n1067 VDD.n1064 75.5806
R17494 VDD.n1040 VDD.n1037 75.5806
R17495 VDD.n1020 VDD.n1017 75.5806
R17496 VDD.n1010 VDD.n1007 75.5806
R17497 VDD.n847 VDD.n844 75.5806
R17498 VDD.n837 VDD.n834 75.5806
R17499 VDD.n817 VDD.n814 75.5806
R17500 VDD.n807 VDD.n804 75.5806
R17501 VDD.n780 VDD.n777 75.5806
R17502 VDD.n760 VDD.n757 75.5806
R17503 VDD.n750 VDD.n747 75.5806
R17504 VDD.n587 VDD.n584 75.5806
R17505 VDD.n577 VDD.n574 75.5806
R17506 VDD.n557 VDD.n554 75.5806
R17507 VDD.n547 VDD.n544 75.5806
R17508 VDD.n520 VDD.n517 75.5806
R17509 VDD.n500 VDD.n497 75.5806
R17510 VDD.n490 VDD.n487 75.5806
R17511 VDD.n7503 VDD.n7500 75.5806
R17512 VDD.n7493 VDD.n7490 75.5806
R17513 VDD.n7473 VDD.n7470 75.5806
R17514 VDD.n7463 VDD.n7460 75.5806
R17515 VDD.n7436 VDD.n7433 75.5806
R17516 VDD.n7416 VDD.n7413 75.5806
R17517 VDD.n7406 VDD.n7403 75.5806
R17518 VDD.n7243 VDD.n7240 75.5806
R17519 VDD.n7233 VDD.n7230 75.5806
R17520 VDD.n7213 VDD.n7210 75.5806
R17521 VDD.n1976 VDD.n1975 75.5806
R17522 VDD.n7179 VDD.n7176 75.5806
R17523 VDD.n7159 VDD.n7156 75.5806
R17524 VDD.n7149 VDD.n7146 75.5806
R17525 VDD.n6139 VDD.n6138 75.5806
R17526 VDD.n6131 VDD.n6128 75.5806
R17527 VDD.n6111 VDD.n6108 75.5806
R17528 VDD.n6084 VDD.n6081 75.5806
R17529 VDD.n6074 VDD.n6071 75.5806
R17530 VDD.n6054 VDD.n6051 75.5806
R17531 VDD.n6044 VDD.n6041 75.5806
R17532 VDD.n6262 VDD.n6261 75.5806
R17533 VDD.n6254 VDD.n6251 75.5806
R17534 VDD.n6234 VDD.n6231 75.5806
R17535 VDD.n6207 VDD.n6204 75.5806
R17536 VDD.n6197 VDD.n6194 75.5806
R17537 VDD.n6177 VDD.n6174 75.5806
R17538 VDD.n6167 VDD.n6164 75.5806
R17539 VDD.n6385 VDD.n6384 75.5806
R17540 VDD.n6377 VDD.n6374 75.5806
R17541 VDD.n6357 VDD.n6354 75.5806
R17542 VDD.n6330 VDD.n6327 75.5806
R17543 VDD.n6320 VDD.n6317 75.5806
R17544 VDD.n6300 VDD.n6297 75.5806
R17545 VDD.n6290 VDD.n6287 75.5806
R17546 VDD.n6508 VDD.n6507 75.5806
R17547 VDD.n6500 VDD.n6497 75.5806
R17548 VDD.n6480 VDD.n6477 75.5806
R17549 VDD.n6453 VDD.n6450 75.5806
R17550 VDD.n6443 VDD.n6440 75.5806
R17551 VDD.n6423 VDD.n6420 75.5806
R17552 VDD.n6413 VDD.n6410 75.5806
R17553 VDD.n6631 VDD.n6630 75.5806
R17554 VDD.n6623 VDD.n6620 75.5806
R17555 VDD.n6603 VDD.n6600 75.5806
R17556 VDD.n6576 VDD.n6573 75.5806
R17557 VDD.n6566 VDD.n6563 75.5806
R17558 VDD.n6546 VDD.n6543 75.5806
R17559 VDD.n6536 VDD.n6533 75.5806
R17560 VDD.n6754 VDD.n6753 75.5806
R17561 VDD.n6746 VDD.n6743 75.5806
R17562 VDD.n6726 VDD.n6723 75.5806
R17563 VDD.n6699 VDD.n6696 75.5806
R17564 VDD.n6689 VDD.n6686 75.5806
R17565 VDD.n6669 VDD.n6666 75.5806
R17566 VDD.n6659 VDD.n6656 75.5806
R17567 VDD.n6877 VDD.n6876 75.5806
R17568 VDD.n6869 VDD.n6866 75.5806
R17569 VDD.n6849 VDD.n6846 75.5806
R17570 VDD.n6822 VDD.n6819 75.5806
R17571 VDD.n6812 VDD.n6809 75.5806
R17572 VDD.n6792 VDD.n6789 75.5806
R17573 VDD.n6782 VDD.n6779 75.5806
R17574 VDD.n4961 VDD.n4958 75.5806
R17575 VDD.n4971 VDD.n4968 75.5806
R17576 VDD.n4991 VDD.n4988 75.5806
R17577 VDD.n5018 VDD.n5015 75.5806
R17578 VDD.n5028 VDD.n5025 75.5806
R17579 VDD.n5048 VDD.n5045 75.5806
R17580 VDD.n5058 VDD.n5055 75.5806
R17581 VDD.n4802 VDD.n4799 75.5806
R17582 VDD.n4792 VDD.n4789 75.5806
R17583 VDD.n4772 VDD.n4769 75.5806
R17584 VDD.n2112 VDD.n2111 75.5806
R17585 VDD.n4738 VDD.n4735 75.5806
R17586 VDD.n4718 VDD.n4715 75.5806
R17587 VDD.n4708 VDD.n4705 75.5806
R17588 VDD.n4677 VDD.n4674 75.5806
R17589 VDD.n4667 VDD.n4664 75.5806
R17590 VDD.n4647 VDD.n4644 75.5806
R17591 VDD.n2248 VDD.n2247 75.5806
R17592 VDD.n4613 VDD.n4610 75.5806
R17593 VDD.n4593 VDD.n4590 75.5806
R17594 VDD.n4583 VDD.n4580 75.5806
R17595 VDD.n4552 VDD.n4549 75.5806
R17596 VDD.n4542 VDD.n4539 75.5806
R17597 VDD.n4522 VDD.n4519 75.5806
R17598 VDD.n2384 VDD.n2383 75.5806
R17599 VDD.n4488 VDD.n4485 75.5806
R17600 VDD.n4468 VDD.n4465 75.5806
R17601 VDD.n4458 VDD.n4455 75.5806
R17602 VDD.n4427 VDD.n4424 75.5806
R17603 VDD.n4417 VDD.n4414 75.5806
R17604 VDD.n4397 VDD.n4394 75.5806
R17605 VDD.n2520 VDD.n2519 75.5806
R17606 VDD.n4363 VDD.n4360 75.5806
R17607 VDD.n4343 VDD.n4340 75.5806
R17608 VDD.n4333 VDD.n4330 75.5806
R17609 VDD.n4302 VDD.n4299 75.5806
R17610 VDD.n4292 VDD.n4289 75.5806
R17611 VDD.n4272 VDD.n4269 75.5806
R17612 VDD.n2656 VDD.n2655 75.5806
R17613 VDD.n4238 VDD.n4235 75.5806
R17614 VDD.n4218 VDD.n4215 75.5806
R17615 VDD.n4208 VDD.n4205 75.5806
R17616 VDD.n4177 VDD.n4174 75.5806
R17617 VDD.n4167 VDD.n4164 75.5806
R17618 VDD.n4147 VDD.n4144 75.5806
R17619 VDD.n2792 VDD.n2791 75.5806
R17620 VDD.n4113 VDD.n4110 75.5806
R17621 VDD.n4093 VDD.n4090 75.5806
R17622 VDD.n4083 VDD.n4080 75.5806
R17623 VDD.n4052 VDD.n4049 75.5806
R17624 VDD.n4042 VDD.n4039 75.5806
R17625 VDD.n4022 VDD.n4019 75.5806
R17626 VDD.n2928 VDD.n2927 75.5806
R17627 VDD.n3988 VDD.n3985 75.5806
R17628 VDD.n3968 VDD.n3965 75.5806
R17629 VDD.n3958 VDD.n3955 75.5806
R17630 VDD.n3608 VDD.n3607 75.5806
R17631 VDD.n3600 VDD.n3597 75.5806
R17632 VDD.n3927 VDD.n3924 75.5806
R17633 VDD.n3917 VDD.n3914 75.5806
R17634 VDD.n3897 VDD.n3894 75.5806
R17635 VDD.n3754 VDD.n3753 75.5806
R17636 VDD.n3863 VDD.n3860 75.5806
R17637 VDD.n3843 VDD.n3840 75.5806
R17638 VDD.n3833 VDD.n3830 75.5806
R17639 VDD.n3142 VDD.t1124 73.6406
R17640 VDD.n3158 VDD.t1110 73.6406
R17641 VDD.n3206 VDD.t1154 73.6406
R17642 VDD.n3222 VDD.t1151 73.6406
R17643 VDD.n3103 VDD.t1143 73.6406
R17644 VDD.n3246 VDD.t1133 73.6406
R17645 VDD.n3357 VDD.t1114 73.6406
R17646 VDD.n3623 VDD.t1147 73.6406
R17647 VDD.n3064 VDD.t1157 73.6406
R17648 VDD.n3080 VDD.t1119 73.6406
R17649 VDD.n3651 VDD.t1144 73.6406
R17650 VDD.n3667 VDD.t1109 73.6406
R17651 VDD.n3049 VDD.t1120 73.6406
R17652 VDD.n3038 VDD.t1140 73.6406
R17653 VDD.n3690 VDD.t1150 73.6406
R17654 VDD.n3122 VDD.t1136 73.6406
R17655 VDD.n3177 VDD.t1121 73.6406
R17656 VDD.n3711 VDD.t1123 73.6406
R17657 VDD.n3149 VDD.t1128 73.6304
R17658 VDD.n3138 VDD.t1113 73.6304
R17659 VDD.n3165 VDD.t1141 73.6304
R17660 VDD.n3155 VDD.t1132 73.6304
R17661 VDD.n3213 VDD.t1122 73.6304
R17662 VDD.n3202 VDD.t1156 73.6304
R17663 VDD.n3229 VDD.t1138 73.6304
R17664 VDD.n3219 VDD.t1155 73.6304
R17665 VDD.n3110 VDD.t1111 73.6304
R17666 VDD.n3099 VDD.t1135 73.6304
R17667 VDD.n3253 VDD.t1129 73.6304
R17668 VDD.n3243 VDD.t1130 73.6304
R17669 VDD.n3364 VDD.t1137 73.6304
R17670 VDD.n3353 VDD.t1152 73.6304
R17671 VDD.n3630 VDD.t1146 73.6304
R17672 VDD.n3620 VDD.t1115 73.6304
R17673 VDD.n3071 VDD.t1125 73.6304
R17674 VDD.n3060 VDD.t1126 73.6304
R17675 VDD.n3087 VDD.t1139 73.6304
R17676 VDD.n3077 VDD.t1158 73.6304
R17677 VDD.n3658 VDD.t1145 73.6304
R17678 VDD.n3647 VDD.t1112 73.6304
R17679 VDD.n3674 VDD.t1108 73.6304
R17680 VDD.n3664 VDD.t1131 73.6304
R17681 VDD.n3044 VDD.t1134 73.6304
R17682 VDD.n3697 VDD.t1148 73.6304
R17683 VDD.n3687 VDD.t1117 73.6304
R17684 VDD.n3129 VDD.t1153 73.6304
R17685 VDD.n3118 VDD.t1127 73.6304
R17686 VDD.n3184 VDD.t1116 73.6304
R17687 VDD.n3174 VDD.t1149 73.6304
R17688 VDD.n3718 VDD.t1118 73.6304
R17689 VDD.n3708 VDD.t1142 73.6304
R17690 VDD.n3394 VDD 71.7309
R17691 VDD.n3395 VDD.t781 69.9039
R17692 VDD VDD.t805 69.9004
R17693 VDD.n3405 VDD.t177 69.8804
R17694 VDD.n3400 VDD.t813 69.8804
R17695 VDD.n3489 VDD.t270 69.8804
R17696 VDD.n3500 VDD.t993 69.8804
R17697 VDD.n3495 VDD.t53 69.8804
R17698 VDD.n3583 VDD.t902 69.8804
R17699 VDD.n3342 VDD 63.2179
R17700 VDD.n337 VDD.n336 54.1632
R17701 VDD.n3450 VDD 53.5114
R17702 VDD.n3451 VDD 43.8048
R17703 VDD.n7517 VDD.n7257 42.18
R17704 VDD.n7531 VDD.n7530 37.0005
R17705 VDD.n7530 VDD.t241 37.0005
R17706 VDD.n37 VDD.n36 37.0005
R17707 VDD.n36 VDD.t241 37.0005
R17708 VDD.n7541 VDD.n7540 37.0005
R17709 VDD.n7540 VDD.t603 37.0005
R17710 VDD.n27 VDD.n26 37.0005
R17711 VDD.n26 VDD.t603 37.0005
R17712 VDD.n7551 VDD.n7550 37.0005
R17713 VDD.n7550 VDD.t830 37.0005
R17714 VDD.n14 VDD.n13 37.0005
R17715 VDD.n13 VDD.t830 37.0005
R17716 VDD.n7730 VDD.n7729 37.0005
R17717 VDD.n7729 VDD.t239 37.0005
R17718 VDD.n7560 VDD.n7559 37.0005
R17719 VDD.t239 VDD.n7560 37.0005
R17720 VDD.n7717 VDD.n7716 37.0005
R17721 VDD.n7716 VDD.t224 37.0005
R17722 VDD.n7568 VDD.n7567 37.0005
R17723 VDD.n7567 VDD.t224 37.0005
R17724 VDD.n7707 VDD.n7706 37.0005
R17725 VDD.n7706 VDD.t578 37.0005
R17726 VDD.n7581 VDD.n7580 37.0005
R17727 VDD.n7580 VDD.t578 37.0005
R17728 VDD.n7585 VDD.n7583 37.0005
R17729 VDD.n7583 VDD.t832 37.0005
R17730 VDD.n7698 VDD.n7584 37.0005
R17731 VDD.n7584 VDD.t832 37.0005
R17732 VDD.n7690 VDD.n7689 37.0005
R17733 VDD.n7689 VDD.t580 37.0005
R17734 VDD.n7596 VDD.n7595 37.0005
R17735 VDD.n7595 VDD.t580 37.0005
R17736 VDD.n7680 VDD.n7679 37.0005
R17737 VDD.n7679 VDD.t405 37.0005
R17738 VDD.n7609 VDD.n7608 37.0005
R17739 VDD.n7608 VDD.t405 37.0005
R17740 VDD.n7670 VDD.n7669 37.0005
R17741 VDD.n7669 VDD.t73 37.0005
R17742 VDD.n7620 VDD.n7619 37.0005
R17743 VDD.n7619 VDD.t73 37.0005
R17744 VDD.n7660 VDD.n7659 37.0005
R17745 VDD.n7659 VDD.t403 37.0005
R17746 VDD.n7630 VDD.n7629 37.0005
R17747 VDD.n7629 VDD.t403 37.0005
R17748 VDD.n7650 VDD.n7649 37.0005
R17749 VDD.n7649 VDD.t856 37.0005
R17750 VDD.n7643 VDD.n7642 37.0005
R17751 VDD.n7642 VDD.t856 37.0005
R17752 VDD.n32 VDD.n30 37.0005
R17753 VDD.n30 VDD.t241 37.0005
R17754 VDD.n7531 VDD.n31 37.0005
R17755 VDD.n31 VDD.t241 37.0005
R17756 VDD.n19 VDD.n17 37.0005
R17757 VDD.n17 VDD.t603 37.0005
R17758 VDD.n7541 VDD.n18 37.0005
R17759 VDD.n18 VDD.t603 37.0005
R17760 VDD.n10 VDD.n8 37.0005
R17761 VDD.n8 VDD.t830 37.0005
R17762 VDD.n7551 VDD.n9 37.0005
R17763 VDD.n9 VDD.t830 37.0005
R17764 VDD.n7728 VDD.n7727 37.0005
R17765 VDD.t239 VDD.n7728 37.0005
R17766 VDD.n7730 VDD.n3 37.0005
R17767 VDD.t239 VDD.n3 37.0005
R17768 VDD.n7564 VDD.n7562 37.0005
R17769 VDD.n7562 VDD.t224 37.0005
R17770 VDD.n7717 VDD.n7563 37.0005
R17771 VDD.n7563 VDD.t224 37.0005
R17772 VDD.n7573 VDD.n7571 37.0005
R17773 VDD.n7571 VDD.t578 37.0005
R17774 VDD.n7707 VDD.n7572 37.0005
R17775 VDD.n7572 VDD.t578 37.0005
R17776 VDD.n7589 VDD.n7587 37.0005
R17777 VDD.n7587 VDD.t580 37.0005
R17778 VDD.n7690 VDD.n7588 37.0005
R17779 VDD.n7588 VDD.t580 37.0005
R17780 VDD.n7601 VDD.n7599 37.0005
R17781 VDD.n7599 VDD.t405 37.0005
R17782 VDD.n7680 VDD.n7600 37.0005
R17783 VDD.n7600 VDD.t405 37.0005
R17784 VDD.n7614 VDD.n7612 37.0005
R17785 VDD.n7612 VDD.t73 37.0005
R17786 VDD.n7670 VDD.n7613 37.0005
R17787 VDD.n7613 VDD.t73 37.0005
R17788 VDD.n7625 VDD.n7623 37.0005
R17789 VDD.n7623 VDD.t403 37.0005
R17790 VDD.n7660 VDD.n7624 37.0005
R17791 VDD.n7624 VDD.t403 37.0005
R17792 VDD.n7635 VDD.n7633 37.0005
R17793 VDD.n7633 VDD.t856 37.0005
R17794 VDD.n7650 VDD.n7634 37.0005
R17795 VDD.n7634 VDD.t856 37.0005
R17796 VDD.n41 VDD.n39 37.0005
R17797 VDD.n39 VDD.t867 37.0005
R17798 VDD.n7522 VDD.n40 37.0005
R17799 VDD.n1890 VDD.n1889 37.0005
R17800 VDD.n1889 VDD.t243 37.0005
R17801 VDD.n1657 VDD.n1656 37.0005
R17802 VDD.n1656 VDD.t243 37.0005
R17803 VDD.n1880 VDD.n1879 37.0005
R17804 VDD.n1879 VDD.t599 37.0005
R17805 VDD.n1667 VDD.n1666 37.0005
R17806 VDD.n1666 VDD.t599 37.0005
R17807 VDD.n1870 VDD.n1869 37.0005
R17808 VDD.n1869 VDD.t923 37.0005
R17809 VDD.n1680 VDD.n1679 37.0005
R17810 VDD.n1679 VDD.t923 37.0005
R17811 VDD.n1860 VDD.n1859 37.0005
R17812 VDD.n1859 VDD.t358 37.0005
R17813 VDD.n1691 VDD.n1690 37.0005
R17814 VDD.n1690 VDD.t358 37.0005
R17815 VDD.n1850 VDD.n1849 37.0005
R17816 VDD.n1849 VDD.t567 37.0005
R17817 VDD.n1701 VDD.n1700 37.0005
R17818 VDD.n1700 VDD.t567 37.0005
R17819 VDD.n1840 VDD.n1839 37.0005
R17820 VDD.n1839 VDD.t597 37.0005
R17821 VDD.n1714 VDD.n1713 37.0005
R17822 VDD.n1713 VDD.t597 37.0005
R17823 VDD.n1718 VDD.n1716 37.0005
R17824 VDD.n1716 VDD.t925 37.0005
R17825 VDD.n1831 VDD.n1717 37.0005
R17826 VDD.n1717 VDD.t925 37.0005
R17827 VDD.n1823 VDD.n1822 37.0005
R17828 VDD.n1822 VDD.t595 37.0005
R17829 VDD.n1729 VDD.n1728 37.0005
R17830 VDD.n1728 VDD.t595 37.0005
R17831 VDD.n1813 VDD.n1812 37.0005
R17832 VDD.n1812 VDD.t157 37.0005
R17833 VDD.n1742 VDD.n1741 37.0005
R17834 VDD.n1741 VDD.t157 37.0005
R17835 VDD.n1803 VDD.n1802 37.0005
R17836 VDD.n1802 VDD.t27 37.0005
R17837 VDD.n1753 VDD.n1752 37.0005
R17838 VDD.n1752 VDD.t27 37.0005
R17839 VDD.n1793 VDD.n1792 37.0005
R17840 VDD.n1792 VDD.t422 37.0005
R17841 VDD.n1763 VDD.n1762 37.0005
R17842 VDD.n1762 VDD.t422 37.0005
R17843 VDD.n1783 VDD.n1782 37.0005
R17844 VDD.n1782 VDD.t54 37.0005
R17845 VDD.n1776 VDD.n1775 37.0005
R17846 VDD.n1775 VDD.t54 37.0005
R17847 VDD.n1651 VDD.n1649 37.0005
R17848 VDD.n1649 VDD.t243 37.0005
R17849 VDD.n1890 VDD.n1650 37.0005
R17850 VDD.n1650 VDD.t243 37.0005
R17851 VDD.n1662 VDD.n1660 37.0005
R17852 VDD.n1660 VDD.t599 37.0005
R17853 VDD.n1880 VDD.n1661 37.0005
R17854 VDD.n1661 VDD.t599 37.0005
R17855 VDD.n1672 VDD.n1670 37.0005
R17856 VDD.n1670 VDD.t923 37.0005
R17857 VDD.n1870 VDD.n1671 37.0005
R17858 VDD.n1671 VDD.t923 37.0005
R17859 VDD.n1685 VDD.n1683 37.0005
R17860 VDD.n1683 VDD.t358 37.0005
R17861 VDD.n1860 VDD.n1684 37.0005
R17862 VDD.n1684 VDD.t358 37.0005
R17863 VDD.n1696 VDD.n1694 37.0005
R17864 VDD.n1694 VDD.t567 37.0005
R17865 VDD.n1850 VDD.n1695 37.0005
R17866 VDD.n1695 VDD.t567 37.0005
R17867 VDD.n1706 VDD.n1704 37.0005
R17868 VDD.n1704 VDD.t597 37.0005
R17869 VDD.n1840 VDD.n1705 37.0005
R17870 VDD.n1705 VDD.t597 37.0005
R17871 VDD.n1722 VDD.n1720 37.0005
R17872 VDD.n1720 VDD.t595 37.0005
R17873 VDD.n1823 VDD.n1721 37.0005
R17874 VDD.n1721 VDD.t595 37.0005
R17875 VDD.n1734 VDD.n1732 37.0005
R17876 VDD.n1732 VDD.t157 37.0005
R17877 VDD.n1813 VDD.n1733 37.0005
R17878 VDD.n1733 VDD.t157 37.0005
R17879 VDD.n1747 VDD.n1745 37.0005
R17880 VDD.n1745 VDD.t27 37.0005
R17881 VDD.n1803 VDD.n1746 37.0005
R17882 VDD.n1746 VDD.t27 37.0005
R17883 VDD.n1758 VDD.n1756 37.0005
R17884 VDD.n1756 VDD.t422 37.0005
R17885 VDD.n1793 VDD.n1757 37.0005
R17886 VDD.n1757 VDD.t422 37.0005
R17887 VDD.n1768 VDD.n1766 37.0005
R17888 VDD.n1766 VDD.t54 37.0005
R17889 VDD.n1783 VDD.n1767 37.0005
R17890 VDD.n1767 VDD.t54 37.0005
R17891 VDD.n1645 VDD.n1644 37.0005
R17892 VDD.t863 VDD.n1645 37.0005
R17893 VDD.n1898 VDD.n1643 37.0005
R17894 VDD.n1630 VDD.n1629 37.0005
R17895 VDD.n1629 VDD.t418 37.0005
R17896 VDD.n1397 VDD.n1396 37.0005
R17897 VDD.n1396 VDD.t418 37.0005
R17898 VDD.n1620 VDD.n1619 37.0005
R17899 VDD.n1619 VDD.t806 37.0005
R17900 VDD.n1407 VDD.n1406 37.0005
R17901 VDD.n1406 VDD.t806 37.0005
R17902 VDD.n1610 VDD.n1609 37.0005
R17903 VDD.n1609 VDD.t4 37.0005
R17904 VDD.n1420 VDD.n1419 37.0005
R17905 VDD.n1419 VDD.t4 37.0005
R17906 VDD.n1600 VDD.n1599 37.0005
R17907 VDD.n1599 VDD.t15 37.0005
R17908 VDD.n1431 VDD.n1430 37.0005
R17909 VDD.n1430 VDD.t15 37.0005
R17910 VDD.n1590 VDD.n1589 37.0005
R17911 VDD.n1589 VDD.t93 37.0005
R17912 VDD.n1441 VDD.n1440 37.0005
R17913 VDD.n1440 VDD.t93 37.0005
R17914 VDD.n1580 VDD.n1579 37.0005
R17915 VDD.n1579 VDD.t769 37.0005
R17916 VDD.n1454 VDD.n1453 37.0005
R17917 VDD.n1453 VDD.t769 37.0005
R17918 VDD.n1458 VDD.n1456 37.0005
R17919 VDD.n1456 VDD.t6 37.0005
R17920 VDD.n1571 VDD.n1457 37.0005
R17921 VDD.n1457 VDD.t6 37.0005
R17922 VDD.n1563 VDD.n1562 37.0005
R17923 VDD.n1562 VDD.t771 37.0005
R17924 VDD.n1469 VDD.n1468 37.0005
R17925 VDD.n1468 VDD.t771 37.0005
R17926 VDD.n1553 VDD.n1552 37.0005
R17927 VDD.n1552 VDD.t815 37.0005
R17928 VDD.n1482 VDD.n1481 37.0005
R17929 VDD.n1481 VDD.t815 37.0005
R17930 VDD.n1543 VDD.n1542 37.0005
R17931 VDD.n1542 VDD.t644 37.0005
R17932 VDD.n1493 VDD.n1492 37.0005
R17933 VDD.n1492 VDD.t644 37.0005
R17934 VDD.n1533 VDD.n1532 37.0005
R17935 VDD.n1532 VDD.t298 37.0005
R17936 VDD.n1503 VDD.n1502 37.0005
R17937 VDD.n1502 VDD.t298 37.0005
R17938 VDD.n1523 VDD.n1522 37.0005
R17939 VDD.n1522 VDD.t994 37.0005
R17940 VDD.n1516 VDD.n1515 37.0005
R17941 VDD.n1515 VDD.t994 37.0005
R17942 VDD.n1391 VDD.n1389 37.0005
R17943 VDD.n1389 VDD.t418 37.0005
R17944 VDD.n1630 VDD.n1390 37.0005
R17945 VDD.n1390 VDD.t418 37.0005
R17946 VDD.n1402 VDD.n1400 37.0005
R17947 VDD.n1400 VDD.t806 37.0005
R17948 VDD.n1620 VDD.n1401 37.0005
R17949 VDD.n1401 VDD.t806 37.0005
R17950 VDD.n1412 VDD.n1410 37.0005
R17951 VDD.n1410 VDD.t4 37.0005
R17952 VDD.n1610 VDD.n1411 37.0005
R17953 VDD.n1411 VDD.t4 37.0005
R17954 VDD.n1425 VDD.n1423 37.0005
R17955 VDD.n1423 VDD.t15 37.0005
R17956 VDD.n1600 VDD.n1424 37.0005
R17957 VDD.n1424 VDD.t15 37.0005
R17958 VDD.n1436 VDD.n1434 37.0005
R17959 VDD.n1434 VDD.t93 37.0005
R17960 VDD.n1590 VDD.n1435 37.0005
R17961 VDD.n1435 VDD.t93 37.0005
R17962 VDD.n1446 VDD.n1444 37.0005
R17963 VDD.n1444 VDD.t769 37.0005
R17964 VDD.n1580 VDD.n1445 37.0005
R17965 VDD.n1445 VDD.t769 37.0005
R17966 VDD.n1462 VDD.n1460 37.0005
R17967 VDD.n1460 VDD.t771 37.0005
R17968 VDD.n1563 VDD.n1461 37.0005
R17969 VDD.n1461 VDD.t771 37.0005
R17970 VDD.n1474 VDD.n1472 37.0005
R17971 VDD.n1472 VDD.t815 37.0005
R17972 VDD.n1553 VDD.n1473 37.0005
R17973 VDD.n1473 VDD.t815 37.0005
R17974 VDD.n1487 VDD.n1485 37.0005
R17975 VDD.n1485 VDD.t644 37.0005
R17976 VDD.n1543 VDD.n1486 37.0005
R17977 VDD.n1486 VDD.t644 37.0005
R17978 VDD.n1498 VDD.n1496 37.0005
R17979 VDD.n1496 VDD.t298 37.0005
R17980 VDD.n1533 VDD.n1497 37.0005
R17981 VDD.n1497 VDD.t298 37.0005
R17982 VDD.n1508 VDD.n1506 37.0005
R17983 VDD.n1506 VDD.t994 37.0005
R17984 VDD.n1523 VDD.n1507 37.0005
R17985 VDD.n1507 VDD.t994 37.0005
R17986 VDD.n1385 VDD.n1384 37.0005
R17987 VDD.t609 VDD.n1385 37.0005
R17988 VDD.n1638 VDD.n1383 37.0005
R17989 VDD.n1370 VDD.n1369 37.0005
R17990 VDD.n1369 VDD.t480 37.0005
R17991 VDD.n1137 VDD.n1136 37.0005
R17992 VDD.n1136 VDD.t480 37.0005
R17993 VDD.n1360 VDD.n1359 37.0005
R17994 VDD.n1359 VDD.t393 37.0005
R17995 VDD.n1147 VDD.n1146 37.0005
R17996 VDD.n1146 VDD.t393 37.0005
R17997 VDD.n1350 VDD.n1349 37.0005
R17998 VDD.n1349 VDD.t101 37.0005
R17999 VDD.n1160 VDD.n1159 37.0005
R18000 VDD.n1159 VDD.t101 37.0005
R18001 VDD.n1340 VDD.n1339 37.0005
R18002 VDD.n1339 VDD.t538 37.0005
R18003 VDD.n1171 VDD.n1170 37.0005
R18004 VDD.n1170 VDD.t538 37.0005
R18005 VDD.n1330 VDD.n1329 37.0005
R18006 VDD.n1329 VDD.t412 37.0005
R18007 VDD.n1181 VDD.n1180 37.0005
R18008 VDD.n1180 VDD.t412 37.0005
R18009 VDD.n1320 VDD.n1319 37.0005
R18010 VDD.n1319 VDD.t778 37.0005
R18011 VDD.n1194 VDD.n1193 37.0005
R18012 VDD.n1193 VDD.t778 37.0005
R18013 VDD.n1198 VDD.n1196 37.0005
R18014 VDD.n1196 VDD.t103 37.0005
R18015 VDD.n1311 VDD.n1197 37.0005
R18016 VDD.n1197 VDD.t103 37.0005
R18017 VDD.n1303 VDD.n1302 37.0005
R18018 VDD.n1302 VDD.t191 37.0005
R18019 VDD.n1209 VDD.n1208 37.0005
R18020 VDD.n1208 VDD.t191 37.0005
R18021 VDD.n1293 VDD.n1292 37.0005
R18022 VDD.n1292 VDD.t178 37.0005
R18023 VDD.n1222 VDD.n1221 37.0005
R18024 VDD.n1221 VDD.t178 37.0005
R18025 VDD.n1283 VDD.n1282 37.0005
R18026 VDD.n1282 VDD.t211 37.0005
R18027 VDD.n1233 VDD.n1232 37.0005
R18028 VDD.n1232 VDD.t211 37.0005
R18029 VDD.n1273 VDD.n1272 37.0005
R18030 VDD.n1272 VDD.t360 37.0005
R18031 VDD.n1243 VDD.n1242 37.0005
R18032 VDD.n1242 VDD.t360 37.0005
R18033 VDD.n1263 VDD.n1262 37.0005
R18034 VDD.n1262 VDD.t114 37.0005
R18035 VDD.n1256 VDD.n1255 37.0005
R18036 VDD.n1255 VDD.t114 37.0005
R18037 VDD.n1131 VDD.n1129 37.0005
R18038 VDD.n1129 VDD.t480 37.0005
R18039 VDD.n1370 VDD.n1130 37.0005
R18040 VDD.n1130 VDD.t480 37.0005
R18041 VDD.n1142 VDD.n1140 37.0005
R18042 VDD.n1140 VDD.t393 37.0005
R18043 VDD.n1360 VDD.n1141 37.0005
R18044 VDD.n1141 VDD.t393 37.0005
R18045 VDD.n1152 VDD.n1150 37.0005
R18046 VDD.n1150 VDD.t101 37.0005
R18047 VDD.n1350 VDD.n1151 37.0005
R18048 VDD.n1151 VDD.t101 37.0005
R18049 VDD.n1165 VDD.n1163 37.0005
R18050 VDD.n1163 VDD.t538 37.0005
R18051 VDD.n1340 VDD.n1164 37.0005
R18052 VDD.n1164 VDD.t538 37.0005
R18053 VDD.n1176 VDD.n1174 37.0005
R18054 VDD.n1174 VDD.t412 37.0005
R18055 VDD.n1330 VDD.n1175 37.0005
R18056 VDD.n1175 VDD.t412 37.0005
R18057 VDD.n1186 VDD.n1184 37.0005
R18058 VDD.n1184 VDD.t778 37.0005
R18059 VDD.n1320 VDD.n1185 37.0005
R18060 VDD.n1185 VDD.t778 37.0005
R18061 VDD.n1202 VDD.n1200 37.0005
R18062 VDD.n1200 VDD.t191 37.0005
R18063 VDD.n1303 VDD.n1201 37.0005
R18064 VDD.n1201 VDD.t191 37.0005
R18065 VDD.n1214 VDD.n1212 37.0005
R18066 VDD.n1212 VDD.t178 37.0005
R18067 VDD.n1293 VDD.n1213 37.0005
R18068 VDD.n1213 VDD.t178 37.0005
R18069 VDD.n1227 VDD.n1225 37.0005
R18070 VDD.n1225 VDD.t211 37.0005
R18071 VDD.n1283 VDD.n1226 37.0005
R18072 VDD.n1226 VDD.t211 37.0005
R18073 VDD.n1238 VDD.n1236 37.0005
R18074 VDD.n1236 VDD.t360 37.0005
R18075 VDD.n1273 VDD.n1237 37.0005
R18076 VDD.n1237 VDD.t360 37.0005
R18077 VDD.n1248 VDD.n1246 37.0005
R18078 VDD.n1246 VDD.t114 37.0005
R18079 VDD.n1263 VDD.n1247 37.0005
R18080 VDD.n1247 VDD.t114 37.0005
R18081 VDD.n1125 VDD.n1124 37.0005
R18082 VDD.t961 VDD.n1125 37.0005
R18083 VDD.n1378 VDD.n1123 37.0005
R18084 VDD.n1110 VDD.n1109 37.0005
R18085 VDD.n1109 VDD.t247 37.0005
R18086 VDD.n877 VDD.n876 37.0005
R18087 VDD.n876 VDD.t247 37.0005
R18088 VDD.n1100 VDD.n1099 37.0005
R18089 VDD.n1099 VDD.t601 37.0005
R18090 VDD.n887 VDD.n886 37.0005
R18091 VDD.n886 VDD.t601 37.0005
R18092 VDD.n1090 VDD.n1089 37.0005
R18093 VDD.n1089 VDD.t657 37.0005
R18094 VDD.n900 VDD.n899 37.0005
R18095 VDD.n899 VDD.t657 37.0005
R18096 VDD.n1080 VDD.n1079 37.0005
R18097 VDD.n1079 VDD.t642 37.0005
R18098 VDD.n911 VDD.n910 37.0005
R18099 VDD.n910 VDD.t642 37.0005
R18100 VDD.n1070 VDD.n1069 37.0005
R18101 VDD.n1069 VDD.t429 37.0005
R18102 VDD.n921 VDD.n920 37.0005
R18103 VDD.n920 VDD.t429 37.0005
R18104 VDD.n1060 VDD.n1059 37.0005
R18105 VDD.n1059 VDD.t174 37.0005
R18106 VDD.n934 VDD.n933 37.0005
R18107 VDD.n933 VDD.t174 37.0005
R18108 VDD.n938 VDD.n936 37.0005
R18109 VDD.n936 VDD.t659 37.0005
R18110 VDD.n1051 VDD.n937 37.0005
R18111 VDD.n937 VDD.t659 37.0005
R18112 VDD.n1043 VDD.n1042 37.0005
R18113 VDD.n1042 VDD.t172 37.0005
R18114 VDD.n949 VDD.n948 37.0005
R18115 VDD.n948 VDD.t172 37.0005
R18116 VDD.n1033 VDD.n1032 37.0005
R18117 VDD.n1032 VDD.t346 37.0005
R18118 VDD.n962 VDD.n961 37.0005
R18119 VDD.n961 VDD.t346 37.0005
R18120 VDD.n1023 VDD.n1022 37.0005
R18121 VDD.n1022 VDD.t9 37.0005
R18122 VDD.n973 VDD.n972 37.0005
R18123 VDD.n972 VDD.t9 37.0005
R18124 VDD.n1013 VDD.n1012 37.0005
R18125 VDD.n1012 VDD.t318 37.0005
R18126 VDD.n983 VDD.n982 37.0005
R18127 VDD.n982 VDD.t318 37.0005
R18128 VDD.n1003 VDD.n1002 37.0005
R18129 VDD.n1002 VDD.t808 37.0005
R18130 VDD.n996 VDD.n995 37.0005
R18131 VDD.n995 VDD.t808 37.0005
R18132 VDD.n871 VDD.n869 37.0005
R18133 VDD.n869 VDD.t247 37.0005
R18134 VDD.n1110 VDD.n870 37.0005
R18135 VDD.n870 VDD.t247 37.0005
R18136 VDD.n882 VDD.n880 37.0005
R18137 VDD.n880 VDD.t601 37.0005
R18138 VDD.n1100 VDD.n881 37.0005
R18139 VDD.n881 VDD.t601 37.0005
R18140 VDD.n892 VDD.n890 37.0005
R18141 VDD.n890 VDD.t657 37.0005
R18142 VDD.n1090 VDD.n891 37.0005
R18143 VDD.n891 VDD.t657 37.0005
R18144 VDD.n905 VDD.n903 37.0005
R18145 VDD.n903 VDD.t642 37.0005
R18146 VDD.n1080 VDD.n904 37.0005
R18147 VDD.n904 VDD.t642 37.0005
R18148 VDD.n916 VDD.n914 37.0005
R18149 VDD.n914 VDD.t429 37.0005
R18150 VDD.n1070 VDD.n915 37.0005
R18151 VDD.n915 VDD.t429 37.0005
R18152 VDD.n926 VDD.n924 37.0005
R18153 VDD.n924 VDD.t174 37.0005
R18154 VDD.n1060 VDD.n925 37.0005
R18155 VDD.n925 VDD.t174 37.0005
R18156 VDD.n942 VDD.n940 37.0005
R18157 VDD.n940 VDD.t172 37.0005
R18158 VDD.n1043 VDD.n941 37.0005
R18159 VDD.n941 VDD.t172 37.0005
R18160 VDD.n954 VDD.n952 37.0005
R18161 VDD.n952 VDD.t346 37.0005
R18162 VDD.n1033 VDD.n953 37.0005
R18163 VDD.n953 VDD.t346 37.0005
R18164 VDD.n967 VDD.n965 37.0005
R18165 VDD.n965 VDD.t9 37.0005
R18166 VDD.n1023 VDD.n966 37.0005
R18167 VDD.n966 VDD.t9 37.0005
R18168 VDD.n978 VDD.n976 37.0005
R18169 VDD.n976 VDD.t318 37.0005
R18170 VDD.n1013 VDD.n977 37.0005
R18171 VDD.n977 VDD.t318 37.0005
R18172 VDD.n988 VDD.n986 37.0005
R18173 VDD.n986 VDD.t808 37.0005
R18174 VDD.n1003 VDD.n987 37.0005
R18175 VDD.n987 VDD.t808 37.0005
R18176 VDD.n865 VDD.n864 37.0005
R18177 VDD.t865 VDD.n865 37.0005
R18178 VDD.n1118 VDD.n863 37.0005
R18179 VDD.n850 VDD.n849 37.0005
R18180 VDD.n849 VDD.t353 37.0005
R18181 VDD.n617 VDD.n616 37.0005
R18182 VDD.n616 VDD.t353 37.0005
R18183 VDD.n840 VDD.n839 37.0005
R18184 VDD.n839 VDD.t120 37.0005
R18185 VDD.n627 VDD.n626 37.0005
R18186 VDD.n626 VDD.t120 37.0005
R18187 VDD.n830 VDD.n829 37.0005
R18188 VDD.n829 VDD.t41 37.0005
R18189 VDD.n640 VDD.n639 37.0005
R18190 VDD.n639 VDD.t41 37.0005
R18191 VDD.n820 VDD.n819 37.0005
R18192 VDD.n819 VDD.t384 37.0005
R18193 VDD.n651 VDD.n650 37.0005
R18194 VDD.n650 VDD.t384 37.0005
R18195 VDD.n810 VDD.n809 37.0005
R18196 VDD.n809 VDD.t220 37.0005
R18197 VDD.n661 VDD.n660 37.0005
R18198 VDD.n660 VDD.t220 37.0005
R18199 VDD.n800 VDD.n799 37.0005
R18200 VDD.n799 VDD.t166 37.0005
R18201 VDD.n674 VDD.n673 37.0005
R18202 VDD.n673 VDD.t166 37.0005
R18203 VDD.n678 VDD.n676 37.0005
R18204 VDD.n676 VDD.t43 37.0005
R18205 VDD.n791 VDD.n677 37.0005
R18206 VDD.n677 VDD.t43 37.0005
R18207 VDD.n783 VDD.n782 37.0005
R18208 VDD.n782 VDD.t164 37.0005
R18209 VDD.n689 VDD.n688 37.0005
R18210 VDD.n688 VDD.t164 37.0005
R18211 VDD.n773 VDD.n772 37.0005
R18212 VDD.n772 VDD.t60 37.0005
R18213 VDD.n702 VDD.n701 37.0005
R18214 VDD.n701 VDD.t60 37.0005
R18215 VDD.n763 VDD.n762 37.0005
R18216 VDD.n762 VDD.t356 37.0005
R18217 VDD.n713 VDD.n712 37.0005
R18218 VDD.n712 VDD.t356 37.0005
R18219 VDD.n753 VDD.n752 37.0005
R18220 VDD.n752 VDD.t63 37.0005
R18221 VDD.n723 VDD.n722 37.0005
R18222 VDD.n722 VDD.t63 37.0005
R18223 VDD.n743 VDD.n742 37.0005
R18224 VDD.n742 VDD.t278 37.0005
R18225 VDD.n736 VDD.n735 37.0005
R18226 VDD.n735 VDD.t278 37.0005
R18227 VDD.n611 VDD.n609 37.0005
R18228 VDD.n609 VDD.t353 37.0005
R18229 VDD.n850 VDD.n610 37.0005
R18230 VDD.n610 VDD.t353 37.0005
R18231 VDD.n622 VDD.n620 37.0005
R18232 VDD.n620 VDD.t120 37.0005
R18233 VDD.n840 VDD.n621 37.0005
R18234 VDD.n621 VDD.t120 37.0005
R18235 VDD.n632 VDD.n630 37.0005
R18236 VDD.n630 VDD.t41 37.0005
R18237 VDD.n830 VDD.n631 37.0005
R18238 VDD.n631 VDD.t41 37.0005
R18239 VDD.n645 VDD.n643 37.0005
R18240 VDD.n643 VDD.t384 37.0005
R18241 VDD.n820 VDD.n644 37.0005
R18242 VDD.n644 VDD.t384 37.0005
R18243 VDD.n656 VDD.n654 37.0005
R18244 VDD.n654 VDD.t220 37.0005
R18245 VDD.n810 VDD.n655 37.0005
R18246 VDD.n655 VDD.t220 37.0005
R18247 VDD.n666 VDD.n664 37.0005
R18248 VDD.n664 VDD.t166 37.0005
R18249 VDD.n800 VDD.n665 37.0005
R18250 VDD.n665 VDD.t166 37.0005
R18251 VDD.n682 VDD.n680 37.0005
R18252 VDD.n680 VDD.t164 37.0005
R18253 VDD.n783 VDD.n681 37.0005
R18254 VDD.n681 VDD.t164 37.0005
R18255 VDD.n694 VDD.n692 37.0005
R18256 VDD.n692 VDD.t60 37.0005
R18257 VDD.n773 VDD.n693 37.0005
R18258 VDD.n693 VDD.t60 37.0005
R18259 VDD.n707 VDD.n705 37.0005
R18260 VDD.n705 VDD.t356 37.0005
R18261 VDD.n763 VDD.n706 37.0005
R18262 VDD.n706 VDD.t356 37.0005
R18263 VDD.n718 VDD.n716 37.0005
R18264 VDD.n716 VDD.t63 37.0005
R18265 VDD.n753 VDD.n717 37.0005
R18266 VDD.n717 VDD.t63 37.0005
R18267 VDD.n728 VDD.n726 37.0005
R18268 VDD.n726 VDD.t278 37.0005
R18269 VDD.n743 VDD.n727 37.0005
R18270 VDD.n727 VDD.t278 37.0005
R18271 VDD.n605 VDD.n604 37.0005
R18272 VDD.t605 VDD.n605 37.0005
R18273 VDD.n858 VDD.n603 37.0005
R18274 VDD.n590 VDD.n589 37.0005
R18275 VDD.n589 VDD.t11 37.0005
R18276 VDD.n357 VDD.n356 37.0005
R18277 VDD.n356 VDD.t11 37.0005
R18278 VDD.n580 VDD.n579 37.0005
R18279 VDD.n579 VDD.t333 37.0005
R18280 VDD.n367 VDD.n366 37.0005
R18281 VDD.n366 VDD.t333 37.0005
R18282 VDD.n570 VDD.n569 37.0005
R18283 VDD.n569 VDD.t555 37.0005
R18284 VDD.n380 VDD.n379 37.0005
R18285 VDD.n379 VDD.t555 37.0005
R18286 VDD.n560 VDD.n559 37.0005
R18287 VDD.n559 VDD.t249 37.0005
R18288 VDD.n391 VDD.n390 37.0005
R18289 VDD.n390 VDD.t249 37.0005
R18290 VDD.n550 VDD.n549 37.0005
R18291 VDD.n549 VDD.t75 37.0005
R18292 VDD.n401 VDD.n400 37.0005
R18293 VDD.n400 VDD.t75 37.0005
R18294 VDD.n540 VDD.n539 37.0005
R18295 VDD.n539 VDD.t233 37.0005
R18296 VDD.n414 VDD.n413 37.0005
R18297 VDD.n413 VDD.t233 37.0005
R18298 VDD.n418 VDD.n416 37.0005
R18299 VDD.n416 VDD.t58 37.0005
R18300 VDD.n531 VDD.n417 37.0005
R18301 VDD.n417 VDD.t58 37.0005
R18302 VDD.n523 VDD.n522 37.0005
R18303 VDD.n522 VDD.t204 37.0005
R18304 VDD.n429 VDD.n428 37.0005
R18305 VDD.n428 VDD.t204 37.0005
R18306 VDD.n513 VDD.n512 37.0005
R18307 VDD.n512 VDD.t988 37.0005
R18308 VDD.n442 VDD.n441 37.0005
R18309 VDD.n441 VDD.t988 37.0005
R18310 VDD.n503 VDD.n502 37.0005
R18311 VDD.n502 VDD.t339 37.0005
R18312 VDD.n453 VDD.n452 37.0005
R18313 VDD.n452 VDD.t339 37.0005
R18314 VDD.n493 VDD.n492 37.0005
R18315 VDD.n492 VDD.t335 37.0005
R18316 VDD.n463 VDD.n462 37.0005
R18317 VDD.n462 VDD.t335 37.0005
R18318 VDD.n483 VDD.n482 37.0005
R18319 VDD.n482 VDD.t362 37.0005
R18320 VDD.n476 VDD.n475 37.0005
R18321 VDD.n475 VDD.t362 37.0005
R18322 VDD.n351 VDD.n349 37.0005
R18323 VDD.n349 VDD.t11 37.0005
R18324 VDD.n590 VDD.n350 37.0005
R18325 VDD.n350 VDD.t11 37.0005
R18326 VDD.n362 VDD.n360 37.0005
R18327 VDD.n360 VDD.t333 37.0005
R18328 VDD.n580 VDD.n361 37.0005
R18329 VDD.n361 VDD.t333 37.0005
R18330 VDD.n372 VDD.n370 37.0005
R18331 VDD.n370 VDD.t555 37.0005
R18332 VDD.n570 VDD.n371 37.0005
R18333 VDD.n371 VDD.t555 37.0005
R18334 VDD.n385 VDD.n383 37.0005
R18335 VDD.n383 VDD.t249 37.0005
R18336 VDD.n560 VDD.n384 37.0005
R18337 VDD.n384 VDD.t249 37.0005
R18338 VDD.n396 VDD.n394 37.0005
R18339 VDD.n394 VDD.t75 37.0005
R18340 VDD.n550 VDD.n395 37.0005
R18341 VDD.n395 VDD.t75 37.0005
R18342 VDD.n406 VDD.n404 37.0005
R18343 VDD.n404 VDD.t233 37.0005
R18344 VDD.n540 VDD.n405 37.0005
R18345 VDD.n405 VDD.t233 37.0005
R18346 VDD.n422 VDD.n420 37.0005
R18347 VDD.n420 VDD.t204 37.0005
R18348 VDD.n523 VDD.n421 37.0005
R18349 VDD.n421 VDD.t204 37.0005
R18350 VDD.n434 VDD.n432 37.0005
R18351 VDD.n432 VDD.t988 37.0005
R18352 VDD.n513 VDD.n433 37.0005
R18353 VDD.n433 VDD.t988 37.0005
R18354 VDD.n447 VDD.n445 37.0005
R18355 VDD.n445 VDD.t339 37.0005
R18356 VDD.n503 VDD.n446 37.0005
R18357 VDD.n446 VDD.t339 37.0005
R18358 VDD.n458 VDD.n456 37.0005
R18359 VDD.n456 VDD.t335 37.0005
R18360 VDD.n493 VDD.n457 37.0005
R18361 VDD.n457 VDD.t335 37.0005
R18362 VDD.n468 VDD.n466 37.0005
R18363 VDD.n466 VDD.t362 37.0005
R18364 VDD.n483 VDD.n467 37.0005
R18365 VDD.n467 VDD.t362 37.0005
R18366 VDD.n345 VDD.n344 37.0005
R18367 VDD.t963 VDD.n345 37.0005
R18368 VDD.n598 VDD.n343 37.0005
R18369 VDD.n292 VDD.n291 37.0005
R18370 VDD.n339 VDD.n338 37.0005
R18371 VDD.n338 VDD.t401 37.0005
R18372 VDD.n333 VDD.n295 37.0005
R18373 VDD.n295 VDD.t786 37.0005
R18374 VDD.n331 VDD.n330 37.0005
R18375 VDD.n330 VDD.t89 37.0005
R18376 VDD.n296 VDD.n294 37.0005
R18377 VDD.n294 VDD.t786 37.0005
R18378 VDD.n328 VDD.n327 37.0005
R18379 VDD.n146 VDD.n143 37.0005
R18380 VDD.n143 VDD.t213 37.0005
R18381 VDD.n150 VDD.n144 37.0005
R18382 VDD.n140 VDD.n139 37.0005
R18383 VDD.t370 VDD.n140 37.0005
R18384 VDD.n157 VDD.n138 37.0005
R18385 VDD.n129 VDD.n127 37.0005
R18386 VDD.n127 VDD.t1072 37.0005
R18387 VDD.n171 VDD.n128 37.0005
R18388 VDD.n128 VDD.t1072 37.0005
R18389 VDD.n160 VDD.n130 37.0005
R18390 VDD.n130 VDD.t654 37.0005
R18391 VDD.n164 VDD.n131 37.0005
R18392 VDD.n124 VDD.n123 37.0005
R18393 VDD.t846 VDD.n124 37.0005
R18394 VDD.n178 VDD.n122 37.0005
R18395 VDD.n181 VDD.n118 37.0005
R18396 VDD.n118 VDD.t619 37.0005
R18397 VDD.n185 VDD.n119 37.0005
R18398 VDD.n115 VDD.n114 37.0005
R18399 VDD.t128 VDD.n115 37.0005
R18400 VDD.n192 VDD.n113 37.0005
R18401 VDD.n104 VDD.n102 37.0005
R18402 VDD.n102 VDD.t1026 37.0005
R18403 VDD.n206 VDD.n103 37.0005
R18404 VDD.n103 VDD.t1026 37.0005
R18405 VDD.n195 VDD.n105 37.0005
R18406 VDD.n105 VDD.t976 37.0005
R18407 VDD.n199 VDD.n106 37.0005
R18408 VDD.n99 VDD.n98 37.0005
R18409 VDD.t170 VDD.n99 37.0005
R18410 VDD.n213 VDD.n97 37.0005
R18411 VDD.n216 VDD.n93 37.0005
R18412 VDD.n93 VDD.t838 37.0005
R18413 VDD.n220 VDD.n94 37.0005
R18414 VDD.n90 VDD.n89 37.0005
R18415 VDD.t921 VDD.n90 37.0005
R18416 VDD.n227 VDD.n88 37.0005
R18417 VDD.n79 VDD.n77 37.0005
R18418 VDD.n77 VDD.t1065 37.0005
R18419 VDD.n241 VDD.n78 37.0005
R18420 VDD.n78 VDD.t1065 37.0005
R18421 VDD.n230 VDD.n80 37.0005
R18422 VDD.n80 VDD.t957 37.0005
R18423 VDD.n234 VDD.n81 37.0005
R18424 VDD.n74 VDD.n73 37.0005
R18425 VDD.t878 VDD.n74 37.0005
R18426 VDD.n248 VDD.n72 37.0005
R18427 VDD.n251 VDD.n68 37.0005
R18428 VDD.n68 VDD.t351 37.0005
R18429 VDD.n255 VDD.n69 37.0005
R18430 VDD.n65 VDD.n64 37.0005
R18431 VDD.t646 VDD.n65 37.0005
R18432 VDD.n262 VDD.n63 37.0005
R18433 VDD.n54 VDD.n52 37.0005
R18434 VDD.n52 VDD.t1089 37.0005
R18435 VDD.n276 VDD.n53 37.0005
R18436 VDD.n53 VDD.t1089 37.0005
R18437 VDD.n265 VDD.n55 37.0005
R18438 VDD.n55 VDD.t77 37.0005
R18439 VDD.n269 VDD.n56 37.0005
R18440 VDD.n49 VDD.n48 37.0005
R18441 VDD.t629 VDD.n49 37.0005
R18442 VDD.n283 VDD.n47 37.0005
R18443 VDD.n7506 VDD.n7505 37.0005
R18444 VDD.n7505 VDD.t155 37.0005
R18445 VDD.n7273 VDD.n7272 37.0005
R18446 VDD.n7272 VDD.t155 37.0005
R18447 VDD.n7496 VDD.n7495 37.0005
R18448 VDD.n7495 VDD.t337 37.0005
R18449 VDD.n7283 VDD.n7282 37.0005
R18450 VDD.n7282 VDD.t337 37.0005
R18451 VDD.n7486 VDD.n7485 37.0005
R18452 VDD.n7485 VDD.t911 37.0005
R18453 VDD.n7296 VDD.n7295 37.0005
R18454 VDD.n7295 VDD.t911 37.0005
R18455 VDD.n7476 VDD.n7475 37.0005
R18456 VDD.n7475 VDD.t13 37.0005
R18457 VDD.n7307 VDD.n7306 37.0005
R18458 VDD.n7306 VDD.t13 37.0005
R18459 VDD.n7466 VDD.n7465 37.0005
R18460 VDD.n7465 VDD.t112 37.0005
R18461 VDD.n7317 VDD.n7316 37.0005
R18462 VDD.n7316 VDD.t112 37.0005
R18463 VDD.n7456 VDD.n7455 37.0005
R18464 VDD.n7455 VDD.t948 37.0005
R18465 VDD.n7330 VDD.n7329 37.0005
R18466 VDD.n7329 VDD.t948 37.0005
R18467 VDD.n7334 VDD.n7332 37.0005
R18468 VDD.n7332 VDD.t913 37.0005
R18469 VDD.n7447 VDD.n7333 37.0005
R18470 VDD.n7333 VDD.t913 37.0005
R18471 VDD.n7439 VDD.n7438 37.0005
R18472 VDD.n7438 VDD.t222 37.0005
R18473 VDD.n7345 VDD.n7344 37.0005
R18474 VDD.n7344 VDD.t222 37.0005
R18475 VDD.n7429 VDD.n7428 37.0005
R18476 VDD.n7428 VDD.t48 37.0005
R18477 VDD.n7358 VDD.n7357 37.0005
R18478 VDD.n7357 VDD.t48 37.0005
R18479 VDD.n7419 VDD.n7418 37.0005
R18480 VDD.n7418 VDD.t639 37.0005
R18481 VDD.n7369 VDD.n7368 37.0005
R18482 VDD.n7368 VDD.t639 37.0005
R18483 VDD.n7409 VDD.n7408 37.0005
R18484 VDD.n7408 VDD.t652 37.0005
R18485 VDD.n7379 VDD.n7378 37.0005
R18486 VDD.n7378 VDD.t652 37.0005
R18487 VDD.n7399 VDD.n7398 37.0005
R18488 VDD.n7398 VDD.t544 37.0005
R18489 VDD.n7392 VDD.n7391 37.0005
R18490 VDD.n7391 VDD.t544 37.0005
R18491 VDD.n7267 VDD.n7265 37.0005
R18492 VDD.n7265 VDD.t155 37.0005
R18493 VDD.n7506 VDD.n7266 37.0005
R18494 VDD.n7266 VDD.t155 37.0005
R18495 VDD.n7278 VDD.n7276 37.0005
R18496 VDD.n7276 VDD.t337 37.0005
R18497 VDD.n7496 VDD.n7277 37.0005
R18498 VDD.n7277 VDD.t337 37.0005
R18499 VDD.n7288 VDD.n7286 37.0005
R18500 VDD.n7286 VDD.t911 37.0005
R18501 VDD.n7486 VDD.n7287 37.0005
R18502 VDD.n7287 VDD.t911 37.0005
R18503 VDD.n7301 VDD.n7299 37.0005
R18504 VDD.n7299 VDD.t13 37.0005
R18505 VDD.n7476 VDD.n7300 37.0005
R18506 VDD.n7300 VDD.t13 37.0005
R18507 VDD.n7312 VDD.n7310 37.0005
R18508 VDD.n7310 VDD.t112 37.0005
R18509 VDD.n7466 VDD.n7311 37.0005
R18510 VDD.n7311 VDD.t112 37.0005
R18511 VDD.n7322 VDD.n7320 37.0005
R18512 VDD.n7320 VDD.t948 37.0005
R18513 VDD.n7456 VDD.n7321 37.0005
R18514 VDD.n7321 VDD.t948 37.0005
R18515 VDD.n7338 VDD.n7336 37.0005
R18516 VDD.n7336 VDD.t222 37.0005
R18517 VDD.n7439 VDD.n7337 37.0005
R18518 VDD.n7337 VDD.t222 37.0005
R18519 VDD.n7350 VDD.n7348 37.0005
R18520 VDD.n7348 VDD.t48 37.0005
R18521 VDD.n7429 VDD.n7349 37.0005
R18522 VDD.n7349 VDD.t48 37.0005
R18523 VDD.n7363 VDD.n7361 37.0005
R18524 VDD.n7361 VDD.t639 37.0005
R18525 VDD.n7419 VDD.n7362 37.0005
R18526 VDD.n7362 VDD.t639 37.0005
R18527 VDD.n7374 VDD.n7372 37.0005
R18528 VDD.n7372 VDD.t652 37.0005
R18529 VDD.n7409 VDD.n7373 37.0005
R18530 VDD.n7373 VDD.t652 37.0005
R18531 VDD.n7384 VDD.n7382 37.0005
R18532 VDD.n7382 VDD.t544 37.0005
R18533 VDD.n7399 VDD.n7383 37.0005
R18534 VDD.n7383 VDD.t544 37.0005
R18535 VDD.n7261 VDD.n7260 37.0005
R18536 VDD.t607 VDD.n7261 37.0005
R18537 VDD.n7514 VDD.n7259 37.0005
R18538 VDD.n7246 VDD.n7245 37.0005
R18539 VDD.n7245 VDD.t439 37.0005
R18540 VDD.n1917 VDD.n1916 37.0005
R18541 VDD.n1916 VDD.t439 37.0005
R18542 VDD.n7236 VDD.n7235 37.0005
R18543 VDD.n7235 VDD.t572 37.0005
R18544 VDD.n1927 VDD.n1926 37.0005
R18545 VDD.n1926 VDD.t572 37.0005
R18546 VDD.n7226 VDD.n7225 37.0005
R18547 VDD.n7225 VDD.t1020 37.0005
R18548 VDD.n1940 VDD.n1939 37.0005
R18549 VDD.n1939 VDD.t1020 37.0005
R18550 VDD.n7216 VDD.n7215 37.0005
R18551 VDD.n7215 VDD.t500 37.0005
R18552 VDD.n1952 VDD.n1951 37.0005
R18553 VDD.n1951 VDD.t500 37.0005
R18554 VDD.n1970 VDD.n1969 37.0005
R18555 VDD.n1969 VDD.t149 37.0005
R18556 VDD.n7202 VDD.n7201 37.0005
R18557 VDD.n7201 VDD.t35 37.0005
R18558 VDD.n1980 VDD.n1979 37.0005
R18559 VDD.t35 VDD.n1980 37.0005
R18560 VDD.n1983 VDD.n1981 37.0005
R18561 VDD.n1981 VDD.t1074 37.0005
R18562 VDD.n7190 VDD.n1982 37.0005
R18563 VDD.n1982 VDD.t1074 37.0005
R18564 VDD.n7182 VDD.n7181 37.0005
R18565 VDD.n7181 VDD.t106 37.0005
R18566 VDD.n1994 VDD.n1993 37.0005
R18567 VDD.n1993 VDD.t106 37.0005
R18568 VDD.n7172 VDD.n7171 37.0005
R18569 VDD.n7171 VDD.t29 37.0005
R18570 VDD.n2007 VDD.n2006 37.0005
R18571 VDD.n2006 VDD.t29 37.0005
R18572 VDD.n7162 VDD.n7161 37.0005
R18573 VDD.n7161 VDD.t522 37.0005
R18574 VDD.n2018 VDD.n2017 37.0005
R18575 VDD.n2017 VDD.t522 37.0005
R18576 VDD.n7152 VDD.n7151 37.0005
R18577 VDD.n7151 VDD.t193 37.0005
R18578 VDD.n2028 VDD.n2027 37.0005
R18579 VDD.n2027 VDD.t193 37.0005
R18580 VDD.n7142 VDD.n7141 37.0005
R18581 VDD.n7141 VDD.t546 37.0005
R18582 VDD.n7135 VDD.n7134 37.0005
R18583 VDD.n7134 VDD.t546 37.0005
R18584 VDD.n1905 VDD.n1904 37.0005
R18585 VDD.t649 VDD.n1905 37.0005
R18586 VDD.n7254 VDD.n1903 37.0005
R18587 VDD.n1911 VDD.n1909 37.0005
R18588 VDD.n1909 VDD.t439 37.0005
R18589 VDD.n7246 VDD.n1910 37.0005
R18590 VDD.n1910 VDD.t439 37.0005
R18591 VDD.n1922 VDD.n1920 37.0005
R18592 VDD.n1920 VDD.t572 37.0005
R18593 VDD.n7236 VDD.n1921 37.0005
R18594 VDD.n1921 VDD.t572 37.0005
R18595 VDD.n1932 VDD.n1930 37.0005
R18596 VDD.n1930 VDD.t1020 37.0005
R18597 VDD.n7226 VDD.n1931 37.0005
R18598 VDD.n1931 VDD.t1020 37.0005
R18599 VDD.n1945 VDD.n1943 37.0005
R18600 VDD.n1943 VDD.t500 37.0005
R18601 VDD.n7216 VDD.n1944 37.0005
R18602 VDD.n1944 VDD.t500 37.0005
R18603 VDD.n7200 VDD.n7199 37.0005
R18604 VDD.t35 VDD.n7200 37.0005
R18605 VDD.n7202 VDD.n1965 37.0005
R18606 VDD.t35 VDD.n1965 37.0005
R18607 VDD.n1987 VDD.n1985 37.0005
R18608 VDD.n1985 VDD.t106 37.0005
R18609 VDD.n7182 VDD.n1986 37.0005
R18610 VDD.n1986 VDD.t106 37.0005
R18611 VDD.n1999 VDD.n1997 37.0005
R18612 VDD.n1997 VDD.t29 37.0005
R18613 VDD.n7172 VDD.n1998 37.0005
R18614 VDD.n1998 VDD.t29 37.0005
R18615 VDD.n2012 VDD.n2010 37.0005
R18616 VDD.n2010 VDD.t522 37.0005
R18617 VDD.n7162 VDD.n2011 37.0005
R18618 VDD.n2011 VDD.t522 37.0005
R18619 VDD.n2023 VDD.n2021 37.0005
R18620 VDD.n2021 VDD.t193 37.0005
R18621 VDD.n7152 VDD.n2022 37.0005
R18622 VDD.n2022 VDD.t193 37.0005
R18623 VDD.n2033 VDD.n2031 37.0005
R18624 VDD.n2031 VDD.t546 37.0005
R18625 VDD.n7142 VDD.n2032 37.0005
R18626 VDD.n2032 VDD.t546 37.0005
R18627 VDD.n1957 VDD.n1955 37.0005
R18628 VDD.n1955 VDD.t149 37.0005
R18629 VDD.n7206 VDD.n1960 37.0005
R18630 VDD.n1960 VDD.t149 37.0005
R18631 VDD.n7206 VDD.n1956 37.0005
R18632 VDD.n1956 VDD.t149 37.0005
R18633 VDD.n6995 VDD.n6992 37.0005
R18634 VDD.n6992 VDD.t939 37.0005
R18635 VDD.n6999 VDD.n6993 37.0005
R18636 VDD.n6989 VDD.n6988 37.0005
R18637 VDD.t968 VDD.n6989 37.0005
R18638 VDD.n7006 VDD.n6987 37.0005
R18639 VDD.n6978 VDD.n6976 37.0005
R18640 VDD.n6976 VDD.t954 37.0005
R18641 VDD.n7020 VDD.n6977 37.0005
R18642 VDD.n6977 VDD.t954 37.0005
R18643 VDD.n7009 VDD.n6979 37.0005
R18644 VDD.n6979 VDD.t1036 37.0005
R18645 VDD.n7013 VDD.n6980 37.0005
R18646 VDD.n6973 VDD.n6972 37.0005
R18647 VDD.t931 VDD.n6973 37.0005
R18648 VDD.n7027 VDD.n6971 37.0005
R18649 VDD.n7030 VDD.n6967 37.0005
R18650 VDD.n6967 VDD.t126 37.0005
R18651 VDD.n7034 VDD.n6968 37.0005
R18652 VDD.n6964 VDD.n6963 37.0005
R18653 VDD.t71 VDD.n6964 37.0005
R18654 VDD.n7041 VDD.n6962 37.0005
R18655 VDD.n6953 VDD.n6951 37.0005
R18656 VDD.n6951 VDD.t420 37.0005
R18657 VDD.n7055 VDD.n6952 37.0005
R18658 VDD.n6952 VDD.t420 37.0005
R18659 VDD.n7044 VDD.n6954 37.0005
R18660 VDD.n6954 VDD.t1012 37.0005
R18661 VDD.n7048 VDD.n6955 37.0005
R18662 VDD.n6948 VDD.n6947 37.0005
R18663 VDD.t189 VDD.n6948 37.0005
R18664 VDD.n7062 VDD.n6946 37.0005
R18665 VDD.n7065 VDD.n6942 37.0005
R18666 VDD.n6942 VDD.t798 37.0005
R18667 VDD.n7069 VDD.n6943 37.0005
R18668 VDD.n6939 VDD.n6938 37.0005
R18669 VDD.t791 VDD.n6939 37.0005
R18670 VDD.n7076 VDD.n6937 37.0005
R18671 VDD.n6928 VDD.n6926 37.0005
R18672 VDD.n6926 VDD.t399 37.0005
R18673 VDD.n7090 VDD.n6927 37.0005
R18674 VDD.n6927 VDD.t399 37.0005
R18675 VDD.n7079 VDD.n6929 37.0005
R18676 VDD.n6929 VDD.t1040 37.0005
R18677 VDD.n7083 VDD.n6930 37.0005
R18678 VDD.n6923 VDD.n6922 37.0005
R18679 VDD.t583 VDD.n6923 37.0005
R18680 VDD.n7097 VDD.n6921 37.0005
R18681 VDD.n7100 VDD.n6917 37.0005
R18682 VDD.n6917 VDD.t773 37.0005
R18683 VDD.n7104 VDD.n6918 37.0005
R18684 VDD.n6914 VDD.n6913 37.0005
R18685 VDD.t276 VDD.n6914 37.0005
R18686 VDD.n7111 VDD.n6912 37.0005
R18687 VDD.n7126 VDD.n7125 37.0005
R18688 VDD.n7125 VDD.t950 37.0005
R18689 VDD.n7124 VDD.n7123 37.0005
R18690 VDD.t950 VDD.n7124 37.0005
R18691 VDD.n7114 VDD.n6907 37.0005
R18692 VDD.n6907 VDD.t1008 37.0005
R18693 VDD.n7118 VDD.n6908 37.0005
R18694 VDD.n6902 VDD.n6896 37.0005
R18695 VDD.n6896 VDD.t301 37.0005
R18696 VDD.n6898 VDD.n6895 37.0005
R18697 VDD.n5902 VDD.n5901 37.0005
R18698 VDD.t245 VDD.n5902 37.0005
R18699 VDD.n6134 VDD.n6133 37.0005
R18700 VDD.n6133 VDD.t37 37.0005
R18701 VDD.n5911 VDD.n5910 37.0005
R18702 VDD.n5910 VDD.t37 37.0005
R18703 VDD.n6124 VDD.n6123 37.0005
R18704 VDD.n6123 VDD.t530 37.0005
R18705 VDD.n5921 VDD.n5920 37.0005
R18706 VDD.n5920 VDD.t530 37.0005
R18707 VDD.n6114 VDD.n6113 37.0005
R18708 VDD.n6113 VDD.t56 37.0005
R18709 VDD.n5932 VDD.n5931 37.0005
R18710 VDD.n5931 VDD.t56 37.0005
R18711 VDD.n6104 VDD.n6103 37.0005
R18712 VDD.n6103 VDD.t322 37.0005
R18713 VDD.n5945 VDD.n5944 37.0005
R18714 VDD.n5944 VDD.t322 37.0005
R18715 VDD.n5949 VDD.n5947 37.0005
R18716 VDD.n5947 VDD.t1024 37.0005
R18717 VDD.n6095 VDD.n5948 37.0005
R18718 VDD.n5948 VDD.t1024 37.0005
R18719 VDD.n6087 VDD.n6086 37.0005
R18720 VDD.n6086 VDD.t324 37.0005
R18721 VDD.n5960 VDD.n5959 37.0005
R18722 VDD.n5959 VDD.t324 37.0005
R18723 VDD.n6077 VDD.n6076 37.0005
R18724 VDD.n6076 VDD.t202 37.0005
R18725 VDD.n5973 VDD.n5972 37.0005
R18726 VDD.n5972 VDD.t202 37.0005
R18727 VDD.n6067 VDD.n6066 37.0005
R18728 VDD.n6066 VDD.t534 37.0005
R18729 VDD.n5983 VDD.n5982 37.0005
R18730 VDD.n5982 VDD.t534 37.0005
R18731 VDD.n6057 VDD.n6056 37.0005
R18732 VDD.n6056 VDD.t1000 37.0005
R18733 VDD.n5994 VDD.n5993 37.0005
R18734 VDD.n5993 VDD.t1000 37.0005
R18735 VDD.n6047 VDD.n6046 37.0005
R18736 VDD.n6046 VDD.t185 37.0005
R18737 VDD.n6007 VDD.n6006 37.0005
R18738 VDD.n6006 VDD.t185 37.0005
R18739 VDD.n6037 VDD.n6036 37.0005
R18740 VDD.n6036 VDD.t494 37.0005
R18741 VDD.n6017 VDD.n6016 37.0005
R18742 VDD.n6016 VDD.t494 37.0005
R18743 VDD.n5906 VDD.n5904 37.0005
R18744 VDD.n5904 VDD.t37 37.0005
R18745 VDD.n6134 VDD.n5905 37.0005
R18746 VDD.n5905 VDD.t37 37.0005
R18747 VDD.n5916 VDD.n5914 37.0005
R18748 VDD.n5914 VDD.t530 37.0005
R18749 VDD.n6124 VDD.n5915 37.0005
R18750 VDD.n5915 VDD.t530 37.0005
R18751 VDD.n5926 VDD.n5924 37.0005
R18752 VDD.n5924 VDD.t56 37.0005
R18753 VDD.n6114 VDD.n5925 37.0005
R18754 VDD.n5925 VDD.t56 37.0005
R18755 VDD.n5937 VDD.n5935 37.0005
R18756 VDD.n5935 VDD.t322 37.0005
R18757 VDD.n6104 VDD.n5936 37.0005
R18758 VDD.n5936 VDD.t322 37.0005
R18759 VDD.n5953 VDD.n5951 37.0005
R18760 VDD.n5951 VDD.t324 37.0005
R18761 VDD.n6087 VDD.n5952 37.0005
R18762 VDD.n5952 VDD.t324 37.0005
R18763 VDD.n5965 VDD.n5963 37.0005
R18764 VDD.n5963 VDD.t202 37.0005
R18765 VDD.n6077 VDD.n5964 37.0005
R18766 VDD.n5964 VDD.t202 37.0005
R18767 VDD.n5978 VDD.n5976 37.0005
R18768 VDD.n5976 VDD.t534 37.0005
R18769 VDD.n6067 VDD.n5977 37.0005
R18770 VDD.n5977 VDD.t534 37.0005
R18771 VDD.n5988 VDD.n5986 37.0005
R18772 VDD.n5986 VDD.t1000 37.0005
R18773 VDD.n6057 VDD.n5987 37.0005
R18774 VDD.n5987 VDD.t1000 37.0005
R18775 VDD.n5999 VDD.n5997 37.0005
R18776 VDD.n5997 VDD.t185 37.0005
R18777 VDD.n6047 VDD.n5998 37.0005
R18778 VDD.n5998 VDD.t185 37.0005
R18779 VDD.n6012 VDD.n6010 37.0005
R18780 VDD.n6010 VDD.t494 37.0005
R18781 VDD.n6037 VDD.n6011 37.0005
R18782 VDD.n6011 VDD.t494 37.0005
R18783 VDD.n6021 VDD.n6019 37.0005
R18784 VDD.n6019 VDD.t888 37.0005
R18785 VDD.n6028 VDD.n6020 37.0005
R18786 VDD.n6145 VDD.n6144 37.0005
R18787 VDD.t245 VDD.n6145 37.0005
R18788 VDD.n6147 VDD.n6146 37.0005
R18789 VDD.n6146 VDD.t245 37.0005
R18790 VDD.n6147 VDD.n5894 37.0005
R18791 VDD.t245 VDD.n5894 37.0005
R18792 VDD.n5766 VDD.n5765 37.0005
R18793 VDD.t141 VDD.n5766 37.0005
R18794 VDD.n6257 VDD.n6256 37.0005
R18795 VDD.n6256 VDD.t263 37.0005
R18796 VDD.n5775 VDD.n5774 37.0005
R18797 VDD.n5774 VDD.t263 37.0005
R18798 VDD.n6247 VDD.n6246 37.0005
R18799 VDD.n6246 VDD.t435 37.0005
R18800 VDD.n5785 VDD.n5784 37.0005
R18801 VDD.n5784 VDD.t435 37.0005
R18802 VDD.n6237 VDD.n6236 37.0005
R18803 VDD.n6236 VDD.t827 37.0005
R18804 VDD.n5796 VDD.n5795 37.0005
R18805 VDD.n5795 VDD.t827 37.0005
R18806 VDD.n6227 VDD.n6226 37.0005
R18807 VDD.n6226 VDD.t944 37.0005
R18808 VDD.n5809 VDD.n5808 37.0005
R18809 VDD.n5808 VDD.t944 37.0005
R18810 VDD.n5813 VDD.n5811 37.0005
R18811 VDD.n5811 VDD.t1079 37.0005
R18812 VDD.n6218 VDD.n5812 37.0005
R18813 VDD.n5812 VDD.t1079 37.0005
R18814 VDD.n6210 VDD.n6209 37.0005
R18815 VDD.n6209 VDD.t632 37.0005
R18816 VDD.n5824 VDD.n5823 37.0005
R18817 VDD.n5823 VDD.t632 37.0005
R18818 VDD.n6200 VDD.n6199 37.0005
R18819 VDD.n6199 VDD.t187 37.0005
R18820 VDD.n5837 VDD.n5836 37.0005
R18821 VDD.n5836 VDD.t187 37.0005
R18822 VDD.n6190 VDD.n6189 37.0005
R18823 VDD.n6189 VDD.t471 37.0005
R18824 VDD.n5847 VDD.n5846 37.0005
R18825 VDD.n5846 VDD.t471 37.0005
R18826 VDD.n6180 VDD.n6179 37.0005
R18827 VDD.n6179 VDD.t1056 37.0005
R18828 VDD.n5858 VDD.n5857 37.0005
R18829 VDD.n5857 VDD.t1056 37.0005
R18830 VDD.n6170 VDD.n6169 37.0005
R18831 VDD.n6169 VDD.t341 37.0005
R18832 VDD.n5871 VDD.n5870 37.0005
R18833 VDD.n5870 VDD.t341 37.0005
R18834 VDD.n6160 VDD.n6159 37.0005
R18835 VDD.n6159 VDD.t516 37.0005
R18836 VDD.n5881 VDD.n5880 37.0005
R18837 VDD.n5880 VDD.t516 37.0005
R18838 VDD.n5770 VDD.n5768 37.0005
R18839 VDD.n5768 VDD.t263 37.0005
R18840 VDD.n6257 VDD.n5769 37.0005
R18841 VDD.n5769 VDD.t263 37.0005
R18842 VDD.n5780 VDD.n5778 37.0005
R18843 VDD.n5778 VDD.t435 37.0005
R18844 VDD.n6247 VDD.n5779 37.0005
R18845 VDD.n5779 VDD.t435 37.0005
R18846 VDD.n5790 VDD.n5788 37.0005
R18847 VDD.n5788 VDD.t827 37.0005
R18848 VDD.n6237 VDD.n5789 37.0005
R18849 VDD.n5789 VDD.t827 37.0005
R18850 VDD.n5801 VDD.n5799 37.0005
R18851 VDD.n5799 VDD.t944 37.0005
R18852 VDD.n6227 VDD.n5800 37.0005
R18853 VDD.n5800 VDD.t944 37.0005
R18854 VDD.n5817 VDD.n5815 37.0005
R18855 VDD.n5815 VDD.t632 37.0005
R18856 VDD.n6210 VDD.n5816 37.0005
R18857 VDD.n5816 VDD.t632 37.0005
R18858 VDD.n5829 VDD.n5827 37.0005
R18859 VDD.n5827 VDD.t187 37.0005
R18860 VDD.n6200 VDD.n5828 37.0005
R18861 VDD.n5828 VDD.t187 37.0005
R18862 VDD.n5842 VDD.n5840 37.0005
R18863 VDD.n5840 VDD.t471 37.0005
R18864 VDD.n6190 VDD.n5841 37.0005
R18865 VDD.n5841 VDD.t471 37.0005
R18866 VDD.n5852 VDD.n5850 37.0005
R18867 VDD.n5850 VDD.t1056 37.0005
R18868 VDD.n6180 VDD.n5851 37.0005
R18869 VDD.n5851 VDD.t1056 37.0005
R18870 VDD.n5863 VDD.n5861 37.0005
R18871 VDD.n5861 VDD.t341 37.0005
R18872 VDD.n6170 VDD.n5862 37.0005
R18873 VDD.n5862 VDD.t341 37.0005
R18874 VDD.n5876 VDD.n5874 37.0005
R18875 VDD.n5874 VDD.t516 37.0005
R18876 VDD.n6160 VDD.n5875 37.0005
R18877 VDD.n5875 VDD.t516 37.0005
R18878 VDD.n5885 VDD.n5883 37.0005
R18879 VDD.n5883 VDD.t881 37.0005
R18880 VDD.n6151 VDD.n5884 37.0005
R18881 VDD.n6268 VDD.n6267 37.0005
R18882 VDD.t141 VDD.n6268 37.0005
R18883 VDD.n6270 VDD.n6269 37.0005
R18884 VDD.n6269 VDD.t141 37.0005
R18885 VDD.n6270 VDD.n5758 37.0005
R18886 VDD.t141 VDD.n5758 37.0005
R18887 VDD.n5630 VDD.n5629 37.0005
R18888 VDD.t364 VDD.n5630 37.0005
R18889 VDD.n6380 VDD.n6379 37.0005
R18890 VDD.n6379 VDD.t109 37.0005
R18891 VDD.n5639 VDD.n5638 37.0005
R18892 VDD.n5638 VDD.t109 37.0005
R18893 VDD.n6370 VDD.n6369 37.0005
R18894 VDD.n6369 VDD.t506 37.0005
R18895 VDD.n5649 VDD.n5648 37.0005
R18896 VDD.n5648 VDD.t506 37.0005
R18897 VDD.n6360 VDD.n6359 37.0005
R18898 VDD.n6359 VDD.t552 37.0005
R18899 VDD.n5660 VDD.n5659 37.0005
R18900 VDD.n5659 VDD.t552 37.0005
R18901 VDD.n6350 VDD.n6349 37.0005
R18902 VDD.n6349 VDD.t145 37.0005
R18903 VDD.n5673 VDD.n5672 37.0005
R18904 VDD.n5672 VDD.t145 37.0005
R18905 VDD.n5677 VDD.n5675 37.0005
R18906 VDD.n5675 VDD.t1054 37.0005
R18907 VDD.n6341 VDD.n5676 37.0005
R18908 VDD.n5676 VDD.t1054 37.0005
R18909 VDD.n6333 VDD.n6332 37.0005
R18910 VDD.n6332 VDD.t147 37.0005
R18911 VDD.n5688 VDD.n5687 37.0005
R18912 VDD.n5687 VDD.t147 37.0005
R18913 VDD.n6323 VDD.n6322 37.0005
R18914 VDD.n6322 VDD.t116 37.0005
R18915 VDD.n5701 VDD.n5700 37.0005
R18916 VDD.n5700 VDD.t116 37.0005
R18917 VDD.n6313 VDD.n6312 37.0005
R18918 VDD.n6312 VDD.t453 37.0005
R18919 VDD.n5711 VDD.n5710 37.0005
R18920 VDD.n5710 VDD.t453 37.0005
R18921 VDD.n6303 VDD.n6302 37.0005
R18922 VDD.n6302 VDD.t1028 37.0005
R18923 VDD.n5722 VDD.n5721 37.0005
R18924 VDD.n5721 VDD.t1028 37.0005
R18925 VDD.n6293 VDD.n6292 37.0005
R18926 VDD.n6292 VDD.t368 37.0005
R18927 VDD.n5735 VDD.n5734 37.0005
R18928 VDD.n5734 VDD.t368 37.0005
R18929 VDD.n6283 VDD.n6282 37.0005
R18930 VDD.n6282 VDD.t463 37.0005
R18931 VDD.n5745 VDD.n5744 37.0005
R18932 VDD.n5744 VDD.t463 37.0005
R18933 VDD.n5634 VDD.n5632 37.0005
R18934 VDD.n5632 VDD.t109 37.0005
R18935 VDD.n6380 VDD.n5633 37.0005
R18936 VDD.n5633 VDD.t109 37.0005
R18937 VDD.n5644 VDD.n5642 37.0005
R18938 VDD.n5642 VDD.t506 37.0005
R18939 VDD.n6370 VDD.n5643 37.0005
R18940 VDD.n5643 VDD.t506 37.0005
R18941 VDD.n5654 VDD.n5652 37.0005
R18942 VDD.n5652 VDD.t552 37.0005
R18943 VDD.n6360 VDD.n5653 37.0005
R18944 VDD.n5653 VDD.t552 37.0005
R18945 VDD.n5665 VDD.n5663 37.0005
R18946 VDD.n5663 VDD.t145 37.0005
R18947 VDD.n6350 VDD.n5664 37.0005
R18948 VDD.n5664 VDD.t145 37.0005
R18949 VDD.n5681 VDD.n5679 37.0005
R18950 VDD.n5679 VDD.t147 37.0005
R18951 VDD.n6333 VDD.n5680 37.0005
R18952 VDD.n5680 VDD.t147 37.0005
R18953 VDD.n5693 VDD.n5691 37.0005
R18954 VDD.n5691 VDD.t116 37.0005
R18955 VDD.n6323 VDD.n5692 37.0005
R18956 VDD.n5692 VDD.t116 37.0005
R18957 VDD.n5706 VDD.n5704 37.0005
R18958 VDD.n5704 VDD.t453 37.0005
R18959 VDD.n6313 VDD.n5705 37.0005
R18960 VDD.n5705 VDD.t453 37.0005
R18961 VDD.n5716 VDD.n5714 37.0005
R18962 VDD.n5714 VDD.t1028 37.0005
R18963 VDD.n6303 VDD.n5715 37.0005
R18964 VDD.n5715 VDD.t1028 37.0005
R18965 VDD.n5727 VDD.n5725 37.0005
R18966 VDD.n5725 VDD.t368 37.0005
R18967 VDD.n6293 VDD.n5726 37.0005
R18968 VDD.n5726 VDD.t368 37.0005
R18969 VDD.n5740 VDD.n5738 37.0005
R18970 VDD.n5738 VDD.t463 37.0005
R18971 VDD.n6283 VDD.n5739 37.0005
R18972 VDD.n5739 VDD.t463 37.0005
R18973 VDD.n5749 VDD.n5747 37.0005
R18974 VDD.n5747 VDD.t916 37.0005
R18975 VDD.n6274 VDD.n5748 37.0005
R18976 VDD.n6391 VDD.n6390 37.0005
R18977 VDD.t364 VDD.n6391 37.0005
R18978 VDD.n6393 VDD.n6392 37.0005
R18979 VDD.n6392 VDD.t364 37.0005
R18980 VDD.n6393 VDD.n5622 37.0005
R18981 VDD.t364 VDD.n5622 37.0005
R18982 VDD.n5494 VDD.n5493 37.0005
R18983 VDD.t46 VDD.n5494 37.0005
R18984 VDD.n6503 VDD.n6502 37.0005
R18985 VDD.n6502 VDD.t253 37.0005
R18986 VDD.n5503 VDD.n5502 37.0005
R18987 VDD.n5502 VDD.t253 37.0005
R18988 VDD.n6493 VDD.n6492 37.0005
R18989 VDD.n6492 VDD.t459 37.0005
R18990 VDD.n5513 VDD.n5512 37.0005
R18991 VDD.n5512 VDD.t459 37.0005
R18992 VDD.n6483 VDD.n6482 37.0005
R18993 VDD.n6482 VDD.t237 37.0005
R18994 VDD.n5524 VDD.n5523 37.0005
R18995 VDD.n5523 VDD.t237 37.0005
R18996 VDD.n6473 VDD.n6472 37.0005
R18997 VDD.n6472 VDD.t257 37.0005
R18998 VDD.n5537 VDD.n5536 37.0005
R18999 VDD.n5536 VDD.t257 37.0005
R19000 VDD.n5541 VDD.n5539 37.0005
R19001 VDD.n5539 VDD.t1096 37.0005
R19002 VDD.n6464 VDD.n5540 37.0005
R19003 VDD.n5540 VDD.t1096 37.0005
R19004 VDD.n6456 VDD.n6455 37.0005
R19005 VDD.n6455 VDD.t135 37.0005
R19006 VDD.n5552 VDD.n5551 37.0005
R19007 VDD.n5551 VDD.t135 37.0005
R19008 VDD.n6446 VDD.n6445 37.0005
R19009 VDD.n6445 VDD.t794 37.0005
R19010 VDD.n5565 VDD.n5564 37.0005
R19011 VDD.n5564 VDD.t794 37.0005
R19012 VDD.n6436 VDD.n6435 37.0005
R19013 VDD.n6435 VDD.t490 37.0005
R19014 VDD.n5575 VDD.n5574 37.0005
R19015 VDD.n5574 VDD.t490 37.0005
R19016 VDD.n6426 VDD.n6425 37.0005
R19017 VDD.n6425 VDD.t1002 37.0005
R19018 VDD.n5586 VDD.n5585 37.0005
R19019 VDD.n5585 VDD.t1002 37.0005
R19020 VDD.n6416 VDD.n6415 37.0005
R19021 VDD.n6415 VDD.t871 37.0005
R19022 VDD.n5599 VDD.n5598 37.0005
R19023 VDD.n5598 VDD.t871 37.0005
R19024 VDD.n6406 VDD.n6405 37.0005
R19025 VDD.n6405 VDD.t443 37.0005
R19026 VDD.n5609 VDD.n5608 37.0005
R19027 VDD.n5608 VDD.t443 37.0005
R19028 VDD.n5498 VDD.n5496 37.0005
R19029 VDD.n5496 VDD.t253 37.0005
R19030 VDD.n6503 VDD.n5497 37.0005
R19031 VDD.n5497 VDD.t253 37.0005
R19032 VDD.n5508 VDD.n5506 37.0005
R19033 VDD.n5506 VDD.t459 37.0005
R19034 VDD.n6493 VDD.n5507 37.0005
R19035 VDD.n5507 VDD.t459 37.0005
R19036 VDD.n5518 VDD.n5516 37.0005
R19037 VDD.n5516 VDD.t237 37.0005
R19038 VDD.n6483 VDD.n5517 37.0005
R19039 VDD.n5517 VDD.t237 37.0005
R19040 VDD.n5529 VDD.n5527 37.0005
R19041 VDD.n5527 VDD.t257 37.0005
R19042 VDD.n6473 VDD.n5528 37.0005
R19043 VDD.n5528 VDD.t257 37.0005
R19044 VDD.n5545 VDD.n5543 37.0005
R19045 VDD.n5543 VDD.t135 37.0005
R19046 VDD.n6456 VDD.n5544 37.0005
R19047 VDD.n5544 VDD.t135 37.0005
R19048 VDD.n5557 VDD.n5555 37.0005
R19049 VDD.n5555 VDD.t794 37.0005
R19050 VDD.n6446 VDD.n5556 37.0005
R19051 VDD.n5556 VDD.t794 37.0005
R19052 VDD.n5570 VDD.n5568 37.0005
R19053 VDD.n5568 VDD.t490 37.0005
R19054 VDD.n6436 VDD.n5569 37.0005
R19055 VDD.n5569 VDD.t490 37.0005
R19056 VDD.n5580 VDD.n5578 37.0005
R19057 VDD.n5578 VDD.t1002 37.0005
R19058 VDD.n6426 VDD.n5579 37.0005
R19059 VDD.n5579 VDD.t1002 37.0005
R19060 VDD.n5591 VDD.n5589 37.0005
R19061 VDD.n5589 VDD.t871 37.0005
R19062 VDD.n6416 VDD.n5590 37.0005
R19063 VDD.n5590 VDD.t871 37.0005
R19064 VDD.n5604 VDD.n5602 37.0005
R19065 VDD.n5602 VDD.t443 37.0005
R19066 VDD.n6406 VDD.n5603 37.0005
R19067 VDD.n5603 VDD.t443 37.0005
R19068 VDD.n5613 VDD.n5611 37.0005
R19069 VDD.n5611 VDD.t621 37.0005
R19070 VDD.n6397 VDD.n5612 37.0005
R19071 VDD.n6514 VDD.n6513 37.0005
R19072 VDD.t46 VDD.n6514 37.0005
R19073 VDD.n6516 VDD.n6515 37.0005
R19074 VDD.n6515 VDD.t46 37.0005
R19075 VDD.n6516 VDD.n5486 37.0005
R19076 VDD.t46 VDD.n5486 37.0005
R19077 VDD.n5358 VDD.n5357 37.0005
R19078 VDD.t312 VDD.n5358 37.0005
R19079 VDD.n6626 VDD.n6625 37.0005
R19080 VDD.n6625 VDD.t33 37.0005
R19081 VDD.n5367 VDD.n5366 37.0005
R19082 VDD.n5366 VDD.t33 37.0005
R19083 VDD.n6616 VDD.n6615 37.0005
R19084 VDD.n6615 VDD.t492 37.0005
R19085 VDD.n5377 VDD.n5376 37.0005
R19086 VDD.n5376 VDD.t492 37.0005
R19087 VDD.n6606 VDD.n6605 37.0005
R19088 VDD.n6605 VDD.t139 37.0005
R19089 VDD.n5388 VDD.n5387 37.0005
R19090 VDD.n5387 VDD.t139 37.0005
R19091 VDD.n6596 VDD.n6595 37.0005
R19092 VDD.n6595 VDD.t208 37.0005
R19093 VDD.n5401 VDD.n5400 37.0005
R19094 VDD.n5400 VDD.t208 37.0005
R19095 VDD.n5405 VDD.n5403 37.0005
R19096 VDD.n5403 VDD.t1084 37.0005
R19097 VDD.n6587 VDD.n5404 37.0005
R19098 VDD.n5404 VDD.t1084 37.0005
R19099 VDD.n6579 VDD.n6578 37.0005
R19100 VDD.n6578 VDD.t280 37.0005
R19101 VDD.n5416 VDD.n5415 37.0005
R19102 VDD.n5415 VDD.t280 37.0005
R19103 VDD.n6569 VDD.n6568 37.0005
R19104 VDD.n6568 VDD.t17 37.0005
R19105 VDD.n5429 VDD.n5428 37.0005
R19106 VDD.n5428 VDD.t17 37.0005
R19107 VDD.n6559 VDD.n6558 37.0005
R19108 VDD.n6558 VDD.t475 37.0005
R19109 VDD.n5439 VDD.n5438 37.0005
R19110 VDD.n5438 VDD.t475 37.0005
R19111 VDD.n6549 VDD.n6548 37.0005
R19112 VDD.n6548 VDD.t1060 37.0005
R19113 VDD.n5450 VDD.n5449 37.0005
R19114 VDD.n5449 VDD.t1060 37.0005
R19115 VDD.n6539 VDD.n6538 37.0005
R19116 VDD.n6538 VDD.t425 37.0005
R19117 VDD.n5463 VDD.n5462 37.0005
R19118 VDD.n5462 VDD.t425 37.0005
R19119 VDD.n6529 VDD.n6528 37.0005
R19120 VDD.n6528 VDD.t478 37.0005
R19121 VDD.n5473 VDD.n5472 37.0005
R19122 VDD.n5472 VDD.t478 37.0005
R19123 VDD.n5362 VDD.n5360 37.0005
R19124 VDD.n5360 VDD.t33 37.0005
R19125 VDD.n6626 VDD.n5361 37.0005
R19126 VDD.n5361 VDD.t33 37.0005
R19127 VDD.n5372 VDD.n5370 37.0005
R19128 VDD.n5370 VDD.t492 37.0005
R19129 VDD.n6616 VDD.n5371 37.0005
R19130 VDD.n5371 VDD.t492 37.0005
R19131 VDD.n5382 VDD.n5380 37.0005
R19132 VDD.n5380 VDD.t139 37.0005
R19133 VDD.n6606 VDD.n5381 37.0005
R19134 VDD.n5381 VDD.t139 37.0005
R19135 VDD.n5393 VDD.n5391 37.0005
R19136 VDD.n5391 VDD.t208 37.0005
R19137 VDD.n6596 VDD.n5392 37.0005
R19138 VDD.n5392 VDD.t208 37.0005
R19139 VDD.n5409 VDD.n5407 37.0005
R19140 VDD.n5407 VDD.t280 37.0005
R19141 VDD.n6579 VDD.n5408 37.0005
R19142 VDD.n5408 VDD.t280 37.0005
R19143 VDD.n5421 VDD.n5419 37.0005
R19144 VDD.n5419 VDD.t17 37.0005
R19145 VDD.n6569 VDD.n5420 37.0005
R19146 VDD.n5420 VDD.t17 37.0005
R19147 VDD.n5434 VDD.n5432 37.0005
R19148 VDD.n5432 VDD.t475 37.0005
R19149 VDD.n6559 VDD.n5433 37.0005
R19150 VDD.n5433 VDD.t475 37.0005
R19151 VDD.n5444 VDD.n5442 37.0005
R19152 VDD.n5442 VDD.t1060 37.0005
R19153 VDD.n6549 VDD.n5443 37.0005
R19154 VDD.n5443 VDD.t1060 37.0005
R19155 VDD.n5455 VDD.n5453 37.0005
R19156 VDD.n5453 VDD.t425 37.0005
R19157 VDD.n6539 VDD.n5454 37.0005
R19158 VDD.n5454 VDD.t425 37.0005
R19159 VDD.n5468 VDD.n5466 37.0005
R19160 VDD.n5466 VDD.t478 37.0005
R19161 VDD.n6529 VDD.n5467 37.0005
R19162 VDD.n5467 VDD.t478 37.0005
R19163 VDD.n5477 VDD.n5475 37.0005
R19164 VDD.n5475 VDD.t23 37.0005
R19165 VDD.n6520 VDD.n5476 37.0005
R19166 VDD.n6637 VDD.n6636 37.0005
R19167 VDD.t312 VDD.n6637 37.0005
R19168 VDD.n6639 VDD.n6638 37.0005
R19169 VDD.n6638 VDD.t312 37.0005
R19170 VDD.n6639 VDD.n5350 37.0005
R19171 VDD.t312 VDD.n5350 37.0005
R19172 VDD.n5222 VDD.n5221 37.0005
R19173 VDD.t305 VDD.n5222 37.0005
R19174 VDD.n6749 VDD.n6748 37.0005
R19175 VDD.n6748 VDD.t320 37.0005
R19176 VDD.n5231 VDD.n5230 37.0005
R19177 VDD.n5230 VDD.t320 37.0005
R19178 VDD.n6739 VDD.n6738 37.0005
R19179 VDD.n6738 VDD.t482 37.0005
R19180 VDD.n5241 VDD.n5240 37.0005
R19181 VDD.n5240 VDD.t482 37.0005
R19182 VDD.n6729 VDD.n6728 37.0005
R19183 VDD.n6728 VDD.t378 37.0005
R19184 VDD.n5252 VDD.n5251 37.0005
R19185 VDD.n5251 VDD.t378 37.0005
R19186 VDD.n6719 VDD.n6718 37.0005
R19187 VDD.n6718 VDD.t316 37.0005
R19188 VDD.n5265 VDD.n5264 37.0005
R19189 VDD.n5264 VDD.t316 37.0005
R19190 VDD.n5269 VDD.n5267 37.0005
R19191 VDD.n5267 VDD.t1058 37.0005
R19192 VDD.n6710 VDD.n5268 37.0005
R19193 VDD.n5268 VDD.t1058 37.0005
R19194 VDD.n6702 VDD.n6701 37.0005
R19195 VDD.n6701 VDD.t314 37.0005
R19196 VDD.n5280 VDD.n5279 37.0005
R19197 VDD.n5279 VDD.t314 37.0005
R19198 VDD.n6692 VDD.n6691 37.0005
R19199 VDD.n6691 VDD.t366 37.0005
R19200 VDD.n5293 VDD.n5292 37.0005
R19201 VDD.n5292 VDD.t366 37.0005
R19202 VDD.n6682 VDD.n6681 37.0005
R19203 VDD.n6681 VDD.t520 37.0005
R19204 VDD.n5303 VDD.n5302 37.0005
R19205 VDD.n5302 VDD.t520 37.0005
R19206 VDD.n6672 VDD.n6671 37.0005
R19207 VDD.n6671 VDD.t1032 37.0005
R19208 VDD.n5314 VDD.n5313 37.0005
R19209 VDD.n5313 VDD.t1032 37.0005
R19210 VDD.n6662 VDD.n6661 37.0005
R19211 VDD.n6661 VDD.t835 37.0005
R19212 VDD.n5327 VDD.n5326 37.0005
R19213 VDD.n5326 VDD.t835 37.0005
R19214 VDD.n6652 VDD.n6651 37.0005
R19215 VDD.n6651 VDD.t465 37.0005
R19216 VDD.n5337 VDD.n5336 37.0005
R19217 VDD.n5336 VDD.t465 37.0005
R19218 VDD.n5226 VDD.n5224 37.0005
R19219 VDD.n5224 VDD.t320 37.0005
R19220 VDD.n6749 VDD.n5225 37.0005
R19221 VDD.n5225 VDD.t320 37.0005
R19222 VDD.n5236 VDD.n5234 37.0005
R19223 VDD.n5234 VDD.t482 37.0005
R19224 VDD.n6739 VDD.n5235 37.0005
R19225 VDD.n5235 VDD.t482 37.0005
R19226 VDD.n5246 VDD.n5244 37.0005
R19227 VDD.n5244 VDD.t378 37.0005
R19228 VDD.n6729 VDD.n5245 37.0005
R19229 VDD.n5245 VDD.t378 37.0005
R19230 VDD.n5257 VDD.n5255 37.0005
R19231 VDD.n5255 VDD.t316 37.0005
R19232 VDD.n6719 VDD.n5256 37.0005
R19233 VDD.n5256 VDD.t316 37.0005
R19234 VDD.n5273 VDD.n5271 37.0005
R19235 VDD.n5271 VDD.t314 37.0005
R19236 VDD.n6702 VDD.n5272 37.0005
R19237 VDD.n5272 VDD.t314 37.0005
R19238 VDD.n5285 VDD.n5283 37.0005
R19239 VDD.n5283 VDD.t366 37.0005
R19240 VDD.n6692 VDD.n5284 37.0005
R19241 VDD.n5284 VDD.t366 37.0005
R19242 VDD.n5298 VDD.n5296 37.0005
R19243 VDD.n5296 VDD.t520 37.0005
R19244 VDD.n6682 VDD.n5297 37.0005
R19245 VDD.n5297 VDD.t520 37.0005
R19246 VDD.n5308 VDD.n5306 37.0005
R19247 VDD.n5306 VDD.t1032 37.0005
R19248 VDD.n6672 VDD.n5307 37.0005
R19249 VDD.n5307 VDD.t1032 37.0005
R19250 VDD.n5319 VDD.n5317 37.0005
R19251 VDD.n5317 VDD.t835 37.0005
R19252 VDD.n6662 VDD.n5318 37.0005
R19253 VDD.n5318 VDD.t835 37.0005
R19254 VDD.n5332 VDD.n5330 37.0005
R19255 VDD.n5330 VDD.t465 37.0005
R19256 VDD.n6652 VDD.n5331 37.0005
R19257 VDD.n5331 VDD.t465 37.0005
R19258 VDD.n5341 VDD.n5339 37.0005
R19259 VDD.n5339 VDD.t840 37.0005
R19260 VDD.n6643 VDD.n5340 37.0005
R19261 VDD.n6760 VDD.n6759 37.0005
R19262 VDD.t305 VDD.n6760 37.0005
R19263 VDD.n6762 VDD.n6761 37.0005
R19264 VDD.n6761 VDD.t305 37.0005
R19265 VDD.n6762 VDD.n5214 37.0005
R19266 VDD.t305 VDD.n5214 37.0005
R19267 VDD.n5086 VDD.n5085 37.0005
R19268 VDD.t349 VDD.n5086 37.0005
R19269 VDD.n6872 VDD.n6871 37.0005
R19270 VDD.n6871 VDD.t431 37.0005
R19271 VDD.n5095 VDD.n5094 37.0005
R19272 VDD.n5094 VDD.t431 37.0005
R19273 VDD.n6862 VDD.n6861 37.0005
R19274 VDD.n6861 VDD.t433 37.0005
R19275 VDD.n5105 VDD.n5104 37.0005
R19276 VDD.n5104 VDD.t433 37.0005
R19277 VDD.n6852 VDD.n6851 37.0005
R19278 VDD.n6851 VDD.t330 37.0005
R19279 VDD.n5116 VDD.n5115 37.0005
R19280 VDD.n5115 VDD.t330 37.0005
R19281 VDD.n6842 VDD.n6841 37.0005
R19282 VDD.n6841 VDD.t228 37.0005
R19283 VDD.n5129 VDD.n5128 37.0005
R19284 VDD.n5128 VDD.t228 37.0005
R19285 VDD.n5133 VDD.n5131 37.0005
R19286 VDD.n5131 VDD.t1076 37.0005
R19287 VDD.n6833 VDD.n5132 37.0005
R19288 VDD.n5132 VDD.t1076 37.0005
R19289 VDD.n6825 VDD.n6824 37.0005
R19290 VDD.n6824 VDD.t226 37.0005
R19291 VDD.n5144 VDD.n5143 37.0005
R19292 VDD.n5143 VDD.t226 37.0005
R19293 VDD.n6815 VDD.n6814 37.0005
R19294 VDD.n6814 VDD.t162 37.0005
R19295 VDD.n5157 VDD.n5156 37.0005
R19296 VDD.n5156 VDD.t162 37.0005
R19297 VDD.n6805 VDD.n6804 37.0005
R19298 VDD.n6804 VDD.t510 37.0005
R19299 VDD.n5167 VDD.n5166 37.0005
R19300 VDD.n5166 VDD.t510 37.0005
R19301 VDD.n6795 VDD.n6794 37.0005
R19302 VDD.n6794 VDD.t1030 37.0005
R19303 VDD.n5178 VDD.n5177 37.0005
R19304 VDD.n5177 VDD.t1030 37.0005
R19305 VDD.n6785 VDD.n6784 37.0005
R19306 VDD.n6784 VDD.t390 37.0005
R19307 VDD.n5191 VDD.n5190 37.0005
R19308 VDD.n5190 VDD.t390 37.0005
R19309 VDD.n6775 VDD.n6774 37.0005
R19310 VDD.n6774 VDD.t457 37.0005
R19311 VDD.n5201 VDD.n5200 37.0005
R19312 VDD.n5200 VDD.t457 37.0005
R19313 VDD.n5090 VDD.n5088 37.0005
R19314 VDD.n5088 VDD.t431 37.0005
R19315 VDD.n6872 VDD.n5089 37.0005
R19316 VDD.n5089 VDD.t431 37.0005
R19317 VDD.n5100 VDD.n5098 37.0005
R19318 VDD.n5098 VDD.t433 37.0005
R19319 VDD.n6862 VDD.n5099 37.0005
R19320 VDD.n5099 VDD.t433 37.0005
R19321 VDD.n5110 VDD.n5108 37.0005
R19322 VDD.n5108 VDD.t330 37.0005
R19323 VDD.n6852 VDD.n5109 37.0005
R19324 VDD.n5109 VDD.t330 37.0005
R19325 VDD.n5121 VDD.n5119 37.0005
R19326 VDD.n5119 VDD.t228 37.0005
R19327 VDD.n6842 VDD.n5120 37.0005
R19328 VDD.n5120 VDD.t228 37.0005
R19329 VDD.n5137 VDD.n5135 37.0005
R19330 VDD.n5135 VDD.t226 37.0005
R19331 VDD.n6825 VDD.n5136 37.0005
R19332 VDD.n5136 VDD.t226 37.0005
R19333 VDD.n5149 VDD.n5147 37.0005
R19334 VDD.n5147 VDD.t162 37.0005
R19335 VDD.n6815 VDD.n5148 37.0005
R19336 VDD.n5148 VDD.t162 37.0005
R19337 VDD.n5162 VDD.n5160 37.0005
R19338 VDD.n5160 VDD.t510 37.0005
R19339 VDD.n6805 VDD.n5161 37.0005
R19340 VDD.n5161 VDD.t510 37.0005
R19341 VDD.n5172 VDD.n5170 37.0005
R19342 VDD.n5170 VDD.t1030 37.0005
R19343 VDD.n6795 VDD.n5171 37.0005
R19344 VDD.n5171 VDD.t1030 37.0005
R19345 VDD.n5183 VDD.n5181 37.0005
R19346 VDD.n5181 VDD.t390 37.0005
R19347 VDD.n6785 VDD.n5182 37.0005
R19348 VDD.n5182 VDD.t390 37.0005
R19349 VDD.n5196 VDD.n5194 37.0005
R19350 VDD.n5194 VDD.t457 37.0005
R19351 VDD.n6775 VDD.n5195 37.0005
R19352 VDD.n5195 VDD.t457 37.0005
R19353 VDD.n5205 VDD.n5203 37.0005
R19354 VDD.n5203 VDD.t919 37.0005
R19355 VDD.n6766 VDD.n5204 37.0005
R19356 VDD.n6883 VDD.n6882 37.0005
R19357 VDD.t349 VDD.n6883 37.0005
R19358 VDD.n6885 VDD.n6884 37.0005
R19359 VDD.n6884 VDD.t349 37.0005
R19360 VDD.n6885 VDD.n5078 37.0005
R19361 VDD.t349 VDD.n5078 37.0005
R19362 VDD.n4944 VDD.n4943 37.0005
R19363 VDD.n4943 VDD.t183 37.0005
R19364 VDD.n4964 VDD.n4963 37.0005
R19365 VDD.n4963 VDD.t181 37.0005
R19366 VDD.n4935 VDD.n4934 37.0005
R19367 VDD.n4934 VDD.t181 37.0005
R19368 VDD.n4974 VDD.n4973 37.0005
R19369 VDD.n4973 VDD.t512 37.0005
R19370 VDD.n4925 VDD.n4924 37.0005
R19371 VDD.n4924 VDD.t512 37.0005
R19372 VDD.n4984 VDD.n4983 37.0005
R19373 VDD.n4983 VDD.t380 37.0005
R19374 VDD.n4914 VDD.n4913 37.0005
R19375 VDD.n4913 VDD.t380 37.0005
R19376 VDD.n4994 VDD.n4993 37.0005
R19377 VDD.n4993 VDD.t118 37.0005
R19378 VDD.n4901 VDD.n4900 37.0005
R19379 VDD.n4900 VDD.t118 37.0005
R19380 VDD.n4890 VDD.n4888 37.0005
R19381 VDD.n4888 VDD.t1052 37.0005
R19382 VDD.n5002 VDD.n4889 37.0005
R19383 VDD.n4889 VDD.t1052 37.0005
R19384 VDD.n5011 VDD.n5010 37.0005
R19385 VDD.n5010 VDD.t84 37.0005
R19386 VDD.n4886 VDD.n4885 37.0005
R19387 VDD.n4885 VDD.t84 37.0005
R19388 VDD.n5021 VDD.n5020 37.0005
R19389 VDD.n5020 VDD.t259 37.0005
R19390 VDD.n4873 VDD.n4872 37.0005
R19391 VDD.n4872 VDD.t259 37.0005
R19392 VDD.n5031 VDD.n5030 37.0005
R19393 VDD.n5030 VDD.t486 37.0005
R19394 VDD.n4863 VDD.n4862 37.0005
R19395 VDD.n4862 VDD.t486 37.0005
R19396 VDD.n5041 VDD.n5040 37.0005
R19397 VDD.n5040 VDD.t1004 37.0005
R19398 VDD.n4852 VDD.n4851 37.0005
R19399 VDD.n4851 VDD.t1004 37.0005
R19400 VDD.n5051 VDD.n5050 37.0005
R19401 VDD.n5050 VDD.t289 37.0005
R19402 VDD.n4839 VDD.n4838 37.0005
R19403 VDD.n4838 VDD.t289 37.0005
R19404 VDD.n5061 VDD.n5060 37.0005
R19405 VDD.n5060 VDD.t496 37.0005
R19406 VDD.n4829 VDD.n4828 37.0005
R19407 VDD.n4828 VDD.t496 37.0005
R19408 VDD.n4930 VDD.n4928 37.0005
R19409 VDD.n4928 VDD.t181 37.0005
R19410 VDD.n4964 VDD.n4929 37.0005
R19411 VDD.n4929 VDD.t181 37.0005
R19412 VDD.n4919 VDD.n4917 37.0005
R19413 VDD.n4917 VDD.t512 37.0005
R19414 VDD.n4974 VDD.n4918 37.0005
R19415 VDD.n4918 VDD.t512 37.0005
R19416 VDD.n4906 VDD.n4904 37.0005
R19417 VDD.n4904 VDD.t380 37.0005
R19418 VDD.n4984 VDD.n4905 37.0005
R19419 VDD.n4905 VDD.t380 37.0005
R19420 VDD.n4894 VDD.n4892 37.0005
R19421 VDD.n4892 VDD.t118 37.0005
R19422 VDD.n4994 VDD.n4893 37.0005
R19423 VDD.n4893 VDD.t118 37.0005
R19424 VDD.n4878 VDD.n4876 37.0005
R19425 VDD.n4876 VDD.t84 37.0005
R19426 VDD.n5011 VDD.n4877 37.0005
R19427 VDD.n4877 VDD.t84 37.0005
R19428 VDD.n4868 VDD.n4866 37.0005
R19429 VDD.n4866 VDD.t259 37.0005
R19430 VDD.n5021 VDD.n4867 37.0005
R19431 VDD.n4867 VDD.t259 37.0005
R19432 VDD.n4857 VDD.n4855 37.0005
R19433 VDD.n4855 VDD.t486 37.0005
R19434 VDD.n5031 VDD.n4856 37.0005
R19435 VDD.n4856 VDD.t486 37.0005
R19436 VDD.n4844 VDD.n4842 37.0005
R19437 VDD.n4842 VDD.t1004 37.0005
R19438 VDD.n5041 VDD.n4843 37.0005
R19439 VDD.n4843 VDD.t1004 37.0005
R19440 VDD.n4834 VDD.n4832 37.0005
R19441 VDD.n4832 VDD.t289 37.0005
R19442 VDD.n5051 VDD.n4833 37.0005
R19443 VDD.n4833 VDD.t289 37.0005
R19444 VDD.n4823 VDD.n4821 37.0005
R19445 VDD.n4821 VDD.t496 37.0005
R19446 VDD.n5061 VDD.n4822 37.0005
R19447 VDD.n4822 VDD.t496 37.0005
R19448 VDD.n4819 VDD.n4818 37.0005
R19449 VDD.t574 VDD.n4819 37.0005
R19450 VDD.n5071 VDD.n4817 37.0005
R19451 VDD.n4940 VDD.n4938 37.0005
R19452 VDD.n4938 VDD.t183 37.0005
R19453 VDD.n4954 VDD.n4950 37.0005
R19454 VDD.n4950 VDD.t183 37.0005
R19455 VDD.n4954 VDD.n4939 37.0005
R19456 VDD.n4939 VDD.t183 37.0005
R19457 VDD.n4805 VDD.n4804 37.0005
R19458 VDD.n4804 VDD.t461 37.0005
R19459 VDD.n2053 VDD.n2052 37.0005
R19460 VDD.n2052 VDD.t461 37.0005
R19461 VDD.n4795 VDD.n4794 37.0005
R19462 VDD.n4794 VDD.t415 37.0005
R19463 VDD.n2063 VDD.n2062 37.0005
R19464 VDD.n2062 VDD.t415 37.0005
R19465 VDD.n4785 VDD.n4784 37.0005
R19466 VDD.n4784 VDD.t1016 37.0005
R19467 VDD.n2076 VDD.n2075 37.0005
R19468 VDD.n2075 VDD.t1016 37.0005
R19469 VDD.n4775 VDD.n4774 37.0005
R19470 VDD.n4774 VDD.t526 37.0005
R19471 VDD.n2088 VDD.n2087 37.0005
R19472 VDD.n2087 VDD.t526 37.0005
R19473 VDD.n2106 VDD.n2105 37.0005
R19474 VDD.n2105 VDD.t261 37.0005
R19475 VDD.n4761 VDD.n4760 37.0005
R19476 VDD.n4760 VDD.t562 37.0005
R19477 VDD.n2116 VDD.n2115 37.0005
R19478 VDD.t562 VDD.n2116 37.0005
R19479 VDD.n2119 VDD.n2117 37.0005
R19480 VDD.n2117 VDD.t1068 37.0005
R19481 VDD.n4749 VDD.n2118 37.0005
R19482 VDD.n2118 VDD.t1068 37.0005
R19483 VDD.n4741 VDD.n4740 37.0005
R19484 VDD.n4740 VDD.t564 37.0005
R19485 VDD.n2130 VDD.n2129 37.0005
R19486 VDD.n2129 VDD.t564 37.0005
R19487 VDD.n4731 VDD.n4730 37.0005
R19488 VDD.n4730 VDD.t848 37.0005
R19489 VDD.n2143 VDD.n2142 37.0005
R19490 VDD.n2142 VDD.t848 37.0005
R19491 VDD.n4721 VDD.n4720 37.0005
R19492 VDD.n4720 VDD.t467 37.0005
R19493 VDD.n2154 VDD.n2153 37.0005
R19494 VDD.n2153 VDD.t467 37.0005
R19495 VDD.n4711 VDD.n4710 37.0005
R19496 VDD.n4710 VDD.t634 37.0005
R19497 VDD.n2164 VDD.n2163 37.0005
R19498 VDD.n2163 VDD.t634 37.0005
R19499 VDD.n4701 VDD.n4700 37.0005
R19500 VDD.n4700 VDD.t548 37.0005
R19501 VDD.n4694 VDD.n4693 37.0005
R19502 VDD.n4693 VDD.t548 37.0005
R19503 VDD.n2041 VDD.n2040 37.0005
R19504 VDD.t303 VDD.n2041 37.0005
R19505 VDD.n4813 VDD.n2039 37.0005
R19506 VDD.n2047 VDD.n2045 37.0005
R19507 VDD.n2045 VDD.t461 37.0005
R19508 VDD.n4805 VDD.n2046 37.0005
R19509 VDD.n2046 VDD.t461 37.0005
R19510 VDD.n2058 VDD.n2056 37.0005
R19511 VDD.n2056 VDD.t415 37.0005
R19512 VDD.n4795 VDD.n2057 37.0005
R19513 VDD.n2057 VDD.t415 37.0005
R19514 VDD.n2068 VDD.n2066 37.0005
R19515 VDD.n2066 VDD.t1016 37.0005
R19516 VDD.n4785 VDD.n2067 37.0005
R19517 VDD.n2067 VDD.t1016 37.0005
R19518 VDD.n2081 VDD.n2079 37.0005
R19519 VDD.n2079 VDD.t526 37.0005
R19520 VDD.n4775 VDD.n2080 37.0005
R19521 VDD.n2080 VDD.t526 37.0005
R19522 VDD.n4759 VDD.n4758 37.0005
R19523 VDD.t562 VDD.n4759 37.0005
R19524 VDD.n4761 VDD.n2101 37.0005
R19525 VDD.t562 VDD.n2101 37.0005
R19526 VDD.n2123 VDD.n2121 37.0005
R19527 VDD.n2121 VDD.t564 37.0005
R19528 VDD.n4741 VDD.n2122 37.0005
R19529 VDD.n2122 VDD.t564 37.0005
R19530 VDD.n2135 VDD.n2133 37.0005
R19531 VDD.n2133 VDD.t848 37.0005
R19532 VDD.n4731 VDD.n2134 37.0005
R19533 VDD.n2134 VDD.t848 37.0005
R19534 VDD.n2148 VDD.n2146 37.0005
R19535 VDD.n2146 VDD.t467 37.0005
R19536 VDD.n4721 VDD.n2147 37.0005
R19537 VDD.n2147 VDD.t467 37.0005
R19538 VDD.n2159 VDD.n2157 37.0005
R19539 VDD.n2157 VDD.t634 37.0005
R19540 VDD.n4711 VDD.n2158 37.0005
R19541 VDD.n2158 VDD.t634 37.0005
R19542 VDD.n2169 VDD.n2167 37.0005
R19543 VDD.n2167 VDD.t548 37.0005
R19544 VDD.n4701 VDD.n2168 37.0005
R19545 VDD.n2168 VDD.t548 37.0005
R19546 VDD.n2093 VDD.n2091 37.0005
R19547 VDD.n2091 VDD.t261 37.0005
R19548 VDD.n4765 VDD.n2096 37.0005
R19549 VDD.n2096 VDD.t261 37.0005
R19550 VDD.n4765 VDD.n2092 37.0005
R19551 VDD.n2092 VDD.t261 37.0005
R19552 VDD.n4680 VDD.n4679 37.0005
R19553 VDD.n4679 VDD.t498 37.0005
R19554 VDD.n2189 VDD.n2188 37.0005
R19555 VDD.n2188 VDD.t498 37.0005
R19556 VDD.n4670 VDD.n4669 37.0005
R19557 VDD.n4669 VDD.t396 37.0005
R19558 VDD.n2199 VDD.n2198 37.0005
R19559 VDD.n2198 VDD.t396 37.0005
R19560 VDD.n4660 VDD.n4659 37.0005
R19561 VDD.n4659 VDD.t1042 37.0005
R19562 VDD.n2212 VDD.n2211 37.0005
R19563 VDD.n2211 VDD.t1042 37.0005
R19564 VDD.n4650 VDD.n4649 37.0005
R19565 VDD.n4649 VDD.t449 37.0005
R19566 VDD.n2224 VDD.n2223 37.0005
R19567 VDD.n2223 VDD.t449 37.0005
R19568 VDD.n2242 VDD.n2241 37.0005
R19569 VDD.n2241 VDD.t133 37.0005
R19570 VDD.n4636 VDD.n4635 37.0005
R19571 VDD.n4635 VDD.t95 37.0005
R19572 VDD.n2252 VDD.n2251 37.0005
R19573 VDD.t95 VDD.n2252 37.0005
R19574 VDD.n2255 VDD.n2253 37.0005
R19575 VDD.n2253 VDD.t1082 37.0005
R19576 VDD.n4624 VDD.n2254 37.0005
R19577 VDD.n2254 VDD.t1082 37.0005
R19578 VDD.n4616 VDD.n4615 37.0005
R19579 VDD.n4615 VDD.t97 37.0005
R19580 VDD.n2266 VDD.n2265 37.0005
R19581 VDD.n2265 VDD.t97 37.0005
R19582 VDD.n4606 VDD.n4605 37.0005
R19583 VDD.n4605 VDD.t143 37.0005
R19584 VDD.n2279 VDD.n2278 37.0005
R19585 VDD.n2278 VDD.t143 37.0005
R19586 VDD.n4596 VDD.n4595 37.0005
R19587 VDD.n4595 VDD.t473 37.0005
R19588 VDD.n2290 VDD.n2289 37.0005
R19589 VDD.n2289 VDD.t473 37.0005
R19590 VDD.n4586 VDD.n4585 37.0005
R19591 VDD.n4585 VDD.t541 37.0005
R19592 VDD.n2300 VDD.n2299 37.0005
R19593 VDD.n2299 VDD.t541 37.0005
R19594 VDD.n4576 VDD.n4575 37.0005
R19595 VDD.n4575 VDD.t788 37.0005
R19596 VDD.n4569 VDD.n4568 37.0005
R19597 VDD.n4568 VDD.t788 37.0005
R19598 VDD.n2177 VDD.n2176 37.0005
R19599 VDD.t65 VDD.n2177 37.0005
R19600 VDD.n4688 VDD.n2175 37.0005
R19601 VDD.n2183 VDD.n2181 37.0005
R19602 VDD.n2181 VDD.t498 37.0005
R19603 VDD.n4680 VDD.n2182 37.0005
R19604 VDD.n2182 VDD.t498 37.0005
R19605 VDD.n2194 VDD.n2192 37.0005
R19606 VDD.n2192 VDD.t396 37.0005
R19607 VDD.n4670 VDD.n2193 37.0005
R19608 VDD.n2193 VDD.t396 37.0005
R19609 VDD.n2204 VDD.n2202 37.0005
R19610 VDD.n2202 VDD.t1042 37.0005
R19611 VDD.n4660 VDD.n2203 37.0005
R19612 VDD.n2203 VDD.t1042 37.0005
R19613 VDD.n2217 VDD.n2215 37.0005
R19614 VDD.n2215 VDD.t449 37.0005
R19615 VDD.n4650 VDD.n2216 37.0005
R19616 VDD.n2216 VDD.t449 37.0005
R19617 VDD.n4634 VDD.n4633 37.0005
R19618 VDD.t95 VDD.n4634 37.0005
R19619 VDD.n4636 VDD.n2237 37.0005
R19620 VDD.t95 VDD.n2237 37.0005
R19621 VDD.n2259 VDD.n2257 37.0005
R19622 VDD.n2257 VDD.t97 37.0005
R19623 VDD.n4616 VDD.n2258 37.0005
R19624 VDD.n2258 VDD.t97 37.0005
R19625 VDD.n2271 VDD.n2269 37.0005
R19626 VDD.n2269 VDD.t143 37.0005
R19627 VDD.n4606 VDD.n2270 37.0005
R19628 VDD.n2270 VDD.t143 37.0005
R19629 VDD.n2284 VDD.n2282 37.0005
R19630 VDD.n2282 VDD.t473 37.0005
R19631 VDD.n4596 VDD.n2283 37.0005
R19632 VDD.n2283 VDD.t473 37.0005
R19633 VDD.n2295 VDD.n2293 37.0005
R19634 VDD.n2293 VDD.t541 37.0005
R19635 VDD.n4586 VDD.n2294 37.0005
R19636 VDD.n2294 VDD.t541 37.0005
R19637 VDD.n2305 VDD.n2303 37.0005
R19638 VDD.n2303 VDD.t788 37.0005
R19639 VDD.n4576 VDD.n2304 37.0005
R19640 VDD.n2304 VDD.t788 37.0005
R19641 VDD.n2229 VDD.n2227 37.0005
R19642 VDD.n2227 VDD.t133 37.0005
R19643 VDD.n4640 VDD.n2232 37.0005
R19644 VDD.n2232 VDD.t133 37.0005
R19645 VDD.n4640 VDD.n2228 37.0005
R19646 VDD.n2228 VDD.t133 37.0005
R19647 VDD.n4555 VDD.n4554 37.0005
R19648 VDD.n4554 VDD.t508 37.0005
R19649 VDD.n2325 VDD.n2324 37.0005
R19650 VDD.n2324 VDD.t508 37.0005
R19651 VDD.n4545 VDD.n4544 37.0005
R19652 VDD.n4544 VDD.t858 37.0005
R19653 VDD.n2335 VDD.n2334 37.0005
R19654 VDD.n2334 VDD.t858 37.0005
R19655 VDD.n4535 VDD.n4534 37.0005
R19656 VDD.n4534 VDD.t1050 37.0005
R19657 VDD.n2348 VDD.n2347 37.0005
R19658 VDD.n2347 VDD.t1050 37.0005
R19659 VDD.n4525 VDD.n4524 37.0005
R19660 VDD.n4524 VDD.t518 37.0005
R19661 VDD.n2360 VDD.n2359 37.0005
R19662 VDD.n2359 VDD.t518 37.0005
R19663 VDD.n2378 VDD.n2377 37.0005
R19664 VDD.n2377 VDD.t266 37.0005
R19665 VDD.n4511 VDD.n4510 37.0005
R19666 VDD.n4510 VDD.t215 37.0005
R19667 VDD.n2388 VDD.n2387 37.0005
R19668 VDD.t215 VDD.n2388 37.0005
R19669 VDD.n2391 VDD.n2389 37.0005
R19670 VDD.n2389 VDD.t1010 37.0005
R19671 VDD.n4499 VDD.n2390 37.0005
R19672 VDD.n2390 VDD.t1010 37.0005
R19673 VDD.n4491 VDD.n4490 37.0005
R19674 VDD.n4490 VDD.t217 37.0005
R19675 VDD.n2402 VDD.n2401 37.0005
R19676 VDD.n2401 VDD.t217 37.0005
R19677 VDD.n4481 VDD.n4480 37.0005
R19678 VDD.n4480 VDD.t91 37.0005
R19679 VDD.n2415 VDD.n2414 37.0005
R19680 VDD.n2414 VDD.t91 37.0005
R19681 VDD.n4471 VDD.n4470 37.0005
R19682 VDD.n4470 VDD.t532 37.0005
R19683 VDD.n2426 VDD.n2425 37.0005
R19684 VDD.n2425 VDD.t532 37.0005
R19685 VDD.n4461 VDD.n4460 37.0005
R19686 VDD.n4460 VDD.t160 37.0005
R19687 VDD.n2436 VDD.n2435 37.0005
R19688 VDD.n2435 VDD.t160 37.0005
R19689 VDD.n4451 VDD.n4450 37.0005
R19690 VDD.n4450 VDD.t590 37.0005
R19691 VDD.n4444 VDD.n4443 37.0005
R19692 VDD.n4443 VDD.t590 37.0005
R19693 VDD.n2313 VDD.n2312 37.0005
R19694 VDD.t25 VDD.n2313 37.0005
R19695 VDD.n4563 VDD.n2311 37.0005
R19696 VDD.n2319 VDD.n2317 37.0005
R19697 VDD.n2317 VDD.t508 37.0005
R19698 VDD.n4555 VDD.n2318 37.0005
R19699 VDD.n2318 VDD.t508 37.0005
R19700 VDD.n2330 VDD.n2328 37.0005
R19701 VDD.n2328 VDD.t858 37.0005
R19702 VDD.n4545 VDD.n2329 37.0005
R19703 VDD.n2329 VDD.t858 37.0005
R19704 VDD.n2340 VDD.n2338 37.0005
R19705 VDD.n2338 VDD.t1050 37.0005
R19706 VDD.n4535 VDD.n2339 37.0005
R19707 VDD.n2339 VDD.t1050 37.0005
R19708 VDD.n2353 VDD.n2351 37.0005
R19709 VDD.n2351 VDD.t518 37.0005
R19710 VDD.n4525 VDD.n2352 37.0005
R19711 VDD.n2352 VDD.t518 37.0005
R19712 VDD.n4509 VDD.n4508 37.0005
R19713 VDD.t215 VDD.n4509 37.0005
R19714 VDD.n4511 VDD.n2373 37.0005
R19715 VDD.t215 VDD.n2373 37.0005
R19716 VDD.n2395 VDD.n2393 37.0005
R19717 VDD.n2393 VDD.t217 37.0005
R19718 VDD.n4491 VDD.n2394 37.0005
R19719 VDD.n2394 VDD.t217 37.0005
R19720 VDD.n2407 VDD.n2405 37.0005
R19721 VDD.n2405 VDD.t91 37.0005
R19722 VDD.n4481 VDD.n2406 37.0005
R19723 VDD.n2406 VDD.t91 37.0005
R19724 VDD.n2420 VDD.n2418 37.0005
R19725 VDD.n2418 VDD.t532 37.0005
R19726 VDD.n4471 VDD.n2419 37.0005
R19727 VDD.n2419 VDD.t532 37.0005
R19728 VDD.n2431 VDD.n2429 37.0005
R19729 VDD.n2429 VDD.t160 37.0005
R19730 VDD.n4461 VDD.n2430 37.0005
R19731 VDD.n2430 VDD.t160 37.0005
R19732 VDD.n2441 VDD.n2439 37.0005
R19733 VDD.n2439 VDD.t590 37.0005
R19734 VDD.n4451 VDD.n2440 37.0005
R19735 VDD.n2440 VDD.t590 37.0005
R19736 VDD.n2365 VDD.n2363 37.0005
R19737 VDD.n2363 VDD.t266 37.0005
R19738 VDD.n4515 VDD.n2368 37.0005
R19739 VDD.n2368 VDD.t266 37.0005
R19740 VDD.n4515 VDD.n2364 37.0005
R19741 VDD.n2364 VDD.t266 37.0005
R19742 VDD.n4430 VDD.n4429 37.0005
R19743 VDD.n4429 VDD.t504 37.0005
R19744 VDD.n2461 VDD.n2460 37.0005
R19745 VDD.n2460 VDD.t504 37.0005
R19746 VDD.n4420 VDD.n4419 37.0005
R19747 VDD.n4419 VDD.t800 37.0005
R19748 VDD.n2471 VDD.n2470 37.0005
R19749 VDD.n2470 VDD.t800 37.0005
R19750 VDD.n4410 VDD.n4409 37.0005
R19751 VDD.n4409 VDD.t1048 37.0005
R19752 VDD.n2484 VDD.n2483 37.0005
R19753 VDD.n2483 VDD.t1048 37.0005
R19754 VDD.n4400 VDD.n4399 37.0005
R19755 VDD.n4399 VDD.t441 37.0005
R19756 VDD.n2496 VDD.n2495 37.0005
R19757 VDD.n2495 VDD.t441 37.0005
R19758 VDD.n2514 VDD.n2513 37.0005
R19759 VDD.n2513 VDD.t328 37.0005
R19760 VDD.n4386 VDD.n4385 37.0005
R19761 VDD.n4385 VDD.t19 37.0005
R19762 VDD.n2524 VDD.n2523 37.0005
R19763 VDD.t19 VDD.n2524 37.0005
R19764 VDD.n2527 VDD.n2525 37.0005
R19765 VDD.n2525 VDD.t1038 37.0005
R19766 VDD.n4374 VDD.n2526 37.0005
R19767 VDD.n2526 VDD.t1038 37.0005
R19768 VDD.n4366 VDD.n4365 37.0005
R19769 VDD.n4365 VDD.t593 37.0005
R19770 VDD.n2538 VDD.n2537 37.0005
R19771 VDD.n2537 VDD.t593 37.0005
R19772 VDD.n4356 VDD.n4355 37.0005
R19773 VDD.n4355 VDD.t199 37.0005
R19774 VDD.n2551 VDD.n2550 37.0005
R19775 VDD.n2550 VDD.t199 37.0005
R19776 VDD.n4346 VDD.n4345 37.0005
R19777 VDD.n4345 VDD.t451 37.0005
R19778 VDD.n2562 VDD.n2561 37.0005
R19779 VDD.n2561 VDD.t451 37.0005
R19780 VDD.n4336 VDD.n4335 37.0005
R19781 VDD.n4335 VDD.t39 37.0005
R19782 VDD.n2572 VDD.n2571 37.0005
R19783 VDD.n2571 VDD.t39 37.0005
R19784 VDD.n4326 VDD.n4325 37.0005
R19785 VDD.n4325 VDD.t69 37.0005
R19786 VDD.n4319 VDD.n4318 37.0005
R19787 VDD.n4318 VDD.t69 37.0005
R19788 VDD.n2449 VDD.n2448 37.0005
R19789 VDD.t796 VDD.n2449 37.0005
R19790 VDD.n4438 VDD.n2447 37.0005
R19791 VDD.n2455 VDD.n2453 37.0005
R19792 VDD.n2453 VDD.t504 37.0005
R19793 VDD.n4430 VDD.n2454 37.0005
R19794 VDD.n2454 VDD.t504 37.0005
R19795 VDD.n2466 VDD.n2464 37.0005
R19796 VDD.n2464 VDD.t800 37.0005
R19797 VDD.n4420 VDD.n2465 37.0005
R19798 VDD.n2465 VDD.t800 37.0005
R19799 VDD.n2476 VDD.n2474 37.0005
R19800 VDD.n2474 VDD.t1048 37.0005
R19801 VDD.n4410 VDD.n2475 37.0005
R19802 VDD.n2475 VDD.t1048 37.0005
R19803 VDD.n2489 VDD.n2487 37.0005
R19804 VDD.n2487 VDD.t441 37.0005
R19805 VDD.n4400 VDD.n2488 37.0005
R19806 VDD.n2488 VDD.t441 37.0005
R19807 VDD.n4384 VDD.n4383 37.0005
R19808 VDD.t19 VDD.n4384 37.0005
R19809 VDD.n4386 VDD.n2509 37.0005
R19810 VDD.t19 VDD.n2509 37.0005
R19811 VDD.n2531 VDD.n2529 37.0005
R19812 VDD.n2529 VDD.t593 37.0005
R19813 VDD.n4366 VDD.n2530 37.0005
R19814 VDD.n2530 VDD.t593 37.0005
R19815 VDD.n2543 VDD.n2541 37.0005
R19816 VDD.n2541 VDD.t199 37.0005
R19817 VDD.n4356 VDD.n2542 37.0005
R19818 VDD.n2542 VDD.t199 37.0005
R19819 VDD.n2556 VDD.n2554 37.0005
R19820 VDD.n2554 VDD.t451 37.0005
R19821 VDD.n4346 VDD.n2555 37.0005
R19822 VDD.n2555 VDD.t451 37.0005
R19823 VDD.n2567 VDD.n2565 37.0005
R19824 VDD.n2565 VDD.t39 37.0005
R19825 VDD.n4336 VDD.n2566 37.0005
R19826 VDD.n2566 VDD.t39 37.0005
R19827 VDD.n2577 VDD.n2575 37.0005
R19828 VDD.n2575 VDD.t69 37.0005
R19829 VDD.n4326 VDD.n2576 37.0005
R19830 VDD.n2576 VDD.t69 37.0005
R19831 VDD.n2501 VDD.n2499 37.0005
R19832 VDD.n2499 VDD.t328 37.0005
R19833 VDD.n4390 VDD.n2504 37.0005
R19834 VDD.n2504 VDD.t328 37.0005
R19835 VDD.n4390 VDD.n2500 37.0005
R19836 VDD.n2500 VDD.t328 37.0005
R19837 VDD.n4305 VDD.n4304 37.0005
R19838 VDD.n4304 VDD.t536 37.0005
R19839 VDD.n2597 VDD.n2596 37.0005
R19840 VDD.n2596 VDD.t536 37.0005
R19841 VDD.n4295 VDD.n4294 37.0005
R19842 VDD.n4294 VDD.t67 37.0005
R19843 VDD.n2607 VDD.n2606 37.0005
R19844 VDD.n2606 VDD.t67 37.0005
R19845 VDD.n4285 VDD.n4284 37.0005
R19846 VDD.n4284 VDD.t1022 37.0005
R19847 VDD.n2620 VDD.n2619 37.0005
R19848 VDD.n2619 VDD.t1022 37.0005
R19849 VDD.n4275 VDD.n4274 37.0005
R19850 VDD.n4274 VDD.t488 37.0005
R19851 VDD.n2632 VDD.n2631 37.0005
R19852 VDD.n2631 VDD.t488 37.0005
R19853 VDD.n2650 VDD.n2649 37.0005
R19854 VDD.n2649 VDD.t31 37.0005
R19855 VDD.n4261 VDD.n4260 37.0005
R19856 VDD.n4260 VDD.t386 37.0005
R19857 VDD.n2660 VDD.n2659 37.0005
R19858 VDD.t386 VDD.n2660 37.0005
R19859 VDD.n2663 VDD.n2661 37.0005
R19860 VDD.n2661 VDD.t1062 37.0005
R19861 VDD.n4249 VDD.n2662 37.0005
R19862 VDD.n2662 VDD.t1062 37.0005
R19863 VDD.n4241 VDD.n4240 37.0005
R19864 VDD.n4240 VDD.t388 37.0005
R19865 VDD.n2674 VDD.n2673 37.0005
R19866 VDD.n2673 VDD.t388 37.0005
R19867 VDD.n4231 VDD.n4230 37.0005
R19868 VDD.n4230 VDD.t344 37.0005
R19869 VDD.n2687 VDD.n2686 37.0005
R19870 VDD.n2686 VDD.t344 37.0005
R19871 VDD.n4221 VDD.n4220 37.0005
R19872 VDD.n4220 VDD.t469 37.0005
R19873 VDD.n2698 VDD.n2697 37.0005
R19874 VDD.n2697 VDD.t469 37.0005
R19875 VDD.n4211 VDD.n4210 37.0005
R19876 VDD.n4210 VDD.t892 37.0005
R19877 VDD.n2708 VDD.n2707 37.0005
R19878 VDD.n2707 VDD.t892 37.0005
R19879 VDD.n4201 VDD.n4200 37.0005
R19880 VDD.n4200 VDD.t2 37.0005
R19881 VDD.n4194 VDD.n4193 37.0005
R19882 VDD.n4193 VDD.t2 37.0005
R19883 VDD.n2585 VDD.n2584 37.0005
R19884 VDD.t764 VDD.n2585 37.0005
R19885 VDD.n4313 VDD.n2583 37.0005
R19886 VDD.n2591 VDD.n2589 37.0005
R19887 VDD.n2589 VDD.t536 37.0005
R19888 VDD.n4305 VDD.n2590 37.0005
R19889 VDD.n2590 VDD.t536 37.0005
R19890 VDD.n2602 VDD.n2600 37.0005
R19891 VDD.n2600 VDD.t67 37.0005
R19892 VDD.n4295 VDD.n2601 37.0005
R19893 VDD.n2601 VDD.t67 37.0005
R19894 VDD.n2612 VDD.n2610 37.0005
R19895 VDD.n2610 VDD.t1022 37.0005
R19896 VDD.n4285 VDD.n2611 37.0005
R19897 VDD.n2611 VDD.t1022 37.0005
R19898 VDD.n2625 VDD.n2623 37.0005
R19899 VDD.n2623 VDD.t488 37.0005
R19900 VDD.n4275 VDD.n2624 37.0005
R19901 VDD.n2624 VDD.t488 37.0005
R19902 VDD.n4259 VDD.n4258 37.0005
R19903 VDD.t386 VDD.n4259 37.0005
R19904 VDD.n4261 VDD.n2645 37.0005
R19905 VDD.t386 VDD.n2645 37.0005
R19906 VDD.n2667 VDD.n2665 37.0005
R19907 VDD.n2665 VDD.t388 37.0005
R19908 VDD.n4241 VDD.n2666 37.0005
R19909 VDD.n2666 VDD.t388 37.0005
R19910 VDD.n2679 VDD.n2677 37.0005
R19911 VDD.n2677 VDD.t344 37.0005
R19912 VDD.n4231 VDD.n2678 37.0005
R19913 VDD.n2678 VDD.t344 37.0005
R19914 VDD.n2692 VDD.n2690 37.0005
R19915 VDD.n2690 VDD.t469 37.0005
R19916 VDD.n4221 VDD.n2691 37.0005
R19917 VDD.n2691 VDD.t469 37.0005
R19918 VDD.n2703 VDD.n2701 37.0005
R19919 VDD.n2701 VDD.t892 37.0005
R19920 VDD.n4211 VDD.n2702 37.0005
R19921 VDD.n2702 VDD.t892 37.0005
R19922 VDD.n2713 VDD.n2711 37.0005
R19923 VDD.n2711 VDD.t2 37.0005
R19924 VDD.n4201 VDD.n2712 37.0005
R19925 VDD.n2712 VDD.t2 37.0005
R19926 VDD.n2637 VDD.n2635 37.0005
R19927 VDD.n2635 VDD.t31 37.0005
R19928 VDD.n4265 VDD.n2640 37.0005
R19929 VDD.n2640 VDD.t31 37.0005
R19930 VDD.n4265 VDD.n2636 37.0005
R19931 VDD.n2636 VDD.t31 37.0005
R19932 VDD.n4180 VDD.n4179 37.0005
R19933 VDD.n4179 VDD.t455 37.0005
R19934 VDD.n2733 VDD.n2732 37.0005
R19935 VDD.n2732 VDD.t455 37.0005
R19936 VDD.n4170 VDD.n4169 37.0005
R19937 VDD.n4169 VDD.t0 37.0005
R19938 VDD.n2743 VDD.n2742 37.0005
R19939 VDD.n2742 VDD.t0 37.0005
R19940 VDD.n4160 VDD.n4159 37.0005
R19941 VDD.n4159 VDD.t1018 37.0005
R19942 VDD.n2756 VDD.n2755 37.0005
R19943 VDD.n2755 VDD.t1018 37.0005
R19944 VDD.n4150 VDD.n4149 37.0005
R19945 VDD.n4149 VDD.t514 37.0005
R19946 VDD.n2768 VDD.n2767 37.0005
R19947 VDD.n2767 VDD.t514 37.0005
R19948 VDD.n2786 VDD.n2785 37.0005
R19949 VDD.n2785 VDD.t373 37.0005
R19950 VDD.n4136 VDD.n4135 37.0005
R19951 VDD.n4135 VDD.t80 37.0005
R19952 VDD.n2796 VDD.n2795 37.0005
R19953 VDD.t80 VDD.n2796 37.0005
R19954 VDD.n2799 VDD.n2797 37.0005
R19955 VDD.n2797 VDD.t1006 37.0005
R19956 VDD.n4124 VDD.n2798 37.0005
R19957 VDD.n2798 VDD.t1006 37.0005
R19958 VDD.n4116 VDD.n4115 37.0005
R19959 VDD.n4115 VDD.t82 37.0005
R19960 VDD.n2810 VDD.n2809 37.0005
R19961 VDD.n2809 VDD.t82 37.0005
R19962 VDD.n4106 VDD.n4105 37.0005
R19963 VDD.n4105 VDD.t168 37.0005
R19964 VDD.n2823 VDD.n2822 37.0005
R19965 VDD.n2822 VDD.t168 37.0005
R19966 VDD.n4096 VDD.n4095 37.0005
R19967 VDD.n4095 VDD.t524 37.0005
R19968 VDD.n2834 VDD.n2833 37.0005
R19969 VDD.n2833 VDD.t524 37.0005
R19970 VDD.n4086 VDD.n4085 37.0005
R19971 VDD.n4085 VDD.t99 37.0005
R19972 VDD.n2844 VDD.n2843 37.0005
R19973 VDD.n2843 VDD.t99 37.0005
R19974 VDD.n4076 VDD.n4075 37.0005
R19975 VDD.n4075 VDD.t292 37.0005
R19976 VDD.n4069 VDD.n4068 37.0005
R19977 VDD.n4068 VDD.t292 37.0005
R19978 VDD.n2721 VDD.n2720 37.0005
R19979 VDD.t124 VDD.n2721 37.0005
R19980 VDD.n4188 VDD.n2719 37.0005
R19981 VDD.n2727 VDD.n2725 37.0005
R19982 VDD.n2725 VDD.t455 37.0005
R19983 VDD.n4180 VDD.n2726 37.0005
R19984 VDD.n2726 VDD.t455 37.0005
R19985 VDD.n2738 VDD.n2736 37.0005
R19986 VDD.n2736 VDD.t0 37.0005
R19987 VDD.n4170 VDD.n2737 37.0005
R19988 VDD.n2737 VDD.t0 37.0005
R19989 VDD.n2748 VDD.n2746 37.0005
R19990 VDD.n2746 VDD.t1018 37.0005
R19991 VDD.n4160 VDD.n2747 37.0005
R19992 VDD.n2747 VDD.t1018 37.0005
R19993 VDD.n2761 VDD.n2759 37.0005
R19994 VDD.n2759 VDD.t514 37.0005
R19995 VDD.n4150 VDD.n2760 37.0005
R19996 VDD.n2760 VDD.t514 37.0005
R19997 VDD.n4134 VDD.n4133 37.0005
R19998 VDD.t80 VDD.n4134 37.0005
R19999 VDD.n4136 VDD.n2781 37.0005
R20000 VDD.t80 VDD.n2781 37.0005
R20001 VDD.n2803 VDD.n2801 37.0005
R20002 VDD.n2801 VDD.t82 37.0005
R20003 VDD.n4116 VDD.n2802 37.0005
R20004 VDD.n2802 VDD.t82 37.0005
R20005 VDD.n2815 VDD.n2813 37.0005
R20006 VDD.n2813 VDD.t168 37.0005
R20007 VDD.n4106 VDD.n2814 37.0005
R20008 VDD.n2814 VDD.t168 37.0005
R20009 VDD.n2828 VDD.n2826 37.0005
R20010 VDD.n2826 VDD.t524 37.0005
R20011 VDD.n4096 VDD.n2827 37.0005
R20012 VDD.n2827 VDD.t524 37.0005
R20013 VDD.n2839 VDD.n2837 37.0005
R20014 VDD.n2837 VDD.t99 37.0005
R20015 VDD.n4086 VDD.n2838 37.0005
R20016 VDD.n2838 VDD.t99 37.0005
R20017 VDD.n2849 VDD.n2847 37.0005
R20018 VDD.n2847 VDD.t292 37.0005
R20019 VDD.n4076 VDD.n2848 37.0005
R20020 VDD.n2848 VDD.t292 37.0005
R20021 VDD.n2773 VDD.n2771 37.0005
R20022 VDD.n2771 VDD.t373 37.0005
R20023 VDD.n4140 VDD.n2776 37.0005
R20024 VDD.n2776 VDD.t373 37.0005
R20025 VDD.n4140 VDD.n2772 37.0005
R20026 VDD.n2772 VDD.t373 37.0005
R20027 VDD.n4055 VDD.n4054 37.0005
R20028 VDD.n4054 VDD.t502 37.0005
R20029 VDD.n2869 VDD.n2868 37.0005
R20030 VDD.n2868 VDD.t502 37.0005
R20031 VDD.n4045 VDD.n4044 37.0005
R20032 VDD.n4044 VDD.t934 37.0005
R20033 VDD.n2879 VDD.n2878 37.0005
R20034 VDD.n2878 VDD.t934 37.0005
R20035 VDD.n4035 VDD.n4034 37.0005
R20036 VDD.n4034 VDD.t1045 37.0005
R20037 VDD.n2892 VDD.n2891 37.0005
R20038 VDD.n2891 VDD.t1045 37.0005
R20039 VDD.n4025 VDD.n4024 37.0005
R20040 VDD.n4024 VDD.t437 37.0005
R20041 VDD.n2904 VDD.n2903 37.0005
R20042 VDD.n2903 VDD.t437 37.0005
R20043 VDD.n2922 VDD.n2921 37.0005
R20044 VDD.n2921 VDD.t821 37.0005
R20045 VDD.n4011 VDD.n4010 37.0005
R20046 VDD.n4010 VDD.t310 37.0005
R20047 VDD.n2932 VDD.n2931 37.0005
R20048 VDD.t310 VDD.n2932 37.0005
R20049 VDD.n2935 VDD.n2933 37.0005
R20050 VDD.n2933 VDD.t1034 37.0005
R20051 VDD.n3999 VDD.n2934 37.0005
R20052 VDD.n2934 VDD.t1034 37.0005
R20053 VDD.n3991 VDD.n3990 37.0005
R20054 VDD.n3990 VDD.t308 37.0005
R20055 VDD.n2946 VDD.n2945 37.0005
R20056 VDD.n2945 VDD.t308 37.0005
R20057 VDD.n3981 VDD.n3980 37.0005
R20058 VDD.n3980 VDD.t196 37.0005
R20059 VDD.n2959 VDD.n2958 37.0005
R20060 VDD.n2958 VDD.t196 37.0005
R20061 VDD.n3971 VDD.n3970 37.0005
R20062 VDD.n3970 VDD.t447 37.0005
R20063 VDD.n2970 VDD.n2969 37.0005
R20064 VDD.n2969 VDD.t447 37.0005
R20065 VDD.n3961 VDD.n3960 37.0005
R20066 VDD.n3960 VDD.t296 37.0005
R20067 VDD.n2980 VDD.n2979 37.0005
R20068 VDD.n2979 VDD.t296 37.0005
R20069 VDD.n3951 VDD.n3950 37.0005
R20070 VDD.n3950 VDD.t626 37.0005
R20071 VDD.n3944 VDD.n3943 37.0005
R20072 VDD.n3943 VDD.t626 37.0005
R20073 VDD.n2857 VDD.n2856 37.0005
R20074 VDD.t153 VDD.n2857 37.0005
R20075 VDD.n4063 VDD.n2855 37.0005
R20076 VDD.n2863 VDD.n2861 37.0005
R20077 VDD.n2861 VDD.t502 37.0005
R20078 VDD.n4055 VDD.n2862 37.0005
R20079 VDD.n2862 VDD.t502 37.0005
R20080 VDD.n2874 VDD.n2872 37.0005
R20081 VDD.n2872 VDD.t934 37.0005
R20082 VDD.n4045 VDD.n2873 37.0005
R20083 VDD.n2873 VDD.t934 37.0005
R20084 VDD.n2884 VDD.n2882 37.0005
R20085 VDD.n2882 VDD.t1045 37.0005
R20086 VDD.n4035 VDD.n2883 37.0005
R20087 VDD.n2883 VDD.t1045 37.0005
R20088 VDD.n2897 VDD.n2895 37.0005
R20089 VDD.n2895 VDD.t437 37.0005
R20090 VDD.n4025 VDD.n2896 37.0005
R20091 VDD.n2896 VDD.t437 37.0005
R20092 VDD.n4009 VDD.n4008 37.0005
R20093 VDD.t310 VDD.n4009 37.0005
R20094 VDD.n4011 VDD.n2917 37.0005
R20095 VDD.t310 VDD.n2917 37.0005
R20096 VDD.n2939 VDD.n2937 37.0005
R20097 VDD.n2937 VDD.t308 37.0005
R20098 VDD.n3991 VDD.n2938 37.0005
R20099 VDD.n2938 VDD.t308 37.0005
R20100 VDD.n2951 VDD.n2949 37.0005
R20101 VDD.n2949 VDD.t196 37.0005
R20102 VDD.n3981 VDD.n2950 37.0005
R20103 VDD.n2950 VDD.t196 37.0005
R20104 VDD.n2964 VDD.n2962 37.0005
R20105 VDD.n2962 VDD.t447 37.0005
R20106 VDD.n3971 VDD.n2963 37.0005
R20107 VDD.n2963 VDD.t447 37.0005
R20108 VDD.n2975 VDD.n2973 37.0005
R20109 VDD.n2973 VDD.t296 37.0005
R20110 VDD.n3961 VDD.n2974 37.0005
R20111 VDD.n2974 VDD.t296 37.0005
R20112 VDD.n2985 VDD.n2983 37.0005
R20113 VDD.n2983 VDD.t626 37.0005
R20114 VDD.n3951 VDD.n2984 37.0005
R20115 VDD.n2984 VDD.t626 37.0005
R20116 VDD.n2909 VDD.n2907 37.0005
R20117 VDD.n2907 VDD.t821 37.0005
R20118 VDD.n4015 VDD.n2912 37.0005
R20119 VDD.n2912 VDD.t821 37.0005
R20120 VDD.n4015 VDD.n2908 37.0005
R20121 VDD.n2908 VDD.t821 37.0005
R20122 VDD.n3616 VDD.n3615 37.0005
R20123 VDD.n3615 VDD.t86 37.0005
R20124 VDD.n3275 VDD.n3274 37.0005
R20125 VDD.t86 VDD.n3275 37.0005
R20126 VDD.n3603 VDD.n3602 37.0005
R20127 VDD.n3602 VDD.t88 37.0005
R20128 VDD.n3284 VDD.n3283 37.0005
R20129 VDD.n3283 VDD.t88 37.0005
R20130 VDD.n3293 VDD.n3292 37.0005
R20131 VDD.n3292 VDD.t21 37.0005
R20132 VDD.n3614 VDD.n3613 37.0005
R20133 VDD.t86 VDD.n3614 37.0005
R20134 VDD.n3616 VDD.n3267 37.0005
R20135 VDD.t86 VDD.n3267 37.0005
R20136 VDD.n3279 VDD.n3277 37.0005
R20137 VDD.n3277 VDD.t88 37.0005
R20138 VDD.n3603 VDD.n3278 37.0005
R20139 VDD.n3278 VDD.t88 37.0005
R20140 VDD.n3289 VDD.n3287 37.0005
R20141 VDD.n3287 VDD.t21 37.0005
R20142 VDD.n3593 VDD.n3299 37.0005
R20143 VDD.n3299 VDD.t21 37.0005
R20144 VDD.n3593 VDD.n3288 37.0005
R20145 VDD.n3288 VDD.t21 37.0005
R20146 VDD.n3349 VDD.n3347 37.0005
R20147 VDD.n3347 VDD.t176 37.0005
R20148 VDD.n3439 VDD.n3348 37.0005
R20149 VDD.n3348 VDD.t176 37.0005
R20150 VDD.n3346 VDD.n3345 37.0005
R20151 VDD.t985 VDD.n3346 37.0005
R20152 VDD.n3448 VDD.n3344 37.0005
R20153 VDD.n3426 VDD.n3425 37.0005
R20154 VDD.t854 VDD.n3426 37.0005
R20155 VDD.n3434 VDD.n3424 37.0005
R20156 VDD.n3458 VDD.n3456 37.0005
R20157 VDD.n3456 VDD.t812 37.0005
R20158 VDD.n3476 VDD.n3457 37.0005
R20159 VDD.n3457 VDD.t812 37.0005
R20160 VDD.n3455 VDD.n3454 37.0005
R20161 VDD.t131 VDD.n3455 37.0005
R20162 VDD.n3485 VDD.n3453 37.0005
R20163 VDD.n3464 VDD.n3463 37.0005
R20164 VDD.t810 VDD.n3464 37.0005
R20165 VDD.n3472 VDD.n3462 37.0005
R20166 VDD.n3324 VDD.n3322 37.0005
R20167 VDD.n3322 VDD.t256 37.0005
R20168 VDD.n3505 VDD.n3323 37.0005
R20169 VDD.n3323 VDD.t256 37.0005
R20170 VDD.n3329 VDD.n3328 37.0005
R20171 VDD.t884 VDD.n3329 37.0005
R20172 VDD.n3337 VDD.n3327 37.0005
R20173 VDD.n3319 VDD.n3318 37.0005
R20174 VDD.t271 VDD.n3319 37.0005
R20175 VDD.n3512 VDD.n3317 37.0005
R20176 VDD.n3312 VDD.n3310 37.0005
R20177 VDD.n3310 VDD.t998 37.0005
R20178 VDD.n3534 VDD.n3311 37.0005
R20179 VDD.n3311 VDD.t998 37.0005
R20180 VDD.n3309 VDD.n3308 37.0005
R20181 VDD.t122 VDD.n3309 37.0005
R20182 VDD.n3543 VDD.n3307 37.0005
R20183 VDD.n3521 VDD.n3520 37.0005
R20184 VDD.t996 VDD.n3521 37.0005
R20185 VDD.n3529 VDD.n3519 37.0005
R20186 VDD.n3552 VDD.n3550 37.0005
R20187 VDD.n3550 VDD.t410 37.0005
R20188 VDD.n3570 VDD.n3551 37.0005
R20189 VDD.n3551 VDD.t410 37.0005
R20190 VDD.n3549 VDD.n3548 37.0005
R20191 VDD.t137 VDD.n3549 37.0005
R20192 VDD.n3579 VDD.n3547 37.0005
R20193 VDD.n3558 VDD.n3557 37.0005
R20194 VDD.t408 VDD.n3558 37.0005
R20195 VDD.n3566 VDD.n3556 37.0005
R20196 VDD.n3380 VDD.n3378 37.0005
R20197 VDD.n3378 VDD.t784 37.0005
R20198 VDD.n3410 VDD.n3379 37.0005
R20199 VDD.n3379 VDD.t784 37.0005
R20200 VDD.n3385 VDD.n3384 37.0005
R20201 VDD.t206 VDD.n3385 37.0005
R20202 VDD.n3393 VDD.n3383 37.0005
R20203 VDD.n3375 VDD.n3374 37.0005
R20204 VDD.t782 VDD.n3375 37.0005
R20205 VDD.n3417 VDD.n3373 37.0005
R20206 VDD.n3930 VDD.n3929 37.0005
R20207 VDD.n3929 VDD.t528 37.0005
R20208 VDD.n3005 VDD.n3004 37.0005
R20209 VDD.n3004 VDD.t528 37.0005
R20210 VDD.n3920 VDD.n3919 37.0005
R20211 VDD.n3919 VDD.t151 37.0005
R20212 VDD.n3015 VDD.n3014 37.0005
R20213 VDD.n3014 VDD.t151 37.0005
R20214 VDD.n3910 VDD.n3909 37.0005
R20215 VDD.n3909 VDD.t1014 37.0005
R20216 VDD.n3028 VDD.n3027 37.0005
R20217 VDD.n3027 VDD.t1014 37.0005
R20218 VDD.n3900 VDD.n3899 37.0005
R20219 VDD.n3899 VDD.t484 37.0005
R20220 VDD.n3730 VDD.n3729 37.0005
R20221 VDD.n3729 VDD.t484 37.0005
R20222 VDD.n3748 VDD.n3747 37.0005
R20223 VDD.n3747 VDD.t51 37.0005
R20224 VDD.n3886 VDD.n3885 37.0005
R20225 VDD.n3885 VDD.t231 37.0005
R20226 VDD.n3758 VDD.n3757 37.0005
R20227 VDD.t231 VDD.n3758 37.0005
R20228 VDD.n3761 VDD.n3759 37.0005
R20229 VDD.n3759 VDD.t1091 37.0005
R20230 VDD.n3874 VDD.n3760 37.0005
R20231 VDD.n3760 VDD.t1091 37.0005
R20232 VDD.n3866 VDD.n3865 37.0005
R20233 VDD.n3865 VDD.t284 37.0005
R20234 VDD.n3772 VDD.n3771 37.0005
R20235 VDD.n3771 VDD.t284 37.0005
R20236 VDD.n3856 VDD.n3855 37.0005
R20237 VDD.n3855 VDD.t558 37.0005
R20238 VDD.n3785 VDD.n3784 37.0005
R20239 VDD.n3784 VDD.t558 37.0005
R20240 VDD.n3846 VDD.n3845 37.0005
R20241 VDD.n3845 VDD.t445 37.0005
R20242 VDD.n3796 VDD.n3795 37.0005
R20243 VDD.n3795 VDD.t445 37.0005
R20244 VDD.n3836 VDD.n3835 37.0005
R20245 VDD.n3835 VDD.t427 37.0005
R20246 VDD.n3806 VDD.n3805 37.0005
R20247 VDD.n3805 VDD.t427 37.0005
R20248 VDD.n3826 VDD.n3825 37.0005
R20249 VDD.n3825 VDD.t235 37.0005
R20250 VDD.n3819 VDD.n3818 37.0005
R20251 VDD.n3818 VDD.t235 37.0005
R20252 VDD.n2993 VDD.n2992 37.0005
R20253 VDD.t941 VDD.n2993 37.0005
R20254 VDD.n3938 VDD.n2991 37.0005
R20255 VDD.n2999 VDD.n2997 37.0005
R20256 VDD.n2997 VDD.t528 37.0005
R20257 VDD.n3930 VDD.n2998 37.0005
R20258 VDD.n2998 VDD.t528 37.0005
R20259 VDD.n3010 VDD.n3008 37.0005
R20260 VDD.n3008 VDD.t151 37.0005
R20261 VDD.n3920 VDD.n3009 37.0005
R20262 VDD.n3009 VDD.t151 37.0005
R20263 VDD.n3020 VDD.n3018 37.0005
R20264 VDD.n3018 VDD.t1014 37.0005
R20265 VDD.n3910 VDD.n3019 37.0005
R20266 VDD.n3019 VDD.t1014 37.0005
R20267 VDD.n3033 VDD.n3031 37.0005
R20268 VDD.n3031 VDD.t484 37.0005
R20269 VDD.n3900 VDD.n3032 37.0005
R20270 VDD.n3032 VDD.t484 37.0005
R20271 VDD.n3884 VDD.n3883 37.0005
R20272 VDD.t231 VDD.n3884 37.0005
R20273 VDD.n3886 VDD.n3743 37.0005
R20274 VDD.t231 VDD.n3743 37.0005
R20275 VDD.n3765 VDD.n3763 37.0005
R20276 VDD.n3763 VDD.t284 37.0005
R20277 VDD.n3866 VDD.n3764 37.0005
R20278 VDD.n3764 VDD.t284 37.0005
R20279 VDD.n3777 VDD.n3775 37.0005
R20280 VDD.n3775 VDD.t558 37.0005
R20281 VDD.n3856 VDD.n3776 37.0005
R20282 VDD.n3776 VDD.t558 37.0005
R20283 VDD.n3790 VDD.n3788 37.0005
R20284 VDD.n3788 VDD.t445 37.0005
R20285 VDD.n3846 VDD.n3789 37.0005
R20286 VDD.n3789 VDD.t445 37.0005
R20287 VDD.n3801 VDD.n3799 37.0005
R20288 VDD.n3799 VDD.t427 37.0005
R20289 VDD.n3836 VDD.n3800 37.0005
R20290 VDD.n3800 VDD.t427 37.0005
R20291 VDD.n3811 VDD.n3809 37.0005
R20292 VDD.n3809 VDD.t235 37.0005
R20293 VDD.n3826 VDD.n3810 37.0005
R20294 VDD.n3810 VDD.t235 37.0005
R20295 VDD.n3735 VDD.n3733 37.0005
R20296 VDD.n3733 VDD.t51 37.0005
R20297 VDD.n3890 VDD.n3738 37.0005
R20298 VDD.n3738 VDD.t51 37.0005
R20299 VDD.n3890 VDD.n3734 37.0005
R20300 VDD.n3734 VDD.t51 37.0005
R20301 VDD.n329 VDD.n328 36.7882
R20302 VDD.n3726 VDD.n3707 34.7977
R20303 VDD.n341 VDD.n285 34.146
R20304 VDD.n7130 VDD.n6887 33.6641
R20305 VDD.n3686 VDD.n3685 33.3344
R20306 VDD.n3199 VDD.n3135 33.3344
R20307 VDD.n42 VDD.n40 31.6493
R20308 VDD.n1647 VDD.n1643 31.6493
R20309 VDD.n1387 VDD.n1383 31.6493
R20310 VDD.n1127 VDD.n1123 31.6493
R20311 VDD.n867 VDD.n863 31.6493
R20312 VDD.n607 VDD.n603 31.6493
R20313 VDD.n347 VDD.n343 31.6493
R20314 VDD.n7263 VDD.n7259 31.6493
R20315 VDD.n1907 VDD.n1903 31.6493
R20316 VDD.n6022 VDD.n6020 31.6493
R20317 VDD.n5886 VDD.n5884 31.6493
R20318 VDD.n5750 VDD.n5748 31.6493
R20319 VDD.n5614 VDD.n5612 31.6493
R20320 VDD.n5478 VDD.n5476 31.6493
R20321 VDD.n5342 VDD.n5340 31.6493
R20322 VDD.n5206 VDD.n5204 31.6493
R20323 VDD.n5068 VDD.n4817 31.6493
R20324 VDD.n2043 VDD.n2039 31.6493
R20325 VDD.n2179 VDD.n2175 31.6493
R20326 VDD.n2315 VDD.n2311 31.6493
R20327 VDD.n2451 VDD.n2447 31.6493
R20328 VDD.n2587 VDD.n2583 31.6493
R20329 VDD.n2723 VDD.n2719 31.6493
R20330 VDD.n2859 VDD.n2855 31.6493
R20331 VDD.n2995 VDD.n2991 31.6493
R20332 VDD.n324 VDD.n323 31.0857
R20333 VDD.n3685 VDD.n3644 29.9244
R20334 VDD.n3644 VDD.n3057 29.9244
R20335 VDD.n3241 VDD.n3057 29.9244
R20336 VDD.n3241 VDD.n3240 29.9244
R20337 VDD.n3240 VDD.n3199 29.9244
R20338 VDD.n3196 VDD.n3096 29.9244
R20339 VDD.n3263 VDD.n3096 29.9244
R20340 VDD.n3640 VDD.n3263 29.9244
R20341 VDD.n3641 VDD.n3640 29.9244
R20342 VDD.n3641 VDD.n3037 29.9244
R20343 VDD.n3707 VDD.n3037 29.9244
R20344 VDD.n3195 VDD.n3194 29.7994
R20345 VDD.n147 VDD.n144 28.7118
R20346 VDD.n142 VDD.n138 28.7118
R20347 VDD.n161 VDD.n131 28.7118
R20348 VDD.n126 VDD.n122 28.7118
R20349 VDD.n182 VDD.n119 28.7118
R20350 VDD.n117 VDD.n113 28.7118
R20351 VDD.n196 VDD.n106 28.7118
R20352 VDD.n101 VDD.n97 28.7118
R20353 VDD.n217 VDD.n94 28.7118
R20354 VDD.n92 VDD.n88 28.7118
R20355 VDD.n231 VDD.n81 28.7118
R20356 VDD.n76 VDD.n72 28.7118
R20357 VDD.n252 VDD.n69 28.7118
R20358 VDD.n67 VDD.n63 28.7118
R20359 VDD.n266 VDD.n56 28.7118
R20360 VDD.n51 VDD.n47 28.7118
R20361 VDD.n6996 VDD.n6993 28.7118
R20362 VDD.n6991 VDD.n6987 28.7118
R20363 VDD.n7010 VDD.n6980 28.7118
R20364 VDD.n6975 VDD.n6971 28.7118
R20365 VDD.n7031 VDD.n6968 28.7118
R20366 VDD.n6966 VDD.n6962 28.7118
R20367 VDD.n7045 VDD.n6955 28.7118
R20368 VDD.n6950 VDD.n6946 28.7118
R20369 VDD.n7066 VDD.n6943 28.7118
R20370 VDD.n6941 VDD.n6937 28.7118
R20371 VDD.n7080 VDD.n6930 28.7118
R20372 VDD.n6925 VDD.n6921 28.7118
R20373 VDD.n7101 VDD.n6918 28.7118
R20374 VDD.n6916 VDD.n6912 28.7118
R20375 VDD.n7115 VDD.n6908 28.7118
R20376 VDD.n6899 VDD.n6895 28.7118
R20377 VDD.n3445 VDD.n3344 28.7118
R20378 VDD.n3428 VDD.n3424 28.7118
R20379 VDD.n3482 VDD.n3453 28.7118
R20380 VDD.n3466 VDD.n3462 28.7118
R20381 VDD.n3334 VDD.n3327 28.7118
R20382 VDD.n3321 VDD.n3317 28.7118
R20383 VDD.n3540 VDD.n3307 28.7118
R20384 VDD.n3523 VDD.n3519 28.7118
R20385 VDD.n3576 VDD.n3547 28.7118
R20386 VDD.n3560 VDD.n3556 28.7118
R20387 VDD.n3390 VDD.n3383 28.7118
R20388 VDD.n3377 VDD.n3373 28.7118
R20389 VDD VDD.n263 26.3103
R20390 VDD VDD.n249 26.3103
R20391 VDD VDD.n228 26.3103
R20392 VDD VDD.n214 26.3103
R20393 VDD VDD.n193 26.3103
R20394 VDD VDD.n179 26.3103
R20395 VDD VDD.n158 26.3103
R20396 VDD VDD.n7112 26.3103
R20397 VDD VDD.n7098 26.3103
R20398 VDD VDD.n7077 26.3103
R20399 VDD VDD.n7063 26.3103
R20400 VDD VDD.n7042 26.3103
R20401 VDD VDD.n7028 26.3103
R20402 VDD VDD.n7007 26.3103
R20403 VDD.n3198 VDD.n3197 25.8669
R20404 VDD.n3239 VDD.n3238 25.8669
R20405 VDD.n3262 VDD.n3242 25.8669
R20406 VDD.n3643 VDD.n3642 25.8669
R20407 VDD.n3684 VDD.n3683 25.8669
R20408 VDD.n3706 VDD.n3686 25.8669
R20409 VDD.n3193 VDD.n3135 25.8669
R20410 VDD.n329 VDD.n299 24.6676
R20411 VDD.n3305 VDD 24.3918
R20412 VDD.t89 VDD.n301 23.5846
R20413 VDD.n301 VDD.t786 23.5846
R20414 VDD.n336 VDD.t786 23.5846
R20415 VDD.t401 VDD.n337 23.5846
R20416 VDD.n7529 VDD.n38 23.1255
R20417 VDD.n7529 VDD.n7528 23.1255
R20418 VDD.n33 VDD.n29 23.1255
R20419 VDD.n7535 VDD.n29 23.1255
R20420 VDD.n7539 VDD.n28 23.1255
R20421 VDD.n7539 VDD.n7538 23.1255
R20422 VDD.n20 VDD.n16 23.1255
R20423 VDD.n7545 VDD.n16 23.1255
R20424 VDD.n7549 VDD.n15 23.1255
R20425 VDD.n7549 VDD.n7548 23.1255
R20426 VDD.n11 VDD.n7 23.1255
R20427 VDD.n7555 VDD.n7 23.1255
R20428 VDD.n7557 VDD.n5 23.1255
R20429 VDD.n7556 VDD.n5 23.1255
R20430 VDD.n7558 VDD.n6 23.1255
R20431 VDD.n7722 VDD.n6 23.1255
R20432 VDD.n7565 VDD.n7561 23.1255
R20433 VDD.n7721 VDD.n7561 23.1255
R20434 VDD.n7715 VDD.n7569 23.1255
R20435 VDD.n7715 VDD.n7714 23.1255
R20436 VDD.n7574 VDD.n7570 23.1255
R20437 VDD.n7711 VDD.n7570 23.1255
R20438 VDD.n7705 VDD.n7582 23.1255
R20439 VDD.n7705 VDD.n7704 23.1255
R20440 VDD.n7700 VDD.n7699 23.1255
R20441 VDD.n7701 VDD.n7700 23.1255
R20442 VDD.n7697 VDD.n7696 23.1255
R20443 VDD.n7696 VDD.n7695 23.1255
R20444 VDD.n7590 VDD.n7586 23.1255
R20445 VDD.n7694 VDD.n7586 23.1255
R20446 VDD.n7688 VDD.n7597 23.1255
R20447 VDD.n7688 VDD.n7687 23.1255
R20448 VDD.n7602 VDD.n7598 23.1255
R20449 VDD.n7684 VDD.n7598 23.1255
R20450 VDD.n7678 VDD.n7610 23.1255
R20451 VDD.n7678 VDD.n7677 23.1255
R20452 VDD.n7615 VDD.n7611 23.1255
R20453 VDD.n7674 VDD.n7611 23.1255
R20454 VDD.n7668 VDD.n7621 23.1255
R20455 VDD.n7668 VDD.n7667 23.1255
R20456 VDD.n7626 VDD.n7622 23.1255
R20457 VDD.n7664 VDD.n7622 23.1255
R20458 VDD.n7658 VDD.n7631 23.1255
R20459 VDD.n7658 VDD.n7657 23.1255
R20460 VDD.n7636 VDD.n7632 23.1255
R20461 VDD.n7654 VDD.n7632 23.1255
R20462 VDD.n7648 VDD.n7644 23.1255
R20463 VDD.n7648 VDD.n7647 23.1255
R20464 VDD.n7527 VDD.n7526 23.1255
R20465 VDD.n7528 VDD.n7527 23.1255
R20466 VDD.n7534 VDD.n7533 23.1255
R20467 VDD.n7535 VDD.n7534 23.1255
R20468 VDD.n7537 VDD.n7536 23.1255
R20469 VDD.n7538 VDD.n7537 23.1255
R20470 VDD.n7544 VDD.n7543 23.1255
R20471 VDD.n7545 VDD.n7544 23.1255
R20472 VDD.n7547 VDD.n7546 23.1255
R20473 VDD.n7548 VDD.n7547 23.1255
R20474 VDD.n7554 VDD.n7553 23.1255
R20475 VDD.n7555 VDD.n7554 23.1255
R20476 VDD.n7725 VDD.n7723 23.1255
R20477 VDD.n7723 VDD.n7556 23.1255
R20478 VDD.n7726 VDD.n7724 23.1255
R20479 VDD.n7724 VDD.n7722 23.1255
R20480 VDD.n7720 VDD.n7719 23.1255
R20481 VDD.n7721 VDD.n7720 23.1255
R20482 VDD.n7713 VDD.n7712 23.1255
R20483 VDD.n7714 VDD.n7713 23.1255
R20484 VDD.n7710 VDD.n7709 23.1255
R20485 VDD.n7711 VDD.n7710 23.1255
R20486 VDD.n7703 VDD.n7702 23.1255
R20487 VDD.n7704 VDD.n7703 23.1255
R20488 VDD.n7693 VDD.n7692 23.1255
R20489 VDD.n7694 VDD.n7693 23.1255
R20490 VDD.n7686 VDD.n7685 23.1255
R20491 VDD.n7687 VDD.n7686 23.1255
R20492 VDD.n7683 VDD.n7682 23.1255
R20493 VDD.n7684 VDD.n7683 23.1255
R20494 VDD.n7676 VDD.n7675 23.1255
R20495 VDD.n7677 VDD.n7676 23.1255
R20496 VDD.n7673 VDD.n7672 23.1255
R20497 VDD.n7674 VDD.n7673 23.1255
R20498 VDD.n7666 VDD.n7665 23.1255
R20499 VDD.n7667 VDD.n7666 23.1255
R20500 VDD.n7663 VDD.n7662 23.1255
R20501 VDD.n7664 VDD.n7663 23.1255
R20502 VDD.n7656 VDD.n7655 23.1255
R20503 VDD.n7657 VDD.n7656 23.1255
R20504 VDD.n7653 VDD.n7652 23.1255
R20505 VDD.n7654 VDD.n7653 23.1255
R20506 VDD.n7646 VDD.n7645 23.1255
R20507 VDD.n7647 VDD.n7646 23.1255
R20508 VDD.n7524 VDD.n7523 23.1255
R20509 VDD.n7525 VDD.n7524 23.1255
R20510 VDD.n44 VDD.n43 23.1255
R20511 VDD.n1652 VDD.n1648 23.1255
R20512 VDD.n1894 VDD.n1648 23.1255
R20513 VDD.n1888 VDD.n1658 23.1255
R20514 VDD.n1888 VDD.n1887 23.1255
R20515 VDD.n1663 VDD.n1659 23.1255
R20516 VDD.n1884 VDD.n1659 23.1255
R20517 VDD.n1878 VDD.n1668 23.1255
R20518 VDD.n1878 VDD.n1877 23.1255
R20519 VDD.n1673 VDD.n1669 23.1255
R20520 VDD.n1874 VDD.n1669 23.1255
R20521 VDD.n1868 VDD.n1681 23.1255
R20522 VDD.n1868 VDD.n1867 23.1255
R20523 VDD.n1686 VDD.n1682 23.1255
R20524 VDD.n1864 VDD.n1682 23.1255
R20525 VDD.n1858 VDD.n1692 23.1255
R20526 VDD.n1858 VDD.n1857 23.1255
R20527 VDD.n1697 VDD.n1693 23.1255
R20528 VDD.n1854 VDD.n1693 23.1255
R20529 VDD.n1848 VDD.n1702 23.1255
R20530 VDD.n1848 VDD.n1847 23.1255
R20531 VDD.n1707 VDD.n1703 23.1255
R20532 VDD.n1844 VDD.n1703 23.1255
R20533 VDD.n1838 VDD.n1715 23.1255
R20534 VDD.n1838 VDD.n1837 23.1255
R20535 VDD.n1833 VDD.n1832 23.1255
R20536 VDD.n1834 VDD.n1833 23.1255
R20537 VDD.n1830 VDD.n1829 23.1255
R20538 VDD.n1829 VDD.n1828 23.1255
R20539 VDD.n1723 VDD.n1719 23.1255
R20540 VDD.n1827 VDD.n1719 23.1255
R20541 VDD.n1821 VDD.n1730 23.1255
R20542 VDD.n1821 VDD.n1820 23.1255
R20543 VDD.n1735 VDD.n1731 23.1255
R20544 VDD.n1817 VDD.n1731 23.1255
R20545 VDD.n1811 VDD.n1743 23.1255
R20546 VDD.n1811 VDD.n1810 23.1255
R20547 VDD.n1748 VDD.n1744 23.1255
R20548 VDD.n1807 VDD.n1744 23.1255
R20549 VDD.n1801 VDD.n1754 23.1255
R20550 VDD.n1801 VDD.n1800 23.1255
R20551 VDD.n1759 VDD.n1755 23.1255
R20552 VDD.n1797 VDD.n1755 23.1255
R20553 VDD.n1791 VDD.n1764 23.1255
R20554 VDD.n1791 VDD.n1790 23.1255
R20555 VDD.n1769 VDD.n1765 23.1255
R20556 VDD.n1787 VDD.n1765 23.1255
R20557 VDD.n1781 VDD.n1777 23.1255
R20558 VDD.n1781 VDD.n1780 23.1255
R20559 VDD.n1893 VDD.n1892 23.1255
R20560 VDD.n1894 VDD.n1893 23.1255
R20561 VDD.n1886 VDD.n1885 23.1255
R20562 VDD.n1887 VDD.n1886 23.1255
R20563 VDD.n1883 VDD.n1882 23.1255
R20564 VDD.n1884 VDD.n1883 23.1255
R20565 VDD.n1876 VDD.n1875 23.1255
R20566 VDD.n1877 VDD.n1876 23.1255
R20567 VDD.n1873 VDD.n1872 23.1255
R20568 VDD.n1874 VDD.n1873 23.1255
R20569 VDD.n1866 VDD.n1865 23.1255
R20570 VDD.n1867 VDD.n1866 23.1255
R20571 VDD.n1863 VDD.n1862 23.1255
R20572 VDD.n1864 VDD.n1863 23.1255
R20573 VDD.n1856 VDD.n1855 23.1255
R20574 VDD.n1857 VDD.n1856 23.1255
R20575 VDD.n1853 VDD.n1852 23.1255
R20576 VDD.n1854 VDD.n1853 23.1255
R20577 VDD.n1846 VDD.n1845 23.1255
R20578 VDD.n1847 VDD.n1846 23.1255
R20579 VDD.n1843 VDD.n1842 23.1255
R20580 VDD.n1844 VDD.n1843 23.1255
R20581 VDD.n1836 VDD.n1835 23.1255
R20582 VDD.n1837 VDD.n1836 23.1255
R20583 VDD.n1826 VDD.n1825 23.1255
R20584 VDD.n1827 VDD.n1826 23.1255
R20585 VDD.n1819 VDD.n1818 23.1255
R20586 VDD.n1820 VDD.n1819 23.1255
R20587 VDD.n1816 VDD.n1815 23.1255
R20588 VDD.n1817 VDD.n1816 23.1255
R20589 VDD.n1809 VDD.n1808 23.1255
R20590 VDD.n1810 VDD.n1809 23.1255
R20591 VDD.n1806 VDD.n1805 23.1255
R20592 VDD.n1807 VDD.n1806 23.1255
R20593 VDD.n1799 VDD.n1798 23.1255
R20594 VDD.n1800 VDD.n1799 23.1255
R20595 VDD.n1796 VDD.n1795 23.1255
R20596 VDD.n1797 VDD.n1796 23.1255
R20597 VDD.n1789 VDD.n1788 23.1255
R20598 VDD.n1790 VDD.n1789 23.1255
R20599 VDD.n1786 VDD.n1785 23.1255
R20600 VDD.n1787 VDD.n1786 23.1255
R20601 VDD.n1779 VDD.n1778 23.1255
R20602 VDD.n1780 VDD.n1779 23.1255
R20603 VDD.n1897 VDD.n1896 23.1255
R20604 VDD.n1896 VDD.n1895 23.1255
R20605 VDD.n1646 VDD.n1642 23.1255
R20606 VDD.n1392 VDD.n1388 23.1255
R20607 VDD.n1634 VDD.n1388 23.1255
R20608 VDD.n1628 VDD.n1398 23.1255
R20609 VDD.n1628 VDD.n1627 23.1255
R20610 VDD.n1403 VDD.n1399 23.1255
R20611 VDD.n1624 VDD.n1399 23.1255
R20612 VDD.n1618 VDD.n1408 23.1255
R20613 VDD.n1618 VDD.n1617 23.1255
R20614 VDD.n1413 VDD.n1409 23.1255
R20615 VDD.n1614 VDD.n1409 23.1255
R20616 VDD.n1608 VDD.n1421 23.1255
R20617 VDD.n1608 VDD.n1607 23.1255
R20618 VDD.n1426 VDD.n1422 23.1255
R20619 VDD.n1604 VDD.n1422 23.1255
R20620 VDD.n1598 VDD.n1432 23.1255
R20621 VDD.n1598 VDD.n1597 23.1255
R20622 VDD.n1437 VDD.n1433 23.1255
R20623 VDD.n1594 VDD.n1433 23.1255
R20624 VDD.n1588 VDD.n1442 23.1255
R20625 VDD.n1588 VDD.n1587 23.1255
R20626 VDD.n1447 VDD.n1443 23.1255
R20627 VDD.n1584 VDD.n1443 23.1255
R20628 VDD.n1578 VDD.n1455 23.1255
R20629 VDD.n1578 VDD.n1577 23.1255
R20630 VDD.n1573 VDD.n1572 23.1255
R20631 VDD.n1574 VDD.n1573 23.1255
R20632 VDD.n1570 VDD.n1569 23.1255
R20633 VDD.n1569 VDD.n1568 23.1255
R20634 VDD.n1463 VDD.n1459 23.1255
R20635 VDD.n1567 VDD.n1459 23.1255
R20636 VDD.n1561 VDD.n1470 23.1255
R20637 VDD.n1561 VDD.n1560 23.1255
R20638 VDD.n1475 VDD.n1471 23.1255
R20639 VDD.n1557 VDD.n1471 23.1255
R20640 VDD.n1551 VDD.n1483 23.1255
R20641 VDD.n1551 VDD.n1550 23.1255
R20642 VDD.n1488 VDD.n1484 23.1255
R20643 VDD.n1547 VDD.n1484 23.1255
R20644 VDD.n1541 VDD.n1494 23.1255
R20645 VDD.n1541 VDD.n1540 23.1255
R20646 VDD.n1499 VDD.n1495 23.1255
R20647 VDD.n1537 VDD.n1495 23.1255
R20648 VDD.n1531 VDD.n1504 23.1255
R20649 VDD.n1531 VDD.n1530 23.1255
R20650 VDD.n1509 VDD.n1505 23.1255
R20651 VDD.n1527 VDD.n1505 23.1255
R20652 VDD.n1521 VDD.n1517 23.1255
R20653 VDD.n1521 VDD.n1520 23.1255
R20654 VDD.n1633 VDD.n1632 23.1255
R20655 VDD.n1634 VDD.n1633 23.1255
R20656 VDD.n1626 VDD.n1625 23.1255
R20657 VDD.n1627 VDD.n1626 23.1255
R20658 VDD.n1623 VDD.n1622 23.1255
R20659 VDD.n1624 VDD.n1623 23.1255
R20660 VDD.n1616 VDD.n1615 23.1255
R20661 VDD.n1617 VDD.n1616 23.1255
R20662 VDD.n1613 VDD.n1612 23.1255
R20663 VDD.n1614 VDD.n1613 23.1255
R20664 VDD.n1606 VDD.n1605 23.1255
R20665 VDD.n1607 VDD.n1606 23.1255
R20666 VDD.n1603 VDD.n1602 23.1255
R20667 VDD.n1604 VDD.n1603 23.1255
R20668 VDD.n1596 VDD.n1595 23.1255
R20669 VDD.n1597 VDD.n1596 23.1255
R20670 VDD.n1593 VDD.n1592 23.1255
R20671 VDD.n1594 VDD.n1593 23.1255
R20672 VDD.n1586 VDD.n1585 23.1255
R20673 VDD.n1587 VDD.n1586 23.1255
R20674 VDD.n1583 VDD.n1582 23.1255
R20675 VDD.n1584 VDD.n1583 23.1255
R20676 VDD.n1576 VDD.n1575 23.1255
R20677 VDD.n1577 VDD.n1576 23.1255
R20678 VDD.n1566 VDD.n1565 23.1255
R20679 VDD.n1567 VDD.n1566 23.1255
R20680 VDD.n1559 VDD.n1558 23.1255
R20681 VDD.n1560 VDD.n1559 23.1255
R20682 VDD.n1556 VDD.n1555 23.1255
R20683 VDD.n1557 VDD.n1556 23.1255
R20684 VDD.n1549 VDD.n1548 23.1255
R20685 VDD.n1550 VDD.n1549 23.1255
R20686 VDD.n1546 VDD.n1545 23.1255
R20687 VDD.n1547 VDD.n1546 23.1255
R20688 VDD.n1539 VDD.n1538 23.1255
R20689 VDD.n1540 VDD.n1539 23.1255
R20690 VDD.n1536 VDD.n1535 23.1255
R20691 VDD.n1537 VDD.n1536 23.1255
R20692 VDD.n1529 VDD.n1528 23.1255
R20693 VDD.n1530 VDD.n1529 23.1255
R20694 VDD.n1526 VDD.n1525 23.1255
R20695 VDD.n1527 VDD.n1526 23.1255
R20696 VDD.n1519 VDD.n1518 23.1255
R20697 VDD.n1520 VDD.n1519 23.1255
R20698 VDD.n1637 VDD.n1636 23.1255
R20699 VDD.n1636 VDD.n1635 23.1255
R20700 VDD.n1386 VDD.n1382 23.1255
R20701 VDD.n1132 VDD.n1128 23.1255
R20702 VDD.n1374 VDD.n1128 23.1255
R20703 VDD.n1368 VDD.n1138 23.1255
R20704 VDD.n1368 VDD.n1367 23.1255
R20705 VDD.n1143 VDD.n1139 23.1255
R20706 VDD.n1364 VDD.n1139 23.1255
R20707 VDD.n1358 VDD.n1148 23.1255
R20708 VDD.n1358 VDD.n1357 23.1255
R20709 VDD.n1153 VDD.n1149 23.1255
R20710 VDD.n1354 VDD.n1149 23.1255
R20711 VDD.n1348 VDD.n1161 23.1255
R20712 VDD.n1348 VDD.n1347 23.1255
R20713 VDD.n1166 VDD.n1162 23.1255
R20714 VDD.n1344 VDD.n1162 23.1255
R20715 VDD.n1338 VDD.n1172 23.1255
R20716 VDD.n1338 VDD.n1337 23.1255
R20717 VDD.n1177 VDD.n1173 23.1255
R20718 VDD.n1334 VDD.n1173 23.1255
R20719 VDD.n1328 VDD.n1182 23.1255
R20720 VDD.n1328 VDD.n1327 23.1255
R20721 VDD.n1187 VDD.n1183 23.1255
R20722 VDD.n1324 VDD.n1183 23.1255
R20723 VDD.n1318 VDD.n1195 23.1255
R20724 VDD.n1318 VDD.n1317 23.1255
R20725 VDD.n1313 VDD.n1312 23.1255
R20726 VDD.n1314 VDD.n1313 23.1255
R20727 VDD.n1310 VDD.n1309 23.1255
R20728 VDD.n1309 VDD.n1308 23.1255
R20729 VDD.n1203 VDD.n1199 23.1255
R20730 VDD.n1307 VDD.n1199 23.1255
R20731 VDD.n1301 VDD.n1210 23.1255
R20732 VDD.n1301 VDD.n1300 23.1255
R20733 VDD.n1215 VDD.n1211 23.1255
R20734 VDD.n1297 VDD.n1211 23.1255
R20735 VDD.n1291 VDD.n1223 23.1255
R20736 VDD.n1291 VDD.n1290 23.1255
R20737 VDD.n1228 VDD.n1224 23.1255
R20738 VDD.n1287 VDD.n1224 23.1255
R20739 VDD.n1281 VDD.n1234 23.1255
R20740 VDD.n1281 VDD.n1280 23.1255
R20741 VDD.n1239 VDD.n1235 23.1255
R20742 VDD.n1277 VDD.n1235 23.1255
R20743 VDD.n1271 VDD.n1244 23.1255
R20744 VDD.n1271 VDD.n1270 23.1255
R20745 VDD.n1249 VDD.n1245 23.1255
R20746 VDD.n1267 VDD.n1245 23.1255
R20747 VDD.n1261 VDD.n1257 23.1255
R20748 VDD.n1261 VDD.n1260 23.1255
R20749 VDD.n1373 VDD.n1372 23.1255
R20750 VDD.n1374 VDD.n1373 23.1255
R20751 VDD.n1366 VDD.n1365 23.1255
R20752 VDD.n1367 VDD.n1366 23.1255
R20753 VDD.n1363 VDD.n1362 23.1255
R20754 VDD.n1364 VDD.n1363 23.1255
R20755 VDD.n1356 VDD.n1355 23.1255
R20756 VDD.n1357 VDD.n1356 23.1255
R20757 VDD.n1353 VDD.n1352 23.1255
R20758 VDD.n1354 VDD.n1353 23.1255
R20759 VDD.n1346 VDD.n1345 23.1255
R20760 VDD.n1347 VDD.n1346 23.1255
R20761 VDD.n1343 VDD.n1342 23.1255
R20762 VDD.n1344 VDD.n1343 23.1255
R20763 VDD.n1336 VDD.n1335 23.1255
R20764 VDD.n1337 VDD.n1336 23.1255
R20765 VDD.n1333 VDD.n1332 23.1255
R20766 VDD.n1334 VDD.n1333 23.1255
R20767 VDD.n1326 VDD.n1325 23.1255
R20768 VDD.n1327 VDD.n1326 23.1255
R20769 VDD.n1323 VDD.n1322 23.1255
R20770 VDD.n1324 VDD.n1323 23.1255
R20771 VDD.n1316 VDD.n1315 23.1255
R20772 VDD.n1317 VDD.n1316 23.1255
R20773 VDD.n1306 VDD.n1305 23.1255
R20774 VDD.n1307 VDD.n1306 23.1255
R20775 VDD.n1299 VDD.n1298 23.1255
R20776 VDD.n1300 VDD.n1299 23.1255
R20777 VDD.n1296 VDD.n1295 23.1255
R20778 VDD.n1297 VDD.n1296 23.1255
R20779 VDD.n1289 VDD.n1288 23.1255
R20780 VDD.n1290 VDD.n1289 23.1255
R20781 VDD.n1286 VDD.n1285 23.1255
R20782 VDD.n1287 VDD.n1286 23.1255
R20783 VDD.n1279 VDD.n1278 23.1255
R20784 VDD.n1280 VDD.n1279 23.1255
R20785 VDD.n1276 VDD.n1275 23.1255
R20786 VDD.n1277 VDD.n1276 23.1255
R20787 VDD.n1269 VDD.n1268 23.1255
R20788 VDD.n1270 VDD.n1269 23.1255
R20789 VDD.n1266 VDD.n1265 23.1255
R20790 VDD.n1267 VDD.n1266 23.1255
R20791 VDD.n1259 VDD.n1258 23.1255
R20792 VDD.n1260 VDD.n1259 23.1255
R20793 VDD.n1377 VDD.n1376 23.1255
R20794 VDD.n1376 VDD.n1375 23.1255
R20795 VDD.n1126 VDD.n1122 23.1255
R20796 VDD.n872 VDD.n868 23.1255
R20797 VDD.n1114 VDD.n868 23.1255
R20798 VDD.n1108 VDD.n878 23.1255
R20799 VDD.n1108 VDD.n1107 23.1255
R20800 VDD.n883 VDD.n879 23.1255
R20801 VDD.n1104 VDD.n879 23.1255
R20802 VDD.n1098 VDD.n888 23.1255
R20803 VDD.n1098 VDD.n1097 23.1255
R20804 VDD.n893 VDD.n889 23.1255
R20805 VDD.n1094 VDD.n889 23.1255
R20806 VDD.n1088 VDD.n901 23.1255
R20807 VDD.n1088 VDD.n1087 23.1255
R20808 VDD.n906 VDD.n902 23.1255
R20809 VDD.n1084 VDD.n902 23.1255
R20810 VDD.n1078 VDD.n912 23.1255
R20811 VDD.n1078 VDD.n1077 23.1255
R20812 VDD.n917 VDD.n913 23.1255
R20813 VDD.n1074 VDD.n913 23.1255
R20814 VDD.n1068 VDD.n922 23.1255
R20815 VDD.n1068 VDD.n1067 23.1255
R20816 VDD.n927 VDD.n923 23.1255
R20817 VDD.n1064 VDD.n923 23.1255
R20818 VDD.n1058 VDD.n935 23.1255
R20819 VDD.n1058 VDD.n1057 23.1255
R20820 VDD.n1053 VDD.n1052 23.1255
R20821 VDD.n1054 VDD.n1053 23.1255
R20822 VDD.n1050 VDD.n1049 23.1255
R20823 VDD.n1049 VDD.n1048 23.1255
R20824 VDD.n943 VDD.n939 23.1255
R20825 VDD.n1047 VDD.n939 23.1255
R20826 VDD.n1041 VDD.n950 23.1255
R20827 VDD.n1041 VDD.n1040 23.1255
R20828 VDD.n955 VDD.n951 23.1255
R20829 VDD.n1037 VDD.n951 23.1255
R20830 VDD.n1031 VDD.n963 23.1255
R20831 VDD.n1031 VDD.n1030 23.1255
R20832 VDD.n968 VDD.n964 23.1255
R20833 VDD.n1027 VDD.n964 23.1255
R20834 VDD.n1021 VDD.n974 23.1255
R20835 VDD.n1021 VDD.n1020 23.1255
R20836 VDD.n979 VDD.n975 23.1255
R20837 VDD.n1017 VDD.n975 23.1255
R20838 VDD.n1011 VDD.n984 23.1255
R20839 VDD.n1011 VDD.n1010 23.1255
R20840 VDD.n989 VDD.n985 23.1255
R20841 VDD.n1007 VDD.n985 23.1255
R20842 VDD.n1001 VDD.n997 23.1255
R20843 VDD.n1001 VDD.n1000 23.1255
R20844 VDD.n1113 VDD.n1112 23.1255
R20845 VDD.n1114 VDD.n1113 23.1255
R20846 VDD.n1106 VDD.n1105 23.1255
R20847 VDD.n1107 VDD.n1106 23.1255
R20848 VDD.n1103 VDD.n1102 23.1255
R20849 VDD.n1104 VDD.n1103 23.1255
R20850 VDD.n1096 VDD.n1095 23.1255
R20851 VDD.n1097 VDD.n1096 23.1255
R20852 VDD.n1093 VDD.n1092 23.1255
R20853 VDD.n1094 VDD.n1093 23.1255
R20854 VDD.n1086 VDD.n1085 23.1255
R20855 VDD.n1087 VDD.n1086 23.1255
R20856 VDD.n1083 VDD.n1082 23.1255
R20857 VDD.n1084 VDD.n1083 23.1255
R20858 VDD.n1076 VDD.n1075 23.1255
R20859 VDD.n1077 VDD.n1076 23.1255
R20860 VDD.n1073 VDD.n1072 23.1255
R20861 VDD.n1074 VDD.n1073 23.1255
R20862 VDD.n1066 VDD.n1065 23.1255
R20863 VDD.n1067 VDD.n1066 23.1255
R20864 VDD.n1063 VDD.n1062 23.1255
R20865 VDD.n1064 VDD.n1063 23.1255
R20866 VDD.n1056 VDD.n1055 23.1255
R20867 VDD.n1057 VDD.n1056 23.1255
R20868 VDD.n1046 VDD.n1045 23.1255
R20869 VDD.n1047 VDD.n1046 23.1255
R20870 VDD.n1039 VDD.n1038 23.1255
R20871 VDD.n1040 VDD.n1039 23.1255
R20872 VDD.n1036 VDD.n1035 23.1255
R20873 VDD.n1037 VDD.n1036 23.1255
R20874 VDD.n1029 VDD.n1028 23.1255
R20875 VDD.n1030 VDD.n1029 23.1255
R20876 VDD.n1026 VDD.n1025 23.1255
R20877 VDD.n1027 VDD.n1026 23.1255
R20878 VDD.n1019 VDD.n1018 23.1255
R20879 VDD.n1020 VDD.n1019 23.1255
R20880 VDD.n1016 VDD.n1015 23.1255
R20881 VDD.n1017 VDD.n1016 23.1255
R20882 VDD.n1009 VDD.n1008 23.1255
R20883 VDD.n1010 VDD.n1009 23.1255
R20884 VDD.n1006 VDD.n1005 23.1255
R20885 VDD.n1007 VDD.n1006 23.1255
R20886 VDD.n999 VDD.n998 23.1255
R20887 VDD.n1000 VDD.n999 23.1255
R20888 VDD.n1117 VDD.n1116 23.1255
R20889 VDD.n1116 VDD.n1115 23.1255
R20890 VDD.n866 VDD.n862 23.1255
R20891 VDD.n612 VDD.n608 23.1255
R20892 VDD.n854 VDD.n608 23.1255
R20893 VDD.n848 VDD.n618 23.1255
R20894 VDD.n848 VDD.n847 23.1255
R20895 VDD.n623 VDD.n619 23.1255
R20896 VDD.n844 VDD.n619 23.1255
R20897 VDD.n838 VDD.n628 23.1255
R20898 VDD.n838 VDD.n837 23.1255
R20899 VDD.n633 VDD.n629 23.1255
R20900 VDD.n834 VDD.n629 23.1255
R20901 VDD.n828 VDD.n641 23.1255
R20902 VDD.n828 VDD.n827 23.1255
R20903 VDD.n646 VDD.n642 23.1255
R20904 VDD.n824 VDD.n642 23.1255
R20905 VDD.n818 VDD.n652 23.1255
R20906 VDD.n818 VDD.n817 23.1255
R20907 VDD.n657 VDD.n653 23.1255
R20908 VDD.n814 VDD.n653 23.1255
R20909 VDD.n808 VDD.n662 23.1255
R20910 VDD.n808 VDD.n807 23.1255
R20911 VDD.n667 VDD.n663 23.1255
R20912 VDD.n804 VDD.n663 23.1255
R20913 VDD.n798 VDD.n675 23.1255
R20914 VDD.n798 VDD.n797 23.1255
R20915 VDD.n793 VDD.n792 23.1255
R20916 VDD.n794 VDD.n793 23.1255
R20917 VDD.n790 VDD.n789 23.1255
R20918 VDD.n789 VDD.n788 23.1255
R20919 VDD.n683 VDD.n679 23.1255
R20920 VDD.n787 VDD.n679 23.1255
R20921 VDD.n781 VDD.n690 23.1255
R20922 VDD.n781 VDD.n780 23.1255
R20923 VDD.n695 VDD.n691 23.1255
R20924 VDD.n777 VDD.n691 23.1255
R20925 VDD.n771 VDD.n703 23.1255
R20926 VDD.n771 VDD.n770 23.1255
R20927 VDD.n708 VDD.n704 23.1255
R20928 VDD.n767 VDD.n704 23.1255
R20929 VDD.n761 VDD.n714 23.1255
R20930 VDD.n761 VDD.n760 23.1255
R20931 VDD.n719 VDD.n715 23.1255
R20932 VDD.n757 VDD.n715 23.1255
R20933 VDD.n751 VDD.n724 23.1255
R20934 VDD.n751 VDD.n750 23.1255
R20935 VDD.n729 VDD.n725 23.1255
R20936 VDD.n747 VDD.n725 23.1255
R20937 VDD.n741 VDD.n737 23.1255
R20938 VDD.n741 VDD.n740 23.1255
R20939 VDD.n853 VDD.n852 23.1255
R20940 VDD.n854 VDD.n853 23.1255
R20941 VDD.n846 VDD.n845 23.1255
R20942 VDD.n847 VDD.n846 23.1255
R20943 VDD.n843 VDD.n842 23.1255
R20944 VDD.n844 VDD.n843 23.1255
R20945 VDD.n836 VDD.n835 23.1255
R20946 VDD.n837 VDD.n836 23.1255
R20947 VDD.n833 VDD.n832 23.1255
R20948 VDD.n834 VDD.n833 23.1255
R20949 VDD.n826 VDD.n825 23.1255
R20950 VDD.n827 VDD.n826 23.1255
R20951 VDD.n823 VDD.n822 23.1255
R20952 VDD.n824 VDD.n823 23.1255
R20953 VDD.n816 VDD.n815 23.1255
R20954 VDD.n817 VDD.n816 23.1255
R20955 VDD.n813 VDD.n812 23.1255
R20956 VDD.n814 VDD.n813 23.1255
R20957 VDD.n806 VDD.n805 23.1255
R20958 VDD.n807 VDD.n806 23.1255
R20959 VDD.n803 VDD.n802 23.1255
R20960 VDD.n804 VDD.n803 23.1255
R20961 VDD.n796 VDD.n795 23.1255
R20962 VDD.n797 VDD.n796 23.1255
R20963 VDD.n786 VDD.n785 23.1255
R20964 VDD.n787 VDD.n786 23.1255
R20965 VDD.n779 VDD.n778 23.1255
R20966 VDD.n780 VDD.n779 23.1255
R20967 VDD.n776 VDD.n775 23.1255
R20968 VDD.n777 VDD.n776 23.1255
R20969 VDD.n769 VDD.n768 23.1255
R20970 VDD.n770 VDD.n769 23.1255
R20971 VDD.n766 VDD.n765 23.1255
R20972 VDD.n767 VDD.n766 23.1255
R20973 VDD.n759 VDD.n758 23.1255
R20974 VDD.n760 VDD.n759 23.1255
R20975 VDD.n756 VDD.n755 23.1255
R20976 VDD.n757 VDD.n756 23.1255
R20977 VDD.n749 VDD.n748 23.1255
R20978 VDD.n750 VDD.n749 23.1255
R20979 VDD.n746 VDD.n745 23.1255
R20980 VDD.n747 VDD.n746 23.1255
R20981 VDD.n739 VDD.n738 23.1255
R20982 VDD.n740 VDD.n739 23.1255
R20983 VDD.n857 VDD.n856 23.1255
R20984 VDD.n856 VDD.n855 23.1255
R20985 VDD.n606 VDD.n602 23.1255
R20986 VDD.n352 VDD.n348 23.1255
R20987 VDD.n594 VDD.n348 23.1255
R20988 VDD.n588 VDD.n358 23.1255
R20989 VDD.n588 VDD.n587 23.1255
R20990 VDD.n363 VDD.n359 23.1255
R20991 VDD.n584 VDD.n359 23.1255
R20992 VDD.n578 VDD.n368 23.1255
R20993 VDD.n578 VDD.n577 23.1255
R20994 VDD.n373 VDD.n369 23.1255
R20995 VDD.n574 VDD.n369 23.1255
R20996 VDD.n568 VDD.n381 23.1255
R20997 VDD.n568 VDD.n567 23.1255
R20998 VDD.n386 VDD.n382 23.1255
R20999 VDD.n564 VDD.n382 23.1255
R21000 VDD.n558 VDD.n392 23.1255
R21001 VDD.n558 VDD.n557 23.1255
R21002 VDD.n397 VDD.n393 23.1255
R21003 VDD.n554 VDD.n393 23.1255
R21004 VDD.n548 VDD.n402 23.1255
R21005 VDD.n548 VDD.n547 23.1255
R21006 VDD.n407 VDD.n403 23.1255
R21007 VDD.n544 VDD.n403 23.1255
R21008 VDD.n538 VDD.n415 23.1255
R21009 VDD.n538 VDD.n537 23.1255
R21010 VDD.n533 VDD.n532 23.1255
R21011 VDD.n534 VDD.n533 23.1255
R21012 VDD.n530 VDD.n529 23.1255
R21013 VDD.n529 VDD.n528 23.1255
R21014 VDD.n423 VDD.n419 23.1255
R21015 VDD.n527 VDD.n419 23.1255
R21016 VDD.n521 VDD.n430 23.1255
R21017 VDD.n521 VDD.n520 23.1255
R21018 VDD.n435 VDD.n431 23.1255
R21019 VDD.n517 VDD.n431 23.1255
R21020 VDD.n511 VDD.n443 23.1255
R21021 VDD.n511 VDD.n510 23.1255
R21022 VDD.n448 VDD.n444 23.1255
R21023 VDD.n507 VDD.n444 23.1255
R21024 VDD.n501 VDD.n454 23.1255
R21025 VDD.n501 VDD.n500 23.1255
R21026 VDD.n459 VDD.n455 23.1255
R21027 VDD.n497 VDD.n455 23.1255
R21028 VDD.n491 VDD.n464 23.1255
R21029 VDD.n491 VDD.n490 23.1255
R21030 VDD.n469 VDD.n465 23.1255
R21031 VDD.n487 VDD.n465 23.1255
R21032 VDD.n481 VDD.n477 23.1255
R21033 VDD.n481 VDD.n480 23.1255
R21034 VDD.n593 VDD.n592 23.1255
R21035 VDD.n594 VDD.n593 23.1255
R21036 VDD.n586 VDD.n585 23.1255
R21037 VDD.n587 VDD.n586 23.1255
R21038 VDD.n583 VDD.n582 23.1255
R21039 VDD.n584 VDD.n583 23.1255
R21040 VDD.n576 VDD.n575 23.1255
R21041 VDD.n577 VDD.n576 23.1255
R21042 VDD.n573 VDD.n572 23.1255
R21043 VDD.n574 VDD.n573 23.1255
R21044 VDD.n566 VDD.n565 23.1255
R21045 VDD.n567 VDD.n566 23.1255
R21046 VDD.n563 VDD.n562 23.1255
R21047 VDD.n564 VDD.n563 23.1255
R21048 VDD.n556 VDD.n555 23.1255
R21049 VDD.n557 VDD.n556 23.1255
R21050 VDD.n553 VDD.n552 23.1255
R21051 VDD.n554 VDD.n553 23.1255
R21052 VDD.n546 VDD.n545 23.1255
R21053 VDD.n547 VDD.n546 23.1255
R21054 VDD.n543 VDD.n542 23.1255
R21055 VDD.n544 VDD.n543 23.1255
R21056 VDD.n536 VDD.n535 23.1255
R21057 VDD.n537 VDD.n536 23.1255
R21058 VDD.n526 VDD.n525 23.1255
R21059 VDD.n527 VDD.n526 23.1255
R21060 VDD.n519 VDD.n518 23.1255
R21061 VDD.n520 VDD.n519 23.1255
R21062 VDD.n516 VDD.n515 23.1255
R21063 VDD.n517 VDD.n516 23.1255
R21064 VDD.n509 VDD.n508 23.1255
R21065 VDD.n510 VDD.n509 23.1255
R21066 VDD.n506 VDD.n505 23.1255
R21067 VDD.n507 VDD.n506 23.1255
R21068 VDD.n499 VDD.n498 23.1255
R21069 VDD.n500 VDD.n499 23.1255
R21070 VDD.n496 VDD.n495 23.1255
R21071 VDD.n497 VDD.n496 23.1255
R21072 VDD.n489 VDD.n488 23.1255
R21073 VDD.n490 VDD.n489 23.1255
R21074 VDD.n486 VDD.n485 23.1255
R21075 VDD.n487 VDD.n486 23.1255
R21076 VDD.n479 VDD.n478 23.1255
R21077 VDD.n480 VDD.n479 23.1255
R21078 VDD.n597 VDD.n596 23.1255
R21079 VDD.n596 VDD.n595 23.1255
R21080 VDD.n346 VDD.n342 23.1255
R21081 VDD.n152 VDD.n151 23.1255
R21082 VDD.n153 VDD.n152 23.1255
R21083 VDD.n149 VDD.n148 23.1255
R21084 VDD.n156 VDD.n155 23.1255
R21085 VDD.n155 VDD.n154 23.1255
R21086 VDD.n141 VDD.n137 23.1255
R21087 VDD.n173 VDD.n172 23.1255
R21088 VDD.n174 VDD.n173 23.1255
R21089 VDD.n170 VDD.n169 23.1255
R21090 VDD.n169 VDD.n168 23.1255
R21091 VDD.n166 VDD.n165 23.1255
R21092 VDD.n167 VDD.n166 23.1255
R21093 VDD.n163 VDD.n162 23.1255
R21094 VDD.n177 VDD.n176 23.1255
R21095 VDD.n176 VDD.n175 23.1255
R21096 VDD.n125 VDD.n121 23.1255
R21097 VDD.n187 VDD.n186 23.1255
R21098 VDD.n188 VDD.n187 23.1255
R21099 VDD.n184 VDD.n183 23.1255
R21100 VDD.n191 VDD.n190 23.1255
R21101 VDD.n190 VDD.n189 23.1255
R21102 VDD.n116 VDD.n112 23.1255
R21103 VDD.n208 VDD.n207 23.1255
R21104 VDD.n209 VDD.n208 23.1255
R21105 VDD.n205 VDD.n204 23.1255
R21106 VDD.n204 VDD.n203 23.1255
R21107 VDD.n201 VDD.n200 23.1255
R21108 VDD.n202 VDD.n201 23.1255
R21109 VDD.n198 VDD.n197 23.1255
R21110 VDD.n212 VDD.n211 23.1255
R21111 VDD.n211 VDD.n210 23.1255
R21112 VDD.n100 VDD.n96 23.1255
R21113 VDD.n222 VDD.n221 23.1255
R21114 VDD.n223 VDD.n222 23.1255
R21115 VDD.n219 VDD.n218 23.1255
R21116 VDD.n226 VDD.n225 23.1255
R21117 VDD.n225 VDD.n224 23.1255
R21118 VDD.n91 VDD.n87 23.1255
R21119 VDD.n243 VDD.n242 23.1255
R21120 VDD.n244 VDD.n243 23.1255
R21121 VDD.n240 VDD.n239 23.1255
R21122 VDD.n239 VDD.n238 23.1255
R21123 VDD.n236 VDD.n235 23.1255
R21124 VDD.n237 VDD.n236 23.1255
R21125 VDD.n233 VDD.n232 23.1255
R21126 VDD.n247 VDD.n246 23.1255
R21127 VDD.n246 VDD.n245 23.1255
R21128 VDD.n75 VDD.n71 23.1255
R21129 VDD.n257 VDD.n256 23.1255
R21130 VDD.n258 VDD.n257 23.1255
R21131 VDD.n254 VDD.n253 23.1255
R21132 VDD.n261 VDD.n260 23.1255
R21133 VDD.n260 VDD.n259 23.1255
R21134 VDD.n66 VDD.n62 23.1255
R21135 VDD.n278 VDD.n277 23.1255
R21136 VDD.n279 VDD.n278 23.1255
R21137 VDD.n275 VDD.n274 23.1255
R21138 VDD.n274 VDD.n273 23.1255
R21139 VDD.n271 VDD.n270 23.1255
R21140 VDD.n272 VDD.n271 23.1255
R21141 VDD.n268 VDD.n267 23.1255
R21142 VDD.n282 VDD.n281 23.1255
R21143 VDD.n281 VDD.n280 23.1255
R21144 VDD.n50 VDD.n46 23.1255
R21145 VDD.n7268 VDD.n7264 23.1255
R21146 VDD.n7510 VDD.n7264 23.1255
R21147 VDD.n7504 VDD.n7274 23.1255
R21148 VDD.n7504 VDD.n7503 23.1255
R21149 VDD.n7279 VDD.n7275 23.1255
R21150 VDD.n7500 VDD.n7275 23.1255
R21151 VDD.n7494 VDD.n7284 23.1255
R21152 VDD.n7494 VDD.n7493 23.1255
R21153 VDD.n7289 VDD.n7285 23.1255
R21154 VDD.n7490 VDD.n7285 23.1255
R21155 VDD.n7484 VDD.n7297 23.1255
R21156 VDD.n7484 VDD.n7483 23.1255
R21157 VDD.n7302 VDD.n7298 23.1255
R21158 VDD.n7480 VDD.n7298 23.1255
R21159 VDD.n7474 VDD.n7308 23.1255
R21160 VDD.n7474 VDD.n7473 23.1255
R21161 VDD.n7313 VDD.n7309 23.1255
R21162 VDD.n7470 VDD.n7309 23.1255
R21163 VDD.n7464 VDD.n7318 23.1255
R21164 VDD.n7464 VDD.n7463 23.1255
R21165 VDD.n7323 VDD.n7319 23.1255
R21166 VDD.n7460 VDD.n7319 23.1255
R21167 VDD.n7454 VDD.n7331 23.1255
R21168 VDD.n7454 VDD.n7453 23.1255
R21169 VDD.n7449 VDD.n7448 23.1255
R21170 VDD.n7450 VDD.n7449 23.1255
R21171 VDD.n7446 VDD.n7445 23.1255
R21172 VDD.n7445 VDD.n7444 23.1255
R21173 VDD.n7339 VDD.n7335 23.1255
R21174 VDD.n7443 VDD.n7335 23.1255
R21175 VDD.n7437 VDD.n7346 23.1255
R21176 VDD.n7437 VDD.n7436 23.1255
R21177 VDD.n7351 VDD.n7347 23.1255
R21178 VDD.n7433 VDD.n7347 23.1255
R21179 VDD.n7427 VDD.n7359 23.1255
R21180 VDD.n7427 VDD.n7426 23.1255
R21181 VDD.n7364 VDD.n7360 23.1255
R21182 VDD.n7423 VDD.n7360 23.1255
R21183 VDD.n7417 VDD.n7370 23.1255
R21184 VDD.n7417 VDD.n7416 23.1255
R21185 VDD.n7375 VDD.n7371 23.1255
R21186 VDD.n7413 VDD.n7371 23.1255
R21187 VDD.n7407 VDD.n7380 23.1255
R21188 VDD.n7407 VDD.n7406 23.1255
R21189 VDD.n7385 VDD.n7381 23.1255
R21190 VDD.n7403 VDD.n7381 23.1255
R21191 VDD.n7397 VDD.n7393 23.1255
R21192 VDD.n7397 VDD.n7396 23.1255
R21193 VDD.n7509 VDD.n7508 23.1255
R21194 VDD.n7510 VDD.n7509 23.1255
R21195 VDD.n7502 VDD.n7501 23.1255
R21196 VDD.n7503 VDD.n7502 23.1255
R21197 VDD.n7499 VDD.n7498 23.1255
R21198 VDD.n7500 VDD.n7499 23.1255
R21199 VDD.n7492 VDD.n7491 23.1255
R21200 VDD.n7493 VDD.n7492 23.1255
R21201 VDD.n7489 VDD.n7488 23.1255
R21202 VDD.n7490 VDD.n7489 23.1255
R21203 VDD.n7482 VDD.n7481 23.1255
R21204 VDD.n7483 VDD.n7482 23.1255
R21205 VDD.n7479 VDD.n7478 23.1255
R21206 VDD.n7480 VDD.n7479 23.1255
R21207 VDD.n7472 VDD.n7471 23.1255
R21208 VDD.n7473 VDD.n7472 23.1255
R21209 VDD.n7469 VDD.n7468 23.1255
R21210 VDD.n7470 VDD.n7469 23.1255
R21211 VDD.n7462 VDD.n7461 23.1255
R21212 VDD.n7463 VDD.n7462 23.1255
R21213 VDD.n7459 VDD.n7458 23.1255
R21214 VDD.n7460 VDD.n7459 23.1255
R21215 VDD.n7452 VDD.n7451 23.1255
R21216 VDD.n7453 VDD.n7452 23.1255
R21217 VDD.n7442 VDD.n7441 23.1255
R21218 VDD.n7443 VDD.n7442 23.1255
R21219 VDD.n7435 VDD.n7434 23.1255
R21220 VDD.n7436 VDD.n7435 23.1255
R21221 VDD.n7432 VDD.n7431 23.1255
R21222 VDD.n7433 VDD.n7432 23.1255
R21223 VDD.n7425 VDD.n7424 23.1255
R21224 VDD.n7426 VDD.n7425 23.1255
R21225 VDD.n7422 VDD.n7421 23.1255
R21226 VDD.n7423 VDD.n7422 23.1255
R21227 VDD.n7415 VDD.n7414 23.1255
R21228 VDD.n7416 VDD.n7415 23.1255
R21229 VDD.n7412 VDD.n7411 23.1255
R21230 VDD.n7413 VDD.n7412 23.1255
R21231 VDD.n7405 VDD.n7404 23.1255
R21232 VDD.n7406 VDD.n7405 23.1255
R21233 VDD.n7402 VDD.n7401 23.1255
R21234 VDD.n7403 VDD.n7402 23.1255
R21235 VDD.n7395 VDD.n7394 23.1255
R21236 VDD.n7396 VDD.n7395 23.1255
R21237 VDD.n7513 VDD.n7512 23.1255
R21238 VDD.n7512 VDD.n7511 23.1255
R21239 VDD.n7262 VDD.n7258 23.1255
R21240 VDD.n1912 VDD.n1908 23.1255
R21241 VDD.n7250 VDD.n1908 23.1255
R21242 VDD.n7244 VDD.n1918 23.1255
R21243 VDD.n7244 VDD.n7243 23.1255
R21244 VDD.n1923 VDD.n1919 23.1255
R21245 VDD.n7240 VDD.n1919 23.1255
R21246 VDD.n7234 VDD.n1928 23.1255
R21247 VDD.n7234 VDD.n7233 23.1255
R21248 VDD.n1933 VDD.n1929 23.1255
R21249 VDD.n7230 VDD.n1929 23.1255
R21250 VDD.n7224 VDD.n1941 23.1255
R21251 VDD.n7224 VDD.n7223 23.1255
R21252 VDD.n1946 VDD.n1942 23.1255
R21253 VDD.n7220 VDD.n1942 23.1255
R21254 VDD.n7214 VDD.n1953 23.1255
R21255 VDD.n7214 VDD.n7213 23.1255
R21256 VDD.n1958 VDD.n1954 23.1255
R21257 VDD.n7210 VDD.n1954 23.1255
R21258 VDD.n1972 VDD.n1971 23.1255
R21259 VDD.n1975 VDD.n1972 23.1255
R21260 VDD.n1977 VDD.n1967 23.1255
R21261 VDD.n1976 VDD.n1967 23.1255
R21262 VDD.n1978 VDD.n1968 23.1255
R21263 VDD.n7194 VDD.n1968 23.1255
R21264 VDD.n7192 VDD.n7191 23.1255
R21265 VDD.n7193 VDD.n7192 23.1255
R21266 VDD.n7189 VDD.n7188 23.1255
R21267 VDD.n7188 VDD.n7187 23.1255
R21268 VDD.n1988 VDD.n1984 23.1255
R21269 VDD.n7186 VDD.n1984 23.1255
R21270 VDD.n7180 VDD.n1995 23.1255
R21271 VDD.n7180 VDD.n7179 23.1255
R21272 VDD.n2000 VDD.n1996 23.1255
R21273 VDD.n7176 VDD.n1996 23.1255
R21274 VDD.n7170 VDD.n2008 23.1255
R21275 VDD.n7170 VDD.n7169 23.1255
R21276 VDD.n2013 VDD.n2009 23.1255
R21277 VDD.n7166 VDD.n2009 23.1255
R21278 VDD.n7160 VDD.n2019 23.1255
R21279 VDD.n7160 VDD.n7159 23.1255
R21280 VDD.n2024 VDD.n2020 23.1255
R21281 VDD.n7156 VDD.n2020 23.1255
R21282 VDD.n7150 VDD.n2029 23.1255
R21283 VDD.n7150 VDD.n7149 23.1255
R21284 VDD.n2034 VDD.n2030 23.1255
R21285 VDD.n7146 VDD.n2030 23.1255
R21286 VDD.n7140 VDD.n7136 23.1255
R21287 VDD.n7140 VDD.n7139 23.1255
R21288 VDD.n1906 VDD.n1902 23.1255
R21289 VDD.n7253 VDD.n7252 23.1255
R21290 VDD.n7252 VDD.n7251 23.1255
R21291 VDD.n7249 VDD.n7248 23.1255
R21292 VDD.n7250 VDD.n7249 23.1255
R21293 VDD.n7242 VDD.n7241 23.1255
R21294 VDD.n7243 VDD.n7242 23.1255
R21295 VDD.n7239 VDD.n7238 23.1255
R21296 VDD.n7240 VDD.n7239 23.1255
R21297 VDD.n7232 VDD.n7231 23.1255
R21298 VDD.n7233 VDD.n7232 23.1255
R21299 VDD.n7229 VDD.n7228 23.1255
R21300 VDD.n7230 VDD.n7229 23.1255
R21301 VDD.n7222 VDD.n7221 23.1255
R21302 VDD.n7223 VDD.n7222 23.1255
R21303 VDD.n7219 VDD.n7218 23.1255
R21304 VDD.n7220 VDD.n7219 23.1255
R21305 VDD.n7212 VDD.n7211 23.1255
R21306 VDD.n7213 VDD.n7212 23.1255
R21307 VDD.n7197 VDD.n7195 23.1255
R21308 VDD.n7195 VDD.n1976 23.1255
R21309 VDD.n7198 VDD.n7196 23.1255
R21310 VDD.n7196 VDD.n7194 23.1255
R21311 VDD.n7185 VDD.n7184 23.1255
R21312 VDD.n7186 VDD.n7185 23.1255
R21313 VDD.n7178 VDD.n7177 23.1255
R21314 VDD.n7179 VDD.n7178 23.1255
R21315 VDD.n7175 VDD.n7174 23.1255
R21316 VDD.n7176 VDD.n7175 23.1255
R21317 VDD.n7168 VDD.n7167 23.1255
R21318 VDD.n7169 VDD.n7168 23.1255
R21319 VDD.n7165 VDD.n7164 23.1255
R21320 VDD.n7166 VDD.n7165 23.1255
R21321 VDD.n7158 VDD.n7157 23.1255
R21322 VDD.n7159 VDD.n7158 23.1255
R21323 VDD.n7155 VDD.n7154 23.1255
R21324 VDD.n7156 VDD.n7155 23.1255
R21325 VDD.n7148 VDD.n7147 23.1255
R21326 VDD.n7149 VDD.n7148 23.1255
R21327 VDD.n7145 VDD.n7144 23.1255
R21328 VDD.n7146 VDD.n7145 23.1255
R21329 VDD.n7138 VDD.n7137 23.1255
R21330 VDD.n7139 VDD.n7138 23.1255
R21331 VDD.n1974 VDD.n1973 23.1255
R21332 VDD.n1975 VDD.n1974 23.1255
R21333 VDD.n7209 VDD.n7208 23.1255
R21334 VDD.n7210 VDD.n7209 23.1255
R21335 VDD.n7001 VDD.n7000 23.1255
R21336 VDD.n7002 VDD.n7001 23.1255
R21337 VDD.n6998 VDD.n6997 23.1255
R21338 VDD.n7005 VDD.n7004 23.1255
R21339 VDD.n7004 VDD.n7003 23.1255
R21340 VDD.n6990 VDD.n6986 23.1255
R21341 VDD.n7022 VDD.n7021 23.1255
R21342 VDD.n7023 VDD.n7022 23.1255
R21343 VDD.n7019 VDD.n7018 23.1255
R21344 VDD.n7018 VDD.n7017 23.1255
R21345 VDD.n7015 VDD.n7014 23.1255
R21346 VDD.n7016 VDD.n7015 23.1255
R21347 VDD.n7012 VDD.n7011 23.1255
R21348 VDD.n7026 VDD.n7025 23.1255
R21349 VDD.n7025 VDD.n7024 23.1255
R21350 VDD.n6974 VDD.n6970 23.1255
R21351 VDD.n7036 VDD.n7035 23.1255
R21352 VDD.n7037 VDD.n7036 23.1255
R21353 VDD.n7033 VDD.n7032 23.1255
R21354 VDD.n7040 VDD.n7039 23.1255
R21355 VDD.n7039 VDD.n7038 23.1255
R21356 VDD.n6965 VDD.n6961 23.1255
R21357 VDD.n7057 VDD.n7056 23.1255
R21358 VDD.n7058 VDD.n7057 23.1255
R21359 VDD.n7054 VDD.n7053 23.1255
R21360 VDD.n7053 VDD.n7052 23.1255
R21361 VDD.n7050 VDD.n7049 23.1255
R21362 VDD.n7051 VDD.n7050 23.1255
R21363 VDD.n7047 VDD.n7046 23.1255
R21364 VDD.n7061 VDD.n7060 23.1255
R21365 VDD.n7060 VDD.n7059 23.1255
R21366 VDD.n6949 VDD.n6945 23.1255
R21367 VDD.n7071 VDD.n7070 23.1255
R21368 VDD.n7072 VDD.n7071 23.1255
R21369 VDD.n7068 VDD.n7067 23.1255
R21370 VDD.n7075 VDD.n7074 23.1255
R21371 VDD.n7074 VDD.n7073 23.1255
R21372 VDD.n6940 VDD.n6936 23.1255
R21373 VDD.n7092 VDD.n7091 23.1255
R21374 VDD.n7093 VDD.n7092 23.1255
R21375 VDD.n7089 VDD.n7088 23.1255
R21376 VDD.n7088 VDD.n7087 23.1255
R21377 VDD.n7085 VDD.n7084 23.1255
R21378 VDD.n7086 VDD.n7085 23.1255
R21379 VDD.n7082 VDD.n7081 23.1255
R21380 VDD.n7096 VDD.n7095 23.1255
R21381 VDD.n7095 VDD.n7094 23.1255
R21382 VDD.n6924 VDD.n6920 23.1255
R21383 VDD.n7106 VDD.n7105 23.1255
R21384 VDD.n7107 VDD.n7106 23.1255
R21385 VDD.n7103 VDD.n7102 23.1255
R21386 VDD.n7110 VDD.n7109 23.1255
R21387 VDD.n7109 VDD.n7108 23.1255
R21388 VDD.n6915 VDD.n6911 23.1255
R21389 VDD.n6893 VDD.n6891 23.1255
R21390 VDD.n6906 VDD.n6893 23.1255
R21391 VDD.n6894 VDD.n6892 23.1255
R21392 VDD.n7122 VDD.n6894 23.1255
R21393 VDD.n7120 VDD.n7119 23.1255
R21394 VDD.n7121 VDD.n7120 23.1255
R21395 VDD.n7117 VDD.n7116 23.1255
R21396 VDD.n6904 VDD.n6903 23.1255
R21397 VDD.n6905 VDD.n6904 23.1255
R21398 VDD.n6901 VDD.n6900 23.1255
R21399 VDD.n5899 VDD.n5896 23.1255
R21400 VDD.n5898 VDD.n5896 23.1255
R21401 VDD.n5900 VDD.n5897 23.1255
R21402 VDD.n6139 VDD.n5897 23.1255
R21403 VDD.n5907 VDD.n5903 23.1255
R21404 VDD.n6138 VDD.n5903 23.1255
R21405 VDD.n6132 VDD.n5912 23.1255
R21406 VDD.n6132 VDD.n6131 23.1255
R21407 VDD.n5917 VDD.n5913 23.1255
R21408 VDD.n6128 VDD.n5913 23.1255
R21409 VDD.n6122 VDD.n5922 23.1255
R21410 VDD.n6122 VDD.n6121 23.1255
R21411 VDD.n5927 VDD.n5923 23.1255
R21412 VDD.n6118 VDD.n5923 23.1255
R21413 VDD.n6112 VDD.n5933 23.1255
R21414 VDD.n6112 VDD.n6111 23.1255
R21415 VDD.n5938 VDD.n5934 23.1255
R21416 VDD.n6108 VDD.n5934 23.1255
R21417 VDD.n6102 VDD.n5946 23.1255
R21418 VDD.n6102 VDD.n6101 23.1255
R21419 VDD.n6097 VDD.n6096 23.1255
R21420 VDD.n6098 VDD.n6097 23.1255
R21421 VDD.n6094 VDD.n6093 23.1255
R21422 VDD.n6093 VDD.n6092 23.1255
R21423 VDD.n5954 VDD.n5950 23.1255
R21424 VDD.n6091 VDD.n5950 23.1255
R21425 VDD.n6085 VDD.n5961 23.1255
R21426 VDD.n6085 VDD.n6084 23.1255
R21427 VDD.n5966 VDD.n5962 23.1255
R21428 VDD.n6081 VDD.n5962 23.1255
R21429 VDD.n6075 VDD.n5974 23.1255
R21430 VDD.n6075 VDD.n6074 23.1255
R21431 VDD.n5979 VDD.n5975 23.1255
R21432 VDD.n6071 VDD.n5975 23.1255
R21433 VDD.n6065 VDD.n5984 23.1255
R21434 VDD.n6065 VDD.n6064 23.1255
R21435 VDD.n5989 VDD.n5985 23.1255
R21436 VDD.n6061 VDD.n5985 23.1255
R21437 VDD.n6055 VDD.n5995 23.1255
R21438 VDD.n6055 VDD.n6054 23.1255
R21439 VDD.n6000 VDD.n5996 23.1255
R21440 VDD.n6051 VDD.n5996 23.1255
R21441 VDD.n6045 VDD.n6008 23.1255
R21442 VDD.n6045 VDD.n6044 23.1255
R21443 VDD.n6013 VDD.n6009 23.1255
R21444 VDD.n6041 VDD.n6009 23.1255
R21445 VDD.n6035 VDD.n6018 23.1255
R21446 VDD.n6035 VDD.n6034 23.1255
R21447 VDD.n6137 VDD.n6136 23.1255
R21448 VDD.n6138 VDD.n6137 23.1255
R21449 VDD.n6130 VDD.n6129 23.1255
R21450 VDD.n6131 VDD.n6130 23.1255
R21451 VDD.n6127 VDD.n6126 23.1255
R21452 VDD.n6128 VDD.n6127 23.1255
R21453 VDD.n6120 VDD.n6119 23.1255
R21454 VDD.n6121 VDD.n6120 23.1255
R21455 VDD.n6117 VDD.n6116 23.1255
R21456 VDD.n6118 VDD.n6117 23.1255
R21457 VDD.n6110 VDD.n6109 23.1255
R21458 VDD.n6111 VDD.n6110 23.1255
R21459 VDD.n6107 VDD.n6106 23.1255
R21460 VDD.n6108 VDD.n6107 23.1255
R21461 VDD.n6100 VDD.n6099 23.1255
R21462 VDD.n6101 VDD.n6100 23.1255
R21463 VDD.n6090 VDD.n6089 23.1255
R21464 VDD.n6091 VDD.n6090 23.1255
R21465 VDD.n6083 VDD.n6082 23.1255
R21466 VDD.n6084 VDD.n6083 23.1255
R21467 VDD.n6080 VDD.n6079 23.1255
R21468 VDD.n6081 VDD.n6080 23.1255
R21469 VDD.n6073 VDD.n6072 23.1255
R21470 VDD.n6074 VDD.n6073 23.1255
R21471 VDD.n6070 VDD.n6069 23.1255
R21472 VDD.n6071 VDD.n6070 23.1255
R21473 VDD.n6063 VDD.n6062 23.1255
R21474 VDD.n6064 VDD.n6063 23.1255
R21475 VDD.n6060 VDD.n6059 23.1255
R21476 VDD.n6061 VDD.n6060 23.1255
R21477 VDD.n6053 VDD.n6052 23.1255
R21478 VDD.n6054 VDD.n6053 23.1255
R21479 VDD.n6050 VDD.n6049 23.1255
R21480 VDD.n6051 VDD.n6050 23.1255
R21481 VDD.n6043 VDD.n6042 23.1255
R21482 VDD.n6044 VDD.n6043 23.1255
R21483 VDD.n6040 VDD.n6039 23.1255
R21484 VDD.n6041 VDD.n6040 23.1255
R21485 VDD.n6033 VDD.n6032 23.1255
R21486 VDD.n6034 VDD.n6033 23.1255
R21487 VDD.n6030 VDD.n6029 23.1255
R21488 VDD.n6031 VDD.n6030 23.1255
R21489 VDD.n6024 VDD.n6023 23.1255
R21490 VDD.n6143 VDD.n6141 23.1255
R21491 VDD.n6141 VDD.n6139 23.1255
R21492 VDD.n6142 VDD.n6140 23.1255
R21493 VDD.n6140 VDD.n5898 23.1255
R21494 VDD.n5763 VDD.n5760 23.1255
R21495 VDD.n5762 VDD.n5760 23.1255
R21496 VDD.n5764 VDD.n5761 23.1255
R21497 VDD.n6262 VDD.n5761 23.1255
R21498 VDD.n5771 VDD.n5767 23.1255
R21499 VDD.n6261 VDD.n5767 23.1255
R21500 VDD.n6255 VDD.n5776 23.1255
R21501 VDD.n6255 VDD.n6254 23.1255
R21502 VDD.n5781 VDD.n5777 23.1255
R21503 VDD.n6251 VDD.n5777 23.1255
R21504 VDD.n6245 VDD.n5786 23.1255
R21505 VDD.n6245 VDD.n6244 23.1255
R21506 VDD.n5791 VDD.n5787 23.1255
R21507 VDD.n6241 VDD.n5787 23.1255
R21508 VDD.n6235 VDD.n5797 23.1255
R21509 VDD.n6235 VDD.n6234 23.1255
R21510 VDD.n5802 VDD.n5798 23.1255
R21511 VDD.n6231 VDD.n5798 23.1255
R21512 VDD.n6225 VDD.n5810 23.1255
R21513 VDD.n6225 VDD.n6224 23.1255
R21514 VDD.n6220 VDD.n6219 23.1255
R21515 VDD.n6221 VDD.n6220 23.1255
R21516 VDD.n6217 VDD.n6216 23.1255
R21517 VDD.n6216 VDD.n6215 23.1255
R21518 VDD.n5818 VDD.n5814 23.1255
R21519 VDD.n6214 VDD.n5814 23.1255
R21520 VDD.n6208 VDD.n5825 23.1255
R21521 VDD.n6208 VDD.n6207 23.1255
R21522 VDD.n5830 VDD.n5826 23.1255
R21523 VDD.n6204 VDD.n5826 23.1255
R21524 VDD.n6198 VDD.n5838 23.1255
R21525 VDD.n6198 VDD.n6197 23.1255
R21526 VDD.n5843 VDD.n5839 23.1255
R21527 VDD.n6194 VDD.n5839 23.1255
R21528 VDD.n6188 VDD.n5848 23.1255
R21529 VDD.n6188 VDD.n6187 23.1255
R21530 VDD.n5853 VDD.n5849 23.1255
R21531 VDD.n6184 VDD.n5849 23.1255
R21532 VDD.n6178 VDD.n5859 23.1255
R21533 VDD.n6178 VDD.n6177 23.1255
R21534 VDD.n5864 VDD.n5860 23.1255
R21535 VDD.n6174 VDD.n5860 23.1255
R21536 VDD.n6168 VDD.n5872 23.1255
R21537 VDD.n6168 VDD.n6167 23.1255
R21538 VDD.n5877 VDD.n5873 23.1255
R21539 VDD.n6164 VDD.n5873 23.1255
R21540 VDD.n6158 VDD.n5882 23.1255
R21541 VDD.n6158 VDD.n6157 23.1255
R21542 VDD.n6260 VDD.n6259 23.1255
R21543 VDD.n6261 VDD.n6260 23.1255
R21544 VDD.n6253 VDD.n6252 23.1255
R21545 VDD.n6254 VDD.n6253 23.1255
R21546 VDD.n6250 VDD.n6249 23.1255
R21547 VDD.n6251 VDD.n6250 23.1255
R21548 VDD.n6243 VDD.n6242 23.1255
R21549 VDD.n6244 VDD.n6243 23.1255
R21550 VDD.n6240 VDD.n6239 23.1255
R21551 VDD.n6241 VDD.n6240 23.1255
R21552 VDD.n6233 VDD.n6232 23.1255
R21553 VDD.n6234 VDD.n6233 23.1255
R21554 VDD.n6230 VDD.n6229 23.1255
R21555 VDD.n6231 VDD.n6230 23.1255
R21556 VDD.n6223 VDD.n6222 23.1255
R21557 VDD.n6224 VDD.n6223 23.1255
R21558 VDD.n6213 VDD.n6212 23.1255
R21559 VDD.n6214 VDD.n6213 23.1255
R21560 VDD.n6206 VDD.n6205 23.1255
R21561 VDD.n6207 VDD.n6206 23.1255
R21562 VDD.n6203 VDD.n6202 23.1255
R21563 VDD.n6204 VDD.n6203 23.1255
R21564 VDD.n6196 VDD.n6195 23.1255
R21565 VDD.n6197 VDD.n6196 23.1255
R21566 VDD.n6193 VDD.n6192 23.1255
R21567 VDD.n6194 VDD.n6193 23.1255
R21568 VDD.n6186 VDD.n6185 23.1255
R21569 VDD.n6187 VDD.n6186 23.1255
R21570 VDD.n6183 VDD.n6182 23.1255
R21571 VDD.n6184 VDD.n6183 23.1255
R21572 VDD.n6176 VDD.n6175 23.1255
R21573 VDD.n6177 VDD.n6176 23.1255
R21574 VDD.n6173 VDD.n6172 23.1255
R21575 VDD.n6174 VDD.n6173 23.1255
R21576 VDD.n6166 VDD.n6165 23.1255
R21577 VDD.n6167 VDD.n6166 23.1255
R21578 VDD.n6163 VDD.n6162 23.1255
R21579 VDD.n6164 VDD.n6163 23.1255
R21580 VDD.n6156 VDD.n6155 23.1255
R21581 VDD.n6157 VDD.n6156 23.1255
R21582 VDD.n6153 VDD.n6152 23.1255
R21583 VDD.n6154 VDD.n6153 23.1255
R21584 VDD.n5888 VDD.n5887 23.1255
R21585 VDD.n6266 VDD.n6264 23.1255
R21586 VDD.n6264 VDD.n6262 23.1255
R21587 VDD.n6265 VDD.n6263 23.1255
R21588 VDD.n6263 VDD.n5762 23.1255
R21589 VDD.n5627 VDD.n5624 23.1255
R21590 VDD.n5626 VDD.n5624 23.1255
R21591 VDD.n5628 VDD.n5625 23.1255
R21592 VDD.n6385 VDD.n5625 23.1255
R21593 VDD.n5635 VDD.n5631 23.1255
R21594 VDD.n6384 VDD.n5631 23.1255
R21595 VDD.n6378 VDD.n5640 23.1255
R21596 VDD.n6378 VDD.n6377 23.1255
R21597 VDD.n5645 VDD.n5641 23.1255
R21598 VDD.n6374 VDD.n5641 23.1255
R21599 VDD.n6368 VDD.n5650 23.1255
R21600 VDD.n6368 VDD.n6367 23.1255
R21601 VDD.n5655 VDD.n5651 23.1255
R21602 VDD.n6364 VDD.n5651 23.1255
R21603 VDD.n6358 VDD.n5661 23.1255
R21604 VDD.n6358 VDD.n6357 23.1255
R21605 VDD.n5666 VDD.n5662 23.1255
R21606 VDD.n6354 VDD.n5662 23.1255
R21607 VDD.n6348 VDD.n5674 23.1255
R21608 VDD.n6348 VDD.n6347 23.1255
R21609 VDD.n6343 VDD.n6342 23.1255
R21610 VDD.n6344 VDD.n6343 23.1255
R21611 VDD.n6340 VDD.n6339 23.1255
R21612 VDD.n6339 VDD.n6338 23.1255
R21613 VDD.n5682 VDD.n5678 23.1255
R21614 VDD.n6337 VDD.n5678 23.1255
R21615 VDD.n6331 VDD.n5689 23.1255
R21616 VDD.n6331 VDD.n6330 23.1255
R21617 VDD.n5694 VDD.n5690 23.1255
R21618 VDD.n6327 VDD.n5690 23.1255
R21619 VDD.n6321 VDD.n5702 23.1255
R21620 VDD.n6321 VDD.n6320 23.1255
R21621 VDD.n5707 VDD.n5703 23.1255
R21622 VDD.n6317 VDD.n5703 23.1255
R21623 VDD.n6311 VDD.n5712 23.1255
R21624 VDD.n6311 VDD.n6310 23.1255
R21625 VDD.n5717 VDD.n5713 23.1255
R21626 VDD.n6307 VDD.n5713 23.1255
R21627 VDD.n6301 VDD.n5723 23.1255
R21628 VDD.n6301 VDD.n6300 23.1255
R21629 VDD.n5728 VDD.n5724 23.1255
R21630 VDD.n6297 VDD.n5724 23.1255
R21631 VDD.n6291 VDD.n5736 23.1255
R21632 VDD.n6291 VDD.n6290 23.1255
R21633 VDD.n5741 VDD.n5737 23.1255
R21634 VDD.n6287 VDD.n5737 23.1255
R21635 VDD.n6281 VDD.n5746 23.1255
R21636 VDD.n6281 VDD.n6280 23.1255
R21637 VDD.n6383 VDD.n6382 23.1255
R21638 VDD.n6384 VDD.n6383 23.1255
R21639 VDD.n6376 VDD.n6375 23.1255
R21640 VDD.n6377 VDD.n6376 23.1255
R21641 VDD.n6373 VDD.n6372 23.1255
R21642 VDD.n6374 VDD.n6373 23.1255
R21643 VDD.n6366 VDD.n6365 23.1255
R21644 VDD.n6367 VDD.n6366 23.1255
R21645 VDD.n6363 VDD.n6362 23.1255
R21646 VDD.n6364 VDD.n6363 23.1255
R21647 VDD.n6356 VDD.n6355 23.1255
R21648 VDD.n6357 VDD.n6356 23.1255
R21649 VDD.n6353 VDD.n6352 23.1255
R21650 VDD.n6354 VDD.n6353 23.1255
R21651 VDD.n6346 VDD.n6345 23.1255
R21652 VDD.n6347 VDD.n6346 23.1255
R21653 VDD.n6336 VDD.n6335 23.1255
R21654 VDD.n6337 VDD.n6336 23.1255
R21655 VDD.n6329 VDD.n6328 23.1255
R21656 VDD.n6330 VDD.n6329 23.1255
R21657 VDD.n6326 VDD.n6325 23.1255
R21658 VDD.n6327 VDD.n6326 23.1255
R21659 VDD.n6319 VDD.n6318 23.1255
R21660 VDD.n6320 VDD.n6319 23.1255
R21661 VDD.n6316 VDD.n6315 23.1255
R21662 VDD.n6317 VDD.n6316 23.1255
R21663 VDD.n6309 VDD.n6308 23.1255
R21664 VDD.n6310 VDD.n6309 23.1255
R21665 VDD.n6306 VDD.n6305 23.1255
R21666 VDD.n6307 VDD.n6306 23.1255
R21667 VDD.n6299 VDD.n6298 23.1255
R21668 VDD.n6300 VDD.n6299 23.1255
R21669 VDD.n6296 VDD.n6295 23.1255
R21670 VDD.n6297 VDD.n6296 23.1255
R21671 VDD.n6289 VDD.n6288 23.1255
R21672 VDD.n6290 VDD.n6289 23.1255
R21673 VDD.n6286 VDD.n6285 23.1255
R21674 VDD.n6287 VDD.n6286 23.1255
R21675 VDD.n6279 VDD.n6278 23.1255
R21676 VDD.n6280 VDD.n6279 23.1255
R21677 VDD.n6276 VDD.n6275 23.1255
R21678 VDD.n6277 VDD.n6276 23.1255
R21679 VDD.n5752 VDD.n5751 23.1255
R21680 VDD.n6389 VDD.n6387 23.1255
R21681 VDD.n6387 VDD.n6385 23.1255
R21682 VDD.n6388 VDD.n6386 23.1255
R21683 VDD.n6386 VDD.n5626 23.1255
R21684 VDD.n5491 VDD.n5488 23.1255
R21685 VDD.n5490 VDD.n5488 23.1255
R21686 VDD.n5492 VDD.n5489 23.1255
R21687 VDD.n6508 VDD.n5489 23.1255
R21688 VDD.n5499 VDD.n5495 23.1255
R21689 VDD.n6507 VDD.n5495 23.1255
R21690 VDD.n6501 VDD.n5504 23.1255
R21691 VDD.n6501 VDD.n6500 23.1255
R21692 VDD.n5509 VDD.n5505 23.1255
R21693 VDD.n6497 VDD.n5505 23.1255
R21694 VDD.n6491 VDD.n5514 23.1255
R21695 VDD.n6491 VDD.n6490 23.1255
R21696 VDD.n5519 VDD.n5515 23.1255
R21697 VDD.n6487 VDD.n5515 23.1255
R21698 VDD.n6481 VDD.n5525 23.1255
R21699 VDD.n6481 VDD.n6480 23.1255
R21700 VDD.n5530 VDD.n5526 23.1255
R21701 VDD.n6477 VDD.n5526 23.1255
R21702 VDD.n6471 VDD.n5538 23.1255
R21703 VDD.n6471 VDD.n6470 23.1255
R21704 VDD.n6466 VDD.n6465 23.1255
R21705 VDD.n6467 VDD.n6466 23.1255
R21706 VDD.n6463 VDD.n6462 23.1255
R21707 VDD.n6462 VDD.n6461 23.1255
R21708 VDD.n5546 VDD.n5542 23.1255
R21709 VDD.n6460 VDD.n5542 23.1255
R21710 VDD.n6454 VDD.n5553 23.1255
R21711 VDD.n6454 VDD.n6453 23.1255
R21712 VDD.n5558 VDD.n5554 23.1255
R21713 VDD.n6450 VDD.n5554 23.1255
R21714 VDD.n6444 VDD.n5566 23.1255
R21715 VDD.n6444 VDD.n6443 23.1255
R21716 VDD.n5571 VDD.n5567 23.1255
R21717 VDD.n6440 VDD.n5567 23.1255
R21718 VDD.n6434 VDD.n5576 23.1255
R21719 VDD.n6434 VDD.n6433 23.1255
R21720 VDD.n5581 VDD.n5577 23.1255
R21721 VDD.n6430 VDD.n5577 23.1255
R21722 VDD.n6424 VDD.n5587 23.1255
R21723 VDD.n6424 VDD.n6423 23.1255
R21724 VDD.n5592 VDD.n5588 23.1255
R21725 VDD.n6420 VDD.n5588 23.1255
R21726 VDD.n6414 VDD.n5600 23.1255
R21727 VDD.n6414 VDD.n6413 23.1255
R21728 VDD.n5605 VDD.n5601 23.1255
R21729 VDD.n6410 VDD.n5601 23.1255
R21730 VDD.n6404 VDD.n5610 23.1255
R21731 VDD.n6404 VDD.n6403 23.1255
R21732 VDD.n6506 VDD.n6505 23.1255
R21733 VDD.n6507 VDD.n6506 23.1255
R21734 VDD.n6499 VDD.n6498 23.1255
R21735 VDD.n6500 VDD.n6499 23.1255
R21736 VDD.n6496 VDD.n6495 23.1255
R21737 VDD.n6497 VDD.n6496 23.1255
R21738 VDD.n6489 VDD.n6488 23.1255
R21739 VDD.n6490 VDD.n6489 23.1255
R21740 VDD.n6486 VDD.n6485 23.1255
R21741 VDD.n6487 VDD.n6486 23.1255
R21742 VDD.n6479 VDD.n6478 23.1255
R21743 VDD.n6480 VDD.n6479 23.1255
R21744 VDD.n6476 VDD.n6475 23.1255
R21745 VDD.n6477 VDD.n6476 23.1255
R21746 VDD.n6469 VDD.n6468 23.1255
R21747 VDD.n6470 VDD.n6469 23.1255
R21748 VDD.n6459 VDD.n6458 23.1255
R21749 VDD.n6460 VDD.n6459 23.1255
R21750 VDD.n6452 VDD.n6451 23.1255
R21751 VDD.n6453 VDD.n6452 23.1255
R21752 VDD.n6449 VDD.n6448 23.1255
R21753 VDD.n6450 VDD.n6449 23.1255
R21754 VDD.n6442 VDD.n6441 23.1255
R21755 VDD.n6443 VDD.n6442 23.1255
R21756 VDD.n6439 VDD.n6438 23.1255
R21757 VDD.n6440 VDD.n6439 23.1255
R21758 VDD.n6432 VDD.n6431 23.1255
R21759 VDD.n6433 VDD.n6432 23.1255
R21760 VDD.n6429 VDD.n6428 23.1255
R21761 VDD.n6430 VDD.n6429 23.1255
R21762 VDD.n6422 VDD.n6421 23.1255
R21763 VDD.n6423 VDD.n6422 23.1255
R21764 VDD.n6419 VDD.n6418 23.1255
R21765 VDD.n6420 VDD.n6419 23.1255
R21766 VDD.n6412 VDD.n6411 23.1255
R21767 VDD.n6413 VDD.n6412 23.1255
R21768 VDD.n6409 VDD.n6408 23.1255
R21769 VDD.n6410 VDD.n6409 23.1255
R21770 VDD.n6402 VDD.n6401 23.1255
R21771 VDD.n6403 VDD.n6402 23.1255
R21772 VDD.n6399 VDD.n6398 23.1255
R21773 VDD.n6400 VDD.n6399 23.1255
R21774 VDD.n5616 VDD.n5615 23.1255
R21775 VDD.n6512 VDD.n6510 23.1255
R21776 VDD.n6510 VDD.n6508 23.1255
R21777 VDD.n6511 VDD.n6509 23.1255
R21778 VDD.n6509 VDD.n5490 23.1255
R21779 VDD.n5355 VDD.n5352 23.1255
R21780 VDD.n5354 VDD.n5352 23.1255
R21781 VDD.n5356 VDD.n5353 23.1255
R21782 VDD.n6631 VDD.n5353 23.1255
R21783 VDD.n5363 VDD.n5359 23.1255
R21784 VDD.n6630 VDD.n5359 23.1255
R21785 VDD.n6624 VDD.n5368 23.1255
R21786 VDD.n6624 VDD.n6623 23.1255
R21787 VDD.n5373 VDD.n5369 23.1255
R21788 VDD.n6620 VDD.n5369 23.1255
R21789 VDD.n6614 VDD.n5378 23.1255
R21790 VDD.n6614 VDD.n6613 23.1255
R21791 VDD.n5383 VDD.n5379 23.1255
R21792 VDD.n6610 VDD.n5379 23.1255
R21793 VDD.n6604 VDD.n5389 23.1255
R21794 VDD.n6604 VDD.n6603 23.1255
R21795 VDD.n5394 VDD.n5390 23.1255
R21796 VDD.n6600 VDD.n5390 23.1255
R21797 VDD.n6594 VDD.n5402 23.1255
R21798 VDD.n6594 VDD.n6593 23.1255
R21799 VDD.n6589 VDD.n6588 23.1255
R21800 VDD.n6590 VDD.n6589 23.1255
R21801 VDD.n6586 VDD.n6585 23.1255
R21802 VDD.n6585 VDD.n6584 23.1255
R21803 VDD.n5410 VDD.n5406 23.1255
R21804 VDD.n6583 VDD.n5406 23.1255
R21805 VDD.n6577 VDD.n5417 23.1255
R21806 VDD.n6577 VDD.n6576 23.1255
R21807 VDD.n5422 VDD.n5418 23.1255
R21808 VDD.n6573 VDD.n5418 23.1255
R21809 VDD.n6567 VDD.n5430 23.1255
R21810 VDD.n6567 VDD.n6566 23.1255
R21811 VDD.n5435 VDD.n5431 23.1255
R21812 VDD.n6563 VDD.n5431 23.1255
R21813 VDD.n6557 VDD.n5440 23.1255
R21814 VDD.n6557 VDD.n6556 23.1255
R21815 VDD.n5445 VDD.n5441 23.1255
R21816 VDD.n6553 VDD.n5441 23.1255
R21817 VDD.n6547 VDD.n5451 23.1255
R21818 VDD.n6547 VDD.n6546 23.1255
R21819 VDD.n5456 VDD.n5452 23.1255
R21820 VDD.n6543 VDD.n5452 23.1255
R21821 VDD.n6537 VDD.n5464 23.1255
R21822 VDD.n6537 VDD.n6536 23.1255
R21823 VDD.n5469 VDD.n5465 23.1255
R21824 VDD.n6533 VDD.n5465 23.1255
R21825 VDD.n6527 VDD.n5474 23.1255
R21826 VDD.n6527 VDD.n6526 23.1255
R21827 VDD.n6629 VDD.n6628 23.1255
R21828 VDD.n6630 VDD.n6629 23.1255
R21829 VDD.n6622 VDD.n6621 23.1255
R21830 VDD.n6623 VDD.n6622 23.1255
R21831 VDD.n6619 VDD.n6618 23.1255
R21832 VDD.n6620 VDD.n6619 23.1255
R21833 VDD.n6612 VDD.n6611 23.1255
R21834 VDD.n6613 VDD.n6612 23.1255
R21835 VDD.n6609 VDD.n6608 23.1255
R21836 VDD.n6610 VDD.n6609 23.1255
R21837 VDD.n6602 VDD.n6601 23.1255
R21838 VDD.n6603 VDD.n6602 23.1255
R21839 VDD.n6599 VDD.n6598 23.1255
R21840 VDD.n6600 VDD.n6599 23.1255
R21841 VDD.n6592 VDD.n6591 23.1255
R21842 VDD.n6593 VDD.n6592 23.1255
R21843 VDD.n6582 VDD.n6581 23.1255
R21844 VDD.n6583 VDD.n6582 23.1255
R21845 VDD.n6575 VDD.n6574 23.1255
R21846 VDD.n6576 VDD.n6575 23.1255
R21847 VDD.n6572 VDD.n6571 23.1255
R21848 VDD.n6573 VDD.n6572 23.1255
R21849 VDD.n6565 VDD.n6564 23.1255
R21850 VDD.n6566 VDD.n6565 23.1255
R21851 VDD.n6562 VDD.n6561 23.1255
R21852 VDD.n6563 VDD.n6562 23.1255
R21853 VDD.n6555 VDD.n6554 23.1255
R21854 VDD.n6556 VDD.n6555 23.1255
R21855 VDD.n6552 VDD.n6551 23.1255
R21856 VDD.n6553 VDD.n6552 23.1255
R21857 VDD.n6545 VDD.n6544 23.1255
R21858 VDD.n6546 VDD.n6545 23.1255
R21859 VDD.n6542 VDD.n6541 23.1255
R21860 VDD.n6543 VDD.n6542 23.1255
R21861 VDD.n6535 VDD.n6534 23.1255
R21862 VDD.n6536 VDD.n6535 23.1255
R21863 VDD.n6532 VDD.n6531 23.1255
R21864 VDD.n6533 VDD.n6532 23.1255
R21865 VDD.n6525 VDD.n6524 23.1255
R21866 VDD.n6526 VDD.n6525 23.1255
R21867 VDD.n6522 VDD.n6521 23.1255
R21868 VDD.n6523 VDD.n6522 23.1255
R21869 VDD.n5480 VDD.n5479 23.1255
R21870 VDD.n6635 VDD.n6633 23.1255
R21871 VDD.n6633 VDD.n6631 23.1255
R21872 VDD.n6634 VDD.n6632 23.1255
R21873 VDD.n6632 VDD.n5354 23.1255
R21874 VDD.n5219 VDD.n5216 23.1255
R21875 VDD.n5218 VDD.n5216 23.1255
R21876 VDD.n5220 VDD.n5217 23.1255
R21877 VDD.n6754 VDD.n5217 23.1255
R21878 VDD.n5227 VDD.n5223 23.1255
R21879 VDD.n6753 VDD.n5223 23.1255
R21880 VDD.n6747 VDD.n5232 23.1255
R21881 VDD.n6747 VDD.n6746 23.1255
R21882 VDD.n5237 VDD.n5233 23.1255
R21883 VDD.n6743 VDD.n5233 23.1255
R21884 VDD.n6737 VDD.n5242 23.1255
R21885 VDD.n6737 VDD.n6736 23.1255
R21886 VDD.n5247 VDD.n5243 23.1255
R21887 VDD.n6733 VDD.n5243 23.1255
R21888 VDD.n6727 VDD.n5253 23.1255
R21889 VDD.n6727 VDD.n6726 23.1255
R21890 VDD.n5258 VDD.n5254 23.1255
R21891 VDD.n6723 VDD.n5254 23.1255
R21892 VDD.n6717 VDD.n5266 23.1255
R21893 VDD.n6717 VDD.n6716 23.1255
R21894 VDD.n6712 VDD.n6711 23.1255
R21895 VDD.n6713 VDD.n6712 23.1255
R21896 VDD.n6709 VDD.n6708 23.1255
R21897 VDD.n6708 VDD.n6707 23.1255
R21898 VDD.n5274 VDD.n5270 23.1255
R21899 VDD.n6706 VDD.n5270 23.1255
R21900 VDD.n6700 VDD.n5281 23.1255
R21901 VDD.n6700 VDD.n6699 23.1255
R21902 VDD.n5286 VDD.n5282 23.1255
R21903 VDD.n6696 VDD.n5282 23.1255
R21904 VDD.n6690 VDD.n5294 23.1255
R21905 VDD.n6690 VDD.n6689 23.1255
R21906 VDD.n5299 VDD.n5295 23.1255
R21907 VDD.n6686 VDD.n5295 23.1255
R21908 VDD.n6680 VDD.n5304 23.1255
R21909 VDD.n6680 VDD.n6679 23.1255
R21910 VDD.n5309 VDD.n5305 23.1255
R21911 VDD.n6676 VDD.n5305 23.1255
R21912 VDD.n6670 VDD.n5315 23.1255
R21913 VDD.n6670 VDD.n6669 23.1255
R21914 VDD.n5320 VDD.n5316 23.1255
R21915 VDD.n6666 VDD.n5316 23.1255
R21916 VDD.n6660 VDD.n5328 23.1255
R21917 VDD.n6660 VDD.n6659 23.1255
R21918 VDD.n5333 VDD.n5329 23.1255
R21919 VDD.n6656 VDD.n5329 23.1255
R21920 VDD.n6650 VDD.n5338 23.1255
R21921 VDD.n6650 VDD.n6649 23.1255
R21922 VDD.n6752 VDD.n6751 23.1255
R21923 VDD.n6753 VDD.n6752 23.1255
R21924 VDD.n6745 VDD.n6744 23.1255
R21925 VDD.n6746 VDD.n6745 23.1255
R21926 VDD.n6742 VDD.n6741 23.1255
R21927 VDD.n6743 VDD.n6742 23.1255
R21928 VDD.n6735 VDD.n6734 23.1255
R21929 VDD.n6736 VDD.n6735 23.1255
R21930 VDD.n6732 VDD.n6731 23.1255
R21931 VDD.n6733 VDD.n6732 23.1255
R21932 VDD.n6725 VDD.n6724 23.1255
R21933 VDD.n6726 VDD.n6725 23.1255
R21934 VDD.n6722 VDD.n6721 23.1255
R21935 VDD.n6723 VDD.n6722 23.1255
R21936 VDD.n6715 VDD.n6714 23.1255
R21937 VDD.n6716 VDD.n6715 23.1255
R21938 VDD.n6705 VDD.n6704 23.1255
R21939 VDD.n6706 VDD.n6705 23.1255
R21940 VDD.n6698 VDD.n6697 23.1255
R21941 VDD.n6699 VDD.n6698 23.1255
R21942 VDD.n6695 VDD.n6694 23.1255
R21943 VDD.n6696 VDD.n6695 23.1255
R21944 VDD.n6688 VDD.n6687 23.1255
R21945 VDD.n6689 VDD.n6688 23.1255
R21946 VDD.n6685 VDD.n6684 23.1255
R21947 VDD.n6686 VDD.n6685 23.1255
R21948 VDD.n6678 VDD.n6677 23.1255
R21949 VDD.n6679 VDD.n6678 23.1255
R21950 VDD.n6675 VDD.n6674 23.1255
R21951 VDD.n6676 VDD.n6675 23.1255
R21952 VDD.n6668 VDD.n6667 23.1255
R21953 VDD.n6669 VDD.n6668 23.1255
R21954 VDD.n6665 VDD.n6664 23.1255
R21955 VDD.n6666 VDD.n6665 23.1255
R21956 VDD.n6658 VDD.n6657 23.1255
R21957 VDD.n6659 VDD.n6658 23.1255
R21958 VDD.n6655 VDD.n6654 23.1255
R21959 VDD.n6656 VDD.n6655 23.1255
R21960 VDD.n6648 VDD.n6647 23.1255
R21961 VDD.n6649 VDD.n6648 23.1255
R21962 VDD.n6645 VDD.n6644 23.1255
R21963 VDD.n6646 VDD.n6645 23.1255
R21964 VDD.n5344 VDD.n5343 23.1255
R21965 VDD.n6758 VDD.n6756 23.1255
R21966 VDD.n6756 VDD.n6754 23.1255
R21967 VDD.n6757 VDD.n6755 23.1255
R21968 VDD.n6755 VDD.n5218 23.1255
R21969 VDD.n5083 VDD.n5080 23.1255
R21970 VDD.n5082 VDD.n5080 23.1255
R21971 VDD.n5084 VDD.n5081 23.1255
R21972 VDD.n6877 VDD.n5081 23.1255
R21973 VDD.n5091 VDD.n5087 23.1255
R21974 VDD.n6876 VDD.n5087 23.1255
R21975 VDD.n6870 VDD.n5096 23.1255
R21976 VDD.n6870 VDD.n6869 23.1255
R21977 VDD.n5101 VDD.n5097 23.1255
R21978 VDD.n6866 VDD.n5097 23.1255
R21979 VDD.n6860 VDD.n5106 23.1255
R21980 VDD.n6860 VDD.n6859 23.1255
R21981 VDD.n5111 VDD.n5107 23.1255
R21982 VDD.n6856 VDD.n5107 23.1255
R21983 VDD.n6850 VDD.n5117 23.1255
R21984 VDD.n6850 VDD.n6849 23.1255
R21985 VDD.n5122 VDD.n5118 23.1255
R21986 VDD.n6846 VDD.n5118 23.1255
R21987 VDD.n6840 VDD.n5130 23.1255
R21988 VDD.n6840 VDD.n6839 23.1255
R21989 VDD.n6835 VDD.n6834 23.1255
R21990 VDD.n6836 VDD.n6835 23.1255
R21991 VDD.n6832 VDD.n6831 23.1255
R21992 VDD.n6831 VDD.n6830 23.1255
R21993 VDD.n5138 VDD.n5134 23.1255
R21994 VDD.n6829 VDD.n5134 23.1255
R21995 VDD.n6823 VDD.n5145 23.1255
R21996 VDD.n6823 VDD.n6822 23.1255
R21997 VDD.n5150 VDD.n5146 23.1255
R21998 VDD.n6819 VDD.n5146 23.1255
R21999 VDD.n6813 VDD.n5158 23.1255
R22000 VDD.n6813 VDD.n6812 23.1255
R22001 VDD.n5163 VDD.n5159 23.1255
R22002 VDD.n6809 VDD.n5159 23.1255
R22003 VDD.n6803 VDD.n5168 23.1255
R22004 VDD.n6803 VDD.n6802 23.1255
R22005 VDD.n5173 VDD.n5169 23.1255
R22006 VDD.n6799 VDD.n5169 23.1255
R22007 VDD.n6793 VDD.n5179 23.1255
R22008 VDD.n6793 VDD.n6792 23.1255
R22009 VDD.n5184 VDD.n5180 23.1255
R22010 VDD.n6789 VDD.n5180 23.1255
R22011 VDD.n6783 VDD.n5192 23.1255
R22012 VDD.n6783 VDD.n6782 23.1255
R22013 VDD.n5197 VDD.n5193 23.1255
R22014 VDD.n6779 VDD.n5193 23.1255
R22015 VDD.n6773 VDD.n5202 23.1255
R22016 VDD.n6773 VDD.n6772 23.1255
R22017 VDD.n6875 VDD.n6874 23.1255
R22018 VDD.n6876 VDD.n6875 23.1255
R22019 VDD.n6868 VDD.n6867 23.1255
R22020 VDD.n6869 VDD.n6868 23.1255
R22021 VDD.n6865 VDD.n6864 23.1255
R22022 VDD.n6866 VDD.n6865 23.1255
R22023 VDD.n6858 VDD.n6857 23.1255
R22024 VDD.n6859 VDD.n6858 23.1255
R22025 VDD.n6855 VDD.n6854 23.1255
R22026 VDD.n6856 VDD.n6855 23.1255
R22027 VDD.n6848 VDD.n6847 23.1255
R22028 VDD.n6849 VDD.n6848 23.1255
R22029 VDD.n6845 VDD.n6844 23.1255
R22030 VDD.n6846 VDD.n6845 23.1255
R22031 VDD.n6838 VDD.n6837 23.1255
R22032 VDD.n6839 VDD.n6838 23.1255
R22033 VDD.n6828 VDD.n6827 23.1255
R22034 VDD.n6829 VDD.n6828 23.1255
R22035 VDD.n6821 VDD.n6820 23.1255
R22036 VDD.n6822 VDD.n6821 23.1255
R22037 VDD.n6818 VDD.n6817 23.1255
R22038 VDD.n6819 VDD.n6818 23.1255
R22039 VDD.n6811 VDD.n6810 23.1255
R22040 VDD.n6812 VDD.n6811 23.1255
R22041 VDD.n6808 VDD.n6807 23.1255
R22042 VDD.n6809 VDD.n6808 23.1255
R22043 VDD.n6801 VDD.n6800 23.1255
R22044 VDD.n6802 VDD.n6801 23.1255
R22045 VDD.n6798 VDD.n6797 23.1255
R22046 VDD.n6799 VDD.n6798 23.1255
R22047 VDD.n6791 VDD.n6790 23.1255
R22048 VDD.n6792 VDD.n6791 23.1255
R22049 VDD.n6788 VDD.n6787 23.1255
R22050 VDD.n6789 VDD.n6788 23.1255
R22051 VDD.n6781 VDD.n6780 23.1255
R22052 VDD.n6782 VDD.n6781 23.1255
R22053 VDD.n6778 VDD.n6777 23.1255
R22054 VDD.n6779 VDD.n6778 23.1255
R22055 VDD.n6771 VDD.n6770 23.1255
R22056 VDD.n6772 VDD.n6771 23.1255
R22057 VDD.n6768 VDD.n6767 23.1255
R22058 VDD.n6769 VDD.n6768 23.1255
R22059 VDD.n5208 VDD.n5207 23.1255
R22060 VDD.n6881 VDD.n6879 23.1255
R22061 VDD.n6879 VDD.n6877 23.1255
R22062 VDD.n6880 VDD.n6878 23.1255
R22063 VDD.n6878 VDD.n5082 23.1255
R22064 VDD.n4949 VDD.n4945 23.1255
R22065 VDD.n4949 VDD.n4948 23.1255
R22066 VDD.n4941 VDD.n4937 23.1255
R22067 VDD.n4958 VDD.n4937 23.1255
R22068 VDD.n4962 VDD.n4936 23.1255
R22069 VDD.n4962 VDD.n4961 23.1255
R22070 VDD.n4931 VDD.n4927 23.1255
R22071 VDD.n4968 VDD.n4927 23.1255
R22072 VDD.n4972 VDD.n4926 23.1255
R22073 VDD.n4972 VDD.n4971 23.1255
R22074 VDD.n4920 VDD.n4916 23.1255
R22075 VDD.n4978 VDD.n4916 23.1255
R22076 VDD.n4982 VDD.n4915 23.1255
R22077 VDD.n4982 VDD.n4981 23.1255
R22078 VDD.n4907 VDD.n4903 23.1255
R22079 VDD.n4988 VDD.n4903 23.1255
R22080 VDD.n4992 VDD.n4902 23.1255
R22081 VDD.n4992 VDD.n4991 23.1255
R22082 VDD.n4895 VDD.n4891 23.1255
R22083 VDD.n4998 VDD.n4891 23.1255
R22084 VDD.n5001 VDD.n5000 23.1255
R22085 VDD.n5000 VDD.n4999 23.1255
R22086 VDD.n5004 VDD.n5003 23.1255
R22087 VDD.n5005 VDD.n5004 23.1255
R22088 VDD.n5009 VDD.n4887 23.1255
R22089 VDD.n5009 VDD.n5008 23.1255
R22090 VDD.n4879 VDD.n4875 23.1255
R22091 VDD.n5015 VDD.n4875 23.1255
R22092 VDD.n5019 VDD.n4874 23.1255
R22093 VDD.n5019 VDD.n5018 23.1255
R22094 VDD.n4869 VDD.n4865 23.1255
R22095 VDD.n5025 VDD.n4865 23.1255
R22096 VDD.n5029 VDD.n4864 23.1255
R22097 VDD.n5029 VDD.n5028 23.1255
R22098 VDD.n4858 VDD.n4854 23.1255
R22099 VDD.n5035 VDD.n4854 23.1255
R22100 VDD.n5039 VDD.n4853 23.1255
R22101 VDD.n5039 VDD.n5038 23.1255
R22102 VDD.n4845 VDD.n4841 23.1255
R22103 VDD.n5045 VDD.n4841 23.1255
R22104 VDD.n5049 VDD.n4840 23.1255
R22105 VDD.n5049 VDD.n5048 23.1255
R22106 VDD.n4835 VDD.n4831 23.1255
R22107 VDD.n5055 VDD.n4831 23.1255
R22108 VDD.n5059 VDD.n4830 23.1255
R22109 VDD.n5059 VDD.n5058 23.1255
R22110 VDD.n4824 VDD.n4820 23.1255
R22111 VDD.n5065 VDD.n4820 23.1255
R22112 VDD.n4960 VDD.n4959 23.1255
R22113 VDD.n4961 VDD.n4960 23.1255
R22114 VDD.n4967 VDD.n4966 23.1255
R22115 VDD.n4968 VDD.n4967 23.1255
R22116 VDD.n4970 VDD.n4969 23.1255
R22117 VDD.n4971 VDD.n4970 23.1255
R22118 VDD.n4977 VDD.n4976 23.1255
R22119 VDD.n4978 VDD.n4977 23.1255
R22120 VDD.n4980 VDD.n4979 23.1255
R22121 VDD.n4981 VDD.n4980 23.1255
R22122 VDD.n4987 VDD.n4986 23.1255
R22123 VDD.n4988 VDD.n4987 23.1255
R22124 VDD.n4990 VDD.n4989 23.1255
R22125 VDD.n4991 VDD.n4990 23.1255
R22126 VDD.n4997 VDD.n4996 23.1255
R22127 VDD.n4998 VDD.n4997 23.1255
R22128 VDD.n5007 VDD.n5006 23.1255
R22129 VDD.n5008 VDD.n5007 23.1255
R22130 VDD.n5014 VDD.n5013 23.1255
R22131 VDD.n5015 VDD.n5014 23.1255
R22132 VDD.n5017 VDD.n5016 23.1255
R22133 VDD.n5018 VDD.n5017 23.1255
R22134 VDD.n5024 VDD.n5023 23.1255
R22135 VDD.n5025 VDD.n5024 23.1255
R22136 VDD.n5027 VDD.n5026 23.1255
R22137 VDD.n5028 VDD.n5027 23.1255
R22138 VDD.n5034 VDD.n5033 23.1255
R22139 VDD.n5035 VDD.n5034 23.1255
R22140 VDD.n5037 VDD.n5036 23.1255
R22141 VDD.n5038 VDD.n5037 23.1255
R22142 VDD.n5044 VDD.n5043 23.1255
R22143 VDD.n5045 VDD.n5044 23.1255
R22144 VDD.n5047 VDD.n5046 23.1255
R22145 VDD.n5048 VDD.n5047 23.1255
R22146 VDD.n5054 VDD.n5053 23.1255
R22147 VDD.n5055 VDD.n5054 23.1255
R22148 VDD.n5057 VDD.n5056 23.1255
R22149 VDD.n5058 VDD.n5057 23.1255
R22150 VDD.n5064 VDD.n5063 23.1255
R22151 VDD.n5065 VDD.n5064 23.1255
R22152 VDD.n5066 VDD.n4816 23.1255
R22153 VDD.n5067 VDD.n5066 23.1255
R22154 VDD.n5070 VDD.n5069 23.1255
R22155 VDD.n4957 VDD.n4956 23.1255
R22156 VDD.n4958 VDD.n4957 23.1255
R22157 VDD.n4947 VDD.n4946 23.1255
R22158 VDD.n4948 VDD.n4947 23.1255
R22159 VDD.n2048 VDD.n2044 23.1255
R22160 VDD.n4809 VDD.n2044 23.1255
R22161 VDD.n4803 VDD.n2054 23.1255
R22162 VDD.n4803 VDD.n4802 23.1255
R22163 VDD.n2059 VDD.n2055 23.1255
R22164 VDD.n4799 VDD.n2055 23.1255
R22165 VDD.n4793 VDD.n2064 23.1255
R22166 VDD.n4793 VDD.n4792 23.1255
R22167 VDD.n2069 VDD.n2065 23.1255
R22168 VDD.n4789 VDD.n2065 23.1255
R22169 VDD.n4783 VDD.n2077 23.1255
R22170 VDD.n4783 VDD.n4782 23.1255
R22171 VDD.n2082 VDD.n2078 23.1255
R22172 VDD.n4779 VDD.n2078 23.1255
R22173 VDD.n4773 VDD.n2089 23.1255
R22174 VDD.n4773 VDD.n4772 23.1255
R22175 VDD.n2094 VDD.n2090 23.1255
R22176 VDD.n4769 VDD.n2090 23.1255
R22177 VDD.n2108 VDD.n2107 23.1255
R22178 VDD.n2111 VDD.n2108 23.1255
R22179 VDD.n2113 VDD.n2103 23.1255
R22180 VDD.n2112 VDD.n2103 23.1255
R22181 VDD.n2114 VDD.n2104 23.1255
R22182 VDD.n4753 VDD.n2104 23.1255
R22183 VDD.n4751 VDD.n4750 23.1255
R22184 VDD.n4752 VDD.n4751 23.1255
R22185 VDD.n4748 VDD.n4747 23.1255
R22186 VDD.n4747 VDD.n4746 23.1255
R22187 VDD.n2124 VDD.n2120 23.1255
R22188 VDD.n4745 VDD.n2120 23.1255
R22189 VDD.n4739 VDD.n2131 23.1255
R22190 VDD.n4739 VDD.n4738 23.1255
R22191 VDD.n2136 VDD.n2132 23.1255
R22192 VDD.n4735 VDD.n2132 23.1255
R22193 VDD.n4729 VDD.n2144 23.1255
R22194 VDD.n4729 VDD.n4728 23.1255
R22195 VDD.n2149 VDD.n2145 23.1255
R22196 VDD.n4725 VDD.n2145 23.1255
R22197 VDD.n4719 VDD.n2155 23.1255
R22198 VDD.n4719 VDD.n4718 23.1255
R22199 VDD.n2160 VDD.n2156 23.1255
R22200 VDD.n4715 VDD.n2156 23.1255
R22201 VDD.n4709 VDD.n2165 23.1255
R22202 VDD.n4709 VDD.n4708 23.1255
R22203 VDD.n2170 VDD.n2166 23.1255
R22204 VDD.n4705 VDD.n2166 23.1255
R22205 VDD.n4699 VDD.n4695 23.1255
R22206 VDD.n4699 VDD.n4698 23.1255
R22207 VDD.n2042 VDD.n2038 23.1255
R22208 VDD.n4812 VDD.n4811 23.1255
R22209 VDD.n4811 VDD.n4810 23.1255
R22210 VDD.n4808 VDD.n4807 23.1255
R22211 VDD.n4809 VDD.n4808 23.1255
R22212 VDD.n4801 VDD.n4800 23.1255
R22213 VDD.n4802 VDD.n4801 23.1255
R22214 VDD.n4798 VDD.n4797 23.1255
R22215 VDD.n4799 VDD.n4798 23.1255
R22216 VDD.n4791 VDD.n4790 23.1255
R22217 VDD.n4792 VDD.n4791 23.1255
R22218 VDD.n4788 VDD.n4787 23.1255
R22219 VDD.n4789 VDD.n4788 23.1255
R22220 VDD.n4781 VDD.n4780 23.1255
R22221 VDD.n4782 VDD.n4781 23.1255
R22222 VDD.n4778 VDD.n4777 23.1255
R22223 VDD.n4779 VDD.n4778 23.1255
R22224 VDD.n4771 VDD.n4770 23.1255
R22225 VDD.n4772 VDD.n4771 23.1255
R22226 VDD.n4756 VDD.n4754 23.1255
R22227 VDD.n4754 VDD.n2112 23.1255
R22228 VDD.n4757 VDD.n4755 23.1255
R22229 VDD.n4755 VDD.n4753 23.1255
R22230 VDD.n4744 VDD.n4743 23.1255
R22231 VDD.n4745 VDD.n4744 23.1255
R22232 VDD.n4737 VDD.n4736 23.1255
R22233 VDD.n4738 VDD.n4737 23.1255
R22234 VDD.n4734 VDD.n4733 23.1255
R22235 VDD.n4735 VDD.n4734 23.1255
R22236 VDD.n4727 VDD.n4726 23.1255
R22237 VDD.n4728 VDD.n4727 23.1255
R22238 VDD.n4724 VDD.n4723 23.1255
R22239 VDD.n4725 VDD.n4724 23.1255
R22240 VDD.n4717 VDD.n4716 23.1255
R22241 VDD.n4718 VDD.n4717 23.1255
R22242 VDD.n4714 VDD.n4713 23.1255
R22243 VDD.n4715 VDD.n4714 23.1255
R22244 VDD.n4707 VDD.n4706 23.1255
R22245 VDD.n4708 VDD.n4707 23.1255
R22246 VDD.n4704 VDD.n4703 23.1255
R22247 VDD.n4705 VDD.n4704 23.1255
R22248 VDD.n4697 VDD.n4696 23.1255
R22249 VDD.n4698 VDD.n4697 23.1255
R22250 VDD.n2110 VDD.n2109 23.1255
R22251 VDD.n2111 VDD.n2110 23.1255
R22252 VDD.n4768 VDD.n4767 23.1255
R22253 VDD.n4769 VDD.n4768 23.1255
R22254 VDD.n2184 VDD.n2180 23.1255
R22255 VDD.n4684 VDD.n2180 23.1255
R22256 VDD.n4678 VDD.n2190 23.1255
R22257 VDD.n4678 VDD.n4677 23.1255
R22258 VDD.n2195 VDD.n2191 23.1255
R22259 VDD.n4674 VDD.n2191 23.1255
R22260 VDD.n4668 VDD.n2200 23.1255
R22261 VDD.n4668 VDD.n4667 23.1255
R22262 VDD.n2205 VDD.n2201 23.1255
R22263 VDD.n4664 VDD.n2201 23.1255
R22264 VDD.n4658 VDD.n2213 23.1255
R22265 VDD.n4658 VDD.n4657 23.1255
R22266 VDD.n2218 VDD.n2214 23.1255
R22267 VDD.n4654 VDD.n2214 23.1255
R22268 VDD.n4648 VDD.n2225 23.1255
R22269 VDD.n4648 VDD.n4647 23.1255
R22270 VDD.n2230 VDD.n2226 23.1255
R22271 VDD.n4644 VDD.n2226 23.1255
R22272 VDD.n2244 VDD.n2243 23.1255
R22273 VDD.n2247 VDD.n2244 23.1255
R22274 VDD.n2249 VDD.n2239 23.1255
R22275 VDD.n2248 VDD.n2239 23.1255
R22276 VDD.n2250 VDD.n2240 23.1255
R22277 VDD.n4628 VDD.n2240 23.1255
R22278 VDD.n4626 VDD.n4625 23.1255
R22279 VDD.n4627 VDD.n4626 23.1255
R22280 VDD.n4623 VDD.n4622 23.1255
R22281 VDD.n4622 VDD.n4621 23.1255
R22282 VDD.n2260 VDD.n2256 23.1255
R22283 VDD.n4620 VDD.n2256 23.1255
R22284 VDD.n4614 VDD.n2267 23.1255
R22285 VDD.n4614 VDD.n4613 23.1255
R22286 VDD.n2272 VDD.n2268 23.1255
R22287 VDD.n4610 VDD.n2268 23.1255
R22288 VDD.n4604 VDD.n2280 23.1255
R22289 VDD.n4604 VDD.n4603 23.1255
R22290 VDD.n2285 VDD.n2281 23.1255
R22291 VDD.n4600 VDD.n2281 23.1255
R22292 VDD.n4594 VDD.n2291 23.1255
R22293 VDD.n4594 VDD.n4593 23.1255
R22294 VDD.n2296 VDD.n2292 23.1255
R22295 VDD.n4590 VDD.n2292 23.1255
R22296 VDD.n4584 VDD.n2301 23.1255
R22297 VDD.n4584 VDD.n4583 23.1255
R22298 VDD.n2306 VDD.n2302 23.1255
R22299 VDD.n4580 VDD.n2302 23.1255
R22300 VDD.n4574 VDD.n4570 23.1255
R22301 VDD.n4574 VDD.n4573 23.1255
R22302 VDD.n2178 VDD.n2174 23.1255
R22303 VDD.n4687 VDD.n4686 23.1255
R22304 VDD.n4686 VDD.n4685 23.1255
R22305 VDD.n4683 VDD.n4682 23.1255
R22306 VDD.n4684 VDD.n4683 23.1255
R22307 VDD.n4676 VDD.n4675 23.1255
R22308 VDD.n4677 VDD.n4676 23.1255
R22309 VDD.n4673 VDD.n4672 23.1255
R22310 VDD.n4674 VDD.n4673 23.1255
R22311 VDD.n4666 VDD.n4665 23.1255
R22312 VDD.n4667 VDD.n4666 23.1255
R22313 VDD.n4663 VDD.n4662 23.1255
R22314 VDD.n4664 VDD.n4663 23.1255
R22315 VDD.n4656 VDD.n4655 23.1255
R22316 VDD.n4657 VDD.n4656 23.1255
R22317 VDD.n4653 VDD.n4652 23.1255
R22318 VDD.n4654 VDD.n4653 23.1255
R22319 VDD.n4646 VDD.n4645 23.1255
R22320 VDD.n4647 VDD.n4646 23.1255
R22321 VDD.n4631 VDD.n4629 23.1255
R22322 VDD.n4629 VDD.n2248 23.1255
R22323 VDD.n4632 VDD.n4630 23.1255
R22324 VDD.n4630 VDD.n4628 23.1255
R22325 VDD.n4619 VDD.n4618 23.1255
R22326 VDD.n4620 VDD.n4619 23.1255
R22327 VDD.n4612 VDD.n4611 23.1255
R22328 VDD.n4613 VDD.n4612 23.1255
R22329 VDD.n4609 VDD.n4608 23.1255
R22330 VDD.n4610 VDD.n4609 23.1255
R22331 VDD.n4602 VDD.n4601 23.1255
R22332 VDD.n4603 VDD.n4602 23.1255
R22333 VDD.n4599 VDD.n4598 23.1255
R22334 VDD.n4600 VDD.n4599 23.1255
R22335 VDD.n4592 VDD.n4591 23.1255
R22336 VDD.n4593 VDD.n4592 23.1255
R22337 VDD.n4589 VDD.n4588 23.1255
R22338 VDD.n4590 VDD.n4589 23.1255
R22339 VDD.n4582 VDD.n4581 23.1255
R22340 VDD.n4583 VDD.n4582 23.1255
R22341 VDD.n4579 VDD.n4578 23.1255
R22342 VDD.n4580 VDD.n4579 23.1255
R22343 VDD.n4572 VDD.n4571 23.1255
R22344 VDD.n4573 VDD.n4572 23.1255
R22345 VDD.n2246 VDD.n2245 23.1255
R22346 VDD.n2247 VDD.n2246 23.1255
R22347 VDD.n4643 VDD.n4642 23.1255
R22348 VDD.n4644 VDD.n4643 23.1255
R22349 VDD.n2320 VDD.n2316 23.1255
R22350 VDD.n4559 VDD.n2316 23.1255
R22351 VDD.n4553 VDD.n2326 23.1255
R22352 VDD.n4553 VDD.n4552 23.1255
R22353 VDD.n2331 VDD.n2327 23.1255
R22354 VDD.n4549 VDD.n2327 23.1255
R22355 VDD.n4543 VDD.n2336 23.1255
R22356 VDD.n4543 VDD.n4542 23.1255
R22357 VDD.n2341 VDD.n2337 23.1255
R22358 VDD.n4539 VDD.n2337 23.1255
R22359 VDD.n4533 VDD.n2349 23.1255
R22360 VDD.n4533 VDD.n4532 23.1255
R22361 VDD.n2354 VDD.n2350 23.1255
R22362 VDD.n4529 VDD.n2350 23.1255
R22363 VDD.n4523 VDD.n2361 23.1255
R22364 VDD.n4523 VDD.n4522 23.1255
R22365 VDD.n2366 VDD.n2362 23.1255
R22366 VDD.n4519 VDD.n2362 23.1255
R22367 VDD.n2380 VDD.n2379 23.1255
R22368 VDD.n2383 VDD.n2380 23.1255
R22369 VDD.n2385 VDD.n2375 23.1255
R22370 VDD.n2384 VDD.n2375 23.1255
R22371 VDD.n2386 VDD.n2376 23.1255
R22372 VDD.n4503 VDD.n2376 23.1255
R22373 VDD.n4501 VDD.n4500 23.1255
R22374 VDD.n4502 VDD.n4501 23.1255
R22375 VDD.n4498 VDD.n4497 23.1255
R22376 VDD.n4497 VDD.n4496 23.1255
R22377 VDD.n2396 VDD.n2392 23.1255
R22378 VDD.n4495 VDD.n2392 23.1255
R22379 VDD.n4489 VDD.n2403 23.1255
R22380 VDD.n4489 VDD.n4488 23.1255
R22381 VDD.n2408 VDD.n2404 23.1255
R22382 VDD.n4485 VDD.n2404 23.1255
R22383 VDD.n4479 VDD.n2416 23.1255
R22384 VDD.n4479 VDD.n4478 23.1255
R22385 VDD.n2421 VDD.n2417 23.1255
R22386 VDD.n4475 VDD.n2417 23.1255
R22387 VDD.n4469 VDD.n2427 23.1255
R22388 VDD.n4469 VDD.n4468 23.1255
R22389 VDD.n2432 VDD.n2428 23.1255
R22390 VDD.n4465 VDD.n2428 23.1255
R22391 VDD.n4459 VDD.n2437 23.1255
R22392 VDD.n4459 VDD.n4458 23.1255
R22393 VDD.n2442 VDD.n2438 23.1255
R22394 VDD.n4455 VDD.n2438 23.1255
R22395 VDD.n4449 VDD.n4445 23.1255
R22396 VDD.n4449 VDD.n4448 23.1255
R22397 VDD.n2314 VDD.n2310 23.1255
R22398 VDD.n4562 VDD.n4561 23.1255
R22399 VDD.n4561 VDD.n4560 23.1255
R22400 VDD.n4558 VDD.n4557 23.1255
R22401 VDD.n4559 VDD.n4558 23.1255
R22402 VDD.n4551 VDD.n4550 23.1255
R22403 VDD.n4552 VDD.n4551 23.1255
R22404 VDD.n4548 VDD.n4547 23.1255
R22405 VDD.n4549 VDD.n4548 23.1255
R22406 VDD.n4541 VDD.n4540 23.1255
R22407 VDD.n4542 VDD.n4541 23.1255
R22408 VDD.n4538 VDD.n4537 23.1255
R22409 VDD.n4539 VDD.n4538 23.1255
R22410 VDD.n4531 VDD.n4530 23.1255
R22411 VDD.n4532 VDD.n4531 23.1255
R22412 VDD.n4528 VDD.n4527 23.1255
R22413 VDD.n4529 VDD.n4528 23.1255
R22414 VDD.n4521 VDD.n4520 23.1255
R22415 VDD.n4522 VDD.n4521 23.1255
R22416 VDD.n4506 VDD.n4504 23.1255
R22417 VDD.n4504 VDD.n2384 23.1255
R22418 VDD.n4507 VDD.n4505 23.1255
R22419 VDD.n4505 VDD.n4503 23.1255
R22420 VDD.n4494 VDD.n4493 23.1255
R22421 VDD.n4495 VDD.n4494 23.1255
R22422 VDD.n4487 VDD.n4486 23.1255
R22423 VDD.n4488 VDD.n4487 23.1255
R22424 VDD.n4484 VDD.n4483 23.1255
R22425 VDD.n4485 VDD.n4484 23.1255
R22426 VDD.n4477 VDD.n4476 23.1255
R22427 VDD.n4478 VDD.n4477 23.1255
R22428 VDD.n4474 VDD.n4473 23.1255
R22429 VDD.n4475 VDD.n4474 23.1255
R22430 VDD.n4467 VDD.n4466 23.1255
R22431 VDD.n4468 VDD.n4467 23.1255
R22432 VDD.n4464 VDD.n4463 23.1255
R22433 VDD.n4465 VDD.n4464 23.1255
R22434 VDD.n4457 VDD.n4456 23.1255
R22435 VDD.n4458 VDD.n4457 23.1255
R22436 VDD.n4454 VDD.n4453 23.1255
R22437 VDD.n4455 VDD.n4454 23.1255
R22438 VDD.n4447 VDD.n4446 23.1255
R22439 VDD.n4448 VDD.n4447 23.1255
R22440 VDD.n2382 VDD.n2381 23.1255
R22441 VDD.n2383 VDD.n2382 23.1255
R22442 VDD.n4518 VDD.n4517 23.1255
R22443 VDD.n4519 VDD.n4518 23.1255
R22444 VDD.n2456 VDD.n2452 23.1255
R22445 VDD.n4434 VDD.n2452 23.1255
R22446 VDD.n4428 VDD.n2462 23.1255
R22447 VDD.n4428 VDD.n4427 23.1255
R22448 VDD.n2467 VDD.n2463 23.1255
R22449 VDD.n4424 VDD.n2463 23.1255
R22450 VDD.n4418 VDD.n2472 23.1255
R22451 VDD.n4418 VDD.n4417 23.1255
R22452 VDD.n2477 VDD.n2473 23.1255
R22453 VDD.n4414 VDD.n2473 23.1255
R22454 VDD.n4408 VDD.n2485 23.1255
R22455 VDD.n4408 VDD.n4407 23.1255
R22456 VDD.n2490 VDD.n2486 23.1255
R22457 VDD.n4404 VDD.n2486 23.1255
R22458 VDD.n4398 VDD.n2497 23.1255
R22459 VDD.n4398 VDD.n4397 23.1255
R22460 VDD.n2502 VDD.n2498 23.1255
R22461 VDD.n4394 VDD.n2498 23.1255
R22462 VDD.n2516 VDD.n2515 23.1255
R22463 VDD.n2519 VDD.n2516 23.1255
R22464 VDD.n2521 VDD.n2511 23.1255
R22465 VDD.n2520 VDD.n2511 23.1255
R22466 VDD.n2522 VDD.n2512 23.1255
R22467 VDD.n4378 VDD.n2512 23.1255
R22468 VDD.n4376 VDD.n4375 23.1255
R22469 VDD.n4377 VDD.n4376 23.1255
R22470 VDD.n4373 VDD.n4372 23.1255
R22471 VDD.n4372 VDD.n4371 23.1255
R22472 VDD.n2532 VDD.n2528 23.1255
R22473 VDD.n4370 VDD.n2528 23.1255
R22474 VDD.n4364 VDD.n2539 23.1255
R22475 VDD.n4364 VDD.n4363 23.1255
R22476 VDD.n2544 VDD.n2540 23.1255
R22477 VDD.n4360 VDD.n2540 23.1255
R22478 VDD.n4354 VDD.n2552 23.1255
R22479 VDD.n4354 VDD.n4353 23.1255
R22480 VDD.n2557 VDD.n2553 23.1255
R22481 VDD.n4350 VDD.n2553 23.1255
R22482 VDD.n4344 VDD.n2563 23.1255
R22483 VDD.n4344 VDD.n4343 23.1255
R22484 VDD.n2568 VDD.n2564 23.1255
R22485 VDD.n4340 VDD.n2564 23.1255
R22486 VDD.n4334 VDD.n2573 23.1255
R22487 VDD.n4334 VDD.n4333 23.1255
R22488 VDD.n2578 VDD.n2574 23.1255
R22489 VDD.n4330 VDD.n2574 23.1255
R22490 VDD.n4324 VDD.n4320 23.1255
R22491 VDD.n4324 VDD.n4323 23.1255
R22492 VDD.n2450 VDD.n2446 23.1255
R22493 VDD.n4437 VDD.n4436 23.1255
R22494 VDD.n4436 VDD.n4435 23.1255
R22495 VDD.n4433 VDD.n4432 23.1255
R22496 VDD.n4434 VDD.n4433 23.1255
R22497 VDD.n4426 VDD.n4425 23.1255
R22498 VDD.n4427 VDD.n4426 23.1255
R22499 VDD.n4423 VDD.n4422 23.1255
R22500 VDD.n4424 VDD.n4423 23.1255
R22501 VDD.n4416 VDD.n4415 23.1255
R22502 VDD.n4417 VDD.n4416 23.1255
R22503 VDD.n4413 VDD.n4412 23.1255
R22504 VDD.n4414 VDD.n4413 23.1255
R22505 VDD.n4406 VDD.n4405 23.1255
R22506 VDD.n4407 VDD.n4406 23.1255
R22507 VDD.n4403 VDD.n4402 23.1255
R22508 VDD.n4404 VDD.n4403 23.1255
R22509 VDD.n4396 VDD.n4395 23.1255
R22510 VDD.n4397 VDD.n4396 23.1255
R22511 VDD.n4381 VDD.n4379 23.1255
R22512 VDD.n4379 VDD.n2520 23.1255
R22513 VDD.n4382 VDD.n4380 23.1255
R22514 VDD.n4380 VDD.n4378 23.1255
R22515 VDD.n4369 VDD.n4368 23.1255
R22516 VDD.n4370 VDD.n4369 23.1255
R22517 VDD.n4362 VDD.n4361 23.1255
R22518 VDD.n4363 VDD.n4362 23.1255
R22519 VDD.n4359 VDD.n4358 23.1255
R22520 VDD.n4360 VDD.n4359 23.1255
R22521 VDD.n4352 VDD.n4351 23.1255
R22522 VDD.n4353 VDD.n4352 23.1255
R22523 VDD.n4349 VDD.n4348 23.1255
R22524 VDD.n4350 VDD.n4349 23.1255
R22525 VDD.n4342 VDD.n4341 23.1255
R22526 VDD.n4343 VDD.n4342 23.1255
R22527 VDD.n4339 VDD.n4338 23.1255
R22528 VDD.n4340 VDD.n4339 23.1255
R22529 VDD.n4332 VDD.n4331 23.1255
R22530 VDD.n4333 VDD.n4332 23.1255
R22531 VDD.n4329 VDD.n4328 23.1255
R22532 VDD.n4330 VDD.n4329 23.1255
R22533 VDD.n4322 VDD.n4321 23.1255
R22534 VDD.n4323 VDD.n4322 23.1255
R22535 VDD.n2518 VDD.n2517 23.1255
R22536 VDD.n2519 VDD.n2518 23.1255
R22537 VDD.n4393 VDD.n4392 23.1255
R22538 VDD.n4394 VDD.n4393 23.1255
R22539 VDD.n2592 VDD.n2588 23.1255
R22540 VDD.n4309 VDD.n2588 23.1255
R22541 VDD.n4303 VDD.n2598 23.1255
R22542 VDD.n4303 VDD.n4302 23.1255
R22543 VDD.n2603 VDD.n2599 23.1255
R22544 VDD.n4299 VDD.n2599 23.1255
R22545 VDD.n4293 VDD.n2608 23.1255
R22546 VDD.n4293 VDD.n4292 23.1255
R22547 VDD.n2613 VDD.n2609 23.1255
R22548 VDD.n4289 VDD.n2609 23.1255
R22549 VDD.n4283 VDD.n2621 23.1255
R22550 VDD.n4283 VDD.n4282 23.1255
R22551 VDD.n2626 VDD.n2622 23.1255
R22552 VDD.n4279 VDD.n2622 23.1255
R22553 VDD.n4273 VDD.n2633 23.1255
R22554 VDD.n4273 VDD.n4272 23.1255
R22555 VDD.n2638 VDD.n2634 23.1255
R22556 VDD.n4269 VDD.n2634 23.1255
R22557 VDD.n2652 VDD.n2651 23.1255
R22558 VDD.n2655 VDD.n2652 23.1255
R22559 VDD.n2657 VDD.n2647 23.1255
R22560 VDD.n2656 VDD.n2647 23.1255
R22561 VDD.n2658 VDD.n2648 23.1255
R22562 VDD.n4253 VDD.n2648 23.1255
R22563 VDD.n4251 VDD.n4250 23.1255
R22564 VDD.n4252 VDD.n4251 23.1255
R22565 VDD.n4248 VDD.n4247 23.1255
R22566 VDD.n4247 VDD.n4246 23.1255
R22567 VDD.n2668 VDD.n2664 23.1255
R22568 VDD.n4245 VDD.n2664 23.1255
R22569 VDD.n4239 VDD.n2675 23.1255
R22570 VDD.n4239 VDD.n4238 23.1255
R22571 VDD.n2680 VDD.n2676 23.1255
R22572 VDD.n4235 VDD.n2676 23.1255
R22573 VDD.n4229 VDD.n2688 23.1255
R22574 VDD.n4229 VDD.n4228 23.1255
R22575 VDD.n2693 VDD.n2689 23.1255
R22576 VDD.n4225 VDD.n2689 23.1255
R22577 VDD.n4219 VDD.n2699 23.1255
R22578 VDD.n4219 VDD.n4218 23.1255
R22579 VDD.n2704 VDD.n2700 23.1255
R22580 VDD.n4215 VDD.n2700 23.1255
R22581 VDD.n4209 VDD.n2709 23.1255
R22582 VDD.n4209 VDD.n4208 23.1255
R22583 VDD.n2714 VDD.n2710 23.1255
R22584 VDD.n4205 VDD.n2710 23.1255
R22585 VDD.n4199 VDD.n4195 23.1255
R22586 VDD.n4199 VDD.n4198 23.1255
R22587 VDD.n2586 VDD.n2582 23.1255
R22588 VDD.n4312 VDD.n4311 23.1255
R22589 VDD.n4311 VDD.n4310 23.1255
R22590 VDD.n4308 VDD.n4307 23.1255
R22591 VDD.n4309 VDD.n4308 23.1255
R22592 VDD.n4301 VDD.n4300 23.1255
R22593 VDD.n4302 VDD.n4301 23.1255
R22594 VDD.n4298 VDD.n4297 23.1255
R22595 VDD.n4299 VDD.n4298 23.1255
R22596 VDD.n4291 VDD.n4290 23.1255
R22597 VDD.n4292 VDD.n4291 23.1255
R22598 VDD.n4288 VDD.n4287 23.1255
R22599 VDD.n4289 VDD.n4288 23.1255
R22600 VDD.n4281 VDD.n4280 23.1255
R22601 VDD.n4282 VDD.n4281 23.1255
R22602 VDD.n4278 VDD.n4277 23.1255
R22603 VDD.n4279 VDD.n4278 23.1255
R22604 VDD.n4271 VDD.n4270 23.1255
R22605 VDD.n4272 VDD.n4271 23.1255
R22606 VDD.n4256 VDD.n4254 23.1255
R22607 VDD.n4254 VDD.n2656 23.1255
R22608 VDD.n4257 VDD.n4255 23.1255
R22609 VDD.n4255 VDD.n4253 23.1255
R22610 VDD.n4244 VDD.n4243 23.1255
R22611 VDD.n4245 VDD.n4244 23.1255
R22612 VDD.n4237 VDD.n4236 23.1255
R22613 VDD.n4238 VDD.n4237 23.1255
R22614 VDD.n4234 VDD.n4233 23.1255
R22615 VDD.n4235 VDD.n4234 23.1255
R22616 VDD.n4227 VDD.n4226 23.1255
R22617 VDD.n4228 VDD.n4227 23.1255
R22618 VDD.n4224 VDD.n4223 23.1255
R22619 VDD.n4225 VDD.n4224 23.1255
R22620 VDD.n4217 VDD.n4216 23.1255
R22621 VDD.n4218 VDD.n4217 23.1255
R22622 VDD.n4214 VDD.n4213 23.1255
R22623 VDD.n4215 VDD.n4214 23.1255
R22624 VDD.n4207 VDD.n4206 23.1255
R22625 VDD.n4208 VDD.n4207 23.1255
R22626 VDD.n4204 VDD.n4203 23.1255
R22627 VDD.n4205 VDD.n4204 23.1255
R22628 VDD.n4197 VDD.n4196 23.1255
R22629 VDD.n4198 VDD.n4197 23.1255
R22630 VDD.n2654 VDD.n2653 23.1255
R22631 VDD.n2655 VDD.n2654 23.1255
R22632 VDD.n4268 VDD.n4267 23.1255
R22633 VDD.n4269 VDD.n4268 23.1255
R22634 VDD.n2728 VDD.n2724 23.1255
R22635 VDD.n4184 VDD.n2724 23.1255
R22636 VDD.n4178 VDD.n2734 23.1255
R22637 VDD.n4178 VDD.n4177 23.1255
R22638 VDD.n2739 VDD.n2735 23.1255
R22639 VDD.n4174 VDD.n2735 23.1255
R22640 VDD.n4168 VDD.n2744 23.1255
R22641 VDD.n4168 VDD.n4167 23.1255
R22642 VDD.n2749 VDD.n2745 23.1255
R22643 VDD.n4164 VDD.n2745 23.1255
R22644 VDD.n4158 VDD.n2757 23.1255
R22645 VDD.n4158 VDD.n4157 23.1255
R22646 VDD.n2762 VDD.n2758 23.1255
R22647 VDD.n4154 VDD.n2758 23.1255
R22648 VDD.n4148 VDD.n2769 23.1255
R22649 VDD.n4148 VDD.n4147 23.1255
R22650 VDD.n2774 VDD.n2770 23.1255
R22651 VDD.n4144 VDD.n2770 23.1255
R22652 VDD.n2788 VDD.n2787 23.1255
R22653 VDD.n2791 VDD.n2788 23.1255
R22654 VDD.n2793 VDD.n2783 23.1255
R22655 VDD.n2792 VDD.n2783 23.1255
R22656 VDD.n2794 VDD.n2784 23.1255
R22657 VDD.n4128 VDD.n2784 23.1255
R22658 VDD.n4126 VDD.n4125 23.1255
R22659 VDD.n4127 VDD.n4126 23.1255
R22660 VDD.n4123 VDD.n4122 23.1255
R22661 VDD.n4122 VDD.n4121 23.1255
R22662 VDD.n2804 VDD.n2800 23.1255
R22663 VDD.n4120 VDD.n2800 23.1255
R22664 VDD.n4114 VDD.n2811 23.1255
R22665 VDD.n4114 VDD.n4113 23.1255
R22666 VDD.n2816 VDD.n2812 23.1255
R22667 VDD.n4110 VDD.n2812 23.1255
R22668 VDD.n4104 VDD.n2824 23.1255
R22669 VDD.n4104 VDD.n4103 23.1255
R22670 VDD.n2829 VDD.n2825 23.1255
R22671 VDD.n4100 VDD.n2825 23.1255
R22672 VDD.n4094 VDD.n2835 23.1255
R22673 VDD.n4094 VDD.n4093 23.1255
R22674 VDD.n2840 VDD.n2836 23.1255
R22675 VDD.n4090 VDD.n2836 23.1255
R22676 VDD.n4084 VDD.n2845 23.1255
R22677 VDD.n4084 VDD.n4083 23.1255
R22678 VDD.n2850 VDD.n2846 23.1255
R22679 VDD.n4080 VDD.n2846 23.1255
R22680 VDD.n4074 VDD.n4070 23.1255
R22681 VDD.n4074 VDD.n4073 23.1255
R22682 VDD.n2722 VDD.n2718 23.1255
R22683 VDD.n4187 VDD.n4186 23.1255
R22684 VDD.n4186 VDD.n4185 23.1255
R22685 VDD.n4183 VDD.n4182 23.1255
R22686 VDD.n4184 VDD.n4183 23.1255
R22687 VDD.n4176 VDD.n4175 23.1255
R22688 VDD.n4177 VDD.n4176 23.1255
R22689 VDD.n4173 VDD.n4172 23.1255
R22690 VDD.n4174 VDD.n4173 23.1255
R22691 VDD.n4166 VDD.n4165 23.1255
R22692 VDD.n4167 VDD.n4166 23.1255
R22693 VDD.n4163 VDD.n4162 23.1255
R22694 VDD.n4164 VDD.n4163 23.1255
R22695 VDD.n4156 VDD.n4155 23.1255
R22696 VDD.n4157 VDD.n4156 23.1255
R22697 VDD.n4153 VDD.n4152 23.1255
R22698 VDD.n4154 VDD.n4153 23.1255
R22699 VDD.n4146 VDD.n4145 23.1255
R22700 VDD.n4147 VDD.n4146 23.1255
R22701 VDD.n4131 VDD.n4129 23.1255
R22702 VDD.n4129 VDD.n2792 23.1255
R22703 VDD.n4132 VDD.n4130 23.1255
R22704 VDD.n4130 VDD.n4128 23.1255
R22705 VDD.n4119 VDD.n4118 23.1255
R22706 VDD.n4120 VDD.n4119 23.1255
R22707 VDD.n4112 VDD.n4111 23.1255
R22708 VDD.n4113 VDD.n4112 23.1255
R22709 VDD.n4109 VDD.n4108 23.1255
R22710 VDD.n4110 VDD.n4109 23.1255
R22711 VDD.n4102 VDD.n4101 23.1255
R22712 VDD.n4103 VDD.n4102 23.1255
R22713 VDD.n4099 VDD.n4098 23.1255
R22714 VDD.n4100 VDD.n4099 23.1255
R22715 VDD.n4092 VDD.n4091 23.1255
R22716 VDD.n4093 VDD.n4092 23.1255
R22717 VDD.n4089 VDD.n4088 23.1255
R22718 VDD.n4090 VDD.n4089 23.1255
R22719 VDD.n4082 VDD.n4081 23.1255
R22720 VDD.n4083 VDD.n4082 23.1255
R22721 VDD.n4079 VDD.n4078 23.1255
R22722 VDD.n4080 VDD.n4079 23.1255
R22723 VDD.n4072 VDD.n4071 23.1255
R22724 VDD.n4073 VDD.n4072 23.1255
R22725 VDD.n2790 VDD.n2789 23.1255
R22726 VDD.n2791 VDD.n2790 23.1255
R22727 VDD.n4143 VDD.n4142 23.1255
R22728 VDD.n4144 VDD.n4143 23.1255
R22729 VDD.n2864 VDD.n2860 23.1255
R22730 VDD.n4059 VDD.n2860 23.1255
R22731 VDD.n4053 VDD.n2870 23.1255
R22732 VDD.n4053 VDD.n4052 23.1255
R22733 VDD.n2875 VDD.n2871 23.1255
R22734 VDD.n4049 VDD.n2871 23.1255
R22735 VDD.n4043 VDD.n2880 23.1255
R22736 VDD.n4043 VDD.n4042 23.1255
R22737 VDD.n2885 VDD.n2881 23.1255
R22738 VDD.n4039 VDD.n2881 23.1255
R22739 VDD.n4033 VDD.n2893 23.1255
R22740 VDD.n4033 VDD.n4032 23.1255
R22741 VDD.n2898 VDD.n2894 23.1255
R22742 VDD.n4029 VDD.n2894 23.1255
R22743 VDD.n4023 VDD.n2905 23.1255
R22744 VDD.n4023 VDD.n4022 23.1255
R22745 VDD.n2910 VDD.n2906 23.1255
R22746 VDD.n4019 VDD.n2906 23.1255
R22747 VDD.n2924 VDD.n2923 23.1255
R22748 VDD.n2927 VDD.n2924 23.1255
R22749 VDD.n2929 VDD.n2919 23.1255
R22750 VDD.n2928 VDD.n2919 23.1255
R22751 VDD.n2930 VDD.n2920 23.1255
R22752 VDD.n4003 VDD.n2920 23.1255
R22753 VDD.n4001 VDD.n4000 23.1255
R22754 VDD.n4002 VDD.n4001 23.1255
R22755 VDD.n3998 VDD.n3997 23.1255
R22756 VDD.n3997 VDD.n3996 23.1255
R22757 VDD.n2940 VDD.n2936 23.1255
R22758 VDD.n3995 VDD.n2936 23.1255
R22759 VDD.n3989 VDD.n2947 23.1255
R22760 VDD.n3989 VDD.n3988 23.1255
R22761 VDD.n2952 VDD.n2948 23.1255
R22762 VDD.n3985 VDD.n2948 23.1255
R22763 VDD.n3979 VDD.n2960 23.1255
R22764 VDD.n3979 VDD.n3978 23.1255
R22765 VDD.n2965 VDD.n2961 23.1255
R22766 VDD.n3975 VDD.n2961 23.1255
R22767 VDD.n3969 VDD.n2971 23.1255
R22768 VDD.n3969 VDD.n3968 23.1255
R22769 VDD.n2976 VDD.n2972 23.1255
R22770 VDD.n3965 VDD.n2972 23.1255
R22771 VDD.n3959 VDD.n2981 23.1255
R22772 VDD.n3959 VDD.n3958 23.1255
R22773 VDD.n2986 VDD.n2982 23.1255
R22774 VDD.n3955 VDD.n2982 23.1255
R22775 VDD.n3949 VDD.n3945 23.1255
R22776 VDD.n3949 VDD.n3948 23.1255
R22777 VDD.n2858 VDD.n2854 23.1255
R22778 VDD.n4062 VDD.n4061 23.1255
R22779 VDD.n4061 VDD.n4060 23.1255
R22780 VDD.n4058 VDD.n4057 23.1255
R22781 VDD.n4059 VDD.n4058 23.1255
R22782 VDD.n4051 VDD.n4050 23.1255
R22783 VDD.n4052 VDD.n4051 23.1255
R22784 VDD.n4048 VDD.n4047 23.1255
R22785 VDD.n4049 VDD.n4048 23.1255
R22786 VDD.n4041 VDD.n4040 23.1255
R22787 VDD.n4042 VDD.n4041 23.1255
R22788 VDD.n4038 VDD.n4037 23.1255
R22789 VDD.n4039 VDD.n4038 23.1255
R22790 VDD.n4031 VDD.n4030 23.1255
R22791 VDD.n4032 VDD.n4031 23.1255
R22792 VDD.n4028 VDD.n4027 23.1255
R22793 VDD.n4029 VDD.n4028 23.1255
R22794 VDD.n4021 VDD.n4020 23.1255
R22795 VDD.n4022 VDD.n4021 23.1255
R22796 VDD.n4006 VDD.n4004 23.1255
R22797 VDD.n4004 VDD.n2928 23.1255
R22798 VDD.n4007 VDD.n4005 23.1255
R22799 VDD.n4005 VDD.n4003 23.1255
R22800 VDD.n3994 VDD.n3993 23.1255
R22801 VDD.n3995 VDD.n3994 23.1255
R22802 VDD.n3987 VDD.n3986 23.1255
R22803 VDD.n3988 VDD.n3987 23.1255
R22804 VDD.n3984 VDD.n3983 23.1255
R22805 VDD.n3985 VDD.n3984 23.1255
R22806 VDD.n3977 VDD.n3976 23.1255
R22807 VDD.n3978 VDD.n3977 23.1255
R22808 VDD.n3974 VDD.n3973 23.1255
R22809 VDD.n3975 VDD.n3974 23.1255
R22810 VDD.n3967 VDD.n3966 23.1255
R22811 VDD.n3968 VDD.n3967 23.1255
R22812 VDD.n3964 VDD.n3963 23.1255
R22813 VDD.n3965 VDD.n3964 23.1255
R22814 VDD.n3957 VDD.n3956 23.1255
R22815 VDD.n3958 VDD.n3957 23.1255
R22816 VDD.n3954 VDD.n3953 23.1255
R22817 VDD.n3955 VDD.n3954 23.1255
R22818 VDD.n3947 VDD.n3946 23.1255
R22819 VDD.n3948 VDD.n3947 23.1255
R22820 VDD.n2926 VDD.n2925 23.1255
R22821 VDD.n2927 VDD.n2926 23.1255
R22822 VDD.n4018 VDD.n4017 23.1255
R22823 VDD.n4019 VDD.n4018 23.1255
R22824 VDD.n3272 VDD.n3269 23.1255
R22825 VDD.n3271 VDD.n3269 23.1255
R22826 VDD.n3273 VDD.n3270 23.1255
R22827 VDD.n3608 VDD.n3270 23.1255
R22828 VDD.n3280 VDD.n3276 23.1255
R22829 VDD.n3607 VDD.n3276 23.1255
R22830 VDD.n3601 VDD.n3285 23.1255
R22831 VDD.n3601 VDD.n3600 23.1255
R22832 VDD.n3290 VDD.n3286 23.1255
R22833 VDD.n3597 VDD.n3286 23.1255
R22834 VDD.n3298 VDD.n3294 23.1255
R22835 VDD.n3298 VDD.n3297 23.1255
R22836 VDD.n3611 VDD.n3609 23.1255
R22837 VDD.n3609 VDD.n3271 23.1255
R22838 VDD.n3612 VDD.n3610 23.1255
R22839 VDD.n3610 VDD.n3608 23.1255
R22840 VDD.n3606 VDD.n3605 23.1255
R22841 VDD.n3607 VDD.n3606 23.1255
R22842 VDD.n3599 VDD.n3598 23.1255
R22843 VDD.n3600 VDD.n3599 23.1255
R22844 VDD.n3296 VDD.n3295 23.1255
R22845 VDD.n3297 VDD.n3296 23.1255
R22846 VDD.n3596 VDD.n3595 23.1255
R22847 VDD.n3597 VDD.n3596 23.1255
R22848 VDD.n3429 VDD.n3350 23.1255
R22849 VDD.n3430 VDD.n3429 23.1255
R22850 VDD.n3441 VDD.n3440 23.1255
R22851 VDD.n3442 VDD.n3441 23.1255
R22852 VDD.n3443 VDD.n3343 23.1255
R22853 VDD.n3444 VDD.n3443 23.1255
R22854 VDD.n3447 VDD.n3446 23.1255
R22855 VDD.n3433 VDD.n3432 23.1255
R22856 VDD.n3432 VDD.n3431 23.1255
R22857 VDD.n3427 VDD.n3423 23.1255
R22858 VDD.n3467 VDD.n3459 23.1255
R22859 VDD.n3468 VDD.n3467 23.1255
R22860 VDD.n3478 VDD.n3477 23.1255
R22861 VDD.n3479 VDD.n3478 23.1255
R22862 VDD.n3480 VDD.n3452 23.1255
R22863 VDD.n3481 VDD.n3480 23.1255
R22864 VDD.n3484 VDD.n3483 23.1255
R22865 VDD.n3471 VDD.n3470 23.1255
R22866 VDD.n3470 VDD.n3469 23.1255
R22867 VDD.n3465 VDD.n3461 23.1255
R22868 VDD.n3507 VDD.n3506 23.1255
R22869 VDD.n3508 VDD.n3507 23.1255
R22870 VDD.n3330 VDD.n3325 23.1255
R22871 VDD.n3331 VDD.n3330 23.1255
R22872 VDD.n3332 VDD.n3326 23.1255
R22873 VDD.n3333 VDD.n3332 23.1255
R22874 VDD.n3336 VDD.n3335 23.1255
R22875 VDD.n3511 VDD.n3510 23.1255
R22876 VDD.n3510 VDD.n3509 23.1255
R22877 VDD.n3320 VDD.n3316 23.1255
R22878 VDD.n3524 VDD.n3313 23.1255
R22879 VDD.n3525 VDD.n3524 23.1255
R22880 VDD.n3536 VDD.n3535 23.1255
R22881 VDD.n3537 VDD.n3536 23.1255
R22882 VDD.n3538 VDD.n3306 23.1255
R22883 VDD.n3539 VDD.n3538 23.1255
R22884 VDD.n3542 VDD.n3541 23.1255
R22885 VDD.n3528 VDD.n3527 23.1255
R22886 VDD.n3527 VDD.n3526 23.1255
R22887 VDD.n3522 VDD.n3518 23.1255
R22888 VDD.n3561 VDD.n3553 23.1255
R22889 VDD.n3562 VDD.n3561 23.1255
R22890 VDD.n3572 VDD.n3571 23.1255
R22891 VDD.n3573 VDD.n3572 23.1255
R22892 VDD.n3574 VDD.n3546 23.1255
R22893 VDD.n3575 VDD.n3574 23.1255
R22894 VDD.n3578 VDD.n3577 23.1255
R22895 VDD.n3565 VDD.n3564 23.1255
R22896 VDD.n3564 VDD.n3563 23.1255
R22897 VDD.n3559 VDD.n3555 23.1255
R22898 VDD.n3412 VDD.n3411 23.1255
R22899 VDD.n3413 VDD.n3412 23.1255
R22900 VDD.n3386 VDD.n3381 23.1255
R22901 VDD.n3387 VDD.n3386 23.1255
R22902 VDD.n3388 VDD.n3382 23.1255
R22903 VDD.n3389 VDD.n3388 23.1255
R22904 VDD.n3392 VDD.n3391 23.1255
R22905 VDD.n3416 VDD.n3415 23.1255
R22906 VDD.n3415 VDD.n3414 23.1255
R22907 VDD.n3376 VDD.n3372 23.1255
R22908 VDD.n3000 VDD.n2996 23.1255
R22909 VDD.n3934 VDD.n2996 23.1255
R22910 VDD.n3928 VDD.n3006 23.1255
R22911 VDD.n3928 VDD.n3927 23.1255
R22912 VDD.n3011 VDD.n3007 23.1255
R22913 VDD.n3924 VDD.n3007 23.1255
R22914 VDD.n3918 VDD.n3016 23.1255
R22915 VDD.n3918 VDD.n3917 23.1255
R22916 VDD.n3021 VDD.n3017 23.1255
R22917 VDD.n3914 VDD.n3017 23.1255
R22918 VDD.n3908 VDD.n3029 23.1255
R22919 VDD.n3908 VDD.n3907 23.1255
R22920 VDD.n3034 VDD.n3030 23.1255
R22921 VDD.n3904 VDD.n3030 23.1255
R22922 VDD.n3898 VDD.n3731 23.1255
R22923 VDD.n3898 VDD.n3897 23.1255
R22924 VDD.n3736 VDD.n3732 23.1255
R22925 VDD.n3894 VDD.n3732 23.1255
R22926 VDD.n3750 VDD.n3749 23.1255
R22927 VDD.n3753 VDD.n3750 23.1255
R22928 VDD.n3755 VDD.n3745 23.1255
R22929 VDD.n3754 VDD.n3745 23.1255
R22930 VDD.n3756 VDD.n3746 23.1255
R22931 VDD.n3878 VDD.n3746 23.1255
R22932 VDD.n3876 VDD.n3875 23.1255
R22933 VDD.n3877 VDD.n3876 23.1255
R22934 VDD.n3873 VDD.n3872 23.1255
R22935 VDD.n3872 VDD.n3871 23.1255
R22936 VDD.n3766 VDD.n3762 23.1255
R22937 VDD.n3870 VDD.n3762 23.1255
R22938 VDD.n3864 VDD.n3773 23.1255
R22939 VDD.n3864 VDD.n3863 23.1255
R22940 VDD.n3778 VDD.n3774 23.1255
R22941 VDD.n3860 VDD.n3774 23.1255
R22942 VDD.n3854 VDD.n3786 23.1255
R22943 VDD.n3854 VDD.n3853 23.1255
R22944 VDD.n3791 VDD.n3787 23.1255
R22945 VDD.n3850 VDD.n3787 23.1255
R22946 VDD.n3844 VDD.n3797 23.1255
R22947 VDD.n3844 VDD.n3843 23.1255
R22948 VDD.n3802 VDD.n3798 23.1255
R22949 VDD.n3840 VDD.n3798 23.1255
R22950 VDD.n3834 VDD.n3807 23.1255
R22951 VDD.n3834 VDD.n3833 23.1255
R22952 VDD.n3812 VDD.n3808 23.1255
R22953 VDD.n3830 VDD.n3808 23.1255
R22954 VDD.n3824 VDD.n3820 23.1255
R22955 VDD.n3824 VDD.n3823 23.1255
R22956 VDD.n2994 VDD.n2990 23.1255
R22957 VDD.n3937 VDD.n3936 23.1255
R22958 VDD.n3936 VDD.n3935 23.1255
R22959 VDD.n3933 VDD.n3932 23.1255
R22960 VDD.n3934 VDD.n3933 23.1255
R22961 VDD.n3926 VDD.n3925 23.1255
R22962 VDD.n3927 VDD.n3926 23.1255
R22963 VDD.n3923 VDD.n3922 23.1255
R22964 VDD.n3924 VDD.n3923 23.1255
R22965 VDD.n3916 VDD.n3915 23.1255
R22966 VDD.n3917 VDD.n3916 23.1255
R22967 VDD.n3913 VDD.n3912 23.1255
R22968 VDD.n3914 VDD.n3913 23.1255
R22969 VDD.n3906 VDD.n3905 23.1255
R22970 VDD.n3907 VDD.n3906 23.1255
R22971 VDD.n3903 VDD.n3902 23.1255
R22972 VDD.n3904 VDD.n3903 23.1255
R22973 VDD.n3896 VDD.n3895 23.1255
R22974 VDD.n3897 VDD.n3896 23.1255
R22975 VDD.n3881 VDD.n3879 23.1255
R22976 VDD.n3879 VDD.n3754 23.1255
R22977 VDD.n3882 VDD.n3880 23.1255
R22978 VDD.n3880 VDD.n3878 23.1255
R22979 VDD.n3869 VDD.n3868 23.1255
R22980 VDD.n3870 VDD.n3869 23.1255
R22981 VDD.n3862 VDD.n3861 23.1255
R22982 VDD.n3863 VDD.n3862 23.1255
R22983 VDD.n3859 VDD.n3858 23.1255
R22984 VDD.n3860 VDD.n3859 23.1255
R22985 VDD.n3852 VDD.n3851 23.1255
R22986 VDD.n3853 VDD.n3852 23.1255
R22987 VDD.n3849 VDD.n3848 23.1255
R22988 VDD.n3850 VDD.n3849 23.1255
R22989 VDD.n3842 VDD.n3841 23.1255
R22990 VDD.n3843 VDD.n3842 23.1255
R22991 VDD.n3839 VDD.n3838 23.1255
R22992 VDD.n3840 VDD.n3839 23.1255
R22993 VDD.n3832 VDD.n3831 23.1255
R22994 VDD.n3833 VDD.n3832 23.1255
R22995 VDD.n3829 VDD.n3828 23.1255
R22996 VDD.n3830 VDD.n3829 23.1255
R22997 VDD.n3822 VDD.n3821 23.1255
R22998 VDD.n3823 VDD.n3822 23.1255
R22999 VDD.n3752 VDD.n3751 23.1255
R23000 VDD.n3753 VDD.n3752 23.1255
R23001 VDD.n3893 VDD.n3892 23.1255
R23002 VDD.n3894 VDD.n3893 23.1255
R23003 VDD.n327 VDD.n326 21.3068
R23004 VDD.n326 VDD.n296 21.3068
R23005 VDD.n286 VDD.t402 20.9643
R23006 VDD.n293 VDD.n290 20.4313
R23007 VDD VDD.n3305 19.2885
R23008 VDD.n3194 VDD 18.5394
R23009 VDD.n304 VDD.t787 18.427
R23010 VDD.n304 VDD.t90 18.427
R23011 VDD.n3169 VDD.n3168 15.5222
R23012 VDD.n3233 VDD.n3232 15.5222
R23013 VDD.n3257 VDD.n3256 15.5222
R23014 VDD.n3634 VDD.n3633 15.5222
R23015 VDD.n3091 VDD.n3090 15.5222
R23016 VDD.n3678 VDD.n3677 15.5222
R23017 VDD.n3701 VDD.n3700 15.5222
R23018 VDD.n3188 VDD.n3187 15.5222
R23019 VDD.n3722 VDD.n3721 15.5222
R23020 VDD.n3545 VDD 14.6853
R23021 VDD.n341 VDD.n340 13.1442
R23022 VDD.n7131 VDD.n7130 10.9545
R23023 VDD VDD.n3300 9.59289
R23024 VDD.n3450 VDD 9.58202
R23025 VDD VDD.n3451 9.58202
R23026 VDD.n3545 VDD 9.58202
R23027 VDD.n1901 VDD.n1900 9.00833
R23028 VDD.n1641 VDD.n1640 9.00833
R23029 VDD.n1381 VDD.n1380 9.00833
R23030 VDD.n1121 VDD.n1120 9.00833
R23031 VDD.n861 VDD.n860 9.00833
R23032 VDD.n601 VDD.n600 9.00833
R23033 VDD.n7517 VDD.n7516 9.00833
R23034 VDD.n7519 VDD.n7518 9.00833
R23035 VDD.n3422 VDD.n3421 8.94311
R23036 VDD.n3460 VDD.n3314 8.94311
R23037 VDD.n3515 VDD.n3514 8.94311
R23038 VDD.n3517 VDD.n3516 8.94311
R23039 VDD.n3554 VDD.n3264 8.94311
R23040 VDD.n3420 VDD.n3419 8.94311
R23041 VDD.n3619 VDD.n3618 8.94311
R23042 VDD.n3154 VDD.n3141 8.48148
R23043 VDD.n3218 VDD.n3205 8.48148
R23044 VDD.n3115 VDD.n3102 8.48148
R23045 VDD.n3369 VDD.n3356 8.48148
R23046 VDD.n3076 VDD.n3063 8.48148
R23047 VDD.n3663 VDD.n3650 8.48148
R23048 VDD.n3056 VDD.n3043 8.48148
R23049 VDD.n3134 VDD.n3121 8.48148
R23050 VDD VDD.n3342 8.38365
R23051 VDD.n3055 VDD.n3048 8.26552
R23052 VDD.n7130 VDD.n7129 7.9105
R23053 VDD.n3401 VDD.n3341 7.9105
R23054 VDD.n3488 VDD.n3487 7.9105
R23055 VDD.n3502 VDD.n3501 7.9105
R23056 VDD.n3496 VDD.n3304 7.9105
R23057 VDD.n3582 VDD.n3581 7.9105
R23058 VDD.n3407 VDD.n3406 7.9105
R23059 VDD.n3591 VDD.n3590 7.9105
R23060 VDD.n3727 VDD.n3726 7.9105
R23061 VDD.n3705 VDD.n2901 7.9105
R23062 VDD.n3682 VDD.n2765 7.9105
R23063 VDD.n3095 VDD.n2629 7.9105
R23064 VDD.n3638 VDD.n2493 7.9105
R23065 VDD.n3261 VDD.n2357 7.9105
R23066 VDD.n3237 VDD.n2221 7.9105
R23067 VDD.n3173 VDD.n2085 7.9105
R23068 VDD.n3192 VDD.n1949 7.9105
R23069 VDD.n3153 VDD 7.85707
R23070 VDD.n3169 VDD 7.85707
R23071 VDD.n3217 VDD 7.85707
R23072 VDD.n3233 VDD 7.85707
R23073 VDD.n3114 VDD 7.85707
R23074 VDD.n3257 VDD 7.85707
R23075 VDD.n3368 VDD 7.85707
R23076 VDD.n3634 VDD 7.85707
R23077 VDD.n3075 VDD 7.85707
R23078 VDD.n3091 VDD 7.85707
R23079 VDD.n3662 VDD 7.85707
R23080 VDD.n3678 VDD 7.85707
R23081 VDD.n3701 VDD 7.85707
R23082 VDD.n3133 VDD 7.85707
R23083 VDD.n3188 VDD 7.85707
R23084 VDD.n3722 VDD 7.85707
R23085 VDD.n7651 VDD.n7650 7.39606
R23086 VDD.n7650 VDD.n7641 7.39606
R23087 VDD.n7661 VDD.n7660 7.39606
R23088 VDD.n7660 VDD.n7628 7.39606
R23089 VDD.n7671 VDD.n7670 7.39606
R23090 VDD.n7670 VDD.n7618 7.39606
R23091 VDD.n7681 VDD.n7680 7.39606
R23092 VDD.n7680 VDD.n7607 7.39606
R23093 VDD.n7691 VDD.n7690 7.39606
R23094 VDD.n7690 VDD.n7594 7.39606
R23095 VDD.n7708 VDD.n7707 7.39606
R23096 VDD.n7707 VDD.n7579 7.39606
R23097 VDD.n7718 VDD.n7717 7.39606
R23098 VDD.n7717 VDD.n7566 7.39606
R23099 VDD.n7730 VDD.n2 7.39606
R23100 VDD.n7730 VDD.n4 7.39606
R23101 VDD.n7551 VDD.n12 7.39606
R23102 VDD.n7552 VDD.n7551 7.39606
R23103 VDD.n7541 VDD.n21 7.39606
R23104 VDD.n7542 VDD.n7541 7.39606
R23105 VDD.n7531 VDD.n34 7.39606
R23106 VDD.n7532 VDD.n7531 7.39606
R23107 VDD.n1784 VDD.n1783 7.39606
R23108 VDD.n1783 VDD.n1774 7.39606
R23109 VDD.n1794 VDD.n1793 7.39606
R23110 VDD.n1793 VDD.n1761 7.39606
R23111 VDD.n1804 VDD.n1803 7.39606
R23112 VDD.n1803 VDD.n1751 7.39606
R23113 VDD.n1814 VDD.n1813 7.39606
R23114 VDD.n1813 VDD.n1740 7.39606
R23115 VDD.n1824 VDD.n1823 7.39606
R23116 VDD.n1823 VDD.n1727 7.39606
R23117 VDD.n1841 VDD.n1840 7.39606
R23118 VDD.n1840 VDD.n1712 7.39606
R23119 VDD.n1851 VDD.n1850 7.39606
R23120 VDD.n1850 VDD.n1699 7.39606
R23121 VDD.n1861 VDD.n1860 7.39606
R23122 VDD.n1860 VDD.n1689 7.39606
R23123 VDD.n1871 VDD.n1870 7.39606
R23124 VDD.n1870 VDD.n1678 7.39606
R23125 VDD.n1881 VDD.n1880 7.39606
R23126 VDD.n1880 VDD.n1665 7.39606
R23127 VDD.n1891 VDD.n1890 7.39606
R23128 VDD.n1890 VDD.n1655 7.39606
R23129 VDD.n1524 VDD.n1523 7.39606
R23130 VDD.n1523 VDD.n1514 7.39606
R23131 VDD.n1534 VDD.n1533 7.39606
R23132 VDD.n1533 VDD.n1501 7.39606
R23133 VDD.n1544 VDD.n1543 7.39606
R23134 VDD.n1543 VDD.n1491 7.39606
R23135 VDD.n1554 VDD.n1553 7.39606
R23136 VDD.n1553 VDD.n1480 7.39606
R23137 VDD.n1564 VDD.n1563 7.39606
R23138 VDD.n1563 VDD.n1467 7.39606
R23139 VDD.n1581 VDD.n1580 7.39606
R23140 VDD.n1580 VDD.n1452 7.39606
R23141 VDD.n1591 VDD.n1590 7.39606
R23142 VDD.n1590 VDD.n1439 7.39606
R23143 VDD.n1601 VDD.n1600 7.39606
R23144 VDD.n1600 VDD.n1429 7.39606
R23145 VDD.n1611 VDD.n1610 7.39606
R23146 VDD.n1610 VDD.n1418 7.39606
R23147 VDD.n1621 VDD.n1620 7.39606
R23148 VDD.n1620 VDD.n1405 7.39606
R23149 VDD.n1631 VDD.n1630 7.39606
R23150 VDD.n1630 VDD.n1395 7.39606
R23151 VDD.n1264 VDD.n1263 7.39606
R23152 VDD.n1263 VDD.n1254 7.39606
R23153 VDD.n1274 VDD.n1273 7.39606
R23154 VDD.n1273 VDD.n1241 7.39606
R23155 VDD.n1284 VDD.n1283 7.39606
R23156 VDD.n1283 VDD.n1231 7.39606
R23157 VDD.n1294 VDD.n1293 7.39606
R23158 VDD.n1293 VDD.n1220 7.39606
R23159 VDD.n1304 VDD.n1303 7.39606
R23160 VDD.n1303 VDD.n1207 7.39606
R23161 VDD.n1321 VDD.n1320 7.39606
R23162 VDD.n1320 VDD.n1192 7.39606
R23163 VDD.n1331 VDD.n1330 7.39606
R23164 VDD.n1330 VDD.n1179 7.39606
R23165 VDD.n1341 VDD.n1340 7.39606
R23166 VDD.n1340 VDD.n1169 7.39606
R23167 VDD.n1351 VDD.n1350 7.39606
R23168 VDD.n1350 VDD.n1158 7.39606
R23169 VDD.n1361 VDD.n1360 7.39606
R23170 VDD.n1360 VDD.n1145 7.39606
R23171 VDD.n1371 VDD.n1370 7.39606
R23172 VDD.n1370 VDD.n1135 7.39606
R23173 VDD.n1004 VDD.n1003 7.39606
R23174 VDD.n1003 VDD.n994 7.39606
R23175 VDD.n1014 VDD.n1013 7.39606
R23176 VDD.n1013 VDD.n981 7.39606
R23177 VDD.n1024 VDD.n1023 7.39606
R23178 VDD.n1023 VDD.n971 7.39606
R23179 VDD.n1034 VDD.n1033 7.39606
R23180 VDD.n1033 VDD.n960 7.39606
R23181 VDD.n1044 VDD.n1043 7.39606
R23182 VDD.n1043 VDD.n947 7.39606
R23183 VDD.n1061 VDD.n1060 7.39606
R23184 VDD.n1060 VDD.n932 7.39606
R23185 VDD.n1071 VDD.n1070 7.39606
R23186 VDD.n1070 VDD.n919 7.39606
R23187 VDD.n1081 VDD.n1080 7.39606
R23188 VDD.n1080 VDD.n909 7.39606
R23189 VDD.n1091 VDD.n1090 7.39606
R23190 VDD.n1090 VDD.n898 7.39606
R23191 VDD.n1101 VDD.n1100 7.39606
R23192 VDD.n1100 VDD.n885 7.39606
R23193 VDD.n1111 VDD.n1110 7.39606
R23194 VDD.n1110 VDD.n875 7.39606
R23195 VDD.n744 VDD.n743 7.39606
R23196 VDD.n743 VDD.n734 7.39606
R23197 VDD.n754 VDD.n753 7.39606
R23198 VDD.n753 VDD.n721 7.39606
R23199 VDD.n764 VDD.n763 7.39606
R23200 VDD.n763 VDD.n711 7.39606
R23201 VDD.n774 VDD.n773 7.39606
R23202 VDD.n773 VDD.n700 7.39606
R23203 VDD.n784 VDD.n783 7.39606
R23204 VDD.n783 VDD.n687 7.39606
R23205 VDD.n801 VDD.n800 7.39606
R23206 VDD.n800 VDD.n672 7.39606
R23207 VDD.n811 VDD.n810 7.39606
R23208 VDD.n810 VDD.n659 7.39606
R23209 VDD.n821 VDD.n820 7.39606
R23210 VDD.n820 VDD.n649 7.39606
R23211 VDD.n831 VDD.n830 7.39606
R23212 VDD.n830 VDD.n638 7.39606
R23213 VDD.n841 VDD.n840 7.39606
R23214 VDD.n840 VDD.n625 7.39606
R23215 VDD.n851 VDD.n850 7.39606
R23216 VDD.n850 VDD.n615 7.39606
R23217 VDD.n484 VDD.n483 7.39606
R23218 VDD.n483 VDD.n474 7.39606
R23219 VDD.n494 VDD.n493 7.39606
R23220 VDD.n493 VDD.n461 7.39606
R23221 VDD.n504 VDD.n503 7.39606
R23222 VDD.n503 VDD.n451 7.39606
R23223 VDD.n514 VDD.n513 7.39606
R23224 VDD.n513 VDD.n440 7.39606
R23225 VDD.n524 VDD.n523 7.39606
R23226 VDD.n523 VDD.n427 7.39606
R23227 VDD.n541 VDD.n540 7.39606
R23228 VDD.n540 VDD.n412 7.39606
R23229 VDD.n551 VDD.n550 7.39606
R23230 VDD.n550 VDD.n399 7.39606
R23231 VDD.n561 VDD.n560 7.39606
R23232 VDD.n560 VDD.n389 7.39606
R23233 VDD.n571 VDD.n570 7.39606
R23234 VDD.n570 VDD.n378 7.39606
R23235 VDD.n581 VDD.n580 7.39606
R23236 VDD.n580 VDD.n365 7.39606
R23237 VDD.n591 VDD.n590 7.39606
R23238 VDD.n590 VDD.n355 7.39606
R23239 VDD.n7400 VDD.n7399 7.39606
R23240 VDD.n7399 VDD.n7390 7.39606
R23241 VDD.n7410 VDD.n7409 7.39606
R23242 VDD.n7409 VDD.n7377 7.39606
R23243 VDD.n7420 VDD.n7419 7.39606
R23244 VDD.n7419 VDD.n7367 7.39606
R23245 VDD.n7430 VDD.n7429 7.39606
R23246 VDD.n7429 VDD.n7356 7.39606
R23247 VDD.n7440 VDD.n7439 7.39606
R23248 VDD.n7439 VDD.n7343 7.39606
R23249 VDD.n7457 VDD.n7456 7.39606
R23250 VDD.n7456 VDD.n7328 7.39606
R23251 VDD.n7467 VDD.n7466 7.39606
R23252 VDD.n7466 VDD.n7315 7.39606
R23253 VDD.n7477 VDD.n7476 7.39606
R23254 VDD.n7476 VDD.n7305 7.39606
R23255 VDD.n7487 VDD.n7486 7.39606
R23256 VDD.n7486 VDD.n7294 7.39606
R23257 VDD.n7497 VDD.n7496 7.39606
R23258 VDD.n7496 VDD.n7281 7.39606
R23259 VDD.n7507 VDD.n7506 7.39606
R23260 VDD.n7506 VDD.n7271 7.39606
R23261 VDD.n7143 VDD.n7142 7.39606
R23262 VDD.n7142 VDD.n7133 7.39606
R23263 VDD.n7153 VDD.n7152 7.39606
R23264 VDD.n7152 VDD.n2026 7.39606
R23265 VDD.n7163 VDD.n7162 7.39606
R23266 VDD.n7162 VDD.n2016 7.39606
R23267 VDD.n7173 VDD.n7172 7.39606
R23268 VDD.n7172 VDD.n2005 7.39606
R23269 VDD.n7183 VDD.n7182 7.39606
R23270 VDD.n7182 VDD.n1992 7.39606
R23271 VDD.n7202 VDD.n1964 7.39606
R23272 VDD.n7202 VDD.n1966 7.39606
R23273 VDD.n7217 VDD.n7216 7.39606
R23274 VDD.n7216 VDD.n1950 7.39606
R23275 VDD.n7227 VDD.n7226 7.39606
R23276 VDD.n7226 VDD.n1938 7.39606
R23277 VDD.n7237 VDD.n7236 7.39606
R23278 VDD.n7236 VDD.n1925 7.39606
R23279 VDD.n7247 VDD.n7246 7.39606
R23280 VDD.n7246 VDD.n1915 7.39606
R23281 VDD.n7207 VDD.n7206 7.39606
R23282 VDD.n7206 VDD.n1959 7.39606
R23283 VDD.n6038 VDD.n6037 7.39606
R23284 VDD.n6037 VDD.n6015 7.39606
R23285 VDD.n6048 VDD.n6047 7.39606
R23286 VDD.n6047 VDD.n6005 7.39606
R23287 VDD.n6058 VDD.n6057 7.39606
R23288 VDD.n6057 VDD.n5992 7.39606
R23289 VDD.n6068 VDD.n6067 7.39606
R23290 VDD.n6067 VDD.n5981 7.39606
R23291 VDD.n6078 VDD.n6077 7.39606
R23292 VDD.n6077 VDD.n5971 7.39606
R23293 VDD.n6088 VDD.n6087 7.39606
R23294 VDD.n6087 VDD.n5958 7.39606
R23295 VDD.n6105 VDD.n6104 7.39606
R23296 VDD.n6104 VDD.n5943 7.39606
R23297 VDD.n6115 VDD.n6114 7.39606
R23298 VDD.n6114 VDD.n5930 7.39606
R23299 VDD.n6125 VDD.n6124 7.39606
R23300 VDD.n6124 VDD.n5919 7.39606
R23301 VDD.n6135 VDD.n6134 7.39606
R23302 VDD.n6134 VDD.n5909 7.39606
R23303 VDD.n6147 VDD.n5893 7.39606
R23304 VDD.n6147 VDD.n5895 7.39606
R23305 VDD.n6161 VDD.n6160 7.39606
R23306 VDD.n6160 VDD.n5879 7.39606
R23307 VDD.n6171 VDD.n6170 7.39606
R23308 VDD.n6170 VDD.n5869 7.39606
R23309 VDD.n6181 VDD.n6180 7.39606
R23310 VDD.n6180 VDD.n5856 7.39606
R23311 VDD.n6191 VDD.n6190 7.39606
R23312 VDD.n6190 VDD.n5845 7.39606
R23313 VDD.n6201 VDD.n6200 7.39606
R23314 VDD.n6200 VDD.n5835 7.39606
R23315 VDD.n6211 VDD.n6210 7.39606
R23316 VDD.n6210 VDD.n5822 7.39606
R23317 VDD.n6228 VDD.n6227 7.39606
R23318 VDD.n6227 VDD.n5807 7.39606
R23319 VDD.n6238 VDD.n6237 7.39606
R23320 VDD.n6237 VDD.n5794 7.39606
R23321 VDD.n6248 VDD.n6247 7.39606
R23322 VDD.n6247 VDD.n5783 7.39606
R23323 VDD.n6258 VDD.n6257 7.39606
R23324 VDD.n6257 VDD.n5773 7.39606
R23325 VDD.n6270 VDD.n5757 7.39606
R23326 VDD.n6270 VDD.n5759 7.39606
R23327 VDD.n6284 VDD.n6283 7.39606
R23328 VDD.n6283 VDD.n5743 7.39606
R23329 VDD.n6294 VDD.n6293 7.39606
R23330 VDD.n6293 VDD.n5733 7.39606
R23331 VDD.n6304 VDD.n6303 7.39606
R23332 VDD.n6303 VDD.n5720 7.39606
R23333 VDD.n6314 VDD.n6313 7.39606
R23334 VDD.n6313 VDD.n5709 7.39606
R23335 VDD.n6324 VDD.n6323 7.39606
R23336 VDD.n6323 VDD.n5699 7.39606
R23337 VDD.n6334 VDD.n6333 7.39606
R23338 VDD.n6333 VDD.n5686 7.39606
R23339 VDD.n6351 VDD.n6350 7.39606
R23340 VDD.n6350 VDD.n5671 7.39606
R23341 VDD.n6361 VDD.n6360 7.39606
R23342 VDD.n6360 VDD.n5658 7.39606
R23343 VDD.n6371 VDD.n6370 7.39606
R23344 VDD.n6370 VDD.n5647 7.39606
R23345 VDD.n6381 VDD.n6380 7.39606
R23346 VDD.n6380 VDD.n5637 7.39606
R23347 VDD.n6393 VDD.n5621 7.39606
R23348 VDD.n6393 VDD.n5623 7.39606
R23349 VDD.n6407 VDD.n6406 7.39606
R23350 VDD.n6406 VDD.n5607 7.39606
R23351 VDD.n6417 VDD.n6416 7.39606
R23352 VDD.n6416 VDD.n5597 7.39606
R23353 VDD.n6427 VDD.n6426 7.39606
R23354 VDD.n6426 VDD.n5584 7.39606
R23355 VDD.n6437 VDD.n6436 7.39606
R23356 VDD.n6436 VDD.n5573 7.39606
R23357 VDD.n6447 VDD.n6446 7.39606
R23358 VDD.n6446 VDD.n5563 7.39606
R23359 VDD.n6457 VDD.n6456 7.39606
R23360 VDD.n6456 VDD.n5550 7.39606
R23361 VDD.n6474 VDD.n6473 7.39606
R23362 VDD.n6473 VDD.n5535 7.39606
R23363 VDD.n6484 VDD.n6483 7.39606
R23364 VDD.n6483 VDD.n5522 7.39606
R23365 VDD.n6494 VDD.n6493 7.39606
R23366 VDD.n6493 VDD.n5511 7.39606
R23367 VDD.n6504 VDD.n6503 7.39606
R23368 VDD.n6503 VDD.n5501 7.39606
R23369 VDD.n6516 VDD.n5485 7.39606
R23370 VDD.n6516 VDD.n5487 7.39606
R23371 VDD.n6530 VDD.n6529 7.39606
R23372 VDD.n6529 VDD.n5471 7.39606
R23373 VDD.n6540 VDD.n6539 7.39606
R23374 VDD.n6539 VDD.n5461 7.39606
R23375 VDD.n6550 VDD.n6549 7.39606
R23376 VDD.n6549 VDD.n5448 7.39606
R23377 VDD.n6560 VDD.n6559 7.39606
R23378 VDD.n6559 VDD.n5437 7.39606
R23379 VDD.n6570 VDD.n6569 7.39606
R23380 VDD.n6569 VDD.n5427 7.39606
R23381 VDD.n6580 VDD.n6579 7.39606
R23382 VDD.n6579 VDD.n5414 7.39606
R23383 VDD.n6597 VDD.n6596 7.39606
R23384 VDD.n6596 VDD.n5399 7.39606
R23385 VDD.n6607 VDD.n6606 7.39606
R23386 VDD.n6606 VDD.n5386 7.39606
R23387 VDD.n6617 VDD.n6616 7.39606
R23388 VDD.n6616 VDD.n5375 7.39606
R23389 VDD.n6627 VDD.n6626 7.39606
R23390 VDD.n6626 VDD.n5365 7.39606
R23391 VDD.n6639 VDD.n5349 7.39606
R23392 VDD.n6639 VDD.n5351 7.39606
R23393 VDD.n6653 VDD.n6652 7.39606
R23394 VDD.n6652 VDD.n5335 7.39606
R23395 VDD.n6663 VDD.n6662 7.39606
R23396 VDD.n6662 VDD.n5325 7.39606
R23397 VDD.n6673 VDD.n6672 7.39606
R23398 VDD.n6672 VDD.n5312 7.39606
R23399 VDD.n6683 VDD.n6682 7.39606
R23400 VDD.n6682 VDD.n5301 7.39606
R23401 VDD.n6693 VDD.n6692 7.39606
R23402 VDD.n6692 VDD.n5291 7.39606
R23403 VDD.n6703 VDD.n6702 7.39606
R23404 VDD.n6702 VDD.n5278 7.39606
R23405 VDD.n6720 VDD.n6719 7.39606
R23406 VDD.n6719 VDD.n5263 7.39606
R23407 VDD.n6730 VDD.n6729 7.39606
R23408 VDD.n6729 VDD.n5250 7.39606
R23409 VDD.n6740 VDD.n6739 7.39606
R23410 VDD.n6739 VDD.n5239 7.39606
R23411 VDD.n6750 VDD.n6749 7.39606
R23412 VDD.n6749 VDD.n5229 7.39606
R23413 VDD.n6762 VDD.n5213 7.39606
R23414 VDD.n6762 VDD.n5215 7.39606
R23415 VDD.n6776 VDD.n6775 7.39606
R23416 VDD.n6775 VDD.n5199 7.39606
R23417 VDD.n6786 VDD.n6785 7.39606
R23418 VDD.n6785 VDD.n5189 7.39606
R23419 VDD.n6796 VDD.n6795 7.39606
R23420 VDD.n6795 VDD.n5176 7.39606
R23421 VDD.n6806 VDD.n6805 7.39606
R23422 VDD.n6805 VDD.n5165 7.39606
R23423 VDD.n6816 VDD.n6815 7.39606
R23424 VDD.n6815 VDD.n5155 7.39606
R23425 VDD.n6826 VDD.n6825 7.39606
R23426 VDD.n6825 VDD.n5142 7.39606
R23427 VDD.n6843 VDD.n6842 7.39606
R23428 VDD.n6842 VDD.n5127 7.39606
R23429 VDD.n6853 VDD.n6852 7.39606
R23430 VDD.n6852 VDD.n5114 7.39606
R23431 VDD.n6863 VDD.n6862 7.39606
R23432 VDD.n6862 VDD.n5103 7.39606
R23433 VDD.n6873 VDD.n6872 7.39606
R23434 VDD.n6872 VDD.n5093 7.39606
R23435 VDD.n6885 VDD.n5077 7.39606
R23436 VDD.n6885 VDD.n5079 7.39606
R23437 VDD.n5061 VDD.n4825 7.39606
R23438 VDD.n5062 VDD.n5061 7.39606
R23439 VDD.n5051 VDD.n4836 7.39606
R23440 VDD.n5052 VDD.n5051 7.39606
R23441 VDD.n5041 VDD.n4846 7.39606
R23442 VDD.n5042 VDD.n5041 7.39606
R23443 VDD.n5031 VDD.n4859 7.39606
R23444 VDD.n5032 VDD.n5031 7.39606
R23445 VDD.n5021 VDD.n4870 7.39606
R23446 VDD.n5022 VDD.n5021 7.39606
R23447 VDD.n5011 VDD.n4880 7.39606
R23448 VDD.n5012 VDD.n5011 7.39606
R23449 VDD.n4994 VDD.n4896 7.39606
R23450 VDD.n4995 VDD.n4994 7.39606
R23451 VDD.n4984 VDD.n4908 7.39606
R23452 VDD.n4985 VDD.n4984 7.39606
R23453 VDD.n4974 VDD.n4921 7.39606
R23454 VDD.n4975 VDD.n4974 7.39606
R23455 VDD.n4964 VDD.n4932 7.39606
R23456 VDD.n4965 VDD.n4964 7.39606
R23457 VDD.n4954 VDD.n4942 7.39606
R23458 VDD.n4955 VDD.n4954 7.39606
R23459 VDD.n4702 VDD.n4701 7.39606
R23460 VDD.n4701 VDD.n4692 7.39606
R23461 VDD.n4712 VDD.n4711 7.39606
R23462 VDD.n4711 VDD.n2162 7.39606
R23463 VDD.n4722 VDD.n4721 7.39606
R23464 VDD.n4721 VDD.n2152 7.39606
R23465 VDD.n4732 VDD.n4731 7.39606
R23466 VDD.n4731 VDD.n2141 7.39606
R23467 VDD.n4742 VDD.n4741 7.39606
R23468 VDD.n4741 VDD.n2128 7.39606
R23469 VDD.n4761 VDD.n2100 7.39606
R23470 VDD.n4761 VDD.n2102 7.39606
R23471 VDD.n4776 VDD.n4775 7.39606
R23472 VDD.n4775 VDD.n2086 7.39606
R23473 VDD.n4786 VDD.n4785 7.39606
R23474 VDD.n4785 VDD.n2074 7.39606
R23475 VDD.n4796 VDD.n4795 7.39606
R23476 VDD.n4795 VDD.n2061 7.39606
R23477 VDD.n4806 VDD.n4805 7.39606
R23478 VDD.n4805 VDD.n2051 7.39606
R23479 VDD.n4766 VDD.n4765 7.39606
R23480 VDD.n4765 VDD.n2095 7.39606
R23481 VDD.n4577 VDD.n4576 7.39606
R23482 VDD.n4576 VDD.n4567 7.39606
R23483 VDD.n4587 VDD.n4586 7.39606
R23484 VDD.n4586 VDD.n2298 7.39606
R23485 VDD.n4597 VDD.n4596 7.39606
R23486 VDD.n4596 VDD.n2288 7.39606
R23487 VDD.n4607 VDD.n4606 7.39606
R23488 VDD.n4606 VDD.n2277 7.39606
R23489 VDD.n4617 VDD.n4616 7.39606
R23490 VDD.n4616 VDD.n2264 7.39606
R23491 VDD.n4636 VDD.n2236 7.39606
R23492 VDD.n4636 VDD.n2238 7.39606
R23493 VDD.n4651 VDD.n4650 7.39606
R23494 VDD.n4650 VDD.n2222 7.39606
R23495 VDD.n4661 VDD.n4660 7.39606
R23496 VDD.n4660 VDD.n2210 7.39606
R23497 VDD.n4671 VDD.n4670 7.39606
R23498 VDD.n4670 VDD.n2197 7.39606
R23499 VDD.n4681 VDD.n4680 7.39606
R23500 VDD.n4680 VDD.n2187 7.39606
R23501 VDD.n4641 VDD.n4640 7.39606
R23502 VDD.n4640 VDD.n2231 7.39606
R23503 VDD.n4452 VDD.n4451 7.39606
R23504 VDD.n4451 VDD.n4442 7.39606
R23505 VDD.n4462 VDD.n4461 7.39606
R23506 VDD.n4461 VDD.n2434 7.39606
R23507 VDD.n4472 VDD.n4471 7.39606
R23508 VDD.n4471 VDD.n2424 7.39606
R23509 VDD.n4482 VDD.n4481 7.39606
R23510 VDD.n4481 VDD.n2413 7.39606
R23511 VDD.n4492 VDD.n4491 7.39606
R23512 VDD.n4491 VDD.n2400 7.39606
R23513 VDD.n4511 VDD.n2372 7.39606
R23514 VDD.n4511 VDD.n2374 7.39606
R23515 VDD.n4526 VDD.n4525 7.39606
R23516 VDD.n4525 VDD.n2358 7.39606
R23517 VDD.n4536 VDD.n4535 7.39606
R23518 VDD.n4535 VDD.n2346 7.39606
R23519 VDD.n4546 VDD.n4545 7.39606
R23520 VDD.n4545 VDD.n2333 7.39606
R23521 VDD.n4556 VDD.n4555 7.39606
R23522 VDD.n4555 VDD.n2323 7.39606
R23523 VDD.n4516 VDD.n4515 7.39606
R23524 VDD.n4515 VDD.n2367 7.39606
R23525 VDD.n4327 VDD.n4326 7.39606
R23526 VDD.n4326 VDD.n4317 7.39606
R23527 VDD.n4337 VDD.n4336 7.39606
R23528 VDD.n4336 VDD.n2570 7.39606
R23529 VDD.n4347 VDD.n4346 7.39606
R23530 VDD.n4346 VDD.n2560 7.39606
R23531 VDD.n4357 VDD.n4356 7.39606
R23532 VDD.n4356 VDD.n2549 7.39606
R23533 VDD.n4367 VDD.n4366 7.39606
R23534 VDD.n4366 VDD.n2536 7.39606
R23535 VDD.n4386 VDD.n2508 7.39606
R23536 VDD.n4386 VDD.n2510 7.39606
R23537 VDD.n4401 VDD.n4400 7.39606
R23538 VDD.n4400 VDD.n2494 7.39606
R23539 VDD.n4411 VDD.n4410 7.39606
R23540 VDD.n4410 VDD.n2482 7.39606
R23541 VDD.n4421 VDD.n4420 7.39606
R23542 VDD.n4420 VDD.n2469 7.39606
R23543 VDD.n4431 VDD.n4430 7.39606
R23544 VDD.n4430 VDD.n2459 7.39606
R23545 VDD.n4391 VDD.n4390 7.39606
R23546 VDD.n4390 VDD.n2503 7.39606
R23547 VDD.n4202 VDD.n4201 7.39606
R23548 VDD.n4201 VDD.n4192 7.39606
R23549 VDD.n4212 VDD.n4211 7.39606
R23550 VDD.n4211 VDD.n2706 7.39606
R23551 VDD.n4222 VDD.n4221 7.39606
R23552 VDD.n4221 VDD.n2696 7.39606
R23553 VDD.n4232 VDD.n4231 7.39606
R23554 VDD.n4231 VDD.n2685 7.39606
R23555 VDD.n4242 VDD.n4241 7.39606
R23556 VDD.n4241 VDD.n2672 7.39606
R23557 VDD.n4261 VDD.n2644 7.39606
R23558 VDD.n4261 VDD.n2646 7.39606
R23559 VDD.n4276 VDD.n4275 7.39606
R23560 VDD.n4275 VDD.n2630 7.39606
R23561 VDD.n4286 VDD.n4285 7.39606
R23562 VDD.n4285 VDD.n2618 7.39606
R23563 VDD.n4296 VDD.n4295 7.39606
R23564 VDD.n4295 VDD.n2605 7.39606
R23565 VDD.n4306 VDD.n4305 7.39606
R23566 VDD.n4305 VDD.n2595 7.39606
R23567 VDD.n4266 VDD.n4265 7.39606
R23568 VDD.n4265 VDD.n2639 7.39606
R23569 VDD.n4077 VDD.n4076 7.39606
R23570 VDD.n4076 VDD.n4067 7.39606
R23571 VDD.n4087 VDD.n4086 7.39606
R23572 VDD.n4086 VDD.n2842 7.39606
R23573 VDD.n4097 VDD.n4096 7.39606
R23574 VDD.n4096 VDD.n2832 7.39606
R23575 VDD.n4107 VDD.n4106 7.39606
R23576 VDD.n4106 VDD.n2821 7.39606
R23577 VDD.n4117 VDD.n4116 7.39606
R23578 VDD.n4116 VDD.n2808 7.39606
R23579 VDD.n4136 VDD.n2780 7.39606
R23580 VDD.n4136 VDD.n2782 7.39606
R23581 VDD.n4151 VDD.n4150 7.39606
R23582 VDD.n4150 VDD.n2766 7.39606
R23583 VDD.n4161 VDD.n4160 7.39606
R23584 VDD.n4160 VDD.n2754 7.39606
R23585 VDD.n4171 VDD.n4170 7.39606
R23586 VDD.n4170 VDD.n2741 7.39606
R23587 VDD.n4181 VDD.n4180 7.39606
R23588 VDD.n4180 VDD.n2731 7.39606
R23589 VDD.n4141 VDD.n4140 7.39606
R23590 VDD.n4140 VDD.n2775 7.39606
R23591 VDD.n3952 VDD.n3951 7.39606
R23592 VDD.n3951 VDD.n3942 7.39606
R23593 VDD.n3962 VDD.n3961 7.39606
R23594 VDD.n3961 VDD.n2978 7.39606
R23595 VDD.n3972 VDD.n3971 7.39606
R23596 VDD.n3971 VDD.n2968 7.39606
R23597 VDD.n3982 VDD.n3981 7.39606
R23598 VDD.n3981 VDD.n2957 7.39606
R23599 VDD.n3992 VDD.n3991 7.39606
R23600 VDD.n3991 VDD.n2944 7.39606
R23601 VDD.n4011 VDD.n2916 7.39606
R23602 VDD.n4011 VDD.n2918 7.39606
R23603 VDD.n4026 VDD.n4025 7.39606
R23604 VDD.n4025 VDD.n2902 7.39606
R23605 VDD.n4036 VDD.n4035 7.39606
R23606 VDD.n4035 VDD.n2890 7.39606
R23607 VDD.n4046 VDD.n4045 7.39606
R23608 VDD.n4045 VDD.n2877 7.39606
R23609 VDD.n4056 VDD.n4055 7.39606
R23610 VDD.n4055 VDD.n2867 7.39606
R23611 VDD.n4016 VDD.n4015 7.39606
R23612 VDD.n4015 VDD.n2911 7.39606
R23613 VDD.n3604 VDD.n3603 7.39606
R23614 VDD.n3603 VDD.n3282 7.39606
R23615 VDD.n3616 VDD.n3266 7.39606
R23616 VDD.n3616 VDD.n3268 7.39606
R23617 VDD.n3594 VDD.n3593 7.39606
R23618 VDD.n3593 VDD.n3291 7.39606
R23619 VDD.n3827 VDD.n3826 7.39606
R23620 VDD.n3826 VDD.n3817 7.39606
R23621 VDD.n3837 VDD.n3836 7.39606
R23622 VDD.n3836 VDD.n3804 7.39606
R23623 VDD.n3847 VDD.n3846 7.39606
R23624 VDD.n3846 VDD.n3794 7.39606
R23625 VDD.n3857 VDD.n3856 7.39606
R23626 VDD.n3856 VDD.n3783 7.39606
R23627 VDD.n3867 VDD.n3866 7.39606
R23628 VDD.n3866 VDD.n3770 7.39606
R23629 VDD.n3886 VDD.n3742 7.39606
R23630 VDD.n3886 VDD.n3744 7.39606
R23631 VDD.n3901 VDD.n3900 7.39606
R23632 VDD.n3900 VDD.n3728 7.39606
R23633 VDD.n3911 VDD.n3910 7.39606
R23634 VDD.n3910 VDD.n3026 7.39606
R23635 VDD.n3921 VDD.n3920 7.39606
R23636 VDD.n3920 VDD.n3013 7.39606
R23637 VDD.n3931 VDD.n3930 7.39606
R23638 VDD.n3930 VDD.n3003 7.39606
R23639 VDD.n3891 VDD.n3890 7.39606
R23640 VDD.n3890 VDD.n3737 7.39606
R23641 VDD.n147 VDD.t213 7.31106
R23642 VDD.t370 VDD.n142 7.31106
R23643 VDD.n161 VDD.t654 7.31106
R23644 VDD.t846 VDD.n126 7.31106
R23645 VDD.n182 VDD.t619 7.31106
R23646 VDD.t128 VDD.n117 7.31106
R23647 VDD.n196 VDD.t976 7.31106
R23648 VDD.t170 VDD.n101 7.31106
R23649 VDD.n217 VDD.t838 7.31106
R23650 VDD.t921 VDD.n92 7.31106
R23651 VDD.n231 VDD.t957 7.31106
R23652 VDD.t878 VDD.n76 7.31106
R23653 VDD.n252 VDD.t351 7.31106
R23654 VDD.t646 VDD.n67 7.31106
R23655 VDD.n266 VDD.t77 7.31106
R23656 VDD.t629 VDD.n51 7.31106
R23657 VDD.n6996 VDD.t939 7.31106
R23658 VDD.t968 VDD.n6991 7.31106
R23659 VDD.n7010 VDD.t1036 7.31106
R23660 VDD.t931 VDD.n6975 7.31106
R23661 VDD.n7031 VDD.t126 7.31106
R23662 VDD.t71 VDD.n6966 7.31106
R23663 VDD.n7045 VDD.t1012 7.31106
R23664 VDD.t189 VDD.n6950 7.31106
R23665 VDD.n7066 VDD.t798 7.31106
R23666 VDD.t791 VDD.n6941 7.31106
R23667 VDD.n7080 VDD.t1040 7.31106
R23668 VDD.t583 VDD.n6925 7.31106
R23669 VDD.n7101 VDD.t773 7.31106
R23670 VDD.t276 VDD.n6916 7.31106
R23671 VDD.n7115 VDD.t1008 7.31106
R23672 VDD.n6899 VDD.t301 7.31106
R23673 VDD.t854 VDD.n3428 7.31106
R23674 VDD.n3445 VDD.t985 7.31106
R23675 VDD.t810 VDD.n3466 7.31106
R23676 VDD.n3482 VDD.t131 7.31106
R23677 VDD.t271 VDD.n3321 7.31106
R23678 VDD.n3334 VDD.t884 7.31106
R23679 VDD.t996 VDD.n3523 7.31106
R23680 VDD.n3540 VDD.t122 7.31106
R23681 VDD.t408 VDD.n3560 7.31106
R23682 VDD.n3576 VDD.t137 7.31106
R23683 VDD.t782 VDD.n3377 7.31106
R23684 VDD.n3390 VDD.t206 7.31106
R23685 VDD VDD.n6763 7.20159
R23686 VDD VDD.n6640 7.20159
R23687 VDD VDD.n6517 7.20159
R23688 VDD VDD.n6394 7.20159
R23689 VDD VDD.n6271 7.20159
R23690 VDD VDD.n6148 7.20159
R23691 VDD.n3154 VDD.n3153 6.96517
R23692 VDD.n3218 VDD.n3217 6.96517
R23693 VDD.n3115 VDD.n3114 6.96517
R23694 VDD.n3369 VDD.n3368 6.96517
R23695 VDD.n3076 VDD.n3075 6.96517
R23696 VDD.n3663 VDD.n3662 6.96517
R23697 VDD.n3056 VDD.n3055 6.96517
R23698 VDD.n3134 VDD.n3133 6.96517
R23699 VDD VDD.n3940 6.79126
R23700 VDD VDD.n4065 6.79126
R23701 VDD VDD.n4190 6.79126
R23702 VDD VDD.n4315 6.79126
R23703 VDD VDD.n4440 6.79126
R23704 VDD VDD.n4565 6.79126
R23705 VDD VDD.n4690 6.79126
R23706 VDD.n322 VDD.n306 6.37981
R23707 VDD.n309 VDD.n306 6.37981
R23708 VDD.n3516 VDD.n3515 5.59193
R23709 VDD.n3686 VDD.n3056 5.50827
R23710 VDD.n3300 VDD 4.96789
R23711 VDD.n6887 VDD.n6886 4.92985
R23712 VDD.n7131 VDD.n4815 4.51952
R23713 VDD.n3153 VDD.n3152 4.5005
R23714 VDD.n3170 VDD.n3169 4.5005
R23715 VDD.n3217 VDD.n3216 4.5005
R23716 VDD.n3234 VDD.n3233 4.5005
R23717 VDD.n3114 VDD.n3113 4.5005
R23718 VDD.n3258 VDD.n3257 4.5005
R23719 VDD.n3368 VDD.n3367 4.5005
R23720 VDD.n3635 VDD.n3634 4.5005
R23721 VDD.n3075 VDD.n3074 4.5005
R23722 VDD.n3092 VDD.n3091 4.5005
R23723 VDD.n3662 VDD.n3661 4.5005
R23724 VDD.n3679 VDD.n3678 4.5005
R23725 VDD.n3055 VDD.n3054 4.5005
R23726 VDD.n3702 VDD.n3701 4.5005
R23727 VDD.n3133 VDD.n3132 4.5005
R23728 VDD.n3189 VDD.n3188 4.5005
R23729 VDD.n3723 VDD.n3722 4.5005
R23730 VDD.n1641 VDD.n1381 4.44435
R23731 VDD.n3501 VDD.n3500 4.44122
R23732 VDD.n3036 VDD 4.43528
R23733 VDD.n2900 VDD 4.43528
R23734 VDD.n2764 VDD 4.43528
R23735 VDD.n2628 VDD 4.43528
R23736 VDD.n2492 VDD 4.43528
R23737 VDD.n2356 VDD 4.43528
R23738 VDD.n2220 VDD 4.43528
R23739 VDD.n2084 VDD 4.43528
R23740 VDD.n1948 VDD 4.43528
R23741 VDD.n42 VDD.t867 4.27344
R23742 VDD.t863 VDD.n1647 4.27344
R23743 VDD.t609 VDD.n1387 4.27344
R23744 VDD.t961 VDD.n1127 4.27344
R23745 VDD.t865 VDD.n867 4.27344
R23746 VDD.t605 VDD.n607 4.27344
R23747 VDD.t963 VDD.n347 4.27344
R23748 VDD.t607 VDD.n7263 4.27344
R23749 VDD.t649 VDD.n1907 4.27344
R23750 VDD.n6022 VDD.t888 4.27344
R23751 VDD.n5886 VDD.t881 4.27344
R23752 VDD.n5750 VDD.t916 4.27344
R23753 VDD.n5614 VDD.t621 4.27344
R23754 VDD.n5478 VDD.t23 4.27344
R23755 VDD.n5342 VDD.t840 4.27344
R23756 VDD.n5206 VDD.t919 4.27344
R23757 VDD.n5068 VDD.t574 4.27344
R23758 VDD.t303 VDD.n2043 4.27344
R23759 VDD.t65 VDD.n2179 4.27344
R23760 VDD.t25 VDD.n2315 4.27344
R23761 VDD.t796 VDD.n2451 4.27344
R23762 VDD.t764 VDD.n2587 4.27344
R23763 VDD.t124 VDD.n2723 4.27344
R23764 VDD.t153 VDD.n2859 4.27344
R23765 VDD.t941 VDD.n2995 4.27344
R23766 VDD.n3198 VDD.n3154 4.23927
R23767 VDD.n3239 VDD.n3218 4.23927
R23768 VDD.n3242 VDD.n3115 4.23927
R23769 VDD.n3370 VDD.n3369 4.23927
R23770 VDD.n3643 VDD.n3076 4.23927
R23771 VDD.n3684 VDD.n3663 4.23927
R23772 VDD.n3135 VDD.n3134 4.23927
R23773 VDD.t401 VDD.n293 4.14288
R23774 VDD.n3422 VDD 3.73292
R23775 VDD.n3460 VDD 3.73292
R23776 VDD.n3514 VDD 3.73292
R23777 VDD.n3517 VDD 3.73292
R23778 VDD.n3554 VDD 3.73292
R23779 VDD.n3419 VDD 3.73292
R23780 VDD.n3618 VDD 3.73292
R23781 VDD.n3420 VDD.n3370 3.53255
R23782 VDD.n3194 VDD.n3193 3.473
R23783 VDD.n3685 VDD.n3684 3.4105
R23784 VDD.n3644 VDD.n3643 3.4105
R23785 VDD.n3370 VDD.n3057 3.4105
R23786 VDD.n3242 VDD.n3241 3.4105
R23787 VDD.n3240 VDD.n3239 3.4105
R23788 VDD.n3199 VDD.n3198 3.4105
R23789 VDD.n3197 VDD.n3196 3.4105
R23790 VDD.n3238 VDD.n3096 3.4105
R23791 VDD.n3263 VDD.n3262 3.4105
R23792 VDD.n3640 VDD.n3639 3.4105
R23793 VDD.n3642 VDD.n3641 3.4105
R23794 VDD.n3683 VDD.n3037 3.4105
R23795 VDD.n3707 VDD.n3706 3.4105
R23796 VDD.n325 VDD.n286 3.29941
R23797 VDD.n4954 VDD.n4953 3.15974
R23798 VDD.n3639 VDD.n3619 3.08605
R23799 VDD.n308 VDD.n307 3.08383
R23800 VDD.n318 VDD.n308 3.08383
R23801 VDD.n3739 VDD 3.063
R23802 VDD.n2913 VDD 3.063
R23803 VDD.n2777 VDD 3.063
R23804 VDD.n2641 VDD 3.063
R23805 VDD.n2505 VDD 3.063
R23806 VDD.n2369 VDD 3.063
R23807 VDD.n2233 VDD 3.063
R23808 VDD.n2097 VDD 3.063
R23809 VDD.n1961 VDD 3.063
R23810 VDD.n3619 VDD.n3264 2.797
R23811 VDD.n3516 VDD.n3264 2.79387
R23812 VDD.n3515 VDD.n3314 2.79387
R23813 VDD.n3421 VDD.n3314 2.79387
R23814 VDD.n861 VDD.n601 2.7876
R23815 VDD.n1121 VDD.n861 2.7876
R23816 VDD.n1381 VDD.n1121 2.7876
R23817 VDD.n1901 VDD.n1641 2.7876
R23818 VDD.n7518 VDD.n1901 2.7876
R23819 VDD.n7518 VDD.n7517 2.7876
R23820 VDD.n6898 VDD.n6897 2.73583
R23821 VDD.n7128 VDD 2.60011
R23822 VDD.n323 VDD.t566 2.59611
R23823 VDD.n3421 VDD.n3420 2.44842
R23824 VDD VDD.n324 2.38637
R23825 VDD.n1899 VDD.n1898 2.3255
R23826 VDD.n1890 VDD.n1654 2.3255
R23827 VDD.n1880 VDD.n1664 2.3255
R23828 VDD.n1870 VDD.n1677 2.3255
R23829 VDD.n1860 VDD.n1688 2.3255
R23830 VDD.n1850 VDD.n1698 2.3255
R23831 VDD.n1840 VDD.n1711 2.3255
R23832 VDD.n1725 VDD.n1718 2.3255
R23833 VDD.n1823 VDD.n1726 2.3255
R23834 VDD.n1813 VDD.n1739 2.3255
R23835 VDD.n1803 VDD.n1750 2.3255
R23836 VDD.n1793 VDD.n1760 2.3255
R23837 VDD.n1783 VDD.n1773 2.3255
R23838 VDD.n1639 VDD.n1638 2.3255
R23839 VDD.n1630 VDD.n1394 2.3255
R23840 VDD.n1620 VDD.n1404 2.3255
R23841 VDD.n1610 VDD.n1417 2.3255
R23842 VDD.n1600 VDD.n1428 2.3255
R23843 VDD.n1590 VDD.n1438 2.3255
R23844 VDD.n1580 VDD.n1451 2.3255
R23845 VDD.n1465 VDD.n1458 2.3255
R23846 VDD.n1563 VDD.n1466 2.3255
R23847 VDD.n1553 VDD.n1479 2.3255
R23848 VDD.n1543 VDD.n1490 2.3255
R23849 VDD.n1533 VDD.n1500 2.3255
R23850 VDD.n1523 VDD.n1513 2.3255
R23851 VDD.n1379 VDD.n1378 2.3255
R23852 VDD.n1370 VDD.n1134 2.3255
R23853 VDD.n1360 VDD.n1144 2.3255
R23854 VDD.n1350 VDD.n1157 2.3255
R23855 VDD.n1340 VDD.n1168 2.3255
R23856 VDD.n1330 VDD.n1178 2.3255
R23857 VDD.n1320 VDD.n1191 2.3255
R23858 VDD.n1205 VDD.n1198 2.3255
R23859 VDD.n1303 VDD.n1206 2.3255
R23860 VDD.n1293 VDD.n1219 2.3255
R23861 VDD.n1283 VDD.n1230 2.3255
R23862 VDD.n1273 VDD.n1240 2.3255
R23863 VDD.n1263 VDD.n1253 2.3255
R23864 VDD.n1119 VDD.n1118 2.3255
R23865 VDD.n1110 VDD.n874 2.3255
R23866 VDD.n1100 VDD.n884 2.3255
R23867 VDD.n1090 VDD.n897 2.3255
R23868 VDD.n1080 VDD.n908 2.3255
R23869 VDD.n1070 VDD.n918 2.3255
R23870 VDD.n1060 VDD.n931 2.3255
R23871 VDD.n945 VDD.n938 2.3255
R23872 VDD.n1043 VDD.n946 2.3255
R23873 VDD.n1033 VDD.n959 2.3255
R23874 VDD.n1023 VDD.n970 2.3255
R23875 VDD.n1013 VDD.n980 2.3255
R23876 VDD.n1003 VDD.n993 2.3255
R23877 VDD.n859 VDD.n858 2.3255
R23878 VDD.n850 VDD.n614 2.3255
R23879 VDD.n840 VDD.n624 2.3255
R23880 VDD.n830 VDD.n637 2.3255
R23881 VDD.n820 VDD.n648 2.3255
R23882 VDD.n810 VDD.n658 2.3255
R23883 VDD.n800 VDD.n671 2.3255
R23884 VDD.n685 VDD.n678 2.3255
R23885 VDD.n783 VDD.n686 2.3255
R23886 VDD.n773 VDD.n699 2.3255
R23887 VDD.n763 VDD.n710 2.3255
R23888 VDD.n753 VDD.n720 2.3255
R23889 VDD.n743 VDD.n733 2.3255
R23890 VDD.n599 VDD.n598 2.3255
R23891 VDD.n590 VDD.n354 2.3255
R23892 VDD.n580 VDD.n364 2.3255
R23893 VDD.n570 VDD.n377 2.3255
R23894 VDD.n560 VDD.n388 2.3255
R23895 VDD.n550 VDD.n398 2.3255
R23896 VDD.n540 VDD.n411 2.3255
R23897 VDD.n425 VDD.n418 2.3255
R23898 VDD.n523 VDD.n426 2.3255
R23899 VDD.n513 VDD.n439 2.3255
R23900 VDD.n503 VDD.n450 2.3255
R23901 VDD.n493 VDD.n460 2.3255
R23902 VDD.n483 VDD.n473 2.3255
R23903 VDD.n284 VDD.n283 2.3255
R23904 VDD.n58 VDD.n54 2.3255
R23905 VDD.n265 VDD.n264 2.3255
R23906 VDD.n263 VDD.n262 2.3255
R23907 VDD.n251 VDD.n250 2.3255
R23908 VDD.n249 VDD.n248 2.3255
R23909 VDD.n83 VDD.n79 2.3255
R23910 VDD.n230 VDD.n229 2.3255
R23911 VDD.n228 VDD.n227 2.3255
R23912 VDD.n216 VDD.n215 2.3255
R23913 VDD.n214 VDD.n213 2.3255
R23914 VDD.n108 VDD.n104 2.3255
R23915 VDD.n195 VDD.n194 2.3255
R23916 VDD.n193 VDD.n192 2.3255
R23917 VDD.n181 VDD.n180 2.3255
R23918 VDD.n179 VDD.n178 2.3255
R23919 VDD.n133 VDD.n129 2.3255
R23920 VDD.n160 VDD.n159 2.3255
R23921 VDD.n158 VDD.n157 2.3255
R23922 VDD.n146 VDD.n145 2.3255
R23923 VDD.n7515 VDD.n7514 2.3255
R23924 VDD.n7506 VDD.n7270 2.3255
R23925 VDD.n7496 VDD.n7280 2.3255
R23926 VDD.n7486 VDD.n7293 2.3255
R23927 VDD.n7476 VDD.n7304 2.3255
R23928 VDD.n7466 VDD.n7314 2.3255
R23929 VDD.n7456 VDD.n7327 2.3255
R23930 VDD.n7341 VDD.n7334 2.3255
R23931 VDD.n7439 VDD.n7342 2.3255
R23932 VDD.n7429 VDD.n7355 2.3255
R23933 VDD.n7419 VDD.n7366 2.3255
R23934 VDD.n7409 VDD.n7376 2.3255
R23935 VDD.n7399 VDD.n7389 2.3255
R23936 VDD.n7114 VDD.n7113 2.3255
R23937 VDD.n7112 VDD.n7111 2.3255
R23938 VDD.n7100 VDD.n7099 2.3255
R23939 VDD.n7098 VDD.n7097 2.3255
R23940 VDD.n6932 VDD.n6928 2.3255
R23941 VDD.n7079 VDD.n7078 2.3255
R23942 VDD.n7077 VDD.n7076 2.3255
R23943 VDD.n7065 VDD.n7064 2.3255
R23944 VDD.n7063 VDD.n7062 2.3255
R23945 VDD.n6957 VDD.n6953 2.3255
R23946 VDD.n7044 VDD.n7043 2.3255
R23947 VDD.n7042 VDD.n7041 2.3255
R23948 VDD.n7030 VDD.n7029 2.3255
R23949 VDD.n7028 VDD.n7027 2.3255
R23950 VDD.n6982 VDD.n6978 2.3255
R23951 VDD.n7009 VDD.n7008 2.3255
R23952 VDD.n7007 VDD.n7006 2.3255
R23953 VDD.n6995 VDD.n6994 2.3255
R23954 VDD.n7127 VDD.n7126 2.3255
R23955 VDD.n6886 VDD.n6885 2.3255
R23956 VDD.n6872 VDD.n5092 2.3255
R23957 VDD.n6862 VDD.n5102 2.3255
R23958 VDD.n6852 VDD.n5113 2.3255
R23959 VDD.n6842 VDD.n5126 2.3255
R23960 VDD.n5139 VDD.n5133 2.3255
R23961 VDD.n6825 VDD.n5141 2.3255
R23962 VDD.n6815 VDD.n5154 2.3255
R23963 VDD.n6805 VDD.n5164 2.3255
R23964 VDD.n6795 VDD.n5175 2.3255
R23965 VDD.n6785 VDD.n5188 2.3255
R23966 VDD.n6775 VDD.n5198 2.3255
R23967 VDD.n6766 VDD.n6765 2.3255
R23968 VDD.n6763 VDD.n6762 2.3255
R23969 VDD.n6749 VDD.n5228 2.3255
R23970 VDD.n6739 VDD.n5238 2.3255
R23971 VDD.n6729 VDD.n5249 2.3255
R23972 VDD.n6719 VDD.n5262 2.3255
R23973 VDD.n5275 VDD.n5269 2.3255
R23974 VDD.n6702 VDD.n5277 2.3255
R23975 VDD.n6692 VDD.n5290 2.3255
R23976 VDD.n6682 VDD.n5300 2.3255
R23977 VDD.n6672 VDD.n5311 2.3255
R23978 VDD.n6662 VDD.n5324 2.3255
R23979 VDD.n6652 VDD.n5334 2.3255
R23980 VDD.n6643 VDD.n6642 2.3255
R23981 VDD.n6640 VDD.n6639 2.3255
R23982 VDD.n6626 VDD.n5364 2.3255
R23983 VDD.n6616 VDD.n5374 2.3255
R23984 VDD.n6606 VDD.n5385 2.3255
R23985 VDD.n6596 VDD.n5398 2.3255
R23986 VDD.n5411 VDD.n5405 2.3255
R23987 VDD.n6579 VDD.n5413 2.3255
R23988 VDD.n6569 VDD.n5426 2.3255
R23989 VDD.n6559 VDD.n5436 2.3255
R23990 VDD.n6549 VDD.n5447 2.3255
R23991 VDD.n6539 VDD.n5460 2.3255
R23992 VDD.n6529 VDD.n5470 2.3255
R23993 VDD.n6520 VDD.n6519 2.3255
R23994 VDD.n6517 VDD.n6516 2.3255
R23995 VDD.n6503 VDD.n5500 2.3255
R23996 VDD.n6493 VDD.n5510 2.3255
R23997 VDD.n6483 VDD.n5521 2.3255
R23998 VDD.n6473 VDD.n5534 2.3255
R23999 VDD.n5547 VDD.n5541 2.3255
R24000 VDD.n6456 VDD.n5549 2.3255
R24001 VDD.n6446 VDD.n5562 2.3255
R24002 VDD.n6436 VDD.n5572 2.3255
R24003 VDD.n6426 VDD.n5583 2.3255
R24004 VDD.n6416 VDD.n5596 2.3255
R24005 VDD.n6406 VDD.n5606 2.3255
R24006 VDD.n6397 VDD.n6396 2.3255
R24007 VDD.n6394 VDD.n6393 2.3255
R24008 VDD.n6380 VDD.n5636 2.3255
R24009 VDD.n6370 VDD.n5646 2.3255
R24010 VDD.n6360 VDD.n5657 2.3255
R24011 VDD.n6350 VDD.n5670 2.3255
R24012 VDD.n5683 VDD.n5677 2.3255
R24013 VDD.n6333 VDD.n5685 2.3255
R24014 VDD.n6323 VDD.n5698 2.3255
R24015 VDD.n6313 VDD.n5708 2.3255
R24016 VDD.n6303 VDD.n5719 2.3255
R24017 VDD.n6293 VDD.n5732 2.3255
R24018 VDD.n6283 VDD.n5742 2.3255
R24019 VDD.n6274 VDD.n6273 2.3255
R24020 VDD.n6271 VDD.n6270 2.3255
R24021 VDD.n6257 VDD.n5772 2.3255
R24022 VDD.n6247 VDD.n5782 2.3255
R24023 VDD.n6237 VDD.n5793 2.3255
R24024 VDD.n6227 VDD.n5806 2.3255
R24025 VDD.n5819 VDD.n5813 2.3255
R24026 VDD.n6210 VDD.n5821 2.3255
R24027 VDD.n6200 VDD.n5834 2.3255
R24028 VDD.n6190 VDD.n5844 2.3255
R24029 VDD.n6180 VDD.n5855 2.3255
R24030 VDD.n6170 VDD.n5868 2.3255
R24031 VDD.n6160 VDD.n5878 2.3255
R24032 VDD.n6151 VDD.n6150 2.3255
R24033 VDD.n6148 VDD.n6147 2.3255
R24034 VDD.n6134 VDD.n5908 2.3255
R24035 VDD.n6124 VDD.n5918 2.3255
R24036 VDD.n6114 VDD.n5929 2.3255
R24037 VDD.n6104 VDD.n5942 2.3255
R24038 VDD.n5955 VDD.n5949 2.3255
R24039 VDD.n6087 VDD.n5957 2.3255
R24040 VDD.n6077 VDD.n5970 2.3255
R24041 VDD.n6067 VDD.n5980 2.3255
R24042 VDD.n6057 VDD.n5991 2.3255
R24043 VDD.n6047 VDD.n6004 2.3255
R24044 VDD.n6037 VDD.n6014 2.3255
R24045 VDD.n6028 VDD.n6027 2.3255
R24046 VDD.n4964 VDD.n4933 2.3255
R24047 VDD.n4974 VDD.n4923 2.3255
R24048 VDD.n4984 VDD.n4912 2.3255
R24049 VDD.n4994 VDD.n4899 2.3255
R24050 VDD.n4898 VDD.n4890 2.3255
R24051 VDD.n5011 VDD.n4884 2.3255
R24052 VDD.n5021 VDD.n4871 2.3255
R24053 VDD.n5031 VDD.n4861 2.3255
R24054 VDD.n5041 VDD.n4850 2.3255
R24055 VDD.n5051 VDD.n4837 2.3255
R24056 VDD.n5061 VDD.n4827 2.3255
R24057 VDD.n5072 VDD.n5071 2.3255
R24058 VDD.n3435 VDD.n3434 2.3255
R24059 VDD.n3439 VDD.n3438 2.3255
R24060 VDD.n3473 VDD.n3472 2.3255
R24061 VDD.n3476 VDD.n3475 2.3255
R24062 VDD.n3513 VDD.n3512 2.3255
R24063 VDD.n3505 VDD.n3504 2.3255
R24064 VDD.n3530 VDD.n3529 2.3255
R24065 VDD.n3534 VDD.n3533 2.3255
R24066 VDD.n3567 VDD.n3566 2.3255
R24067 VDD.n3570 VDD.n3569 2.3255
R24068 VDD.n3418 VDD.n3417 2.3255
R24069 VDD.n3410 VDD.n3409 2.3255
R24070 VDD.n3394 VDD.n3393 2.3255
R24071 VDD.n3449 VDD.n3448 2.3255
R24072 VDD.n3486 VDD.n3485 2.3255
R24073 VDD.n3338 VDD.n3337 2.3255
R24074 VDD.n3544 VDD.n3543 2.3255
R24075 VDD.n3580 VDD.n3579 2.3255
R24076 VDD.n3593 VDD.n3592 2.3255
R24077 VDD.n3617 VDD.n3616 2.3255
R24078 VDD.n3603 VDD.n3281 2.3255
R24079 VDD.n3890 VDD.n3889 2.3255
R24080 VDD.n3887 VDD.n3886 2.3255
R24081 VDD.n3768 VDD.n3761 2.3255
R24082 VDD.n3866 VDD.n3769 2.3255
R24083 VDD.n3856 VDD.n3782 2.3255
R24084 VDD.n3846 VDD.n3793 2.3255
R24085 VDD.n3836 VDD.n3803 2.3255
R24086 VDD.n3826 VDD.n3816 2.3255
R24087 VDD.n3900 VDD.n3727 2.3255
R24088 VDD.n4015 VDD.n4014 2.3255
R24089 VDD.n4012 VDD.n4011 2.3255
R24090 VDD.n2942 VDD.n2935 2.3255
R24091 VDD.n3991 VDD.n2943 2.3255
R24092 VDD.n3981 VDD.n2956 2.3255
R24093 VDD.n3971 VDD.n2967 2.3255
R24094 VDD.n3961 VDD.n2977 2.3255
R24095 VDD.n3951 VDD.n3941 2.3255
R24096 VDD.n3939 VDD.n3938 2.3255
R24097 VDD.n3930 VDD.n3002 2.3255
R24098 VDD.n3920 VDD.n3012 2.3255
R24099 VDD.n3910 VDD.n3025 2.3255
R24100 VDD.n4025 VDD.n2901 2.3255
R24101 VDD.n4140 VDD.n4139 2.3255
R24102 VDD.n4137 VDD.n4136 2.3255
R24103 VDD.n2806 VDD.n2799 2.3255
R24104 VDD.n4116 VDD.n2807 2.3255
R24105 VDD.n4106 VDD.n2820 2.3255
R24106 VDD.n4096 VDD.n2831 2.3255
R24107 VDD.n4086 VDD.n2841 2.3255
R24108 VDD.n4076 VDD.n4066 2.3255
R24109 VDD.n4064 VDD.n4063 2.3255
R24110 VDD.n4055 VDD.n2866 2.3255
R24111 VDD.n4045 VDD.n2876 2.3255
R24112 VDD.n4035 VDD.n2889 2.3255
R24113 VDD.n4150 VDD.n2765 2.3255
R24114 VDD.n4265 VDD.n4264 2.3255
R24115 VDD.n4262 VDD.n4261 2.3255
R24116 VDD.n2670 VDD.n2663 2.3255
R24117 VDD.n4241 VDD.n2671 2.3255
R24118 VDD.n4231 VDD.n2684 2.3255
R24119 VDD.n4221 VDD.n2695 2.3255
R24120 VDD.n4211 VDD.n2705 2.3255
R24121 VDD.n4201 VDD.n4191 2.3255
R24122 VDD.n4189 VDD.n4188 2.3255
R24123 VDD.n4180 VDD.n2730 2.3255
R24124 VDD.n4170 VDD.n2740 2.3255
R24125 VDD.n4160 VDD.n2753 2.3255
R24126 VDD.n4275 VDD.n2629 2.3255
R24127 VDD.n4390 VDD.n4389 2.3255
R24128 VDD.n4387 VDD.n4386 2.3255
R24129 VDD.n2534 VDD.n2527 2.3255
R24130 VDD.n4366 VDD.n2535 2.3255
R24131 VDD.n4356 VDD.n2548 2.3255
R24132 VDD.n4346 VDD.n2559 2.3255
R24133 VDD.n4336 VDD.n2569 2.3255
R24134 VDD.n4326 VDD.n4316 2.3255
R24135 VDD.n4314 VDD.n4313 2.3255
R24136 VDD.n4305 VDD.n2594 2.3255
R24137 VDD.n4295 VDD.n2604 2.3255
R24138 VDD.n4285 VDD.n2617 2.3255
R24139 VDD.n4400 VDD.n2493 2.3255
R24140 VDD.n4515 VDD.n4514 2.3255
R24141 VDD.n4512 VDD.n4511 2.3255
R24142 VDD.n2398 VDD.n2391 2.3255
R24143 VDD.n4491 VDD.n2399 2.3255
R24144 VDD.n4481 VDD.n2412 2.3255
R24145 VDD.n4471 VDD.n2423 2.3255
R24146 VDD.n4461 VDD.n2433 2.3255
R24147 VDD.n4451 VDD.n4441 2.3255
R24148 VDD.n4439 VDD.n4438 2.3255
R24149 VDD.n4430 VDD.n2458 2.3255
R24150 VDD.n4420 VDD.n2468 2.3255
R24151 VDD.n4410 VDD.n2481 2.3255
R24152 VDD.n4525 VDD.n2357 2.3255
R24153 VDD.n4640 VDD.n4639 2.3255
R24154 VDD.n4637 VDD.n4636 2.3255
R24155 VDD.n2262 VDD.n2255 2.3255
R24156 VDD.n4616 VDD.n2263 2.3255
R24157 VDD.n4606 VDD.n2276 2.3255
R24158 VDD.n4596 VDD.n2287 2.3255
R24159 VDD.n4586 VDD.n2297 2.3255
R24160 VDD.n4576 VDD.n4566 2.3255
R24161 VDD.n4564 VDD.n4563 2.3255
R24162 VDD.n4555 VDD.n2322 2.3255
R24163 VDD.n4545 VDD.n2332 2.3255
R24164 VDD.n4535 VDD.n2345 2.3255
R24165 VDD.n4650 VDD.n2221 2.3255
R24166 VDD.n4765 VDD.n4764 2.3255
R24167 VDD.n4762 VDD.n4761 2.3255
R24168 VDD.n2126 VDD.n2119 2.3255
R24169 VDD.n4741 VDD.n2127 2.3255
R24170 VDD.n4731 VDD.n2140 2.3255
R24171 VDD.n4721 VDD.n2151 2.3255
R24172 VDD.n4711 VDD.n2161 2.3255
R24173 VDD.n4701 VDD.n4691 2.3255
R24174 VDD.n4689 VDD.n4688 2.3255
R24175 VDD.n4680 VDD.n2186 2.3255
R24176 VDD.n4670 VDD.n2196 2.3255
R24177 VDD.n4660 VDD.n2209 2.3255
R24178 VDD.n4775 VDD.n2085 2.3255
R24179 VDD.n4814 VDD.n4813 2.3255
R24180 VDD.n4805 VDD.n2050 2.3255
R24181 VDD.n4795 VDD.n2060 2.3255
R24182 VDD.n4785 VDD.n2073 2.3255
R24183 VDD.n7206 VDD.n7205 2.3255
R24184 VDD.n7203 VDD.n7202 2.3255
R24185 VDD.n1990 VDD.n1983 2.3255
R24186 VDD.n7182 VDD.n1991 2.3255
R24187 VDD.n7172 VDD.n2004 2.3255
R24188 VDD.n7162 VDD.n2015 2.3255
R24189 VDD.n7152 VDD.n2025 2.3255
R24190 VDD.n7142 VDD.n7132 2.3255
R24191 VDD.n7216 VDD.n1949 2.3255
R24192 VDD.n7255 VDD.n7254 2.3255
R24193 VDD.n7246 VDD.n1914 2.3255
R24194 VDD.n7236 VDD.n1924 2.3255
R24195 VDD.n7226 VDD.n1937 2.3255
R24196 VDD.n7522 VDD.n7521 2.3255
R24197 VDD.n7531 VDD.n35 2.3255
R24198 VDD.n7541 VDD.n25 2.3255
R24199 VDD.n7551 VDD.n0 2.3255
R24200 VDD.n7731 VDD.n7730 2.3255
R24201 VDD.n7717 VDD.n1 2.3255
R24202 VDD.n7707 VDD.n7578 2.3255
R24203 VDD.n7592 VDD.n7585 2.3255
R24204 VDD.n7690 VDD.n7593 2.3255
R24205 VDD.n7680 VDD.n7606 2.3255
R24206 VDD.n7670 VDD.n7617 2.3255
R24207 VDD.n7660 VDD.n7627 2.3255
R24208 VDD.n7650 VDD.n7640 2.3255
R24209 VDD.n6887 VDD 2.22333
R24210 VDD VDD.n7131 2.22333
R24211 VDD.n314 VDD.n313 2.05606
R24212 VDD.n313 VDD.n310 2.05606
R24213 VDD.n601 VDD.n341 1.71757
R24214 VDD.n324 VDD 1.71534
R24215 VDD.n1664 VDD.n1654 1.66898
R24216 VDD.n1698 VDD.n1688 1.66898
R24217 VDD.n1760 VDD.n1750 1.66898
R24218 VDD.n1404 VDD.n1394 1.66898
R24219 VDD.n1438 VDD.n1428 1.66898
R24220 VDD.n1500 VDD.n1490 1.66898
R24221 VDD.n1144 VDD.n1134 1.66898
R24222 VDD.n1178 VDD.n1168 1.66898
R24223 VDD.n1240 VDD.n1230 1.66898
R24224 VDD.n884 VDD.n874 1.66898
R24225 VDD.n918 VDD.n908 1.66898
R24226 VDD.n980 VDD.n970 1.66898
R24227 VDD.n624 VDD.n614 1.66898
R24228 VDD.n658 VDD.n648 1.66898
R24229 VDD.n720 VDD.n710 1.66898
R24230 VDD.n364 VDD.n354 1.66898
R24231 VDD.n398 VDD.n388 1.66898
R24232 VDD.n460 VDD.n450 1.66898
R24233 VDD.n7280 VDD.n7270 1.66898
R24234 VDD.n7314 VDD.n7304 1.66898
R24235 VDD.n7376 VDD.n7366 1.66898
R24236 VDD.n5102 VDD.n5092 1.66898
R24237 VDD.n5164 VDD.n5154 1.66898
R24238 VDD.n5198 VDD.n5188 1.66898
R24239 VDD.n5238 VDD.n5228 1.66898
R24240 VDD.n5300 VDD.n5290 1.66898
R24241 VDD.n5334 VDD.n5324 1.66898
R24242 VDD.n5374 VDD.n5364 1.66898
R24243 VDD.n5436 VDD.n5426 1.66898
R24244 VDD.n5470 VDD.n5460 1.66898
R24245 VDD.n5510 VDD.n5500 1.66898
R24246 VDD.n5572 VDD.n5562 1.66898
R24247 VDD.n5606 VDD.n5596 1.66898
R24248 VDD.n5646 VDD.n5636 1.66898
R24249 VDD.n5708 VDD.n5698 1.66898
R24250 VDD.n5742 VDD.n5732 1.66898
R24251 VDD.n5782 VDD.n5772 1.66898
R24252 VDD.n5844 VDD.n5834 1.66898
R24253 VDD.n5878 VDD.n5868 1.66898
R24254 VDD.n5918 VDD.n5908 1.66898
R24255 VDD.n5980 VDD.n5970 1.66898
R24256 VDD.n6014 VDD.n6004 1.66898
R24257 VDD.n4933 VDD.n4923 1.66898
R24258 VDD.n4871 VDD.n4861 1.66898
R24259 VDD.n4837 VDD.n4827 1.66898
R24260 VDD.n3803 VDD.n3793 1.66898
R24261 VDD.n2977 VDD.n2967 1.66898
R24262 VDD.n3012 VDD.n3002 1.66898
R24263 VDD.n2841 VDD.n2831 1.66898
R24264 VDD.n2876 VDD.n2866 1.66898
R24265 VDD.n2705 VDD.n2695 1.66898
R24266 VDD.n2740 VDD.n2730 1.66898
R24267 VDD.n2569 VDD.n2559 1.66898
R24268 VDD.n2604 VDD.n2594 1.66898
R24269 VDD.n2433 VDD.n2423 1.66898
R24270 VDD.n2468 VDD.n2458 1.66898
R24271 VDD.n2297 VDD.n2287 1.66898
R24272 VDD.n2332 VDD.n2322 1.66898
R24273 VDD.n2161 VDD.n2151 1.66898
R24274 VDD.n2196 VDD.n2186 1.66898
R24275 VDD.n2060 VDD.n2050 1.66898
R24276 VDD.n2025 VDD.n2015 1.66898
R24277 VDD.n1924 VDD.n1914 1.66898
R24278 VDD.n35 VDD.n25 1.66898
R24279 VDD.n7731 VDD.n1 1.66898
R24280 VDD.n7627 VDD.n7617 1.66898
R24281 VDD.n3583 VDD.n3582 1.64628
R24282 VDD.n3496 VDD.n3495 1.64315
R24283 VDD.n3489 VDD.n3488 1.64315
R24284 VDD.n3401 VDD.n3400 1.64315
R24285 VDD.n3889 VDD.n3739 1.58202
R24286 VDD.n4014 VDD.n2913 1.58202
R24287 VDD.n4139 VDD.n2777 1.58202
R24288 VDD.n4264 VDD.n2641 1.58202
R24289 VDD.n4389 VDD.n2505 1.58202
R24290 VDD.n4514 VDD.n2369 1.58202
R24291 VDD.n4639 VDD.n2233 1.58202
R24292 VDD.n4764 VDD.n2097 1.58202
R24293 VDD.n7205 VDD.n1961 1.58202
R24294 VDD.n3437 VDD 1.53854
R24295 VDD.n3340 VDD 1.53854
R24296 VDD.n3503 VDD 1.53854
R24297 VDD.n3532 VDD 1.53854
R24298 VDD.n3303 VDD 1.53854
R24299 VDD.n3408 VDD 1.53854
R24300 VDD.n3301 VDD 1.53854
R24301 VDD.n3197 VDD.n3173 1.46377
R24302 VDD.n3238 VDD.n3237 1.46377
R24303 VDD.n3262 VDD.n3261 1.46377
R24304 VDD.n3639 VDD.n3638 1.46377
R24305 VDD.n3642 VDD.n3095 1.46377
R24306 VDD.n3683 VDD.n3682 1.46377
R24307 VDD.n3706 VDD.n3705 1.46377
R24308 VDD.n3193 VDD.n3192 1.46377
R24309 VDD.n325 VDD 1.45974
R24310 VDD.n285 VDD 1.33448
R24311 VDD.n7257 VDD 1.33448
R24312 VDD.n3406 VDD.n3405 1.2977
R24313 VDD.n3438 VDD.n3436 1.26409
R24314 VDD.n3475 VDD.n3474 1.26409
R24315 VDD.n3504 VDD.n3315 1.26409
R24316 VDD.n3533 VDD.n3531 1.26409
R24317 VDD.n3569 VDD.n3568 1.26409
R24318 VDD.n3409 VDD.n3371 1.26409
R24319 VDD.n3281 VDD.n3265 1.26409
R24320 VDD.n302 VDD.n297 1.22567
R24321 VDD.n302 VDD.n301 1.22567
R24322 VDD.n335 VDD.n334 1.22567
R24323 VDD.n336 VDD.n335 1.22567
R24324 VDD.n299 VDD.n298 1.22567
R24325 VDD.n3143 VDD.n3142 1.19615
R24326 VDD.n3159 VDD.n3158 1.19615
R24327 VDD.n3207 VDD.n3206 1.19615
R24328 VDD.n3223 VDD.n3222 1.19615
R24329 VDD.n3104 VDD.n3103 1.19615
R24330 VDD.n3247 VDD.n3246 1.19615
R24331 VDD.n3358 VDD.n3357 1.19615
R24332 VDD.n3624 VDD.n3623 1.19615
R24333 VDD.n3065 VDD.n3064 1.19615
R24334 VDD.n3081 VDD.n3080 1.19615
R24335 VDD.n3652 VDD.n3651 1.19615
R24336 VDD.n3668 VDD.n3667 1.19615
R24337 VDD.n3046 VDD.n3045 1.19615
R24338 VDD.n3691 VDD.n3690 1.19615
R24339 VDD.n3123 VDD.n3122 1.19615
R24340 VDD.n3178 VDD.n3177 1.19615
R24341 VDD.n3712 VDD.n3711 1.19615
R24342 VDD.n340 VDD.n339 1.163
R24343 VDD.n3438 VDD.n3437 1.1418
R24344 VDD.n3475 VDD.n3340 1.1418
R24345 VDD.n3504 VDD.n3503 1.1418
R24346 VDD.n3533 VDD.n3532 1.1418
R24347 VDD.n3569 VDD.n3303 1.1418
R24348 VDD.n3409 VDD.n3408 1.1418
R24349 VDD.n3301 VDD.n3281 1.1418
R24350 VDD.n3148 VDD 1.09561
R24351 VDD.n3137 VDD 1.09561
R24352 VDD.n3164 VDD 1.09561
R24353 VDD.n3171 VDD 1.09561
R24354 VDD.n3212 VDD 1.09561
R24355 VDD.n3201 VDD 1.09561
R24356 VDD.n3228 VDD 1.09561
R24357 VDD.n3235 VDD 1.09561
R24358 VDD.n3109 VDD 1.09561
R24359 VDD.n3098 VDD 1.09561
R24360 VDD.n3252 VDD 1.09561
R24361 VDD.n3259 VDD 1.09561
R24362 VDD.n3363 VDD 1.09561
R24363 VDD.n3352 VDD 1.09561
R24364 VDD.n3629 VDD 1.09561
R24365 VDD.n3636 VDD 1.09561
R24366 VDD.n3070 VDD 1.09561
R24367 VDD.n3059 VDD 1.09561
R24368 VDD.n3086 VDD 1.09561
R24369 VDD.n3093 VDD 1.09561
R24370 VDD.n3657 VDD 1.09561
R24371 VDD.n3646 VDD 1.09561
R24372 VDD.n3673 VDD 1.09561
R24373 VDD.n3680 VDD 1.09561
R24374 VDD.n3696 VDD 1.09561
R24375 VDD.n3703 VDD 1.09561
R24376 VDD.n3128 VDD 1.09561
R24377 VDD.n3117 VDD 1.09561
R24378 VDD.n3183 VDD 1.09561
R24379 VDD.n3190 VDD 1.09561
R24380 VDD.n3717 VDD 1.09561
R24381 VDD.n3724 VDD 1.09561
R24382 VDD.n289 VDD.n287 1.02828
R24383 VDD.n337 VDD.n289 1.02828
R24384 VDD.n290 VDD.n288 1.02828
R24385 VDD.n1899 VDD 1.01137
R24386 VDD VDD.n1677 1.01137
R24387 VDD VDD.n1711 1.01137
R24388 VDD VDD.n1725 1.01137
R24389 VDD.n1726 VDD 1.01137
R24390 VDD VDD.n1739 1.01137
R24391 VDD.n1773 VDD 1.01137
R24392 VDD.n1639 VDD 1.01137
R24393 VDD VDD.n1417 1.01137
R24394 VDD VDD.n1451 1.01137
R24395 VDD VDD.n1465 1.01137
R24396 VDD.n1466 VDD 1.01137
R24397 VDD VDD.n1479 1.01137
R24398 VDD.n1513 VDD 1.01137
R24399 VDD.n1379 VDD 1.01137
R24400 VDD VDD.n1157 1.01137
R24401 VDD VDD.n1191 1.01137
R24402 VDD VDD.n1205 1.01137
R24403 VDD.n1206 VDD 1.01137
R24404 VDD VDD.n1219 1.01137
R24405 VDD.n1253 VDD 1.01137
R24406 VDD.n1119 VDD 1.01137
R24407 VDD VDD.n897 1.01137
R24408 VDD VDD.n931 1.01137
R24409 VDD VDD.n945 1.01137
R24410 VDD.n946 VDD 1.01137
R24411 VDD VDD.n959 1.01137
R24412 VDD.n993 VDD 1.01137
R24413 VDD.n859 VDD 1.01137
R24414 VDD VDD.n637 1.01137
R24415 VDD VDD.n671 1.01137
R24416 VDD VDD.n685 1.01137
R24417 VDD.n686 VDD 1.01137
R24418 VDD VDD.n699 1.01137
R24419 VDD.n733 VDD 1.01137
R24420 VDD.n599 VDD 1.01137
R24421 VDD VDD.n377 1.01137
R24422 VDD VDD.n411 1.01137
R24423 VDD VDD.n425 1.01137
R24424 VDD.n426 VDD 1.01137
R24425 VDD VDD.n439 1.01137
R24426 VDD.n473 VDD 1.01137
R24427 VDD.n58 VDD 1.01137
R24428 VDD.n264 VDD 1.01137
R24429 VDD.n250 VDD 1.01137
R24430 VDD.n83 VDD 1.01137
R24431 VDD.n229 VDD 1.01137
R24432 VDD.n215 VDD 1.01137
R24433 VDD.n108 VDD 1.01137
R24434 VDD.n194 VDD 1.01137
R24435 VDD.n180 VDD 1.01137
R24436 VDD.n133 VDD 1.01137
R24437 VDD.n159 VDD 1.01137
R24438 VDD.n145 VDD 1.01137
R24439 VDD.n7515 VDD 1.01137
R24440 VDD VDD.n7293 1.01137
R24441 VDD VDD.n7327 1.01137
R24442 VDD VDD.n7341 1.01137
R24443 VDD.n7342 VDD 1.01137
R24444 VDD VDD.n7355 1.01137
R24445 VDD.n7389 VDD 1.01137
R24446 VDD.n7113 VDD 1.01137
R24447 VDD.n7099 VDD 1.01137
R24448 VDD.n6932 VDD 1.01137
R24449 VDD.n7078 VDD 1.01137
R24450 VDD.n7064 VDD 1.01137
R24451 VDD.n6957 VDD 1.01137
R24452 VDD.n7043 VDD 1.01137
R24453 VDD.n7029 VDD 1.01137
R24454 VDD.n6982 VDD 1.01137
R24455 VDD.n7008 VDD 1.01137
R24456 VDD.n6994 VDD 1.01137
R24457 VDD.n5113 VDD 1.01137
R24458 VDD VDD.n5126 1.01137
R24459 VDD.n5139 VDD 1.01137
R24460 VDD.n5141 VDD 1.01137
R24461 VDD.n5175 VDD 1.01137
R24462 VDD.n6765 VDD 1.01137
R24463 VDD.n5249 VDD 1.01137
R24464 VDD VDD.n5262 1.01137
R24465 VDD.n5275 VDD 1.01137
R24466 VDD.n5277 VDD 1.01137
R24467 VDD.n5311 VDD 1.01137
R24468 VDD.n6642 VDD 1.01137
R24469 VDD.n5385 VDD 1.01137
R24470 VDD VDD.n5398 1.01137
R24471 VDD.n5411 VDD 1.01137
R24472 VDD.n5413 VDD 1.01137
R24473 VDD.n5447 VDD 1.01137
R24474 VDD.n6519 VDD 1.01137
R24475 VDD.n5521 VDD 1.01137
R24476 VDD VDD.n5534 1.01137
R24477 VDD.n5547 VDD 1.01137
R24478 VDD.n5549 VDD 1.01137
R24479 VDD.n5583 VDD 1.01137
R24480 VDD.n6396 VDD 1.01137
R24481 VDD.n5657 VDD 1.01137
R24482 VDD VDD.n5670 1.01137
R24483 VDD.n5683 VDD 1.01137
R24484 VDD.n5685 VDD 1.01137
R24485 VDD.n5719 VDD 1.01137
R24486 VDD.n6273 VDD 1.01137
R24487 VDD.n5793 VDD 1.01137
R24488 VDD VDD.n5806 1.01137
R24489 VDD.n5819 VDD 1.01137
R24490 VDD.n5821 VDD 1.01137
R24491 VDD.n5855 VDD 1.01137
R24492 VDD.n6150 VDD 1.01137
R24493 VDD.n5929 VDD 1.01137
R24494 VDD VDD.n5942 1.01137
R24495 VDD.n5955 VDD 1.01137
R24496 VDD.n5957 VDD 1.01137
R24497 VDD.n5991 VDD 1.01137
R24498 VDD.n6027 VDD 1.01137
R24499 VDD VDD.n4912 1.01137
R24500 VDD.n4899 VDD 1.01137
R24501 VDD VDD.n4898 1.01137
R24502 VDD VDD.n4884 1.01137
R24503 VDD VDD.n4850 1.01137
R24504 VDD.n5072 VDD 1.01137
R24505 VDD.n3887 VDD 1.01137
R24506 VDD VDD.n3768 1.01137
R24507 VDD.n3769 VDD 1.01137
R24508 VDD VDD.n3782 1.01137
R24509 VDD.n3816 VDD 1.01137
R24510 VDD.n4012 VDD 1.01137
R24511 VDD VDD.n2942 1.01137
R24512 VDD.n2943 VDD 1.01137
R24513 VDD VDD.n2956 1.01137
R24514 VDD.n3941 VDD 1.01137
R24515 VDD.n3939 VDD 1.01137
R24516 VDD VDD.n3025 1.01137
R24517 VDD.n4137 VDD 1.01137
R24518 VDD VDD.n2806 1.01137
R24519 VDD.n2807 VDD 1.01137
R24520 VDD VDD.n2820 1.01137
R24521 VDD.n4066 VDD 1.01137
R24522 VDD.n4064 VDD 1.01137
R24523 VDD VDD.n2889 1.01137
R24524 VDD.n4262 VDD 1.01137
R24525 VDD VDD.n2670 1.01137
R24526 VDD.n2671 VDD 1.01137
R24527 VDD VDD.n2684 1.01137
R24528 VDD.n4191 VDD 1.01137
R24529 VDD.n4189 VDD 1.01137
R24530 VDD VDD.n2753 1.01137
R24531 VDD.n4387 VDD 1.01137
R24532 VDD VDD.n2534 1.01137
R24533 VDD.n2535 VDD 1.01137
R24534 VDD VDD.n2548 1.01137
R24535 VDD.n4316 VDD 1.01137
R24536 VDD.n4314 VDD 1.01137
R24537 VDD VDD.n2617 1.01137
R24538 VDD.n4512 VDD 1.01137
R24539 VDD VDD.n2398 1.01137
R24540 VDD.n2399 VDD 1.01137
R24541 VDD VDD.n2412 1.01137
R24542 VDD.n4441 VDD 1.01137
R24543 VDD.n4439 VDD 1.01137
R24544 VDD VDD.n2481 1.01137
R24545 VDD.n4637 VDD 1.01137
R24546 VDD VDD.n2262 1.01137
R24547 VDD.n2263 VDD 1.01137
R24548 VDD VDD.n2276 1.01137
R24549 VDD.n4566 VDD 1.01137
R24550 VDD.n4564 VDD 1.01137
R24551 VDD VDD.n2345 1.01137
R24552 VDD.n4762 VDD 1.01137
R24553 VDD VDD.n2126 1.01137
R24554 VDD.n2127 VDD 1.01137
R24555 VDD VDD.n2140 1.01137
R24556 VDD.n4691 VDD 1.01137
R24557 VDD.n4689 VDD 1.01137
R24558 VDD VDD.n2209 1.01137
R24559 VDD.n4814 VDD 1.01137
R24560 VDD VDD.n2073 1.01137
R24561 VDD.n7203 VDD 1.01137
R24562 VDD VDD.n1990 1.01137
R24563 VDD.n1991 VDD 1.01137
R24564 VDD VDD.n2004 1.01137
R24565 VDD.n7132 VDD 1.01137
R24566 VDD.n7255 VDD 1.01137
R24567 VDD VDD.n1937 1.01137
R24568 VDD.n7521 VDD 1.01137
R24569 VDD VDD.n0 1.01137
R24570 VDD VDD.n7578 1.01137
R24571 VDD VDD.n7592 1.01137
R24572 VDD.n7593 VDD 1.01137
R24573 VDD VDD.n7606 1.01137
R24574 VDD.n7640 VDD 1.01137
R24575 VDD.n3449 VDD 0.980969
R24576 VDD.n3486 VDD 0.980969
R24577 VDD.n3338 VDD 0.980969
R24578 VDD.n3544 VDD 0.980969
R24579 VDD.n3394 VDD 0.980969
R24580 VDD.n3592 VDD 0.980969
R24581 VDD.n3580 VDD 0.965885
R24582 VDD.n7128 VDD.n7127 0.938
R24583 VDD.n285 VDD.n284 0.845609
R24584 VDD.n3435 VDD.n3422 0.845609
R24585 VDD.n3473 VDD.n3460 0.845609
R24586 VDD.n3514 VDD.n3513 0.845609
R24587 VDD.n3530 VDD.n3517 0.845609
R24588 VDD.n3567 VDD.n3554 0.845609
R24589 VDD.n3419 VDD.n3418 0.845609
R24590 VDD.n3618 VDD.n3617 0.845609
R24591 VDD.n1676 VDD.n1664 0.834739
R24592 VDD.n1677 VDD.n1676 0.834739
R24593 VDD.n1710 VDD.n1698 0.834739
R24594 VDD.n1711 VDD.n1710 0.834739
R24595 VDD.n1738 VDD.n1726 0.834739
R24596 VDD.n1739 VDD.n1738 0.834739
R24597 VDD.n1772 VDD.n1760 0.834739
R24598 VDD.n1773 VDD.n1772 0.834739
R24599 VDD.n1416 VDD.n1404 0.834739
R24600 VDD.n1417 VDD.n1416 0.834739
R24601 VDD.n1450 VDD.n1438 0.834739
R24602 VDD.n1451 VDD.n1450 0.834739
R24603 VDD.n1478 VDD.n1466 0.834739
R24604 VDD.n1479 VDD.n1478 0.834739
R24605 VDD.n1512 VDD.n1500 0.834739
R24606 VDD.n1513 VDD.n1512 0.834739
R24607 VDD.n1156 VDD.n1144 0.834739
R24608 VDD.n1157 VDD.n1156 0.834739
R24609 VDD.n1190 VDD.n1178 0.834739
R24610 VDD.n1191 VDD.n1190 0.834739
R24611 VDD.n1218 VDD.n1206 0.834739
R24612 VDD.n1219 VDD.n1218 0.834739
R24613 VDD.n1252 VDD.n1240 0.834739
R24614 VDD.n1253 VDD.n1252 0.834739
R24615 VDD.n896 VDD.n884 0.834739
R24616 VDD.n897 VDD.n896 0.834739
R24617 VDD.n930 VDD.n918 0.834739
R24618 VDD.n931 VDD.n930 0.834739
R24619 VDD.n958 VDD.n946 0.834739
R24620 VDD.n959 VDD.n958 0.834739
R24621 VDD.n992 VDD.n980 0.834739
R24622 VDD.n993 VDD.n992 0.834739
R24623 VDD.n636 VDD.n624 0.834739
R24624 VDD.n637 VDD.n636 0.834739
R24625 VDD.n670 VDD.n658 0.834739
R24626 VDD.n671 VDD.n670 0.834739
R24627 VDD.n698 VDD.n686 0.834739
R24628 VDD.n699 VDD.n698 0.834739
R24629 VDD.n732 VDD.n720 0.834739
R24630 VDD.n733 VDD.n732 0.834739
R24631 VDD.n376 VDD.n364 0.834739
R24632 VDD.n377 VDD.n376 0.834739
R24633 VDD.n410 VDD.n398 0.834739
R24634 VDD.n411 VDD.n410 0.834739
R24635 VDD.n438 VDD.n426 0.834739
R24636 VDD.n439 VDD.n438 0.834739
R24637 VDD.n472 VDD.n460 0.834739
R24638 VDD.n473 VDD.n472 0.834739
R24639 VDD.n59 VDD.n58 0.834739
R24640 VDD.n264 VDD.n59 0.834739
R24641 VDD.n263 VDD.n61 0.834739
R24642 VDD.n250 VDD.n61 0.834739
R24643 VDD.n84 VDD.n83 0.834739
R24644 VDD.n229 VDD.n84 0.834739
R24645 VDD.n228 VDD.n86 0.834739
R24646 VDD.n215 VDD.n86 0.834739
R24647 VDD.n109 VDD.n108 0.834739
R24648 VDD.n194 VDD.n109 0.834739
R24649 VDD.n193 VDD.n111 0.834739
R24650 VDD.n180 VDD.n111 0.834739
R24651 VDD.n134 VDD.n133 0.834739
R24652 VDD.n159 VDD.n134 0.834739
R24653 VDD.n158 VDD.n136 0.834739
R24654 VDD.n145 VDD.n136 0.834739
R24655 VDD.n7292 VDD.n7280 0.834739
R24656 VDD.n7293 VDD.n7292 0.834739
R24657 VDD.n7326 VDD.n7314 0.834739
R24658 VDD.n7327 VDD.n7326 0.834739
R24659 VDD.n7354 VDD.n7342 0.834739
R24660 VDD.n7355 VDD.n7354 0.834739
R24661 VDD.n7388 VDD.n7376 0.834739
R24662 VDD.n7389 VDD.n7388 0.834739
R24663 VDD.n7127 VDD.n6890 0.834739
R24664 VDD.n7113 VDD.n6890 0.834739
R24665 VDD.n7112 VDD.n6910 0.834739
R24666 VDD.n7099 VDD.n6910 0.834739
R24667 VDD.n6933 VDD.n6932 0.834739
R24668 VDD.n7078 VDD.n6933 0.834739
R24669 VDD.n7077 VDD.n6935 0.834739
R24670 VDD.n7064 VDD.n6935 0.834739
R24671 VDD.n6958 VDD.n6957 0.834739
R24672 VDD.n7043 VDD.n6958 0.834739
R24673 VDD.n7042 VDD.n6960 0.834739
R24674 VDD.n7029 VDD.n6960 0.834739
R24675 VDD.n6983 VDD.n6982 0.834739
R24676 VDD.n7008 VDD.n6983 0.834739
R24677 VDD.n7007 VDD.n6985 0.834739
R24678 VDD.n6994 VDD.n6985 0.834739
R24679 VDD.n6886 VDD.n5076 0.834739
R24680 VDD.n5092 VDD.n5076 0.834739
R24681 VDD.n5125 VDD.n5113 0.834739
R24682 VDD.n5126 VDD.n5125 0.834739
R24683 VDD.n5153 VDD.n5141 0.834739
R24684 VDD.n5154 VDD.n5153 0.834739
R24685 VDD.n5187 VDD.n5175 0.834739
R24686 VDD.n5188 VDD.n5187 0.834739
R24687 VDD.n6763 VDD.n5212 0.834739
R24688 VDD.n5228 VDD.n5212 0.834739
R24689 VDD.n5261 VDD.n5249 0.834739
R24690 VDD.n5262 VDD.n5261 0.834739
R24691 VDD.n5289 VDD.n5277 0.834739
R24692 VDD.n5290 VDD.n5289 0.834739
R24693 VDD.n5323 VDD.n5311 0.834739
R24694 VDD.n5324 VDD.n5323 0.834739
R24695 VDD.n6640 VDD.n5348 0.834739
R24696 VDD.n5364 VDD.n5348 0.834739
R24697 VDD.n5397 VDD.n5385 0.834739
R24698 VDD.n5398 VDD.n5397 0.834739
R24699 VDD.n5425 VDD.n5413 0.834739
R24700 VDD.n5426 VDD.n5425 0.834739
R24701 VDD.n5459 VDD.n5447 0.834739
R24702 VDD.n5460 VDD.n5459 0.834739
R24703 VDD.n6517 VDD.n5484 0.834739
R24704 VDD.n5500 VDD.n5484 0.834739
R24705 VDD.n5533 VDD.n5521 0.834739
R24706 VDD.n5534 VDD.n5533 0.834739
R24707 VDD.n5561 VDD.n5549 0.834739
R24708 VDD.n5562 VDD.n5561 0.834739
R24709 VDD.n5595 VDD.n5583 0.834739
R24710 VDD.n5596 VDD.n5595 0.834739
R24711 VDD.n6394 VDD.n5620 0.834739
R24712 VDD.n5636 VDD.n5620 0.834739
R24713 VDD.n5669 VDD.n5657 0.834739
R24714 VDD.n5670 VDD.n5669 0.834739
R24715 VDD.n5697 VDD.n5685 0.834739
R24716 VDD.n5698 VDD.n5697 0.834739
R24717 VDD.n5731 VDD.n5719 0.834739
R24718 VDD.n5732 VDD.n5731 0.834739
R24719 VDD.n6271 VDD.n5756 0.834739
R24720 VDD.n5772 VDD.n5756 0.834739
R24721 VDD.n5805 VDD.n5793 0.834739
R24722 VDD.n5806 VDD.n5805 0.834739
R24723 VDD.n5833 VDD.n5821 0.834739
R24724 VDD.n5834 VDD.n5833 0.834739
R24725 VDD.n5867 VDD.n5855 0.834739
R24726 VDD.n5868 VDD.n5867 0.834739
R24727 VDD.n6148 VDD.n5892 0.834739
R24728 VDD.n5908 VDD.n5892 0.834739
R24729 VDD.n5941 VDD.n5929 0.834739
R24730 VDD.n5942 VDD.n5941 0.834739
R24731 VDD.n5969 VDD.n5957 0.834739
R24732 VDD.n5970 VDD.n5969 0.834739
R24733 VDD.n6003 VDD.n5991 0.834739
R24734 VDD.n6004 VDD.n6003 0.834739
R24735 VDD.n4953 VDD.n4933 0.834739
R24736 VDD.n4912 VDD.n4911 0.834739
R24737 VDD.n4911 VDD.n4899 0.834739
R24738 VDD.n4884 VDD.n4883 0.834739
R24739 VDD.n4883 VDD.n4871 0.834739
R24740 VDD.n4850 VDD.n4849 0.834739
R24741 VDD.n4849 VDD.n4837 0.834739
R24742 VDD.n3889 VDD.n3888 0.834739
R24743 VDD.n3888 VDD.n3887 0.834739
R24744 VDD.n3781 VDD.n3769 0.834739
R24745 VDD.n3782 VDD.n3781 0.834739
R24746 VDD.n3815 VDD.n3803 0.834739
R24747 VDD.n3816 VDD.n3815 0.834739
R24748 VDD.n4014 VDD.n4013 0.834739
R24749 VDD.n4013 VDD.n4012 0.834739
R24750 VDD.n2955 VDD.n2943 0.834739
R24751 VDD.n2956 VDD.n2955 0.834739
R24752 VDD.n2989 VDD.n2977 0.834739
R24753 VDD.n3941 VDD.n2989 0.834739
R24754 VDD.n3024 VDD.n3012 0.834739
R24755 VDD.n3025 VDD.n3024 0.834739
R24756 VDD.n4139 VDD.n4138 0.834739
R24757 VDD.n4138 VDD.n4137 0.834739
R24758 VDD.n2819 VDD.n2807 0.834739
R24759 VDD.n2820 VDD.n2819 0.834739
R24760 VDD.n2853 VDD.n2841 0.834739
R24761 VDD.n4066 VDD.n2853 0.834739
R24762 VDD.n2888 VDD.n2876 0.834739
R24763 VDD.n2889 VDD.n2888 0.834739
R24764 VDD.n4264 VDD.n4263 0.834739
R24765 VDD.n4263 VDD.n4262 0.834739
R24766 VDD.n2683 VDD.n2671 0.834739
R24767 VDD.n2684 VDD.n2683 0.834739
R24768 VDD.n2717 VDD.n2705 0.834739
R24769 VDD.n4191 VDD.n2717 0.834739
R24770 VDD.n2752 VDD.n2740 0.834739
R24771 VDD.n2753 VDD.n2752 0.834739
R24772 VDD.n4389 VDD.n4388 0.834739
R24773 VDD.n4388 VDD.n4387 0.834739
R24774 VDD.n2547 VDD.n2535 0.834739
R24775 VDD.n2548 VDD.n2547 0.834739
R24776 VDD.n2581 VDD.n2569 0.834739
R24777 VDD.n4316 VDD.n2581 0.834739
R24778 VDD.n2616 VDD.n2604 0.834739
R24779 VDD.n2617 VDD.n2616 0.834739
R24780 VDD.n4514 VDD.n4513 0.834739
R24781 VDD.n4513 VDD.n4512 0.834739
R24782 VDD.n2411 VDD.n2399 0.834739
R24783 VDD.n2412 VDD.n2411 0.834739
R24784 VDD.n2445 VDD.n2433 0.834739
R24785 VDD.n4441 VDD.n2445 0.834739
R24786 VDD.n2480 VDD.n2468 0.834739
R24787 VDD.n2481 VDD.n2480 0.834739
R24788 VDD.n4639 VDD.n4638 0.834739
R24789 VDD.n4638 VDD.n4637 0.834739
R24790 VDD.n2275 VDD.n2263 0.834739
R24791 VDD.n2276 VDD.n2275 0.834739
R24792 VDD.n2309 VDD.n2297 0.834739
R24793 VDD.n4566 VDD.n2309 0.834739
R24794 VDD.n2344 VDD.n2332 0.834739
R24795 VDD.n2345 VDD.n2344 0.834739
R24796 VDD.n4764 VDD.n4763 0.834739
R24797 VDD.n4763 VDD.n4762 0.834739
R24798 VDD.n2139 VDD.n2127 0.834739
R24799 VDD.n2140 VDD.n2139 0.834739
R24800 VDD.n2173 VDD.n2161 0.834739
R24801 VDD.n4691 VDD.n2173 0.834739
R24802 VDD.n2208 VDD.n2196 0.834739
R24803 VDD.n2209 VDD.n2208 0.834739
R24804 VDD.n2072 VDD.n2060 0.834739
R24805 VDD.n2073 VDD.n2072 0.834739
R24806 VDD.n7205 VDD.n7204 0.834739
R24807 VDD.n7204 VDD.n7203 0.834739
R24808 VDD.n2003 VDD.n1991 0.834739
R24809 VDD.n2004 VDD.n2003 0.834739
R24810 VDD.n2037 VDD.n2025 0.834739
R24811 VDD.n7132 VDD.n2037 0.834739
R24812 VDD.n1936 VDD.n1924 0.834739
R24813 VDD.n1937 VDD.n1936 0.834739
R24814 VDD.n25 VDD.n24 0.834739
R24815 VDD.n24 VDD.n0 0.834739
R24816 VDD.n7577 VDD.n1 0.834739
R24817 VDD.n7578 VDD.n7577 0.834739
R24818 VDD.n7605 VDD.n7593 0.834739
R24819 VDD.n7606 VDD.n7605 0.834739
R24820 VDD.n7639 VDD.n7627 0.834739
R24821 VDD.n7640 VDD.n7639 0.834739
R24822 VDD.n321 VDD.n320 0.819084
R24823 VDD.n320 VDD.n319 0.819084
R24824 VDD.n1676 VDD.n1674 0.807565
R24825 VDD.n1676 VDD.n1675 0.807565
R24826 VDD.n1710 VDD.n1708 0.807565
R24827 VDD.n1710 VDD.n1709 0.807565
R24828 VDD.n1738 VDD.n1736 0.807565
R24829 VDD.n1738 VDD.n1737 0.807565
R24830 VDD.n1772 VDD.n1770 0.807565
R24831 VDD.n1772 VDD.n1771 0.807565
R24832 VDD.n1416 VDD.n1414 0.807565
R24833 VDD.n1416 VDD.n1415 0.807565
R24834 VDD.n1450 VDD.n1448 0.807565
R24835 VDD.n1450 VDD.n1449 0.807565
R24836 VDD.n1478 VDD.n1476 0.807565
R24837 VDD.n1478 VDD.n1477 0.807565
R24838 VDD.n1512 VDD.n1510 0.807565
R24839 VDD.n1512 VDD.n1511 0.807565
R24840 VDD.n1156 VDD.n1154 0.807565
R24841 VDD.n1156 VDD.n1155 0.807565
R24842 VDD.n1190 VDD.n1188 0.807565
R24843 VDD.n1190 VDD.n1189 0.807565
R24844 VDD.n1218 VDD.n1216 0.807565
R24845 VDD.n1218 VDD.n1217 0.807565
R24846 VDD.n1252 VDD.n1250 0.807565
R24847 VDD.n1252 VDD.n1251 0.807565
R24848 VDD.n896 VDD.n894 0.807565
R24849 VDD.n896 VDD.n895 0.807565
R24850 VDD.n930 VDD.n928 0.807565
R24851 VDD.n930 VDD.n929 0.807565
R24852 VDD.n958 VDD.n956 0.807565
R24853 VDD.n958 VDD.n957 0.807565
R24854 VDD.n992 VDD.n990 0.807565
R24855 VDD.n992 VDD.n991 0.807565
R24856 VDD.n636 VDD.n634 0.807565
R24857 VDD.n636 VDD.n635 0.807565
R24858 VDD.n670 VDD.n668 0.807565
R24859 VDD.n670 VDD.n669 0.807565
R24860 VDD.n698 VDD.n696 0.807565
R24861 VDD.n698 VDD.n697 0.807565
R24862 VDD.n732 VDD.n730 0.807565
R24863 VDD.n732 VDD.n731 0.807565
R24864 VDD.n376 VDD.n374 0.807565
R24865 VDD.n376 VDD.n375 0.807565
R24866 VDD.n410 VDD.n408 0.807565
R24867 VDD.n410 VDD.n409 0.807565
R24868 VDD.n438 VDD.n436 0.807565
R24869 VDD.n438 VDD.n437 0.807565
R24870 VDD.n472 VDD.n470 0.807565
R24871 VDD.n472 VDD.n471 0.807565
R24872 VDD.n325 VDD.n304 0.807565
R24873 VDD.n136 VDD.n135 0.807565
R24874 VDD.n134 VDD.n132 0.807565
R24875 VDD.n111 VDD.n110 0.807565
R24876 VDD.n109 VDD.n107 0.807565
R24877 VDD.n86 VDD.n85 0.807565
R24878 VDD.n84 VDD.n82 0.807565
R24879 VDD.n61 VDD.n60 0.807565
R24880 VDD.n59 VDD.n57 0.807565
R24881 VDD.n7292 VDD.n7290 0.807565
R24882 VDD.n7292 VDD.n7291 0.807565
R24883 VDD.n7326 VDD.n7324 0.807565
R24884 VDD.n7326 VDD.n7325 0.807565
R24885 VDD.n7354 VDD.n7352 0.807565
R24886 VDD.n7354 VDD.n7353 0.807565
R24887 VDD.n7388 VDD.n7386 0.807565
R24888 VDD.n7388 VDD.n7387 0.807565
R24889 VDD.n6985 VDD.n6984 0.807565
R24890 VDD.n6983 VDD.n6981 0.807565
R24891 VDD.n6960 VDD.n6959 0.807565
R24892 VDD.n6958 VDD.n6956 0.807565
R24893 VDD.n6935 VDD.n6934 0.807565
R24894 VDD.n6933 VDD.n6931 0.807565
R24895 VDD.n6910 VDD.n6909 0.807565
R24896 VDD.n6890 VDD.n6889 0.807565
R24897 VDD.n5076 VDD.n5074 0.807565
R24898 VDD.n5076 VDD.n5075 0.807565
R24899 VDD.n5125 VDD.n5123 0.807565
R24900 VDD.n5125 VDD.n5124 0.807565
R24901 VDD.n5153 VDD.n5151 0.807565
R24902 VDD.n5153 VDD.n5152 0.807565
R24903 VDD.n5187 VDD.n5185 0.807565
R24904 VDD.n5187 VDD.n5186 0.807565
R24905 VDD.n5212 VDD.n5210 0.807565
R24906 VDD.n5212 VDD.n5211 0.807565
R24907 VDD.n5261 VDD.n5259 0.807565
R24908 VDD.n5261 VDD.n5260 0.807565
R24909 VDD.n5289 VDD.n5287 0.807565
R24910 VDD.n5289 VDD.n5288 0.807565
R24911 VDD.n5323 VDD.n5321 0.807565
R24912 VDD.n5323 VDD.n5322 0.807565
R24913 VDD.n5348 VDD.n5346 0.807565
R24914 VDD.n5348 VDD.n5347 0.807565
R24915 VDD.n5397 VDD.n5395 0.807565
R24916 VDD.n5397 VDD.n5396 0.807565
R24917 VDD.n5425 VDD.n5423 0.807565
R24918 VDD.n5425 VDD.n5424 0.807565
R24919 VDD.n5459 VDD.n5457 0.807565
R24920 VDD.n5459 VDD.n5458 0.807565
R24921 VDD.n5484 VDD.n5482 0.807565
R24922 VDD.n5484 VDD.n5483 0.807565
R24923 VDD.n5533 VDD.n5531 0.807565
R24924 VDD.n5533 VDD.n5532 0.807565
R24925 VDD.n5561 VDD.n5559 0.807565
R24926 VDD.n5561 VDD.n5560 0.807565
R24927 VDD.n5595 VDD.n5593 0.807565
R24928 VDD.n5595 VDD.n5594 0.807565
R24929 VDD.n5620 VDD.n5618 0.807565
R24930 VDD.n5620 VDD.n5619 0.807565
R24931 VDD.n5669 VDD.n5667 0.807565
R24932 VDD.n5669 VDD.n5668 0.807565
R24933 VDD.n5697 VDD.n5695 0.807565
R24934 VDD.n5697 VDD.n5696 0.807565
R24935 VDD.n5731 VDD.n5729 0.807565
R24936 VDD.n5731 VDD.n5730 0.807565
R24937 VDD.n5756 VDD.n5754 0.807565
R24938 VDD.n5756 VDD.n5755 0.807565
R24939 VDD.n5805 VDD.n5803 0.807565
R24940 VDD.n5805 VDD.n5804 0.807565
R24941 VDD.n5833 VDD.n5831 0.807565
R24942 VDD.n5833 VDD.n5832 0.807565
R24943 VDD.n5867 VDD.n5865 0.807565
R24944 VDD.n5867 VDD.n5866 0.807565
R24945 VDD.n5892 VDD.n5890 0.807565
R24946 VDD.n5892 VDD.n5891 0.807565
R24947 VDD.n5941 VDD.n5939 0.807565
R24948 VDD.n5941 VDD.n5940 0.807565
R24949 VDD.n5969 VDD.n5967 0.807565
R24950 VDD.n5969 VDD.n5968 0.807565
R24951 VDD.n6003 VDD.n6001 0.807565
R24952 VDD.n6003 VDD.n6002 0.807565
R24953 VDD.n4953 VDD.n4951 0.807565
R24954 VDD.n4953 VDD.n4952 0.807565
R24955 VDD.n4911 VDD.n4909 0.807565
R24956 VDD.n4911 VDD.n4910 0.807565
R24957 VDD.n4883 VDD.n4881 0.807565
R24958 VDD.n4883 VDD.n4882 0.807565
R24959 VDD.n4849 VDD.n4847 0.807565
R24960 VDD.n4849 VDD.n4848 0.807565
R24961 VDD.n3888 VDD.n3740 0.807565
R24962 VDD.n3888 VDD.n3741 0.807565
R24963 VDD.n3781 VDD.n3779 0.807565
R24964 VDD.n3781 VDD.n3780 0.807565
R24965 VDD.n3815 VDD.n3813 0.807565
R24966 VDD.n3815 VDD.n3814 0.807565
R24967 VDD.n4013 VDD.n2914 0.807565
R24968 VDD.n4013 VDD.n2915 0.807565
R24969 VDD.n2955 VDD.n2953 0.807565
R24970 VDD.n2955 VDD.n2954 0.807565
R24971 VDD.n2989 VDD.n2987 0.807565
R24972 VDD.n2989 VDD.n2988 0.807565
R24973 VDD.n3024 VDD.n3022 0.807565
R24974 VDD.n3024 VDD.n3023 0.807565
R24975 VDD.n4138 VDD.n2778 0.807565
R24976 VDD.n4138 VDD.n2779 0.807565
R24977 VDD.n2819 VDD.n2817 0.807565
R24978 VDD.n2819 VDD.n2818 0.807565
R24979 VDD.n2853 VDD.n2851 0.807565
R24980 VDD.n2853 VDD.n2852 0.807565
R24981 VDD.n2888 VDD.n2886 0.807565
R24982 VDD.n2888 VDD.n2887 0.807565
R24983 VDD.n4263 VDD.n2642 0.807565
R24984 VDD.n4263 VDD.n2643 0.807565
R24985 VDD.n2683 VDD.n2681 0.807565
R24986 VDD.n2683 VDD.n2682 0.807565
R24987 VDD.n2717 VDD.n2715 0.807565
R24988 VDD.n2717 VDD.n2716 0.807565
R24989 VDD.n2752 VDD.n2750 0.807565
R24990 VDD.n2752 VDD.n2751 0.807565
R24991 VDD.n4388 VDD.n2506 0.807565
R24992 VDD.n4388 VDD.n2507 0.807565
R24993 VDD.n2547 VDD.n2545 0.807565
R24994 VDD.n2547 VDD.n2546 0.807565
R24995 VDD.n2581 VDD.n2579 0.807565
R24996 VDD.n2581 VDD.n2580 0.807565
R24997 VDD.n2616 VDD.n2614 0.807565
R24998 VDD.n2616 VDD.n2615 0.807565
R24999 VDD.n4513 VDD.n2370 0.807565
R25000 VDD.n4513 VDD.n2371 0.807565
R25001 VDD.n2411 VDD.n2409 0.807565
R25002 VDD.n2411 VDD.n2410 0.807565
R25003 VDD.n2445 VDD.n2443 0.807565
R25004 VDD.n2445 VDD.n2444 0.807565
R25005 VDD.n2480 VDD.n2478 0.807565
R25006 VDD.n2480 VDD.n2479 0.807565
R25007 VDD.n4638 VDD.n2234 0.807565
R25008 VDD.n4638 VDD.n2235 0.807565
R25009 VDD.n2275 VDD.n2273 0.807565
R25010 VDD.n2275 VDD.n2274 0.807565
R25011 VDD.n2309 VDD.n2307 0.807565
R25012 VDD.n2309 VDD.n2308 0.807565
R25013 VDD.n2344 VDD.n2342 0.807565
R25014 VDD.n2344 VDD.n2343 0.807565
R25015 VDD.n4763 VDD.n2098 0.807565
R25016 VDD.n4763 VDD.n2099 0.807565
R25017 VDD.n2139 VDD.n2137 0.807565
R25018 VDD.n2139 VDD.n2138 0.807565
R25019 VDD.n2173 VDD.n2171 0.807565
R25020 VDD.n2173 VDD.n2172 0.807565
R25021 VDD.n2208 VDD.n2206 0.807565
R25022 VDD.n2208 VDD.n2207 0.807565
R25023 VDD.n2072 VDD.n2070 0.807565
R25024 VDD.n2072 VDD.n2071 0.807565
R25025 VDD.n7204 VDD.n1962 0.807565
R25026 VDD.n7204 VDD.n1963 0.807565
R25027 VDD.n2003 VDD.n2001 0.807565
R25028 VDD.n2003 VDD.n2002 0.807565
R25029 VDD.n2037 VDD.n2035 0.807565
R25030 VDD.n2037 VDD.n2036 0.807565
R25031 VDD.n1936 VDD.n1934 0.807565
R25032 VDD.n1936 VDD.n1935 0.807565
R25033 VDD.n24 VDD.n22 0.807565
R25034 VDD.n24 VDD.n23 0.807565
R25035 VDD.n7577 VDD.n7575 0.807565
R25036 VDD.n7577 VDD.n7576 0.807565
R25037 VDD.n7605 VDD.n7603 0.807565
R25038 VDD.n7605 VDD.n7604 0.807565
R25039 VDD.n7639 VDD.n7637 0.807565
R25040 VDD.n7639 VDD.n7638 0.807565
R25041 VDD.n3151 VDD.n3150 0.796696
R25042 VDD.n3140 VDD.n3139 0.796696
R25043 VDD.n3167 VDD.n3166 0.796696
R25044 VDD.n3157 VDD.n3156 0.796696
R25045 VDD.n3215 VDD.n3214 0.796696
R25046 VDD.n3204 VDD.n3203 0.796696
R25047 VDD.n3231 VDD.n3230 0.796696
R25048 VDD.n3221 VDD.n3220 0.796696
R25049 VDD.n3112 VDD.n3111 0.796696
R25050 VDD.n3101 VDD.n3100 0.796696
R25051 VDD.n3255 VDD.n3254 0.796696
R25052 VDD.n3245 VDD.n3244 0.796696
R25053 VDD.n3366 VDD.n3365 0.796696
R25054 VDD.n3355 VDD.n3354 0.796696
R25055 VDD.n3632 VDD.n3631 0.796696
R25056 VDD.n3622 VDD.n3621 0.796696
R25057 VDD.n3073 VDD.n3072 0.796696
R25058 VDD.n3062 VDD.n3061 0.796696
R25059 VDD.n3089 VDD.n3088 0.796696
R25060 VDD.n3079 VDD.n3078 0.796696
R25061 VDD.n3660 VDD.n3659 0.796696
R25062 VDD.n3649 VDD.n3648 0.796696
R25063 VDD.n3676 VDD.n3675 0.796696
R25064 VDD.n3666 VDD.n3665 0.796696
R25065 VDD.n3050 VDD.n3049 0.796696
R25066 VDD.n3039 VDD.n3038 0.796696
R25067 VDD.n3699 VDD.n3698 0.796696
R25068 VDD.n3689 VDD.n3688 0.796696
R25069 VDD.n3131 VDD.n3130 0.796696
R25070 VDD.n3120 VDD.n3119 0.796696
R25071 VDD.n3186 VDD.n3185 0.796696
R25072 VDD.n3176 VDD.n3175 0.796696
R25073 VDD.n3720 VDD.n3719 0.796696
R25074 VDD.n3710 VDD.n3709 0.796696
R25075 VDD.n3146 VDD.n3145 0.783833
R25076 VDD.n3162 VDD.n3161 0.783833
R25077 VDD.n3210 VDD.n3209 0.783833
R25078 VDD.n3226 VDD.n3225 0.783833
R25079 VDD.n3107 VDD.n3106 0.783833
R25080 VDD.n3250 VDD.n3249 0.783833
R25081 VDD.n3361 VDD.n3360 0.783833
R25082 VDD.n3627 VDD.n3626 0.783833
R25083 VDD.n3068 VDD.n3067 0.783833
R25084 VDD.n3084 VDD.n3083 0.783833
R25085 VDD.n3655 VDD.n3654 0.783833
R25086 VDD.n3671 VDD.n3670 0.783833
R25087 VDD.n3048 VDD.n3047 0.783833
R25088 VDD.n3694 VDD.n3693 0.783833
R25089 VDD.n3126 VDD.n3125 0.783833
R25090 VDD.n3181 VDD.n3180 0.783833
R25091 VDD.n3715 VDD.n3714 0.783833
R25092 VDD.n316 VDD.n315 0.774559
R25093 VDD.n317 VDD.n316 0.774559
R25094 VDD.n3145 VDD 0.716182
R25095 VDD.n3161 VDD 0.716182
R25096 VDD.n3209 VDD 0.716182
R25097 VDD.n3225 VDD 0.716182
R25098 VDD.n3106 VDD 0.716182
R25099 VDD.n3249 VDD 0.716182
R25100 VDD.n3360 VDD 0.716182
R25101 VDD.n3626 VDD 0.716182
R25102 VDD.n3067 VDD 0.716182
R25103 VDD.n3083 VDD 0.716182
R25104 VDD.n3654 VDD 0.716182
R25105 VDD.n3670 VDD 0.716182
R25106 VDD.n3048 VDD 0.716182
R25107 VDD.n3693 VDD 0.716182
R25108 VDD.n3125 VDD 0.716182
R25109 VDD.n3180 VDD 0.716182
R25110 VDD.n3714 VDD 0.716182
R25111 VDD.n3151 VDD 0.662609
R25112 VDD.n3140 VDD 0.662609
R25113 VDD.n3167 VDD 0.662609
R25114 VDD.n3157 VDD 0.662609
R25115 VDD.n3215 VDD 0.662609
R25116 VDD.n3204 VDD 0.662609
R25117 VDD.n3231 VDD 0.662609
R25118 VDD.n3221 VDD 0.662609
R25119 VDD.n3112 VDD 0.662609
R25120 VDD.n3101 VDD 0.662609
R25121 VDD.n3255 VDD 0.662609
R25122 VDD.n3245 VDD 0.662609
R25123 VDD.n3366 VDD 0.662609
R25124 VDD.n3355 VDD 0.662609
R25125 VDD.n3632 VDD 0.662609
R25126 VDD.n3622 VDD 0.662609
R25127 VDD.n3073 VDD 0.662609
R25128 VDD.n3062 VDD 0.662609
R25129 VDD.n3089 VDD 0.662609
R25130 VDD.n3079 VDD 0.662609
R25131 VDD.n3660 VDD 0.662609
R25132 VDD.n3649 VDD 0.662609
R25133 VDD.n3676 VDD 0.662609
R25134 VDD.n3666 VDD 0.662609
R25135 VDD.n3699 VDD 0.662609
R25136 VDD.n3689 VDD 0.662609
R25137 VDD.n3131 VDD 0.662609
R25138 VDD.n3120 VDD 0.662609
R25139 VDD.n3186 VDD 0.662609
R25140 VDD.n3176 VDD 0.662609
R25141 VDD.n3720 VDD 0.662609
R25142 VDD.n3710 VDD 0.662609
R25143 VDD.n3396 VDD.n3395 0.648317
R25144 VDD.n3588 VDD.n3587 0.648317
R25145 VDD.n3585 VDD.n3584 0.648317
R25146 VDD.n3494 VDD.n3493 0.648317
R25147 VDD.n3499 VDD.n3498 0.648317
R25148 VDD.n3491 VDD.n3490 0.648317
R25149 VDD.n3399 VDD.n3398 0.648317
R25150 VDD.n3404 VDD.n3403 0.648317
R25151 VDD.n326 VDD.n325 0.6205
R25152 VDD.n1653 VDD 0.601043
R25153 VDD.n1687 VDD 0.601043
R25154 VDD.n1724 VDD 0.601043
R25155 VDD.n1749 VDD 0.601043
R25156 VDD.n1393 VDD 0.601043
R25157 VDD.n1427 VDD 0.601043
R25158 VDD.n1464 VDD 0.601043
R25159 VDD.n1489 VDD 0.601043
R25160 VDD.n1133 VDD 0.601043
R25161 VDD.n1167 VDD 0.601043
R25162 VDD.n1204 VDD 0.601043
R25163 VDD.n1229 VDD 0.601043
R25164 VDD.n873 VDD 0.601043
R25165 VDD.n907 VDD 0.601043
R25166 VDD.n944 VDD 0.601043
R25167 VDD.n969 VDD 0.601043
R25168 VDD.n613 VDD 0.601043
R25169 VDD.n647 VDD 0.601043
R25170 VDD.n684 VDD 0.601043
R25171 VDD.n709 VDD 0.601043
R25172 VDD.n353 VDD 0.601043
R25173 VDD.n387 VDD 0.601043
R25174 VDD.n424 VDD 0.601043
R25175 VDD.n449 VDD 0.601043
R25176 VDD VDD.n45 0.601043
R25177 VDD VDD.n70 0.601043
R25178 VDD VDD.n95 0.601043
R25179 VDD VDD.n120 0.601043
R25180 VDD.n7269 VDD 0.601043
R25181 VDD.n7303 VDD 0.601043
R25182 VDD.n7340 VDD 0.601043
R25183 VDD.n7365 VDD 0.601043
R25184 VDD VDD.n6919 0.601043
R25185 VDD VDD.n6944 0.601043
R25186 VDD VDD.n6969 0.601043
R25187 VDD VDD.n5112 0.601043
R25188 VDD VDD.n5140 0.601043
R25189 VDD VDD.n5174 0.601043
R25190 VDD VDD.n5209 0.601043
R25191 VDD.n6764 VDD 0.601043
R25192 VDD VDD.n5248 0.601043
R25193 VDD VDD.n5276 0.601043
R25194 VDD VDD.n5310 0.601043
R25195 VDD VDD.n5345 0.601043
R25196 VDD.n6641 VDD 0.601043
R25197 VDD VDD.n5384 0.601043
R25198 VDD VDD.n5412 0.601043
R25199 VDD VDD.n5446 0.601043
R25200 VDD VDD.n5481 0.601043
R25201 VDD.n6518 VDD 0.601043
R25202 VDD VDD.n5520 0.601043
R25203 VDD VDD.n5548 0.601043
R25204 VDD VDD.n5582 0.601043
R25205 VDD VDD.n5617 0.601043
R25206 VDD.n6395 VDD 0.601043
R25207 VDD VDD.n5656 0.601043
R25208 VDD VDD.n5684 0.601043
R25209 VDD VDD.n5718 0.601043
R25210 VDD VDD.n5753 0.601043
R25211 VDD.n6272 VDD 0.601043
R25212 VDD VDD.n5792 0.601043
R25213 VDD VDD.n5820 0.601043
R25214 VDD VDD.n5854 0.601043
R25215 VDD VDD.n5889 0.601043
R25216 VDD.n6149 VDD 0.601043
R25217 VDD VDD.n5928 0.601043
R25218 VDD VDD.n5956 0.601043
R25219 VDD VDD.n5990 0.601043
R25220 VDD VDD.n6025 0.601043
R25221 VDD.n6026 VDD 0.601043
R25222 VDD.n4922 VDD 0.601043
R25223 VDD.n4897 VDD 0.601043
R25224 VDD.n4860 VDD 0.601043
R25225 VDD.n4826 VDD 0.601043
R25226 VDD VDD.n5073 0.601043
R25227 VDD.n3767 VDD 0.601043
R25228 VDD.n3792 VDD 0.601043
R25229 VDD.n2941 VDD 0.601043
R25230 VDD.n2966 VDD 0.601043
R25231 VDD.n3001 VDD 0.601043
R25232 VDD.n3035 VDD 0.601043
R25233 VDD.n2805 VDD 0.601043
R25234 VDD.n2830 VDD 0.601043
R25235 VDD.n2865 VDD 0.601043
R25236 VDD.n2899 VDD 0.601043
R25237 VDD.n2669 VDD 0.601043
R25238 VDD.n2694 VDD 0.601043
R25239 VDD.n2729 VDD 0.601043
R25240 VDD.n2763 VDD 0.601043
R25241 VDD.n2533 VDD 0.601043
R25242 VDD.n2558 VDD 0.601043
R25243 VDD.n2593 VDD 0.601043
R25244 VDD.n2627 VDD 0.601043
R25245 VDD.n2397 VDD 0.601043
R25246 VDD.n2422 VDD 0.601043
R25247 VDD.n2457 VDD 0.601043
R25248 VDD.n2491 VDD 0.601043
R25249 VDD.n2261 VDD 0.601043
R25250 VDD.n2286 VDD 0.601043
R25251 VDD.n2321 VDD 0.601043
R25252 VDD.n2355 VDD 0.601043
R25253 VDD.n2125 VDD 0.601043
R25254 VDD.n2150 VDD 0.601043
R25255 VDD.n2185 VDD 0.601043
R25256 VDD.n2219 VDD 0.601043
R25257 VDD.n2049 VDD 0.601043
R25258 VDD.n2083 VDD 0.601043
R25259 VDD.n1989 VDD 0.601043
R25260 VDD.n2014 VDD 0.601043
R25261 VDD.n1913 VDD 0.601043
R25262 VDD.n1947 VDD 0.601043
R25263 VDD VDD.n7520 0.601043
R25264 VDD VDD.n7732 0.601043
R25265 VDD.n7591 VDD 0.601043
R25266 VDD.n7616 VDD 0.601043
R25267 VDD.n3395 VDD 0.592985
R25268 VDD.n3588 VDD 0.592985
R25269 VDD.n3584 VDD 0.592985
R25270 VDD.n3494 VDD 0.592985
R25271 VDD.n3499 VDD 0.592985
R25272 VDD.n3490 VDD 0.592985
R25273 VDD.n3399 VDD 0.592985
R25274 VDD.n3404 VDD 0.592985
R25275 VDD.n3050 VDD 0.524957
R25276 VDD.n3039 VDD 0.524957
R25277 VDD.n6897 VDD.n6888 0.5005
R25278 VDD.n340 VDD.n286 0.486913
R25279 VDD.n3147 VDD 0.447191
R25280 VDD.n3136 VDD 0.447191
R25281 VDD.n3163 VDD 0.447191
R25282 VDD.n3172 VDD 0.447191
R25283 VDD.n3211 VDD 0.447191
R25284 VDD.n3200 VDD 0.447191
R25285 VDD.n3227 VDD 0.447191
R25286 VDD.n3236 VDD 0.447191
R25287 VDD.n3108 VDD 0.447191
R25288 VDD.n3097 VDD 0.447191
R25289 VDD.n3251 VDD 0.447191
R25290 VDD.n3260 VDD 0.447191
R25291 VDD.n3362 VDD 0.447191
R25292 VDD.n3351 VDD 0.447191
R25293 VDD.n3628 VDD 0.447191
R25294 VDD.n3637 VDD 0.447191
R25295 VDD.n3069 VDD 0.447191
R25296 VDD.n3058 VDD 0.447191
R25297 VDD.n3085 VDD 0.447191
R25298 VDD.n3094 VDD 0.447191
R25299 VDD.n3656 VDD 0.447191
R25300 VDD.n3645 VDD 0.447191
R25301 VDD.n3672 VDD 0.447191
R25302 VDD.n3681 VDD 0.447191
R25303 VDD.n3046 VDD 0.447191
R25304 VDD.n3695 VDD 0.447191
R25305 VDD.n3704 VDD 0.447191
R25306 VDD.n3127 VDD 0.447191
R25307 VDD.n3116 VDD 0.447191
R25308 VDD.n3182 VDD 0.447191
R25309 VDD.n3191 VDD 0.447191
R25310 VDD.n3716 VDD 0.447191
R25311 VDD.n3725 VDD 0.447191
R25312 VDD.n3406 VDD.n3397 0.447
R25313 VDD.n3590 VDD.n3589 0.447
R25314 VDD.n3590 VDD.n3586 0.447
R25315 VDD.n3497 VDD.n3496 0.447
R25316 VDD.n3501 VDD.n3492 0.447
R25317 VDD.n3488 VDD.n3339 0.447
R25318 VDD.n3402 VDD.n3401 0.447
R25319 VDD.n3582 VDD.n3302 0.446929
R25320 VDD.n7257 VDD.n7256 0.435283
R25321 VDD.n1900 VDD.n1899 0.410826
R25322 VDD.n1654 VDD.n1653 0.410826
R25323 VDD.n1688 VDD.n1687 0.410826
R25324 VDD.n1725 VDD.n1724 0.410826
R25325 VDD.n1750 VDD.n1749 0.410826
R25326 VDD.n1640 VDD.n1639 0.410826
R25327 VDD.n1394 VDD.n1393 0.410826
R25328 VDD.n1428 VDD.n1427 0.410826
R25329 VDD.n1465 VDD.n1464 0.410826
R25330 VDD.n1490 VDD.n1489 0.410826
R25331 VDD.n1380 VDD.n1379 0.410826
R25332 VDD.n1134 VDD.n1133 0.410826
R25333 VDD.n1168 VDD.n1167 0.410826
R25334 VDD.n1205 VDD.n1204 0.410826
R25335 VDD.n1230 VDD.n1229 0.410826
R25336 VDD.n1120 VDD.n1119 0.410826
R25337 VDD.n874 VDD.n873 0.410826
R25338 VDD.n908 VDD.n907 0.410826
R25339 VDD.n945 VDD.n944 0.410826
R25340 VDD.n970 VDD.n969 0.410826
R25341 VDD.n860 VDD.n859 0.410826
R25342 VDD.n614 VDD.n613 0.410826
R25343 VDD.n648 VDD.n647 0.410826
R25344 VDD.n685 VDD.n684 0.410826
R25345 VDD.n710 VDD.n709 0.410826
R25346 VDD.n600 VDD.n599 0.410826
R25347 VDD.n354 VDD.n353 0.410826
R25348 VDD.n388 VDD.n387 0.410826
R25349 VDD.n425 VDD.n424 0.410826
R25350 VDD.n450 VDD.n449 0.410826
R25351 VDD.n284 VDD.n45 0.410826
R25352 VDD.n249 VDD.n70 0.410826
R25353 VDD.n214 VDD.n95 0.410826
R25354 VDD.n179 VDD.n120 0.410826
R25355 VDD.n7516 VDD.n7515 0.410826
R25356 VDD.n7270 VDD.n7269 0.410826
R25357 VDD.n7304 VDD.n7303 0.410826
R25358 VDD.n7341 VDD.n7340 0.410826
R25359 VDD.n7366 VDD.n7365 0.410826
R25360 VDD.n7098 VDD.n6919 0.410826
R25361 VDD.n7063 VDD.n6944 0.410826
R25362 VDD.n7028 VDD.n6969 0.410826
R25363 VDD.n5112 VDD.n5102 0.410826
R25364 VDD.n5140 VDD.n5139 0.410826
R25365 VDD.n5174 VDD.n5164 0.410826
R25366 VDD.n5209 VDD.n5198 0.410826
R25367 VDD.n6765 VDD.n6764 0.410826
R25368 VDD.n5248 VDD.n5238 0.410826
R25369 VDD.n5276 VDD.n5275 0.410826
R25370 VDD.n5310 VDD.n5300 0.410826
R25371 VDD.n5345 VDD.n5334 0.410826
R25372 VDD.n6642 VDD.n6641 0.410826
R25373 VDD.n5384 VDD.n5374 0.410826
R25374 VDD.n5412 VDD.n5411 0.410826
R25375 VDD.n5446 VDD.n5436 0.410826
R25376 VDD.n5481 VDD.n5470 0.410826
R25377 VDD.n6519 VDD.n6518 0.410826
R25378 VDD.n5520 VDD.n5510 0.410826
R25379 VDD.n5548 VDD.n5547 0.410826
R25380 VDD.n5582 VDD.n5572 0.410826
R25381 VDD.n5617 VDD.n5606 0.410826
R25382 VDD.n6396 VDD.n6395 0.410826
R25383 VDD.n5656 VDD.n5646 0.410826
R25384 VDD.n5684 VDD.n5683 0.410826
R25385 VDD.n5718 VDD.n5708 0.410826
R25386 VDD.n5753 VDD.n5742 0.410826
R25387 VDD.n6273 VDD.n6272 0.410826
R25388 VDD.n5792 VDD.n5782 0.410826
R25389 VDD.n5820 VDD.n5819 0.410826
R25390 VDD.n5854 VDD.n5844 0.410826
R25391 VDD.n5889 VDD.n5878 0.410826
R25392 VDD.n6150 VDD.n6149 0.410826
R25393 VDD.n5928 VDD.n5918 0.410826
R25394 VDD.n5956 VDD.n5955 0.410826
R25395 VDD.n5990 VDD.n5980 0.410826
R25396 VDD.n6025 VDD.n6014 0.410826
R25397 VDD.n6027 VDD.n6026 0.410826
R25398 VDD.n4923 VDD.n4922 0.410826
R25399 VDD.n4898 VDD.n4897 0.410826
R25400 VDD.n4861 VDD.n4860 0.410826
R25401 VDD.n4827 VDD.n4826 0.410826
R25402 VDD.n5073 VDD.n5072 0.410826
R25403 VDD.n3768 VDD.n3767 0.410826
R25404 VDD.n3793 VDD.n3792 0.410826
R25405 VDD.n2942 VDD.n2941 0.410826
R25406 VDD.n2967 VDD.n2966 0.410826
R25407 VDD.n3940 VDD.n3939 0.410826
R25408 VDD.n3002 VDD.n3001 0.410826
R25409 VDD.n2806 VDD.n2805 0.410826
R25410 VDD.n2831 VDD.n2830 0.410826
R25411 VDD.n4065 VDD.n4064 0.410826
R25412 VDD.n2866 VDD.n2865 0.410826
R25413 VDD.n2670 VDD.n2669 0.410826
R25414 VDD.n2695 VDD.n2694 0.410826
R25415 VDD.n4190 VDD.n4189 0.410826
R25416 VDD.n2730 VDD.n2729 0.410826
R25417 VDD.n2534 VDD.n2533 0.410826
R25418 VDD.n2559 VDD.n2558 0.410826
R25419 VDD.n4315 VDD.n4314 0.410826
R25420 VDD.n2594 VDD.n2593 0.410826
R25421 VDD.n2398 VDD.n2397 0.410826
R25422 VDD.n2423 VDD.n2422 0.410826
R25423 VDD.n4440 VDD.n4439 0.410826
R25424 VDD.n2458 VDD.n2457 0.410826
R25425 VDD.n2262 VDD.n2261 0.410826
R25426 VDD.n2287 VDD.n2286 0.410826
R25427 VDD.n4565 VDD.n4564 0.410826
R25428 VDD.n2322 VDD.n2321 0.410826
R25429 VDD.n2126 VDD.n2125 0.410826
R25430 VDD.n2151 VDD.n2150 0.410826
R25431 VDD.n4690 VDD.n4689 0.410826
R25432 VDD.n2186 VDD.n2185 0.410826
R25433 VDD.n4815 VDD.n4814 0.410826
R25434 VDD.n2050 VDD.n2049 0.410826
R25435 VDD.n1990 VDD.n1989 0.410826
R25436 VDD.n2015 VDD.n2014 0.410826
R25437 VDD.n7256 VDD.n7255 0.410826
R25438 VDD.n1914 VDD.n1913 0.410826
R25439 VDD.n7521 VDD.n7519 0.410826
R25440 VDD.n7520 VDD.n35 0.410826
R25441 VDD.n7732 VDD.n7731 0.410826
R25442 VDD.n7592 VDD.n7591 0.410826
R25443 VDD.n7617 VDD.n7616 0.410826
R25444 VDD.n3436 VDD.n3435 0.405391
R25445 VDD.n3474 VDD.n3473 0.405391
R25446 VDD.n3513 VDD.n3315 0.405391
R25447 VDD.n3531 VDD.n3530 0.405391
R25448 VDD.n3568 VDD.n3567 0.405391
R25449 VDD.n3418 VDD.n3371 0.405391
R25450 VDD.n3617 VDD.n3265 0.405391
R25451 VDD.n312 VDD.n305 0.397496
R25452 VDD.n312 VDD.n311 0.397496
R25453 VDD.n323 VDD.n322 0.344944
R25454 VDD.n3036 VDD.n3035 0.32387
R25455 VDD.n2900 VDD.n2899 0.32387
R25456 VDD.n2764 VDD.n2763 0.32387
R25457 VDD.n2628 VDD.n2627 0.32387
R25458 VDD.n2492 VDD.n2491 0.32387
R25459 VDD.n2356 VDD.n2355 0.32387
R25460 VDD.n2220 VDD.n2219 0.32387
R25461 VDD.n2084 VDD.n2083 0.32387
R25462 VDD.n1948 VDD.n1947 0.32387
R25463 VDD.n3053 VDD 0.252453
R25464 VDD.n3042 VDD 0.252453
R25465 VDD.n3148 VDD.n3147 0.226043
R25466 VDD.n3137 VDD.n3136 0.226043
R25467 VDD.n3164 VDD.n3163 0.226043
R25468 VDD.n3172 VDD.n3171 0.226043
R25469 VDD.n3212 VDD.n3211 0.226043
R25470 VDD.n3201 VDD.n3200 0.226043
R25471 VDD.n3228 VDD.n3227 0.226043
R25472 VDD.n3236 VDD.n3235 0.226043
R25473 VDD.n3109 VDD.n3108 0.226043
R25474 VDD.n3098 VDD.n3097 0.226043
R25475 VDD.n3252 VDD.n3251 0.226043
R25476 VDD.n3260 VDD.n3259 0.226043
R25477 VDD.n3363 VDD.n3362 0.226043
R25478 VDD.n3352 VDD.n3351 0.226043
R25479 VDD.n3629 VDD.n3628 0.226043
R25480 VDD.n3637 VDD.n3636 0.226043
R25481 VDD.n3070 VDD.n3069 0.226043
R25482 VDD.n3059 VDD.n3058 0.226043
R25483 VDD.n3086 VDD.n3085 0.226043
R25484 VDD.n3094 VDD.n3093 0.226043
R25485 VDD.n3657 VDD.n3656 0.226043
R25486 VDD.n3646 VDD.n3645 0.226043
R25487 VDD.n3673 VDD.n3672 0.226043
R25488 VDD.n3681 VDD.n3680 0.226043
R25489 VDD.n3053 VDD.n3052 0.226043
R25490 VDD.n3042 VDD.n3041 0.226043
R25491 VDD.n3696 VDD.n3695 0.226043
R25492 VDD.n3704 VDD.n3703 0.226043
R25493 VDD.n3128 VDD.n3127 0.226043
R25494 VDD.n3117 VDD.n3116 0.226043
R25495 VDD.n3183 VDD.n3182 0.226043
R25496 VDD.n3191 VDD.n3190 0.226043
R25497 VDD.n3717 VDD.n3716 0.226043
R25498 VDD.n3725 VDD.n3724 0.226043
R25499 VDD.n3142 VDD 0.217464
R25500 VDD.n3158 VDD 0.217464
R25501 VDD.n3206 VDD 0.217464
R25502 VDD.n3222 VDD 0.217464
R25503 VDD.n3103 VDD 0.217464
R25504 VDD.n3246 VDD 0.217464
R25505 VDD.n3357 VDD 0.217464
R25506 VDD.n3623 VDD 0.217464
R25507 VDD.n3064 VDD 0.217464
R25508 VDD.n3080 VDD 0.217464
R25509 VDD.n3651 VDD 0.217464
R25510 VDD.n3667 VDD 0.217464
R25511 VDD.n3049 VDD 0.217464
R25512 VDD.n3038 VDD 0.217464
R25513 VDD.n3690 VDD 0.217464
R25514 VDD.n3122 VDD 0.217464
R25515 VDD.n3177 VDD 0.217464
R25516 VDD.n3711 VDD 0.217464
R25517 VDD.n3150 VDD 0.1255
R25518 VDD.n3143 VDD 0.1255
R25519 VDD.n3139 VDD 0.1255
R25520 VDD.n3166 VDD 0.1255
R25521 VDD.n3159 VDD 0.1255
R25522 VDD.n3156 VDD 0.1255
R25523 VDD.n3214 VDD 0.1255
R25524 VDD.n3207 VDD 0.1255
R25525 VDD.n3203 VDD 0.1255
R25526 VDD.n3230 VDD 0.1255
R25527 VDD.n3223 VDD 0.1255
R25528 VDD.n3220 VDD 0.1255
R25529 VDD.n3111 VDD 0.1255
R25530 VDD.n3104 VDD 0.1255
R25531 VDD.n3100 VDD 0.1255
R25532 VDD.n3254 VDD 0.1255
R25533 VDD.n3247 VDD 0.1255
R25534 VDD.n3244 VDD 0.1255
R25535 VDD.n3365 VDD 0.1255
R25536 VDD.n3358 VDD 0.1255
R25537 VDD.n3354 VDD 0.1255
R25538 VDD.n3631 VDD 0.1255
R25539 VDD.n3624 VDD 0.1255
R25540 VDD.n3621 VDD 0.1255
R25541 VDD.n3072 VDD 0.1255
R25542 VDD.n3065 VDD 0.1255
R25543 VDD.n3061 VDD 0.1255
R25544 VDD.n3088 VDD 0.1255
R25545 VDD.n3081 VDD 0.1255
R25546 VDD.n3078 VDD 0.1255
R25547 VDD.n3659 VDD 0.1255
R25548 VDD.n3652 VDD 0.1255
R25549 VDD.n3648 VDD 0.1255
R25550 VDD.n3675 VDD 0.1255
R25551 VDD.n3668 VDD 0.1255
R25552 VDD.n3665 VDD 0.1255
R25553 VDD.n3052 VDD 0.1255
R25554 VDD.n3045 VDD 0.1255
R25555 VDD.n3041 VDD 0.1255
R25556 VDD.n3698 VDD 0.1255
R25557 VDD.n3691 VDD 0.1255
R25558 VDD.n3688 VDD 0.1255
R25559 VDD.n3130 VDD 0.1255
R25560 VDD.n3123 VDD 0.1255
R25561 VDD.n3119 VDD 0.1255
R25562 VDD.n3185 VDD 0.1255
R25563 VDD.n3178 VDD 0.1255
R25564 VDD.n3175 VDD 0.1255
R25565 VDD.n3719 VDD 0.1255
R25566 VDD.n3712 VDD 0.1255
R25567 VDD.n3709 VDD 0.1255
R25568 VDD.n6888 VDD 0.101043
R25569 VDD.t89 VDD.n329 0.086419
R25570 VDD.n7129 VDD.n6888 0.063
R25571 VDD.n3152 VDD.n3148 0.063
R25572 VDD.n3152 VDD.n3151 0.063
R25573 VDD.n3141 VDD.n3137 0.063
R25574 VDD.n3141 VDD.n3140 0.063
R25575 VDD.n3168 VDD.n3164 0.063
R25576 VDD.n3168 VDD.n3167 0.063
R25577 VDD.n3171 VDD.n3170 0.063
R25578 VDD.n3170 VDD.n3157 0.063
R25579 VDD.n3216 VDD.n3212 0.063
R25580 VDD.n3216 VDD.n3215 0.063
R25581 VDD.n3205 VDD.n3201 0.063
R25582 VDD.n3205 VDD.n3204 0.063
R25583 VDD.n3232 VDD.n3228 0.063
R25584 VDD.n3232 VDD.n3231 0.063
R25585 VDD.n3235 VDD.n3234 0.063
R25586 VDD.n3234 VDD.n3221 0.063
R25587 VDD.n3113 VDD.n3109 0.063
R25588 VDD.n3113 VDD.n3112 0.063
R25589 VDD.n3102 VDD.n3098 0.063
R25590 VDD.n3102 VDD.n3101 0.063
R25591 VDD.n3256 VDD.n3252 0.063
R25592 VDD.n3256 VDD.n3255 0.063
R25593 VDD.n3259 VDD.n3258 0.063
R25594 VDD.n3258 VDD.n3245 0.063
R25595 VDD.n3367 VDD.n3363 0.063
R25596 VDD.n3367 VDD.n3366 0.063
R25597 VDD.n3356 VDD.n3352 0.063
R25598 VDD.n3356 VDD.n3355 0.063
R25599 VDD.n3437 VDD.n3341 0.063
R25600 VDD.n3449 VDD.n3341 0.063
R25601 VDD.n3487 VDD.n3340 0.063
R25602 VDD.n3487 VDD.n3486 0.063
R25603 VDD.n3503 VDD.n3502 0.063
R25604 VDD.n3502 VDD.n3338 0.063
R25605 VDD.n3532 VDD.n3304 0.063
R25606 VDD.n3544 VDD.n3304 0.063
R25607 VDD.n3408 VDD.n3407 0.063
R25608 VDD.n3407 VDD.n3394 0.063
R25609 VDD.n3591 VDD.n3301 0.063
R25610 VDD.n3592 VDD.n3591 0.063
R25611 VDD.n3633 VDD.n3629 0.063
R25612 VDD.n3633 VDD.n3632 0.063
R25613 VDD.n3636 VDD.n3635 0.063
R25614 VDD.n3635 VDD.n3622 0.063
R25615 VDD.n3074 VDD.n3070 0.063
R25616 VDD.n3074 VDD.n3073 0.063
R25617 VDD.n3063 VDD.n3059 0.063
R25618 VDD.n3063 VDD.n3062 0.063
R25619 VDD.n3090 VDD.n3086 0.063
R25620 VDD.n3090 VDD.n3089 0.063
R25621 VDD.n3093 VDD.n3092 0.063
R25622 VDD.n3092 VDD.n3079 0.063
R25623 VDD.n3661 VDD.n3657 0.063
R25624 VDD.n3661 VDD.n3660 0.063
R25625 VDD.n3650 VDD.n3646 0.063
R25626 VDD.n3650 VDD.n3649 0.063
R25627 VDD.n3677 VDD.n3673 0.063
R25628 VDD.n3677 VDD.n3676 0.063
R25629 VDD.n3680 VDD.n3679 0.063
R25630 VDD.n3679 VDD.n3666 0.063
R25631 VDD.n3054 VDD.n3050 0.063
R25632 VDD.n3054 VDD.n3053 0.063
R25633 VDD.n3043 VDD.n3039 0.063
R25634 VDD.n3043 VDD.n3042 0.063
R25635 VDD.n3700 VDD.n3696 0.063
R25636 VDD.n3700 VDD.n3699 0.063
R25637 VDD.n3703 VDD.n3702 0.063
R25638 VDD.n3702 VDD.n3689 0.063
R25639 VDD.n3132 VDD.n3128 0.063
R25640 VDD.n3132 VDD.n3131 0.063
R25641 VDD.n3121 VDD.n3117 0.063
R25642 VDD.n3121 VDD.n3120 0.063
R25643 VDD.n3187 VDD.n3183 0.063
R25644 VDD.n3187 VDD.n3186 0.063
R25645 VDD.n3190 VDD.n3189 0.063
R25646 VDD.n3189 VDD.n3176 0.063
R25647 VDD.n3721 VDD.n3717 0.063
R25648 VDD.n3721 VDD.n3720 0.063
R25649 VDD.n3724 VDD.n3723 0.063
R25650 VDD.n3723 VDD.n3710 0.063
R25651 VDD.n3727 VDD.n3036 0.063
R25652 VDD.n3739 VDD.n3727 0.063
R25653 VDD.n2901 VDD.n2900 0.063
R25654 VDD.n2913 VDD.n2901 0.063
R25655 VDD.n2765 VDD.n2764 0.063
R25656 VDD.n2777 VDD.n2765 0.063
R25657 VDD.n2629 VDD.n2628 0.063
R25658 VDD.n2641 VDD.n2629 0.063
R25659 VDD.n2493 VDD.n2492 0.063
R25660 VDD.n2505 VDD.n2493 0.063
R25661 VDD.n2357 VDD.n2356 0.063
R25662 VDD.n2369 VDD.n2357 0.063
R25663 VDD.n2221 VDD.n2220 0.063
R25664 VDD.n2233 VDD.n2221 0.063
R25665 VDD.n2085 VDD.n2084 0.063
R25666 VDD.n2097 VDD.n2085 0.063
R25667 VDD.n1949 VDD.n1948 0.063
R25668 VDD.n1961 VDD.n1949 0.063
R25669 VDD.n3581 VDD.n3303 0.0620385
R25670 VDD.n3581 VDD.n3580 0.0620385
R25671 VDD VDD.n7128 0.0532344
R25672 VDD.n3196 VDD 0.0477973
R25673 VDD.n3195 VDD 0.0249565
R25674 VDD.n3589 VDD.n3588 0.024
R25675 VDD.n3584 VDD.n3583 0.024
R25676 VDD.n3495 VDD.n3494 0.024
R25677 VDD.n3500 VDD.n3499 0.024
R25678 VDD.n3490 VDD.n3489 0.024
R25679 VDD.n3400 VDD.n3399 0.024
R25680 VDD.n3405 VDD.n3404 0.024
R25681 VDD.n3144 VDD.n3143 0.0216397
R25682 VDD.n3144 VDD 0.0216397
R25683 VDD.n3160 VDD.n3159 0.0216397
R25684 VDD.n3160 VDD 0.0216397
R25685 VDD.n3208 VDD.n3207 0.0216397
R25686 VDD.n3208 VDD 0.0216397
R25687 VDD.n3224 VDD.n3223 0.0216397
R25688 VDD.n3224 VDD 0.0216397
R25689 VDD.n3105 VDD.n3104 0.0216397
R25690 VDD.n3105 VDD 0.0216397
R25691 VDD.n3248 VDD.n3247 0.0216397
R25692 VDD.n3248 VDD 0.0216397
R25693 VDD.n3359 VDD.n3358 0.0216397
R25694 VDD.n3359 VDD 0.0216397
R25695 VDD.n3625 VDD.n3624 0.0216397
R25696 VDD.n3625 VDD 0.0216397
R25697 VDD.n3066 VDD.n3065 0.0216397
R25698 VDD.n3066 VDD 0.0216397
R25699 VDD.n3082 VDD.n3081 0.0216397
R25700 VDD.n3082 VDD 0.0216397
R25701 VDD.n3653 VDD.n3652 0.0216397
R25702 VDD.n3653 VDD 0.0216397
R25703 VDD.n3669 VDD.n3668 0.0216397
R25704 VDD.n3669 VDD 0.0216397
R25705 VDD.n3052 VDD.n3051 0.0216397
R25706 VDD.n3051 VDD 0.0216397
R25707 VDD.n3041 VDD.n3040 0.0216397
R25708 VDD.n3040 VDD 0.0216397
R25709 VDD.n3692 VDD.n3691 0.0216397
R25710 VDD.n3692 VDD 0.0216397
R25711 VDD.n3124 VDD.n3123 0.0216397
R25712 VDD.n3124 VDD 0.0216397
R25713 VDD.n3179 VDD.n3178 0.0216397
R25714 VDD.n3179 VDD 0.0216397
R25715 VDD.n3713 VDD.n3712 0.0216397
R25716 VDD.n3713 VDD 0.0216397
R25717 VDD.n3397 VDD 0.0204394
R25718 VDD.n3586 VDD 0.0204394
R25719 VDD VDD.n3302 0.0204394
R25720 VDD VDD.n3497 0.0204394
R25721 VDD.n3492 VDD 0.0204394
R25722 VDD VDD.n3339 0.0204394
R25723 VDD VDD.n3402 0.0204394
R25724 VDD VDD.n3195 0.0157027
R25725 VDD.n3150 VDD.n3149 0.0107679
R25726 VDD.n3149 VDD 0.0107679
R25727 VDD.n3139 VDD.n3138 0.0107679
R25728 VDD.n3138 VDD 0.0107679
R25729 VDD.n3166 VDD.n3165 0.0107679
R25730 VDD.n3165 VDD 0.0107679
R25731 VDD.n3156 VDD.n3155 0.0107679
R25732 VDD.n3155 VDD 0.0107679
R25733 VDD.n3214 VDD.n3213 0.0107679
R25734 VDD.n3213 VDD 0.0107679
R25735 VDD.n3203 VDD.n3202 0.0107679
R25736 VDD.n3202 VDD 0.0107679
R25737 VDD.n3230 VDD.n3229 0.0107679
R25738 VDD.n3229 VDD 0.0107679
R25739 VDD.n3220 VDD.n3219 0.0107679
R25740 VDD.n3219 VDD 0.0107679
R25741 VDD.n3111 VDD.n3110 0.0107679
R25742 VDD.n3110 VDD 0.0107679
R25743 VDD.n3100 VDD.n3099 0.0107679
R25744 VDD.n3099 VDD 0.0107679
R25745 VDD.n3254 VDD.n3253 0.0107679
R25746 VDD.n3253 VDD 0.0107679
R25747 VDD.n3244 VDD.n3243 0.0107679
R25748 VDD.n3243 VDD 0.0107679
R25749 VDD.n3365 VDD.n3364 0.0107679
R25750 VDD.n3364 VDD 0.0107679
R25751 VDD.n3354 VDD.n3353 0.0107679
R25752 VDD.n3353 VDD 0.0107679
R25753 VDD.n3631 VDD.n3630 0.0107679
R25754 VDD.n3630 VDD 0.0107679
R25755 VDD.n3621 VDD.n3620 0.0107679
R25756 VDD.n3620 VDD 0.0107679
R25757 VDD.n3072 VDD.n3071 0.0107679
R25758 VDD.n3071 VDD 0.0107679
R25759 VDD.n3061 VDD.n3060 0.0107679
R25760 VDD.n3060 VDD 0.0107679
R25761 VDD.n3088 VDD.n3087 0.0107679
R25762 VDD.n3087 VDD 0.0107679
R25763 VDD.n3078 VDD.n3077 0.0107679
R25764 VDD.n3077 VDD 0.0107679
R25765 VDD.n3659 VDD.n3658 0.0107679
R25766 VDD.n3658 VDD 0.0107679
R25767 VDD.n3648 VDD.n3647 0.0107679
R25768 VDD.n3647 VDD 0.0107679
R25769 VDD.n3675 VDD.n3674 0.0107679
R25770 VDD.n3674 VDD 0.0107679
R25771 VDD.n3665 VDD.n3664 0.0107679
R25772 VDD.n3664 VDD 0.0107679
R25773 VDD.n3045 VDD.n3044 0.0107679
R25774 VDD.n3044 VDD 0.0107679
R25775 VDD.n3698 VDD.n3697 0.0107679
R25776 VDD.n3697 VDD 0.0107679
R25777 VDD.n3688 VDD.n3687 0.0107679
R25778 VDD.n3687 VDD 0.0107679
R25779 VDD.n3130 VDD.n3129 0.0107679
R25780 VDD.n3129 VDD 0.0107679
R25781 VDD.n3119 VDD.n3118 0.0107679
R25782 VDD.n3118 VDD 0.0107679
R25783 VDD.n3185 VDD.n3184 0.0107679
R25784 VDD.n3184 VDD 0.0107679
R25785 VDD.n3175 VDD.n3174 0.0107679
R25786 VDD.n3174 VDD 0.0107679
R25787 VDD.n3719 VDD.n3718 0.0107679
R25788 VDD.n3718 VDD 0.0107679
R25789 VDD.n3709 VDD.n3708 0.0107679
R25790 VDD.n3708 VDD 0.0107679
R25791 VDD.n7129 VDD 0.0102656
R25792 VDD.n3394 VDD 0.00534007
R25793 VDD.n3449 VDD.n3342 0.00534007
R25794 VDD VDD.n3449 0.00534007
R25795 VDD.n3486 VDD.n3450 0.00534007
R25796 VDD.n3486 VDD 0.00534007
R25797 VDD.n3451 VDD.n3338 0.00534007
R25798 VDD.n3338 VDD 0.00534007
R25799 VDD.n3544 VDD.n3305 0.00534007
R25800 VDD VDD.n3544 0.00534007
R25801 VDD.n3580 VDD.n3545 0.00534007
R25802 VDD.n3580 VDD 0.00534007
R25803 VDD.n3592 VDD.n3300 0.00534007
R25804 VDD.n3592 VDD 0.00534007
R25805 VDD.n3146 VDD 0.00441667
R25806 VDD.n3162 VDD 0.00441667
R25807 VDD.n3210 VDD 0.00441667
R25808 VDD.n3226 VDD 0.00441667
R25809 VDD.n3107 VDD 0.00441667
R25810 VDD.n3250 VDD 0.00441667
R25811 VDD.n3361 VDD 0.00441667
R25812 VDD.n3396 VDD 0.00441667
R25813 VDD.n3587 VDD 0.00441667
R25814 VDD.n3585 VDD 0.00441667
R25815 VDD.n3493 VDD 0.00441667
R25816 VDD.n3498 VDD 0.00441667
R25817 VDD.n3491 VDD 0.00441667
R25818 VDD.n3398 VDD 0.00441667
R25819 VDD.n3403 VDD 0.00441667
R25820 VDD.n3627 VDD 0.00441667
R25821 VDD.n3068 VDD 0.00441667
R25822 VDD.n3084 VDD 0.00441667
R25823 VDD.n3655 VDD 0.00441667
R25824 VDD.n3671 VDD 0.00441667
R25825 VDD.n3047 VDD 0.00441667
R25826 VDD.n3694 VDD 0.00441667
R25827 VDD.n3126 VDD 0.00441667
R25828 VDD.n3181 VDD 0.00441667
R25829 VDD.n3715 VDD 0.00441667
R25830 VDD VDD.n3146 0.00406061
R25831 VDD VDD.n3162 0.00406061
R25832 VDD VDD.n3210 0.00406061
R25833 VDD VDD.n3226 0.00406061
R25834 VDD VDD.n3107 0.00406061
R25835 VDD VDD.n3250 0.00406061
R25836 VDD VDD.n3361 0.00406061
R25837 VDD VDD.n3396 0.00406061
R25838 VDD.n3587 VDD 0.00406061
R25839 VDD VDD.n3585 0.00406061
R25840 VDD.n3493 VDD 0.00406061
R25841 VDD.n3498 VDD 0.00406061
R25842 VDD VDD.n3491 0.00406061
R25843 VDD.n3398 VDD 0.00406061
R25844 VDD.n3403 VDD 0.00406061
R25845 VDD VDD.n3627 0.00406061
R25846 VDD VDD.n3068 0.00406061
R25847 VDD VDD.n3084 0.00406061
R25848 VDD VDD.n3655 0.00406061
R25849 VDD VDD.n3671 0.00406061
R25850 VDD.n3047 VDD 0.00406061
R25851 VDD VDD.n3694 0.00406061
R25852 VDD VDD.n3126 0.00406061
R25853 VDD VDD.n3181 0.00406061
R25854 VDD VDD.n3715 0.00406061
R25855 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.t1 169.46
R25856 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C.t3 167.809
R25857 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.t0 167.809
R25858 D_FlipFlop_6.3-input-nand_2.C.t5 D_FlipFlop_6.3-input-nand_2.C.n13 167.226
R25859 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C.t7 150.273
R25860 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.t5 150.273
R25861 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C.t6 73.6406
R25862 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C.t4 73.6304
R25863 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C.t2 60.4568
R25864 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C.n7 12.3891
R25865 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.n11 11.4489
R25866 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C 1.68257
R25867 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C.n2 1.38365
R25868 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C.n0 1.19615
R25869 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C.n5 1.1717
R25870 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C 1.08448
R25871 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C 0.932141
R25872 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C 0.720633
R25873 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C.n12 0.280391
R25874 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C 0.217464
R25875 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C 0.1255
R25876 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C 0.1255
R25877 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C 0.1255
R25878 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C.n9 0.0874565
R25879 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C.n6 0.063
R25880 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C 0.063
R25881 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C.n8 0.063
R25882 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C.n3 0.063
R25883 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.n10 0.0435206
R25884 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.n1 0.0216397
R25885 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.C.n14 0.0216397
R25886 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C.n4 0.0107679
R25887 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C 0.0107679
R25888 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 169.46
R25889 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 167.809
R25890 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 167.809
R25891 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 167.226
R25892 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 150.273
R25893 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 150.273
R25894 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 73.6406
R25895 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 73.6304
R25896 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 60.3943
R25897 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 12.3891
R25898 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 11.4489
R25899 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 1.68257
R25900 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 1.38365
R25901 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 1.19615
R25902 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 1.1717
R25903 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 1.08448
R25904 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.932141
R25905 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.720633
R25906 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 0.280391
R25907 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.217464
R25908 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R25909 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R25910 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R25911 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 0.0874565
R25912 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 0.063
R25913 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.063
R25914 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 0.063
R25915 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 0.063
R25916 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 0.0435206
R25917 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 0.0216397
R25918 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 0.0216397
R25919 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 0.0107679
R25920 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.0107679
R25921 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 169.46
R25922 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 168.089
R25923 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 167.809
R25924 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 150.293
R25925 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 73.6304
R25926 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 60.4568
R25927 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 12.0358
R25928 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 11.4489
R25929 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.981478
R25930 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 0.788543
R25931 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.769522
R25932 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 0.720633
R25933 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 0.682565
R25934 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.580578
R25935 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 0.55213
R25936 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 0.470609
R25937 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.447191
R25938 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.428234
R25939 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.1255
R25940 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.1255
R25941 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 0.063
R25942 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 0.063
R25943 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.063
R25944 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 0.063
R25945 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 0.063
R25946 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 0.0435206
R25947 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 0.0107679
R25948 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.0107679
R25949 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z.t3 168.635
R25950 CDAC8_0.switch_8.Z CDAC8_0.switch_8.Z.t0 168.571
R25951 CDAC8_0.switch_8.Z.n0 CDAC8_0.switch_8.Z.t1 60.321
R25952 CDAC8_0.switch_8.Z.n0 CDAC8_0.switch_8.Z.t2 60.321
R25953 CDAC8_0.switch_8.Z.n20 CDAC8_0.switch_8.Z.n19 11.3205
R25954 CDAC8_0.switch_8.Z.n15 CDAC8_0.switch_8.Z.n14 5.49497
R25955 CDAC8_0.switch_8.Z.n19 CDAC8_0.switch_8.Z.n3 2.98587
R25956 CDAC8_0.switch_8.Z.n19 CDAC8_0.switch_8.Z.n18 2.5049
R25957 CDAC8_0.switch_8.Z.n2 CDAC8_0.switch_8.Z 1.36463
R25958 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z.n21 1.04126
R25959 CDAC8_0.switch_8.Z.n21 CDAC8_0.switch_8.Z 0.838391
R25960 CDAC8_0.switch_8.Z.n4 CDAC8_0.switch_8.Z.t4 0.77316
R25961 CDAC8_0.switch_8.Z.n10 CDAC8_0.switch_8.Z.t12 0.77316
R25962 CDAC8_0.switch_8.Z.n3 CDAC8_0.switch_8.Z.t14 0.658247
R25963 CDAC8_0.switch_8.Z.n18 CDAC8_0.switch_8.Z.t6 0.658247
R25964 CDAC8_0.switch_8.Z.n8 CDAC8_0.switch_8.Z.t13 0.611304
R25965 CDAC8_0.switch_8.Z.n9 CDAC8_0.switch_8.Z.t18 0.611304
R25966 CDAC8_0.switch_8.Z.n17 CDAC8_0.switch_8.Z.t5 0.611304
R25967 CDAC8_0.switch_8.Z.n16 CDAC8_0.switch_8.Z.t11 0.611304
R25968 CDAC8_0.switch_8.Z.n7 CDAC8_0.switch_8.Z.t9 0.611304
R25969 CDAC8_0.switch_8.Z.n6 CDAC8_0.switch_8.Z.t15 0.611304
R25970 CDAC8_0.switch_8.Z.n5 CDAC8_0.switch_8.Z.t19 0.611304
R25971 CDAC8_0.switch_8.Z.n4 CDAC8_0.switch_8.Z.t17 0.611304
R25972 CDAC8_0.switch_8.Z.n13 CDAC8_0.switch_8.Z.t16 0.611304
R25973 CDAC8_0.switch_8.Z.n12 CDAC8_0.switch_8.Z.t7 0.611304
R25974 CDAC8_0.switch_8.Z.n11 CDAC8_0.switch_8.Z.t10 0.611304
R25975 CDAC8_0.switch_8.Z.n10 CDAC8_0.switch_8.Z.t8 0.611304
R25976 CDAC8_0.switch_8.Z.n2 CDAC8_0.switch_8.Z.n1 0.405391
R25977 CDAC8_0.switch_8.Z.n1 CDAC8_0.switch_8.Z 0.259656
R25978 CDAC8_0.switch_8.Z.n17 CDAC8_0.switch_8.Z.n16 0.162356
R25979 CDAC8_0.switch_8.Z.n7 CDAC8_0.switch_8.Z.n6 0.162356
R25980 CDAC8_0.switch_8.Z.n6 CDAC8_0.switch_8.Z.n5 0.162356
R25981 CDAC8_0.switch_8.Z.n5 CDAC8_0.switch_8.Z.n4 0.162356
R25982 CDAC8_0.switch_8.Z.n9 CDAC8_0.switch_8.Z.n8 0.162356
R25983 CDAC8_0.switch_8.Z.n13 CDAC8_0.switch_8.Z.n12 0.162356
R25984 CDAC8_0.switch_8.Z.n12 CDAC8_0.switch_8.Z.n11 0.162356
R25985 CDAC8_0.switch_8.Z.n11 CDAC8_0.switch_8.Z.n10 0.162356
R25986 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z 0.1255
R25987 CDAC8_0.switch_8.Z.n18 CDAC8_0.switch_8.Z.n17 0.115412
R25988 CDAC8_0.switch_8.Z.n8 CDAC8_0.switch_8.Z.n3 0.115412
R25989 CDAC8_0.switch_8.Z.n15 CDAC8_0.switch_8.Z.n7 0.0845094
R25990 CDAC8_0.switch_8.Z.n14 CDAC8_0.switch_8.Z.n13 0.0845094
R25991 CDAC8_0.switch_8.Z.n21 CDAC8_0.switch_8.Z.n20 0.0805781
R25992 CDAC8_0.switch_8.Z.n16 CDAC8_0.switch_8.Z.n15 0.0783469
R25993 CDAC8_0.switch_8.Z.n14 CDAC8_0.switch_8.Z.n9 0.0783469
R25994 CDAC8_0.switch_8.Z.n20 CDAC8_0.switch_8.Z.n2 0.063
R25995 CDAC8_0.switch_8.Z CDAC8_0.switch_8.Z.n22 0.063
R25996 CDAC8_0.switch_8.Z.n1 CDAC8_0.switch_8.Z.n0 0.0188121
R25997 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 179.256
R25998 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 168.089
R25999 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 150.293
R26000 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 73.6304
R26001 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 60.4568
R26002 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 12.0358
R26003 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.981478
R26004 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 0.788543
R26005 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.769522
R26006 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.720633
R26007 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 0.682565
R26008 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.580578
R26009 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 0.55213
R26010 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 0.470609
R26011 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.447191
R26012 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.428234
R26013 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1255
R26014 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1255
R26015 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 0.063
R26016 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 0.063
R26017 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 0.063
R26018 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 0.063
R26019 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 0.063
R26020 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 0.0435206
R26021 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 0.0107679
R26022 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.0107679
R26023 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.t2 168.548
R26024 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.t0 168.548
R26025 CDAC8_0.switch_6.Z.n0 CDAC8_0.switch_6.Z.t1 60.321
R26026 CDAC8_0.switch_6.Z.n0 CDAC8_0.switch_6.Z.t3 60.321
R26027 CDAC8_0.switch_6.Z.n102 CDAC8_0.switch_6.Z.n101 22.979
R26028 CDAC8_0.switch_6.Z.n124 CDAC8_0.switch_6.Z.n123 11.3711
R26029 CDAC8_0.switch_6.Z.n123 CDAC8_0.switch_6.Z.n3 11.3479
R26030 CDAC8_0.switch_6.Z.n123 CDAC8_0.switch_6.Z.n122 10.8669
R26031 CDAC8_0.switch_6.Z.n54 CDAC8_0.switch_6.Z.n53 4.99363
R26032 CDAC8_0.switch_6.Z.n57 CDAC8_0.switch_6.Z.n56 4.99363
R26033 CDAC8_0.switch_6.Z.n65 CDAC8_0.switch_6.Z.n64 4.99363
R26034 CDAC8_0.switch_6.Z.n70 CDAC8_0.switch_6.Z.n69 4.99363
R26035 CDAC8_0.switch_6.Z.n73 CDAC8_0.switch_6.Z.n72 4.99363
R26036 CDAC8_0.switch_6.Z.n76 CDAC8_0.switch_6.Z.n75 4.99363
R26037 CDAC8_0.switch_6.Z.n79 CDAC8_0.switch_6.Z.n78 4.99363
R26038 CDAC8_0.switch_6.Z.n83 CDAC8_0.switch_6.Z.n82 4.99363
R26039 CDAC8_0.switch_6.Z.n85 CDAC8_0.switch_6.Z.n43 4.99363
R26040 CDAC8_0.switch_6.Z.n9 CDAC8_0.switch_6.Z.n8 4.99363
R26041 CDAC8_0.switch_6.Z.n12 CDAC8_0.switch_6.Z.n11 4.99363
R26042 CDAC8_0.switch_6.Z.n15 CDAC8_0.switch_6.Z.n14 4.99363
R26043 CDAC8_0.switch_6.Z.n19 CDAC8_0.switch_6.Z.n18 4.99363
R26044 CDAC8_0.switch_6.Z.n119 CDAC8_0.switch_6.Z.n118 4.99363
R26045 CDAC8_0.switch_6.Z.n116 CDAC8_0.switch_6.Z.n115 4.99363
R26046 CDAC8_0.switch_6.Z.n113 CDAC8_0.switch_6.Z.n112 4.99363
R26047 CDAC8_0.switch_6.Z.n110 CDAC8_0.switch_6.Z.n109 4.99363
R26048 CDAC8_0.switch_6.Z.n107 CDAC8_0.switch_6.Z.n106 4.99363
R26049 CDAC8_0.switch_6.Z.n104 CDAC8_0.switch_6.Z.n103 4.99363
R26050 CDAC8_0.switch_6.Z.n41 CDAC8_0.switch_6.Z.n40 4.99363
R26051 CDAC8_0.switch_6.Z.n38 CDAC8_0.switch_6.Z.n37 4.99363
R26052 CDAC8_0.switch_6.Z.n35 CDAC8_0.switch_6.Z.n34 4.99363
R26053 CDAC8_0.switch_6.Z.n32 CDAC8_0.switch_6.Z.n31 4.99363
R26054 CDAC8_0.switch_6.Z.n99 CDAC8_0.switch_6.Z.n98 4.99363
R26055 CDAC8_0.switch_6.Z.n96 CDAC8_0.switch_6.Z.n95 4.99363
R26056 CDAC8_0.switch_6.Z.n93 CDAC8_0.switch_6.Z.n92 4.99363
R26057 CDAC8_0.switch_6.Z.n90 CDAC8_0.switch_6.Z.n89 4.99363
R26058 CDAC8_0.switch_6.Z.n122 CDAC8_0.switch_6.Z.n4 4.61363
R26059 CDAC8_0.switch_6.Z.n62 CDAC8_0.switch_6.Z.n3 4.61363
R26060 CDAC8_0.switch_6.Z.n60 CDAC8_0.switch_6.Z.n59 3.9471
R26061 CDAC8_0.switch_6.Z.n2 CDAC8_0.switch_6.Z.n1 1.58202
R26062 CDAC8_0.switch_6.Z.n32 CDAC8_0.switch_6.Z.t5 0.726216
R26063 CDAC8_0.switch_6.Z.n31 CDAC8_0.switch_6.Z.t37 0.726216
R26064 CDAC8_0.switch_6.Z.n89 CDAC8_0.switch_6.Z.t50 0.726216
R26065 CDAC8_0.switch_6.Z.n90 CDAC8_0.switch_6.Z.t36 0.726216
R26066 CDAC8_0.switch_6.Z.n54 CDAC8_0.switch_6.Z.t31 0.658247
R26067 CDAC8_0.switch_6.Z.n53 CDAC8_0.switch_6.Z.t47 0.658247
R26068 CDAC8_0.switch_6.Z.n8 CDAC8_0.switch_6.Z.t32 0.658247
R26069 CDAC8_0.switch_6.Z.n9 CDAC8_0.switch_6.Z.t63 0.658247
R26070 CDAC8_0.switch_6.Z.n55 CDAC8_0.switch_6.Z.t28 0.611304
R26071 CDAC8_0.switch_6.Z.n51 CDAC8_0.switch_6.Z.t44 0.611304
R26072 CDAC8_0.switch_6.Z.n61 CDAC8_0.switch_6.Z.t40 0.611304
R26073 CDAC8_0.switch_6.Z.n63 CDAC8_0.switch_6.Z.t66 0.611304
R26074 CDAC8_0.switch_6.Z.n49 CDAC8_0.switch_6.Z.t11 0.611304
R26075 CDAC8_0.switch_6.Z.n71 CDAC8_0.switch_6.Z.t8 0.611304
R26076 CDAC8_0.switch_6.Z.n47 CDAC8_0.switch_6.Z.t19 0.611304
R26077 CDAC8_0.switch_6.Z.n77 CDAC8_0.switch_6.Z.t16 0.611304
R26078 CDAC8_0.switch_6.Z.n45 CDAC8_0.switch_6.Z.t48 0.611304
R26079 CDAC8_0.switch_6.Z.n84 CDAC8_0.switch_6.Z.t57 0.611304
R26080 CDAC8_0.switch_6.Z.n86 CDAC8_0.switch_6.Z.t55 0.611304
R26081 CDAC8_0.switch_6.Z.n97 CDAC8_0.switch_6.Z.t64 0.611304
R26082 CDAC8_0.switch_6.Z.n87 CDAC8_0.switch_6.Z.t26 0.611304
R26083 CDAC8_0.switch_6.Z.n91 CDAC8_0.switch_6.Z.t24 0.611304
R26084 CDAC8_0.switch_6.Z.n52 CDAC8_0.switch_6.Z.t43 0.611304
R26085 CDAC8_0.switch_6.Z.n58 CDAC8_0.switch_6.Z.t54 0.611304
R26086 CDAC8_0.switch_6.Z.n50 CDAC8_0.switch_6.Z.t52 0.611304
R26087 CDAC8_0.switch_6.Z.n66 CDAC8_0.switch_6.Z.t14 0.611304
R26088 CDAC8_0.switch_6.Z.n68 CDAC8_0.switch_6.Z.t21 0.611304
R26089 CDAC8_0.switch_6.Z.n48 CDAC8_0.switch_6.Z.t18 0.611304
R26090 CDAC8_0.switch_6.Z.n74 CDAC8_0.switch_6.Z.t35 0.611304
R26091 CDAC8_0.switch_6.Z.n46 CDAC8_0.switch_6.Z.t30 0.611304
R26092 CDAC8_0.switch_6.Z.n80 CDAC8_0.switch_6.Z.t60 0.611304
R26093 CDAC8_0.switch_6.Z.n81 CDAC8_0.switch_6.Z.t6 0.611304
R26094 CDAC8_0.switch_6.Z.n7 CDAC8_0.switch_6.Z.t29 0.611304
R26095 CDAC8_0.switch_6.Z.n13 CDAC8_0.switch_6.Z.t45 0.611304
R26096 CDAC8_0.switch_6.Z.n5 CDAC8_0.switch_6.Z.t41 0.611304
R26097 CDAC8_0.switch_6.Z.n20 CDAC8_0.switch_6.Z.t67 0.611304
R26098 CDAC8_0.switch_6.Z.n120 CDAC8_0.switch_6.Z.t12 0.611304
R26099 CDAC8_0.switch_6.Z.n21 CDAC8_0.switch_6.Z.t9 0.611304
R26100 CDAC8_0.switch_6.Z.n114 CDAC8_0.switch_6.Z.t20 0.611304
R26101 CDAC8_0.switch_6.Z.n24 CDAC8_0.switch_6.Z.t17 0.611304
R26102 CDAC8_0.switch_6.Z.n108 CDAC8_0.switch_6.Z.t49 0.611304
R26103 CDAC8_0.switch_6.Z.n26 CDAC8_0.switch_6.Z.t58 0.611304
R26104 CDAC8_0.switch_6.Z.n42 CDAC8_0.switch_6.Z.t56 0.611304
R26105 CDAC8_0.switch_6.Z.n28 CDAC8_0.switch_6.Z.t65 0.611304
R26106 CDAC8_0.switch_6.Z.n36 CDAC8_0.switch_6.Z.t27 0.611304
R26107 CDAC8_0.switch_6.Z.n30 CDAC8_0.switch_6.Z.t25 0.611304
R26108 CDAC8_0.switch_6.Z.n10 CDAC8_0.switch_6.Z.t62 0.611304
R26109 CDAC8_0.switch_6.Z.n6 CDAC8_0.switch_6.Z.t10 0.611304
R26110 CDAC8_0.switch_6.Z.n16 CDAC8_0.switch_6.Z.t7 0.611304
R26111 CDAC8_0.switch_6.Z.n17 CDAC8_0.switch_6.Z.t34 0.611304
R26112 CDAC8_0.switch_6.Z.n22 CDAC8_0.switch_6.Z.t46 0.611304
R26113 CDAC8_0.switch_6.Z.n117 CDAC8_0.switch_6.Z.t42 0.611304
R26114 CDAC8_0.switch_6.Z.n23 CDAC8_0.switch_6.Z.t53 0.611304
R26115 CDAC8_0.switch_6.Z.n111 CDAC8_0.switch_6.Z.t51 0.611304
R26116 CDAC8_0.switch_6.Z.n25 CDAC8_0.switch_6.Z.t15 0.611304
R26117 CDAC8_0.switch_6.Z.n105 CDAC8_0.switch_6.Z.t23 0.611304
R26118 CDAC8_0.switch_6.Z.n27 CDAC8_0.switch_6.Z.t22 0.611304
R26119 CDAC8_0.switch_6.Z.n39 CDAC8_0.switch_6.Z.t33 0.611304
R26120 CDAC8_0.switch_6.Z.n29 CDAC8_0.switch_6.Z.t61 0.611304
R26121 CDAC8_0.switch_6.Z.n33 CDAC8_0.switch_6.Z.t59 0.611304
R26122 CDAC8_0.switch_6.Z.n100 CDAC8_0.switch_6.Z.t4 0.611304
R26123 CDAC8_0.switch_6.Z.n44 CDAC8_0.switch_6.Z.t13 0.611304
R26124 CDAC8_0.switch_6.Z.n94 CDAC8_0.switch_6.Z.t39 0.611304
R26125 CDAC8_0.switch_6.Z.n88 CDAC8_0.switch_6.Z.t38 0.611304
R26126 CDAC8_0.switch_6.Z.n122 CDAC8_0.switch_6.Z.n121 0.3805
R26127 CDAC8_0.switch_6.Z.n67 CDAC8_0.switch_6.Z.n3 0.3805
R26128 CDAC8_0.switch_6.Z.n1 CDAC8_0.switch_6.Z 0.259656
R26129 CDAC8_0.switch_6.Z.n2 CDAC8_0.switch_6.Z 0.188
R26130 CDAC8_0.switch_6.Z.n10 CDAC8_0.switch_6.Z.n9 0.115412
R26131 CDAC8_0.switch_6.Z.n11 CDAC8_0.switch_6.Z.n6 0.115412
R26132 CDAC8_0.switch_6.Z.n16 CDAC8_0.switch_6.Z.n15 0.115412
R26133 CDAC8_0.switch_6.Z.n18 CDAC8_0.switch_6.Z.n17 0.115412
R26134 CDAC8_0.switch_6.Z.n22 CDAC8_0.switch_6.Z.n4 0.115412
R26135 CDAC8_0.switch_6.Z.n118 CDAC8_0.switch_6.Z.n117 0.115412
R26136 CDAC8_0.switch_6.Z.n116 CDAC8_0.switch_6.Z.n23 0.115412
R26137 CDAC8_0.switch_6.Z.n112 CDAC8_0.switch_6.Z.n111 0.115412
R26138 CDAC8_0.switch_6.Z.n110 CDAC8_0.switch_6.Z.n25 0.115412
R26139 CDAC8_0.switch_6.Z.n106 CDAC8_0.switch_6.Z.n105 0.115412
R26140 CDAC8_0.switch_6.Z.n104 CDAC8_0.switch_6.Z.n27 0.115412
R26141 CDAC8_0.switch_6.Z.n40 CDAC8_0.switch_6.Z.n39 0.115412
R26142 CDAC8_0.switch_6.Z.n38 CDAC8_0.switch_6.Z.n29 0.115412
R26143 CDAC8_0.switch_6.Z.n34 CDAC8_0.switch_6.Z.n33 0.115412
R26144 CDAC8_0.switch_6.Z.n8 CDAC8_0.switch_6.Z.n7 0.115412
R26145 CDAC8_0.switch_6.Z.n13 CDAC8_0.switch_6.Z.n12 0.115412
R26146 CDAC8_0.switch_6.Z.n14 CDAC8_0.switch_6.Z.n5 0.115412
R26147 CDAC8_0.switch_6.Z.n20 CDAC8_0.switch_6.Z.n19 0.115412
R26148 CDAC8_0.switch_6.Z.n121 CDAC8_0.switch_6.Z.n120 0.115412
R26149 CDAC8_0.switch_6.Z.n119 CDAC8_0.switch_6.Z.n21 0.115412
R26150 CDAC8_0.switch_6.Z.n115 CDAC8_0.switch_6.Z.n114 0.115412
R26151 CDAC8_0.switch_6.Z.n113 CDAC8_0.switch_6.Z.n24 0.115412
R26152 CDAC8_0.switch_6.Z.n109 CDAC8_0.switch_6.Z.n108 0.115412
R26153 CDAC8_0.switch_6.Z.n107 CDAC8_0.switch_6.Z.n26 0.115412
R26154 CDAC8_0.switch_6.Z.n41 CDAC8_0.switch_6.Z.n28 0.115412
R26155 CDAC8_0.switch_6.Z.n37 CDAC8_0.switch_6.Z.n36 0.115412
R26156 CDAC8_0.switch_6.Z.n35 CDAC8_0.switch_6.Z.n30 0.115412
R26157 CDAC8_0.switch_6.Z.n53 CDAC8_0.switch_6.Z.n52 0.115412
R26158 CDAC8_0.switch_6.Z.n58 CDAC8_0.switch_6.Z.n57 0.115412
R26159 CDAC8_0.switch_6.Z.n59 CDAC8_0.switch_6.Z.n50 0.115412
R26160 CDAC8_0.switch_6.Z.n66 CDAC8_0.switch_6.Z.n65 0.115412
R26161 CDAC8_0.switch_6.Z.n68 CDAC8_0.switch_6.Z.n67 0.115412
R26162 CDAC8_0.switch_6.Z.n69 CDAC8_0.switch_6.Z.n48 0.115412
R26163 CDAC8_0.switch_6.Z.n74 CDAC8_0.switch_6.Z.n73 0.115412
R26164 CDAC8_0.switch_6.Z.n75 CDAC8_0.switch_6.Z.n46 0.115412
R26165 CDAC8_0.switch_6.Z.n80 CDAC8_0.switch_6.Z.n79 0.115412
R26166 CDAC8_0.switch_6.Z.n82 CDAC8_0.switch_6.Z.n81 0.115412
R26167 CDAC8_0.switch_6.Z.n99 CDAC8_0.switch_6.Z.n44 0.115412
R26168 CDAC8_0.switch_6.Z.n95 CDAC8_0.switch_6.Z.n94 0.115412
R26169 CDAC8_0.switch_6.Z.n93 CDAC8_0.switch_6.Z.n88 0.115412
R26170 CDAC8_0.switch_6.Z.n55 CDAC8_0.switch_6.Z.n54 0.115412
R26171 CDAC8_0.switch_6.Z.n56 CDAC8_0.switch_6.Z.n51 0.115412
R26172 CDAC8_0.switch_6.Z.n61 CDAC8_0.switch_6.Z.n60 0.115412
R26173 CDAC8_0.switch_6.Z.n64 CDAC8_0.switch_6.Z.n63 0.115412
R26174 CDAC8_0.switch_6.Z.n62 CDAC8_0.switch_6.Z.n49 0.115412
R26175 CDAC8_0.switch_6.Z.n71 CDAC8_0.switch_6.Z.n70 0.115412
R26176 CDAC8_0.switch_6.Z.n72 CDAC8_0.switch_6.Z.n47 0.115412
R26177 CDAC8_0.switch_6.Z.n77 CDAC8_0.switch_6.Z.n76 0.115412
R26178 CDAC8_0.switch_6.Z.n78 CDAC8_0.switch_6.Z.n45 0.115412
R26179 CDAC8_0.switch_6.Z.n84 CDAC8_0.switch_6.Z.n83 0.115412
R26180 CDAC8_0.switch_6.Z.n86 CDAC8_0.switch_6.Z.n85 0.115412
R26181 CDAC8_0.switch_6.Z.n98 CDAC8_0.switch_6.Z.n97 0.115412
R26182 CDAC8_0.switch_6.Z.n96 CDAC8_0.switch_6.Z.n87 0.115412
R26183 CDAC8_0.switch_6.Z.n92 CDAC8_0.switch_6.Z.n91 0.115412
R26184 CDAC8_0.switch_6.Z.n102 CDAC8_0.switch_6.Z.n42 0.0845094
R26185 CDAC8_0.switch_6.Z.n101 CDAC8_0.switch_6.Z.n100 0.0845094
R26186 CDAC8_0.switch_6.Z.n124 CDAC8_0.switch_6.Z.n2 0.063
R26187 CDAC8_0.switch_6.Z.n11 CDAC8_0.switch_6.Z.n10 0.0474438
R26188 CDAC8_0.switch_6.Z.n15 CDAC8_0.switch_6.Z.n6 0.0474438
R26189 CDAC8_0.switch_6.Z.n18 CDAC8_0.switch_6.Z.n16 0.0474438
R26190 CDAC8_0.switch_6.Z.n17 CDAC8_0.switch_6.Z.n4 0.0474438
R26191 CDAC8_0.switch_6.Z.n118 CDAC8_0.switch_6.Z.n22 0.0474438
R26192 CDAC8_0.switch_6.Z.n117 CDAC8_0.switch_6.Z.n116 0.0474438
R26193 CDAC8_0.switch_6.Z.n112 CDAC8_0.switch_6.Z.n23 0.0474438
R26194 CDAC8_0.switch_6.Z.n111 CDAC8_0.switch_6.Z.n110 0.0474438
R26195 CDAC8_0.switch_6.Z.n106 CDAC8_0.switch_6.Z.n25 0.0474438
R26196 CDAC8_0.switch_6.Z.n105 CDAC8_0.switch_6.Z.n104 0.0474438
R26197 CDAC8_0.switch_6.Z.n40 CDAC8_0.switch_6.Z.n27 0.0474438
R26198 CDAC8_0.switch_6.Z.n39 CDAC8_0.switch_6.Z.n38 0.0474438
R26199 CDAC8_0.switch_6.Z.n34 CDAC8_0.switch_6.Z.n29 0.0474438
R26200 CDAC8_0.switch_6.Z.n33 CDAC8_0.switch_6.Z.n32 0.0474438
R26201 CDAC8_0.switch_6.Z.n12 CDAC8_0.switch_6.Z.n7 0.0474438
R26202 CDAC8_0.switch_6.Z.n14 CDAC8_0.switch_6.Z.n13 0.0474438
R26203 CDAC8_0.switch_6.Z.n19 CDAC8_0.switch_6.Z.n5 0.0474438
R26204 CDAC8_0.switch_6.Z.n121 CDAC8_0.switch_6.Z.n20 0.0474438
R26205 CDAC8_0.switch_6.Z.n120 CDAC8_0.switch_6.Z.n119 0.0474438
R26206 CDAC8_0.switch_6.Z.n115 CDAC8_0.switch_6.Z.n21 0.0474438
R26207 CDAC8_0.switch_6.Z.n114 CDAC8_0.switch_6.Z.n113 0.0474438
R26208 CDAC8_0.switch_6.Z.n109 CDAC8_0.switch_6.Z.n24 0.0474438
R26209 CDAC8_0.switch_6.Z.n108 CDAC8_0.switch_6.Z.n107 0.0474438
R26210 CDAC8_0.switch_6.Z.n103 CDAC8_0.switch_6.Z.n26 0.0474438
R26211 CDAC8_0.switch_6.Z.n42 CDAC8_0.switch_6.Z.n41 0.0474438
R26212 CDAC8_0.switch_6.Z.n37 CDAC8_0.switch_6.Z.n28 0.0474438
R26213 CDAC8_0.switch_6.Z.n36 CDAC8_0.switch_6.Z.n35 0.0474438
R26214 CDAC8_0.switch_6.Z.n31 CDAC8_0.switch_6.Z.n30 0.0474438
R26215 CDAC8_0.switch_6.Z.n57 CDAC8_0.switch_6.Z.n52 0.0474438
R26216 CDAC8_0.switch_6.Z.n59 CDAC8_0.switch_6.Z.n58 0.0474438
R26217 CDAC8_0.switch_6.Z.n65 CDAC8_0.switch_6.Z.n50 0.0474438
R26218 CDAC8_0.switch_6.Z.n67 CDAC8_0.switch_6.Z.n66 0.0474438
R26219 CDAC8_0.switch_6.Z.n69 CDAC8_0.switch_6.Z.n68 0.0474438
R26220 CDAC8_0.switch_6.Z.n73 CDAC8_0.switch_6.Z.n48 0.0474438
R26221 CDAC8_0.switch_6.Z.n75 CDAC8_0.switch_6.Z.n74 0.0474438
R26222 CDAC8_0.switch_6.Z.n79 CDAC8_0.switch_6.Z.n46 0.0474438
R26223 CDAC8_0.switch_6.Z.n82 CDAC8_0.switch_6.Z.n80 0.0474438
R26224 CDAC8_0.switch_6.Z.n81 CDAC8_0.switch_6.Z.n43 0.0474438
R26225 CDAC8_0.switch_6.Z.n100 CDAC8_0.switch_6.Z.n99 0.0474438
R26226 CDAC8_0.switch_6.Z.n95 CDAC8_0.switch_6.Z.n44 0.0474438
R26227 CDAC8_0.switch_6.Z.n94 CDAC8_0.switch_6.Z.n93 0.0474438
R26228 CDAC8_0.switch_6.Z.n89 CDAC8_0.switch_6.Z.n88 0.0474438
R26229 CDAC8_0.switch_6.Z.n56 CDAC8_0.switch_6.Z.n55 0.0474438
R26230 CDAC8_0.switch_6.Z.n60 CDAC8_0.switch_6.Z.n51 0.0474438
R26231 CDAC8_0.switch_6.Z.n64 CDAC8_0.switch_6.Z.n61 0.0474438
R26232 CDAC8_0.switch_6.Z.n63 CDAC8_0.switch_6.Z.n62 0.0474438
R26233 CDAC8_0.switch_6.Z.n70 CDAC8_0.switch_6.Z.n49 0.0474438
R26234 CDAC8_0.switch_6.Z.n72 CDAC8_0.switch_6.Z.n71 0.0474438
R26235 CDAC8_0.switch_6.Z.n76 CDAC8_0.switch_6.Z.n47 0.0474438
R26236 CDAC8_0.switch_6.Z.n78 CDAC8_0.switch_6.Z.n77 0.0474438
R26237 CDAC8_0.switch_6.Z.n83 CDAC8_0.switch_6.Z.n45 0.0474438
R26238 CDAC8_0.switch_6.Z.n85 CDAC8_0.switch_6.Z.n84 0.0474438
R26239 CDAC8_0.switch_6.Z.n98 CDAC8_0.switch_6.Z.n86 0.0474438
R26240 CDAC8_0.switch_6.Z.n97 CDAC8_0.switch_6.Z.n96 0.0474438
R26241 CDAC8_0.switch_6.Z.n92 CDAC8_0.switch_6.Z.n87 0.0474438
R26242 CDAC8_0.switch_6.Z.n91 CDAC8_0.switch_6.Z.n90 0.0474438
R26243 CDAC8_0.switch_6.Z CDAC8_0.switch_6.Z.n125 0.0454219
R26244 CDAC8_0.switch_6.Z.n103 CDAC8_0.switch_6.Z.n102 0.0314031
R26245 CDAC8_0.switch_6.Z.n101 CDAC8_0.switch_6.Z.n43 0.0314031
R26246 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.n124 0.0278438
R26247 CDAC8_0.switch_6.Z.n1 CDAC8_0.switch_6.Z.n0 0.0188121
R26248 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.t3 169.46
R26249 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout.t2 167.809
R26250 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.t0 167.809
R26251 D_FlipFlop_1.3-input-nand_2.Vout.t4 D_FlipFlop_1.3-input-nand_2.Vout.n11 167.227
R26252 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.t4 150.293
R26253 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.t7 150.273
R26254 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout.t5 73.6406
R26255 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout.t6 73.6304
R26256 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout.t1 60.3809
R26257 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout.n5 12.3891
R26258 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout.n9 11.4489
R26259 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout.n2 1.38365
R26260 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.n1 1.19615
R26261 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.n4 1.1717
R26262 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout 0.848156
R26263 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.Vout.n12 0.447191
R26264 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R26265 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout.n10 0.280391
R26266 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout.n8 0.262643
R26267 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout 0.217464
R26268 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R26269 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R26270 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R26271 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R26272 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout.n7 0.0874565
R26273 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout.n3 0.063
R26274 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout.n6 0.063
R26275 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout 0.063
R26276 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R26277 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout.n0 0.0107679
R26278 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout 0.0107679
R26279 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.t2 169.46
R26280 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.t3 167.809
R26281 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t0 167.809
R26282 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t7 167.226
R26283 D_FlipFlop_1.3-input-nand_2.C.t7 D_FlipFlop_1.3-input-nand_2.C.n10 150.273
R26284 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C.t4 150.273
R26285 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C.t6 73.6406
R26286 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C.t5 73.6304
R26287 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C.t1 60.4568
R26288 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C.n5 12.3891
R26289 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.n12 11.4489
R26290 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C 1.68257
R26291 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C.n0 1.38365
R26292 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C.n8 1.19615
R26293 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C.n3 1.1717
R26294 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C 1.08448
R26295 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C 0.932141
R26296 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.C.n14 0.720633
R26297 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.n11 0.280391
R26298 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C 0.217464
R26299 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C 0.1255
R26300 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C 0.1255
R26301 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C 0.1255
R26302 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.n7 0.0874565
R26303 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C.n4 0.063
R26304 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C 0.063
R26305 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C.n6 0.063
R26306 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C.n1 0.063
R26307 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.n13 0.0435206
R26308 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C.n9 0.0216397
R26309 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C 0.0216397
R26310 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C.n2 0.0107679
R26311 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C 0.0107679
R26312 D_FlipFlop_7.D.n76 D_FlipFlop_7.D.t16 150.273
R26313 D_FlipFlop_7.D.n82 D_FlipFlop_7.D.t7 150.273
R26314 D_FlipFlop_7.D.n62 D_FlipFlop_7.D.t13 150.273
R26315 D_FlipFlop_7.D.n68 D_FlipFlop_7.D.t3 150.273
R26316 D_FlipFlop_7.D.n48 D_FlipFlop_7.D.t29 150.273
R26317 D_FlipFlop_7.D.n54 D_FlipFlop_7.D.t22 150.273
R26318 D_FlipFlop_7.D.n34 D_FlipFlop_7.D.t17 150.273
R26319 D_FlipFlop_7.D.n40 D_FlipFlop_7.D.t8 150.273
R26320 D_FlipFlop_7.D.n20 D_FlipFlop_7.D.t11 150.273
R26321 D_FlipFlop_7.D.n26 D_FlipFlop_7.D.t32 150.273
R26322 D_FlipFlop_7.D.n7 D_FlipFlop_7.D.t30 150.273
R26323 D_FlipFlop_7.D.n13 D_FlipFlop_7.D.t23 150.273
R26324 D_FlipFlop_7.D.n102 D_FlipFlop_7.D.t18 150.273
R26325 D_FlipFlop_7.D.n108 D_FlipFlop_7.D.t9 150.273
R26326 D_FlipFlop_7.D.n89 D_FlipFlop_7.D.t12 150.273
R26327 D_FlipFlop_7.D.n95 D_FlipFlop_7.D.t35 150.273
R26328 D_FlipFlop_7.D.n74 D_FlipFlop_7.D.t5 73.6406
R26329 D_FlipFlop_7.D.n80 D_FlipFlop_7.D.t10 73.6406
R26330 D_FlipFlop_7.D.n60 D_FlipFlop_7.D.t21 73.6406
R26331 D_FlipFlop_7.D.n66 D_FlipFlop_7.D.t28 73.6406
R26332 D_FlipFlop_7.D.n46 D_FlipFlop_7.D.t19 73.6406
R26333 D_FlipFlop_7.D.n52 D_FlipFlop_7.D.t26 73.6406
R26334 D_FlipFlop_7.D.n32 D_FlipFlop_7.D.t14 73.6406
R26335 D_FlipFlop_7.D.n38 D_FlipFlop_7.D.t24 73.6406
R26336 D_FlipFlop_7.D.n18 D_FlipFlop_7.D.t31 73.6406
R26337 D_FlipFlop_7.D.n24 D_FlipFlop_7.D.t4 73.6406
R26338 D_FlipFlop_7.D.n5 D_FlipFlop_7.D.t20 73.6406
R26339 D_FlipFlop_7.D.n11 D_FlipFlop_7.D.t27 73.6406
R26340 D_FlipFlop_7.D.n100 D_FlipFlop_7.D.t15 73.6406
R26341 D_FlipFlop_7.D.n106 D_FlipFlop_7.D.t25 73.6406
R26342 D_FlipFlop_7.D.n87 D_FlipFlop_7.D.t34 73.6406
R26343 D_FlipFlop_7.D.n93 D_FlipFlop_7.D.t6 73.6406
R26344 D_FlipFlop_7.D.n1 D_FlipFlop_7.D.t1 33.6184
R26345 D_FlipFlop_7.D.n1 D_FlipFlop_7.D.t2 28.4497
R26346 D_FlipFlop_7.D.n86 D_FlipFlop_7.D.n85 8.12822
R26347 D_FlipFlop_7.D.n72 D_FlipFlop_7.D.n71 8.12822
R26348 D_FlipFlop_7.D.n58 D_FlipFlop_7.D.n57 8.12822
R26349 D_FlipFlop_7.D.n44 D_FlipFlop_7.D.n43 8.12822
R26350 D_FlipFlop_7.D.n30 D_FlipFlop_7.D.n29 8.12822
R26351 D_FlipFlop_7.D.n17 D_FlipFlop_7.D.n16 8.12822
R26352 D_FlipFlop_7.D.n112 D_FlipFlop_7.D.n111 8.12822
R26353 D_FlipFlop_7.D.n99 D_FlipFlop_7.D.n98 8.12822
R26354 D_FlipFlop_7.D.n31 D_FlipFlop_7.D.n17 6.18977
R26355 D_FlipFlop_7.D.n113 D_FlipFlop_7.D.n99 6.18977
R26356 D_FlipFlop_7.D.n115 D_FlipFlop_7.D.n114 5.69478
R26357 D_FlipFlop_7.D.n86 D_FlipFlop_7.D.n79 4.5005
R26358 D_FlipFlop_7.D.n72 D_FlipFlop_7.D.n65 4.5005
R26359 D_FlipFlop_7.D.n58 D_FlipFlop_7.D.n51 4.5005
R26360 D_FlipFlop_7.D.n44 D_FlipFlop_7.D.n37 4.5005
R26361 D_FlipFlop_7.D.n30 D_FlipFlop_7.D.n23 4.5005
R26362 D_FlipFlop_7.D.n17 D_FlipFlop_7.D.n10 4.5005
R26363 D_FlipFlop_7.D.n112 D_FlipFlop_7.D.n105 4.5005
R26364 D_FlipFlop_7.D.n99 D_FlipFlop_7.D.n92 4.5005
R26365 D_FlipFlop_7.D.n73 D_FlipFlop_7.D.n59 4.43652
R26366 D_FlipFlop_7.D.n4 D_FlipFlop_7.D.n1 3.8456
R26367 D_FlipFlop_7.D.n31 D_FlipFlop_7.D.n30 3.4105
R26368 D_FlipFlop_7.D.n45 D_FlipFlop_7.D.n44 3.4105
R26369 D_FlipFlop_7.D.n59 D_FlipFlop_7.D.n58 3.4105
R26370 D_FlipFlop_7.D.n73 D_FlipFlop_7.D.n72 3.4105
R26371 D_FlipFlop_7.D.n113 D_FlipFlop_7.D.n112 3.4105
R26372 D_FlipFlop_7.D.n114 D_FlipFlop_7.D.n86 3.4105
R26373 D_FlipFlop_7.D.n45 D_FlipFlop_7.D.n31 2.77977
R26374 D_FlipFlop_7.D.n59 D_FlipFlop_7.D.n45 2.77977
R26375 D_FlipFlop_7.D.n114 D_FlipFlop_7.D.n73 2.77977
R26376 D_FlipFlop_7.D.n114 D_FlipFlop_7.D.n113 2.77977
R26377 D_FlipFlop_7.D.n0 D_FlipFlop_7.D.t33 1.13717
R26378 D_FlipFlop_7.D.n3 D_FlipFlop_7.D.n2 0.855396
R26379 D_FlipFlop_7.D.n75 D_FlipFlop_5.Inverter_0.Vin 0.851043
R26380 D_FlipFlop_7.D.n81 D_FlipFlop_5.3-input-nand_0.B 0.851043
R26381 D_FlipFlop_7.D.n61 D_FlipFlop_4.Inverter_0.Vin 0.851043
R26382 D_FlipFlop_7.D.n67 D_FlipFlop_4.3-input-nand_0.B 0.851043
R26383 D_FlipFlop_7.D.n47 D_FlipFlop_1.Inverter_0.Vin 0.851043
R26384 D_FlipFlop_7.D.n53 D_FlipFlop_1.3-input-nand_0.B 0.851043
R26385 D_FlipFlop_7.D.n33 D_FlipFlop_2.Inverter_0.Vin 0.851043
R26386 D_FlipFlop_7.D.n39 D_FlipFlop_2.3-input-nand_0.B 0.851043
R26387 D_FlipFlop_7.D.n19 D_FlipFlop_3.Inverter_0.Vin 0.851043
R26388 D_FlipFlop_7.D.n25 D_FlipFlop_3.3-input-nand_0.B 0.851043
R26389 D_FlipFlop_7.D.n6 D_FlipFlop_0.Inverter_0.Vin 0.851043
R26390 D_FlipFlop_7.D.n12 D_FlipFlop_0.3-input-nand_0.B 0.851043
R26391 D_FlipFlop_7.D.n101 D_FlipFlop_6.Inverter_0.Vin 0.851043
R26392 D_FlipFlop_7.D.n107 D_FlipFlop_6.3-input-nand_0.B 0.851043
R26393 D_FlipFlop_7.D.n88 D_FlipFlop_7.Inverter_0.Vin 0.851043
R26394 D_FlipFlop_7.D.n94 D_FlipFlop_7.3-input-nand_0.B 0.851043
R26395 D_FlipFlop_7.D.n78 D_FlipFlop_7.D.n77 0.55213
R26396 D_FlipFlop_7.D.n84 D_FlipFlop_7.D.n83 0.55213
R26397 D_FlipFlop_7.D.n64 D_FlipFlop_7.D.n63 0.55213
R26398 D_FlipFlop_7.D.n70 D_FlipFlop_7.D.n69 0.55213
R26399 D_FlipFlop_7.D.n50 D_FlipFlop_7.D.n49 0.55213
R26400 D_FlipFlop_7.D.n56 D_FlipFlop_7.D.n55 0.55213
R26401 D_FlipFlop_7.D.n36 D_FlipFlop_7.D.n35 0.55213
R26402 D_FlipFlop_7.D.n42 D_FlipFlop_7.D.n41 0.55213
R26403 D_FlipFlop_7.D.n22 D_FlipFlop_7.D.n21 0.55213
R26404 D_FlipFlop_7.D.n28 D_FlipFlop_7.D.n27 0.55213
R26405 D_FlipFlop_7.D.n9 D_FlipFlop_7.D.n8 0.55213
R26406 D_FlipFlop_7.D.n15 D_FlipFlop_7.D.n14 0.55213
R26407 D_FlipFlop_7.D.n104 D_FlipFlop_7.D.n103 0.55213
R26408 D_FlipFlop_7.D.n110 D_FlipFlop_7.D.n109 0.55213
R26409 D_FlipFlop_7.D.n91 D_FlipFlop_7.D.n90 0.55213
R26410 D_FlipFlop_7.D.n97 D_FlipFlop_7.D.n96 0.55213
R26411 D_FlipFlop_7.D.n78 D_FlipFlop_5.Inverter_0.Vin 0.486828
R26412 D_FlipFlop_7.D.n84 D_FlipFlop_5.3-input-nand_0.B 0.486828
R26413 D_FlipFlop_7.D.n64 D_FlipFlop_4.Inverter_0.Vin 0.486828
R26414 D_FlipFlop_7.D.n70 D_FlipFlop_4.3-input-nand_0.B 0.486828
R26415 D_FlipFlop_7.D.n50 D_FlipFlop_1.Inverter_0.Vin 0.486828
R26416 D_FlipFlop_7.D.n56 D_FlipFlop_1.3-input-nand_0.B 0.486828
R26417 D_FlipFlop_7.D.n36 D_FlipFlop_2.Inverter_0.Vin 0.486828
R26418 D_FlipFlop_7.D.n42 D_FlipFlop_2.3-input-nand_0.B 0.486828
R26419 D_FlipFlop_7.D.n22 D_FlipFlop_3.Inverter_0.Vin 0.486828
R26420 D_FlipFlop_7.D.n28 D_FlipFlop_3.3-input-nand_0.B 0.486828
R26421 D_FlipFlop_7.D.n9 D_FlipFlop_0.Inverter_0.Vin 0.486828
R26422 D_FlipFlop_7.D.n15 D_FlipFlop_0.3-input-nand_0.B 0.486828
R26423 D_FlipFlop_7.D.n104 D_FlipFlop_6.Inverter_0.Vin 0.486828
R26424 D_FlipFlop_7.D.n110 D_FlipFlop_6.3-input-nand_0.B 0.486828
R26425 D_FlipFlop_7.D.n91 D_FlipFlop_7.Inverter_0.Vin 0.486828
R26426 D_FlipFlop_7.D.n97 D_FlipFlop_7.3-input-nand_0.B 0.486828
R26427 D_FlipFlop_7.D.n75 D_FlipFlop_7.D.n74 0.470609
R26428 D_FlipFlop_7.D.n81 D_FlipFlop_7.D.n80 0.470609
R26429 D_FlipFlop_7.D.n61 D_FlipFlop_7.D.n60 0.470609
R26430 D_FlipFlop_7.D.n67 D_FlipFlop_7.D.n66 0.470609
R26431 D_FlipFlop_7.D.n47 D_FlipFlop_7.D.n46 0.470609
R26432 D_FlipFlop_7.D.n53 D_FlipFlop_7.D.n52 0.470609
R26433 D_FlipFlop_7.D.n33 D_FlipFlop_7.D.n32 0.470609
R26434 D_FlipFlop_7.D.n39 D_FlipFlop_7.D.n38 0.470609
R26435 D_FlipFlop_7.D.n19 D_FlipFlop_7.D.n18 0.470609
R26436 D_FlipFlop_7.D.n25 D_FlipFlop_7.D.n24 0.470609
R26437 D_FlipFlop_7.D.n6 D_FlipFlop_7.D.n5 0.470609
R26438 D_FlipFlop_7.D.n12 D_FlipFlop_7.D.n11 0.470609
R26439 D_FlipFlop_7.D.n101 D_FlipFlop_7.D.n100 0.470609
R26440 D_FlipFlop_7.D.n107 D_FlipFlop_7.D.n106 0.470609
R26441 D_FlipFlop_7.D.n88 D_FlipFlop_7.D.n87 0.470609
R26442 D_FlipFlop_7.D.n94 D_FlipFlop_7.D.n93 0.470609
R26443 D_FlipFlop_7.D.n4 D_FlipFlop_7.D.n3 0.3805
R26444 D_FlipFlop_7.D.n115 D_FlipFlop_7.D.n4 0.280803
R26445 D_FlipFlop_7.D.n74 D_FlipFlop_5.Inverter_0.Vin 0.217464
R26446 D_FlipFlop_7.D.n80 D_FlipFlop_5.3-input-nand_0.B 0.217464
R26447 D_FlipFlop_7.D.n60 D_FlipFlop_4.Inverter_0.Vin 0.217464
R26448 D_FlipFlop_7.D.n66 D_FlipFlop_4.3-input-nand_0.B 0.217464
R26449 D_FlipFlop_7.D.n46 D_FlipFlop_1.Inverter_0.Vin 0.217464
R26450 D_FlipFlop_7.D.n52 D_FlipFlop_1.3-input-nand_0.B 0.217464
R26451 D_FlipFlop_7.D.n32 D_FlipFlop_2.Inverter_0.Vin 0.217464
R26452 D_FlipFlop_7.D.n38 D_FlipFlop_2.3-input-nand_0.B 0.217464
R26453 D_FlipFlop_7.D.n18 D_FlipFlop_3.Inverter_0.Vin 0.217464
R26454 D_FlipFlop_7.D.n24 D_FlipFlop_3.3-input-nand_0.B 0.217464
R26455 D_FlipFlop_7.D.n5 D_FlipFlop_0.Inverter_0.Vin 0.217464
R26456 D_FlipFlop_7.D.n11 D_FlipFlop_0.3-input-nand_0.B 0.217464
R26457 D_FlipFlop_7.D.n100 D_FlipFlop_6.Inverter_0.Vin 0.217464
R26458 D_FlipFlop_7.D.n106 D_FlipFlop_6.3-input-nand_0.B 0.217464
R26459 D_FlipFlop_7.D.n87 D_FlipFlop_7.Inverter_0.Vin 0.217464
R26460 D_FlipFlop_7.D.n93 D_FlipFlop_7.3-input-nand_0.B 0.217464
R26461 D_FlipFlop_7.D.n77 D_FlipFlop_5.Inverter_0.Vin 0.1255
R26462 D_FlipFlop_7.D.n83 D_FlipFlop_5.3-input-nand_0.B 0.1255
R26463 D_FlipFlop_7.D.n63 D_FlipFlop_4.Inverter_0.Vin 0.1255
R26464 D_FlipFlop_7.D.n69 D_FlipFlop_4.3-input-nand_0.B 0.1255
R26465 D_FlipFlop_7.D.n49 D_FlipFlop_1.Inverter_0.Vin 0.1255
R26466 D_FlipFlop_7.D.n55 D_FlipFlop_1.3-input-nand_0.B 0.1255
R26467 D_FlipFlop_7.D.n35 D_FlipFlop_2.Inverter_0.Vin 0.1255
R26468 D_FlipFlop_7.D.n41 D_FlipFlop_2.3-input-nand_0.B 0.1255
R26469 D_FlipFlop_7.D.n21 D_FlipFlop_3.Inverter_0.Vin 0.1255
R26470 D_FlipFlop_7.D.n27 D_FlipFlop_3.3-input-nand_0.B 0.1255
R26471 D_FlipFlop_7.D.n8 D_FlipFlop_0.Inverter_0.Vin 0.1255
R26472 D_FlipFlop_7.D.n14 D_FlipFlop_0.3-input-nand_0.B 0.1255
R26473 D_FlipFlop_7.D.n103 D_FlipFlop_6.Inverter_0.Vin 0.1255
R26474 D_FlipFlop_7.D.n109 D_FlipFlop_6.3-input-nand_0.B 0.1255
R26475 D_FlipFlop_7.D.n90 D_FlipFlop_7.Inverter_0.Vin 0.1255
R26476 D_FlipFlop_7.D.n96 D_FlipFlop_7.3-input-nand_0.B 0.1255
R26477 D_FlipFlop_7.D.n116 D_FlipFlop_7.D.n115 0.105716
R26478 D_FlipFlop_7.D.n3 D_FlipFlop_7.D.t0 0.0856875
R26479 D_FlipFlop_7.D.n79 D_FlipFlop_7.D.n75 0.063
R26480 D_FlipFlop_7.D.n79 D_FlipFlop_7.D.n78 0.063
R26481 D_FlipFlop_7.D.n85 D_FlipFlop_7.D.n81 0.063
R26482 D_FlipFlop_7.D.n85 D_FlipFlop_7.D.n84 0.063
R26483 D_FlipFlop_7.D.n65 D_FlipFlop_7.D.n61 0.063
R26484 D_FlipFlop_7.D.n65 D_FlipFlop_7.D.n64 0.063
R26485 D_FlipFlop_7.D.n71 D_FlipFlop_7.D.n67 0.063
R26486 D_FlipFlop_7.D.n71 D_FlipFlop_7.D.n70 0.063
R26487 D_FlipFlop_7.D.n51 D_FlipFlop_7.D.n47 0.063
R26488 D_FlipFlop_7.D.n51 D_FlipFlop_7.D.n50 0.063
R26489 D_FlipFlop_7.D.n57 D_FlipFlop_7.D.n53 0.063
R26490 D_FlipFlop_7.D.n57 D_FlipFlop_7.D.n56 0.063
R26491 D_FlipFlop_7.D.n37 D_FlipFlop_7.D.n33 0.063
R26492 D_FlipFlop_7.D.n37 D_FlipFlop_7.D.n36 0.063
R26493 D_FlipFlop_7.D.n43 D_FlipFlop_7.D.n39 0.063
R26494 D_FlipFlop_7.D.n43 D_FlipFlop_7.D.n42 0.063
R26495 D_FlipFlop_7.D.n23 D_FlipFlop_7.D.n19 0.063
R26496 D_FlipFlop_7.D.n23 D_FlipFlop_7.D.n22 0.063
R26497 D_FlipFlop_7.D.n29 D_FlipFlop_7.D.n25 0.063
R26498 D_FlipFlop_7.D.n29 D_FlipFlop_7.D.n28 0.063
R26499 D_FlipFlop_7.D.n10 D_FlipFlop_7.D.n6 0.063
R26500 D_FlipFlop_7.D.n10 D_FlipFlop_7.D.n9 0.063
R26501 D_FlipFlop_7.D.n16 D_FlipFlop_7.D.n12 0.063
R26502 D_FlipFlop_7.D.n16 D_FlipFlop_7.D.n15 0.063
R26503 D_FlipFlop_7.D.n105 D_FlipFlop_7.D.n101 0.063
R26504 D_FlipFlop_7.D.n105 D_FlipFlop_7.D.n104 0.063
R26505 D_FlipFlop_7.D.n111 D_FlipFlop_7.D.n107 0.063
R26506 D_FlipFlop_7.D.n111 D_FlipFlop_7.D.n110 0.063
R26507 D_FlipFlop_7.D.n92 D_FlipFlop_7.D.n88 0.063
R26508 D_FlipFlop_7.D.n92 D_FlipFlop_7.D.n91 0.063
R26509 D_FlipFlop_7.D.n98 D_FlipFlop_7.D.n94 0.063
R26510 D_FlipFlop_7.D.n98 D_FlipFlop_7.D.n97 0.063
R26511 Comparator_0.Vout D_FlipFlop_7.D.n116 0.0620344
R26512 D_FlipFlop_7.D.n116 D_FlipFlop_7.D.n0 0.0413995
R26513 D_FlipFlop_7.D.n77 D_FlipFlop_7.D.n76 0.0216397
R26514 D_FlipFlop_7.D.n76 D_FlipFlop_5.Inverter_0.Vin 0.0216397
R26515 D_FlipFlop_7.D.n83 D_FlipFlop_7.D.n82 0.0216397
R26516 D_FlipFlop_7.D.n82 D_FlipFlop_5.3-input-nand_0.B 0.0216397
R26517 D_FlipFlop_7.D.n63 D_FlipFlop_7.D.n62 0.0216397
R26518 D_FlipFlop_7.D.n62 D_FlipFlop_4.Inverter_0.Vin 0.0216397
R26519 D_FlipFlop_7.D.n69 D_FlipFlop_7.D.n68 0.0216397
R26520 D_FlipFlop_7.D.n68 D_FlipFlop_4.3-input-nand_0.B 0.0216397
R26521 D_FlipFlop_7.D.n49 D_FlipFlop_7.D.n48 0.0216397
R26522 D_FlipFlop_7.D.n48 D_FlipFlop_1.Inverter_0.Vin 0.0216397
R26523 D_FlipFlop_7.D.n55 D_FlipFlop_7.D.n54 0.0216397
R26524 D_FlipFlop_7.D.n54 D_FlipFlop_1.3-input-nand_0.B 0.0216397
R26525 D_FlipFlop_7.D.n35 D_FlipFlop_7.D.n34 0.0216397
R26526 D_FlipFlop_7.D.n34 D_FlipFlop_2.Inverter_0.Vin 0.0216397
R26527 D_FlipFlop_7.D.n41 D_FlipFlop_7.D.n40 0.0216397
R26528 D_FlipFlop_7.D.n40 D_FlipFlop_2.3-input-nand_0.B 0.0216397
R26529 D_FlipFlop_7.D.n21 D_FlipFlop_7.D.n20 0.0216397
R26530 D_FlipFlop_7.D.n20 D_FlipFlop_3.Inverter_0.Vin 0.0216397
R26531 D_FlipFlop_7.D.n27 D_FlipFlop_7.D.n26 0.0216397
R26532 D_FlipFlop_7.D.n26 D_FlipFlop_3.3-input-nand_0.B 0.0216397
R26533 D_FlipFlop_7.D.n8 D_FlipFlop_7.D.n7 0.0216397
R26534 D_FlipFlop_7.D.n7 D_FlipFlop_0.Inverter_0.Vin 0.0216397
R26535 D_FlipFlop_7.D.n14 D_FlipFlop_7.D.n13 0.0216397
R26536 D_FlipFlop_7.D.n13 D_FlipFlop_0.3-input-nand_0.B 0.0216397
R26537 D_FlipFlop_7.D.n103 D_FlipFlop_7.D.n102 0.0216397
R26538 D_FlipFlop_7.D.n102 D_FlipFlop_6.Inverter_0.Vin 0.0216397
R26539 D_FlipFlop_7.D.n109 D_FlipFlop_7.D.n108 0.0216397
R26540 D_FlipFlop_7.D.n108 D_FlipFlop_6.3-input-nand_0.B 0.0216397
R26541 D_FlipFlop_7.D.n90 D_FlipFlop_7.D.n89 0.0216397
R26542 D_FlipFlop_7.D.n89 D_FlipFlop_7.Inverter_0.Vin 0.0216397
R26543 D_FlipFlop_7.D.n96 D_FlipFlop_7.D.n95 0.0216397
R26544 D_FlipFlop_7.D.n95 D_FlipFlop_7.3-input-nand_0.B 0.0216397
R26545 D_FlipFlop_7.D.n0 Comparator_0.Vout 0.0131087
R26546 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 169.46
R26547 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 168.089
R26548 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 167.809
R26549 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 150.273
R26550 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 73.6406
R26551 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 60.3809
R26552 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 12.0358
R26553 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 11.4489
R26554 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 1.08746
R26555 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.851043
R26556 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.848156
R26557 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 0.788543
R26558 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 0.682565
R26559 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.65675
R26560 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 0.55213
R26561 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.486828
R26562 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 0.470609
R26563 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 0.262643
R26564 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.217464
R26565 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.1255
R26566 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.1255
R26567 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 0.063
R26568 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 0.063
R26569 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 0.063
R26570 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 0.063
R26571 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 0.063
R26572 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 0.0216397
R26573 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.0216397
R26574 Nand_Gate_0.A.n55 Nand_Gate_0.A.t3 169.46
R26575 Nand_Gate_0.A.n57 Nand_Gate_0.A.t2 167.809
R26576 Nand_Gate_0.A.n55 Nand_Gate_0.A.t0 167.809
R26577 Nand_Gate_0.A Nand_Gate_0.A.t13 158.585
R26578 Nand_Gate_0.A Nand_Gate_0.A.t16 158.581
R26579 Nand_Gate_0.A.n42 Nand_Gate_0.A.t11 150.293
R26580 Nand_Gate_0.A.t16 Nand_Gate_0.A.n38 150.293
R26581 Nand_Gate_0.A.t13 Nand_Gate_0.A.n2 150.293
R26582 Nand_Gate_0.A.n29 Nand_Gate_0.A.t10 150.273
R26583 Nand_Gate_0.A.n23 Nand_Gate_0.A.t17 150.273
R26584 Nand_Gate_0.A.n14 Nand_Gate_0.A.t12 150.273
R26585 Nand_Gate_0.A.n8 Nand_Gate_0.A.t8 150.273
R26586 Nand_Gate_0.A.n27 Nand_Gate_0.A.t6 73.6406
R26587 Nand_Gate_0.A.n21 Nand_Gate_0.A.t15 73.6406
R26588 Nand_Gate_0.A.n12 Nand_Gate_0.A.t7 73.6406
R26589 Nand_Gate_0.A.n6 Nand_Gate_0.A.t14 73.6406
R26590 Nand_Gate_0.A.n44 Nand_Gate_0.A.t4 73.6304
R26591 Nand_Gate_0.A.n36 Nand_Gate_0.A.t5 73.6304
R26592 Nand_Gate_0.A.n0 Nand_Gate_0.A.t9 73.6304
R26593 Nand_Gate_0.A.n48 Nand_Gate_0.A.n41 65.2862
R26594 Nand_Gate_0.A.n4 Nand_Gate_0.A.t1 60.3809
R26595 Nand_Gate_0.A.n33 Nand_Gate_0.A.n26 15.5222
R26596 Nand_Gate_0.A.n56 Nand_Gate_0.A.n55 11.4489
R26597 Nand_Gate_0.A.n48 Nand_Gate_0.A.n47 9.57083
R26598 Nand_Gate_0.A.n34 Nand_Gate_0.A.n33 8.26552
R26599 Nand_Gate_0.A.n58 Nand_Gate_0.A.n57 8.21389
R26600 Nand_Gate_0.A.n18 Nand_Gate_0.A.n11 8.1418
R26601 Nand_Gate_0.A.n49 Nand_Gate_0.A.n48 6.58222
R26602 Nand_Gate_0.A.n20 Nand_Gate_0.A.n19 6.47604
R26603 Nand_Gate_0.A.n19 Nand_Gate_0.A 5.35402
R26604 Nand_Gate_0.A.n52 Nand_Gate_0.A 4.55128
R26605 Nand_Gate_0.A.n33 Nand_Gate_0.A.n32 4.5005
R26606 Nand_Gate_0.A.n18 Nand_Gate_0.A.n17 4.5005
R26607 Nand_Gate_0.A.n38 Nand_Gate_0.A.n37 1.19615
R26608 Nand_Gate_0.A.n2 Nand_Gate_0.A.n1 1.19615
R26609 Nand_Gate_0.A.n5 Nand_Gate_0.A 1.08746
R26610 Nand_Gate_0.A.n20 Nand_Gate_0.A 0.973326
R26611 Nand_Gate_0.A.n13 Nand_Gate_0.A 0.851043
R26612 Nand_Gate_0.A.n7 Nand_Gate_0.A 0.851043
R26613 Nand_Gate_0.A.n4 Nand_Gate_0.A 0.848156
R26614 Nand_Gate_0.A.n28 Nand_Gate_0.A.n27 0.796696
R26615 Nand_Gate_0.A.n22 Nand_Gate_0.A.n21 0.796696
R26616 Nand_Gate_0.A.n54 Nand_Gate_0.A.n53 0.788543
R26617 Nand_Gate_0.A.n43 Nand_Gate_0.A 0.769522
R26618 Nand_Gate_0.A.n51 Nand_Gate_0.A.n50 0.755935
R26619 Nand_Gate_0.A.n34 Nand_Gate_0.A 0.716182
R26620 Nand_Gate_0.A.n5 Nand_Gate_0.A.n4 0.682565
R26621 Nand_Gate_0.A.n53 Nand_Gate_0.A 0.65675
R26622 Nand_Gate_0.A.n35 Nand_Gate_0.A.n34 0.556667
R26623 Nand_Gate_0.A.n43 Nand_Gate_0.A.n42 0.55213
R26624 Nand_Gate_0.A.n16 Nand_Gate_0.A.n15 0.55213
R26625 Nand_Gate_0.A.n10 Nand_Gate_0.A.n9 0.55213
R26626 Nand_Gate_0.A.n28 Nand_Gate_0.A 0.524957
R26627 Nand_Gate_0.A.n22 Nand_Gate_0.A 0.524957
R26628 Nand_Gate_0.A.n16 Nand_Gate_0.A 0.486828
R26629 Nand_Gate_0.A.n10 Nand_Gate_0.A 0.486828
R26630 Nand_Gate_0.A.n50 Nand_Gate_0.A 0.48023
R26631 Nand_Gate_0.A.n46 Nand_Gate_0.A.n45 0.470609
R26632 Nand_Gate_0.A.n13 Nand_Gate_0.A.n12 0.470609
R26633 Nand_Gate_0.A.n7 Nand_Gate_0.A.n6 0.470609
R26634 Nand_Gate_0.A.n42 Nand_Gate_0.A 0.447191
R26635 Nand_Gate_0.A.n38 Nand_Gate_0.A 0.447191
R26636 Nand_Gate_0.A.n2 Nand_Gate_0.A 0.447191
R26637 Nand_Gate_0.A.n46 Nand_Gate_0.A 0.428234
R26638 Nand_Gate_0.A.n58 Nand_Gate_0.A.n3 0.425067
R26639 Nand_Gate_0.A Nand_Gate_0.A.n58 0.39003
R26640 Nand_Gate_0.A.n57 Nand_Gate_0.A.n56 0.280391
R26641 Nand_Gate_0.A.n31 Nand_Gate_0.A 0.252453
R26642 Nand_Gate_0.A.n25 Nand_Gate_0.A 0.252453
R26643 Nand_Gate_0.A.n35 Nand_Gate_0.A 0.231583
R26644 Nand_Gate_0.A.n31 Nand_Gate_0.A.n30 0.226043
R26645 Nand_Gate_0.A.n25 Nand_Gate_0.A.n24 0.226043
R26646 Nand_Gate_0.A.n27 Nand_Gate_0.A 0.217464
R26647 Nand_Gate_0.A.n21 Nand_Gate_0.A 0.217464
R26648 Nand_Gate_0.A.n12 Nand_Gate_0.A 0.217464
R26649 Nand_Gate_0.A.n6 Nand_Gate_0.A 0.217464
R26650 Nand_Gate_0.A.n56 Nand_Gate_0.A 0.200143
R26651 Nand_Gate_0.A.n40 Nand_Gate_0.A.n39 0.168133
R26652 Nand_Gate_0.A.n40 Nand_Gate_0.A 0.135934
R26653 Nand_Gate_0.A.n45 Nand_Gate_0.A 0.1255
R26654 Nand_Gate_0.A.n30 Nand_Gate_0.A 0.1255
R26655 Nand_Gate_0.A.n24 Nand_Gate_0.A 0.1255
R26656 Nand_Gate_0.A.n37 Nand_Gate_0.A 0.1255
R26657 Nand_Gate_0.A.n15 Nand_Gate_0.A 0.1255
R26658 Nand_Gate_0.A.n9 Nand_Gate_0.A 0.1255
R26659 Nand_Gate_0.A.n54 Nand_Gate_0.A 0.1255
R26660 Nand_Gate_0.A.n1 Nand_Gate_0.A 0.1255
R26661 Nand_Gate_0.A.n47 Nand_Gate_0.A.n43 0.063
R26662 Nand_Gate_0.A.n47 Nand_Gate_0.A.n46 0.063
R26663 Nand_Gate_0.A.n32 Nand_Gate_0.A.n28 0.063
R26664 Nand_Gate_0.A.n32 Nand_Gate_0.A.n31 0.063
R26665 Nand_Gate_0.A.n26 Nand_Gate_0.A.n22 0.063
R26666 Nand_Gate_0.A.n26 Nand_Gate_0.A.n25 0.063
R26667 Nand_Gate_0.A.n17 Nand_Gate_0.A.n13 0.063
R26668 Nand_Gate_0.A.n17 Nand_Gate_0.A.n16 0.063
R26669 Nand_Gate_0.A.n11 Nand_Gate_0.A.n7 0.063
R26670 Nand_Gate_0.A.n11 Nand_Gate_0.A.n10 0.063
R26671 Nand_Gate_0.A.n19 Nand_Gate_0.A.n18 0.063
R26672 Nand_Gate_0.A.n49 Nand_Gate_0.A.n20 0.063
R26673 Nand_Gate_0.A.n50 Nand_Gate_0.A.n49 0.063
R26674 Nand_Gate_0.A.n52 Nand_Gate_0.A.n5 0.063
R26675 Nand_Gate_0.A.n53 Nand_Gate_0.A.n52 0.063
R26676 Nand_Gate_0.A Nand_Gate_0.A.n54 0.063
R26677 Nand_Gate_0.A.n41 Nand_Gate_0.A.n35 0.024
R26678 Nand_Gate_0.A.n41 Nand_Gate_0.A.n40 0.024
R26679 Nand_Gate_0.A.n30 Nand_Gate_0.A.n29 0.0216397
R26680 Nand_Gate_0.A.n29 Nand_Gate_0.A 0.0216397
R26681 Nand_Gate_0.A.n24 Nand_Gate_0.A.n23 0.0216397
R26682 Nand_Gate_0.A.n23 Nand_Gate_0.A 0.0216397
R26683 Nand_Gate_0.A.n15 Nand_Gate_0.A.n14 0.0216397
R26684 Nand_Gate_0.A.n14 Nand_Gate_0.A 0.0216397
R26685 Nand_Gate_0.A.n9 Nand_Gate_0.A.n8 0.0216397
R26686 Nand_Gate_0.A.n8 Nand_Gate_0.A 0.0216397
R26687 Nand_Gate_0.A.n51 Nand_Gate_0.A 0.0168043
R26688 Nand_Gate_0.A Nand_Gate_0.A.n51 0.0122188
R26689 Nand_Gate_0.A.n45 Nand_Gate_0.A.n44 0.0107679
R26690 Nand_Gate_0.A.n44 Nand_Gate_0.A 0.0107679
R26691 Nand_Gate_0.A.n37 Nand_Gate_0.A.n36 0.0107679
R26692 Nand_Gate_0.A.n36 Nand_Gate_0.A 0.0107679
R26693 Nand_Gate_0.A.n1 Nand_Gate_0.A.n0 0.0107679
R26694 Nand_Gate_0.A.n0 Nand_Gate_0.A 0.0107679
R26695 Nand_Gate_0.A.n39 Nand_Gate_0.A 0.00441667
R26696 Nand_Gate_0.A.n3 Nand_Gate_0.A 0.00441667
R26697 Nand_Gate_0.A.n39 Nand_Gate_0.A 0.00406061
R26698 Nand_Gate_0.A.n3 Nand_Gate_0.A 0.00406061
R26699 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 316.762
R26700 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 168.108
R26701 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 150.293
R26702 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 150.273
R26703 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 73.6406
R26704 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 73.6304
R26705 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 60.3943
R26706 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 12.0358
R26707 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 1.19615
R26708 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.981478
R26709 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 0.788543
R26710 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.769522
R26711 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 0.682565
R26712 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.580578
R26713 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 0.55213
R26714 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 0.484875
R26715 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 0.470609
R26716 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.447191
R26717 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.428234
R26718 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.217464
R26719 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R26720 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R26721 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R26722 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 0.063
R26723 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 0.063
R26724 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.063
R26725 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 0.063
R26726 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 0.063
R26727 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 0.0216397
R26728 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.0216397
R26729 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 0.0107679
R26730 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.0107679
R26731 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 179.256
R26732 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 168.089
R26733 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 150.293
R26734 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 73.6304
R26735 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 60.3943
R26736 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 12.0358
R26737 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.981478
R26738 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 0.788543
R26739 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.769522
R26740 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.720633
R26741 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 0.682565
R26742 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.580578
R26743 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 0.55213
R26744 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 0.470609
R26745 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.447191
R26746 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.428234
R26747 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1255
R26748 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1255
R26749 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 0.063
R26750 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 0.063
R26751 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 0.063
R26752 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 0.063
R26753 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 0.063
R26754 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 0.0435206
R26755 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 0.0107679
R26756 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.0107679
R26757 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 169.46
R26758 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 168.089
R26759 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 167.809
R26760 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 150.293
R26761 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 73.6304
R26762 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 60.3943
R26763 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 12.0358
R26764 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 11.4489
R26765 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.981478
R26766 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 0.788543
R26767 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.769522
R26768 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 0.720633
R26769 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 0.682565
R26770 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.580578
R26771 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 0.55213
R26772 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 0.470609
R26773 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.447191
R26774 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.428234
R26775 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.1255
R26776 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.1255
R26777 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 0.063
R26778 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 0.063
R26779 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.063
R26780 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 0.063
R26781 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 0.063
R26782 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 0.0435206
R26783 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 0.0107679
R26784 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.0107679
R26785 Nand_Gate_2.A.n55 Nand_Gate_2.A.t3 169.46
R26786 Nand_Gate_2.A.n57 Nand_Gate_2.A.t2 167.809
R26787 Nand_Gate_2.A.n55 Nand_Gate_2.A.t0 167.809
R26788 Nand_Gate_2.A Nand_Gate_2.A.t11 158.585
R26789 Nand_Gate_2.A Nand_Gate_2.A.t7 158.581
R26790 Nand_Gate_2.A.n42 Nand_Gate_2.A.t14 150.293
R26791 Nand_Gate_2.A.t7 Nand_Gate_2.A.n38 150.293
R26792 Nand_Gate_2.A.t11 Nand_Gate_2.A.n2 150.293
R26793 Nand_Gate_2.A.n29 Nand_Gate_2.A.t5 150.273
R26794 Nand_Gate_2.A.n23 Nand_Gate_2.A.t9 150.273
R26795 Nand_Gate_2.A.n14 Nand_Gate_2.A.t15 150.273
R26796 Nand_Gate_2.A.n8 Nand_Gate_2.A.t17 150.273
R26797 Nand_Gate_2.A.n27 Nand_Gate_2.A.t10 73.6406
R26798 Nand_Gate_2.A.n21 Nand_Gate_2.A.t6 73.6406
R26799 Nand_Gate_2.A.n12 Nand_Gate_2.A.t4 73.6406
R26800 Nand_Gate_2.A.n6 Nand_Gate_2.A.t16 73.6406
R26801 Nand_Gate_2.A.n44 Nand_Gate_2.A.t12 73.6304
R26802 Nand_Gate_2.A.n36 Nand_Gate_2.A.t13 73.6304
R26803 Nand_Gate_2.A.n0 Nand_Gate_2.A.t8 73.6304
R26804 Nand_Gate_2.A.n4 Nand_Gate_2.A.t1 60.3809
R26805 Nand_Gate_2.A.n48 Nand_Gate_2.A.n41 45.1913
R26806 Nand_Gate_2.A.n33 Nand_Gate_2.A.n26 15.5222
R26807 Nand_Gate_2.A.n56 Nand_Gate_2.A.n55 11.4489
R26808 Nand_Gate_2.A.n48 Nand_Gate_2.A.n47 9.57083
R26809 Nand_Gate_2.A.n34 Nand_Gate_2.A.n33 8.26552
R26810 Nand_Gate_2.A.n58 Nand_Gate_2.A.n57 8.21389
R26811 Nand_Gate_2.A.n18 Nand_Gate_2.A.n11 8.1418
R26812 Nand_Gate_2.A.n49 Nand_Gate_2.A.n48 6.58222
R26813 Nand_Gate_2.A.n20 Nand_Gate_2.A.n19 6.47604
R26814 Nand_Gate_2.A.n19 Nand_Gate_2.A 5.35402
R26815 Nand_Gate_2.A.n52 Nand_Gate_2.A 4.55128
R26816 Nand_Gate_2.A.n33 Nand_Gate_2.A.n32 4.5005
R26817 Nand_Gate_2.A.n18 Nand_Gate_2.A.n17 4.5005
R26818 Nand_Gate_2.A.n38 Nand_Gate_2.A.n37 1.19615
R26819 Nand_Gate_2.A.n2 Nand_Gate_2.A.n1 1.19615
R26820 Nand_Gate_2.A.n5 Nand_Gate_2.A 1.08746
R26821 Nand_Gate_2.A.n20 Nand_Gate_2.A 0.973326
R26822 Nand_Gate_2.A.n13 Nand_Gate_2.A 0.851043
R26823 Nand_Gate_2.A.n7 Nand_Gate_2.A 0.851043
R26824 Nand_Gate_2.A.n4 Nand_Gate_2.A 0.848156
R26825 Nand_Gate_2.A.n28 Nand_Gate_2.A.n27 0.796696
R26826 Nand_Gate_2.A.n22 Nand_Gate_2.A.n21 0.796696
R26827 Nand_Gate_2.A.n54 Nand_Gate_2.A.n53 0.788543
R26828 Nand_Gate_2.A.n43 Nand_Gate_2.A 0.769522
R26829 Nand_Gate_2.A.n51 Nand_Gate_2.A.n50 0.755935
R26830 Nand_Gate_2.A.n34 Nand_Gate_2.A 0.716182
R26831 Nand_Gate_2.A.n5 Nand_Gate_2.A.n4 0.682565
R26832 Nand_Gate_2.A.n53 Nand_Gate_2.A 0.65675
R26833 Nand_Gate_2.A.n43 Nand_Gate_2.A.n42 0.55213
R26834 Nand_Gate_2.A.n16 Nand_Gate_2.A.n15 0.55213
R26835 Nand_Gate_2.A.n10 Nand_Gate_2.A.n9 0.55213
R26836 Nand_Gate_2.A.n35 Nand_Gate_2.A.n34 0.549617
R26837 Nand_Gate_2.A.n28 Nand_Gate_2.A 0.524957
R26838 Nand_Gate_2.A.n22 Nand_Gate_2.A 0.524957
R26839 Nand_Gate_2.A.n16 Nand_Gate_2.A 0.486828
R26840 Nand_Gate_2.A.n10 Nand_Gate_2.A 0.486828
R26841 Nand_Gate_2.A.n50 Nand_Gate_2.A 0.48023
R26842 Nand_Gate_2.A.n46 Nand_Gate_2.A.n45 0.470609
R26843 Nand_Gate_2.A.n13 Nand_Gate_2.A.n12 0.470609
R26844 Nand_Gate_2.A.n7 Nand_Gate_2.A.n6 0.470609
R26845 Nand_Gate_2.A.n42 Nand_Gate_2.A 0.447191
R26846 Nand_Gate_2.A.n38 Nand_Gate_2.A 0.447191
R26847 Nand_Gate_2.A.n2 Nand_Gate_2.A 0.447191
R26848 Nand_Gate_2.A.n46 Nand_Gate_2.A 0.428234
R26849 Nand_Gate_2.A.n58 Nand_Gate_2.A.n3 0.425067
R26850 Nand_Gate_2.A Nand_Gate_2.A.n58 0.39003
R26851 Nand_Gate_2.A.n57 Nand_Gate_2.A.n56 0.280391
R26852 Nand_Gate_2.A.n31 Nand_Gate_2.A 0.252453
R26853 Nand_Gate_2.A.n25 Nand_Gate_2.A 0.252453
R26854 Nand_Gate_2.A.n35 Nand_Gate_2.A 0.238633
R26855 Nand_Gate_2.A.n31 Nand_Gate_2.A.n30 0.226043
R26856 Nand_Gate_2.A.n25 Nand_Gate_2.A.n24 0.226043
R26857 Nand_Gate_2.A.n27 Nand_Gate_2.A 0.217464
R26858 Nand_Gate_2.A.n21 Nand_Gate_2.A 0.217464
R26859 Nand_Gate_2.A.n12 Nand_Gate_2.A 0.217464
R26860 Nand_Gate_2.A.n6 Nand_Gate_2.A 0.217464
R26861 Nand_Gate_2.A.n56 Nand_Gate_2.A 0.200143
R26862 Nand_Gate_2.A.n40 Nand_Gate_2.A.n39 0.175183
R26863 Nand_Gate_2.A.n40 Nand_Gate_2.A 0.1415
R26864 Nand_Gate_2.A.n45 Nand_Gate_2.A 0.1255
R26865 Nand_Gate_2.A.n30 Nand_Gate_2.A 0.1255
R26866 Nand_Gate_2.A.n24 Nand_Gate_2.A 0.1255
R26867 Nand_Gate_2.A.n37 Nand_Gate_2.A 0.1255
R26868 Nand_Gate_2.A.n15 Nand_Gate_2.A 0.1255
R26869 Nand_Gate_2.A.n9 Nand_Gate_2.A 0.1255
R26870 Nand_Gate_2.A.n54 Nand_Gate_2.A 0.1255
R26871 Nand_Gate_2.A.n1 Nand_Gate_2.A 0.1255
R26872 Nand_Gate_2.A.n47 Nand_Gate_2.A.n43 0.063
R26873 Nand_Gate_2.A.n47 Nand_Gate_2.A.n46 0.063
R26874 Nand_Gate_2.A.n32 Nand_Gate_2.A.n28 0.063
R26875 Nand_Gate_2.A.n32 Nand_Gate_2.A.n31 0.063
R26876 Nand_Gate_2.A.n26 Nand_Gate_2.A.n22 0.063
R26877 Nand_Gate_2.A.n26 Nand_Gate_2.A.n25 0.063
R26878 Nand_Gate_2.A.n17 Nand_Gate_2.A.n13 0.063
R26879 Nand_Gate_2.A.n17 Nand_Gate_2.A.n16 0.063
R26880 Nand_Gate_2.A.n11 Nand_Gate_2.A.n7 0.063
R26881 Nand_Gate_2.A.n11 Nand_Gate_2.A.n10 0.063
R26882 Nand_Gate_2.A.n19 Nand_Gate_2.A.n18 0.063
R26883 Nand_Gate_2.A.n49 Nand_Gate_2.A.n20 0.063
R26884 Nand_Gate_2.A.n50 Nand_Gate_2.A.n49 0.063
R26885 Nand_Gate_2.A.n52 Nand_Gate_2.A.n5 0.063
R26886 Nand_Gate_2.A.n53 Nand_Gate_2.A.n52 0.063
R26887 Nand_Gate_2.A Nand_Gate_2.A.n54 0.063
R26888 Nand_Gate_2.A.n41 Nand_Gate_2.A.n35 0.024
R26889 Nand_Gate_2.A.n41 Nand_Gate_2.A.n40 0.024
R26890 Nand_Gate_2.A.n30 Nand_Gate_2.A.n29 0.0216397
R26891 Nand_Gate_2.A.n29 Nand_Gate_2.A 0.0216397
R26892 Nand_Gate_2.A.n24 Nand_Gate_2.A.n23 0.0216397
R26893 Nand_Gate_2.A.n23 Nand_Gate_2.A 0.0216397
R26894 Nand_Gate_2.A.n15 Nand_Gate_2.A.n14 0.0216397
R26895 Nand_Gate_2.A.n14 Nand_Gate_2.A 0.0216397
R26896 Nand_Gate_2.A.n9 Nand_Gate_2.A.n8 0.0216397
R26897 Nand_Gate_2.A.n8 Nand_Gate_2.A 0.0216397
R26898 Nand_Gate_2.A.n51 Nand_Gate_2.A 0.0168043
R26899 Nand_Gate_2.A Nand_Gate_2.A.n51 0.0122188
R26900 Nand_Gate_2.A.n45 Nand_Gate_2.A.n44 0.0107679
R26901 Nand_Gate_2.A.n44 Nand_Gate_2.A 0.0107679
R26902 Nand_Gate_2.A.n37 Nand_Gate_2.A.n36 0.0107679
R26903 Nand_Gate_2.A.n36 Nand_Gate_2.A 0.0107679
R26904 Nand_Gate_2.A.n1 Nand_Gate_2.A.n0 0.0107679
R26905 Nand_Gate_2.A.n0 Nand_Gate_2.A 0.0107679
R26906 Nand_Gate_2.A.n39 Nand_Gate_2.A 0.00441667
R26907 Nand_Gate_2.A.n3 Nand_Gate_2.A 0.00441667
R26908 Nand_Gate_2.A.n39 Nand_Gate_2.A 0.00406061
R26909 Nand_Gate_2.A.n3 Nand_Gate_2.A 0.00406061
R26910 And_Gate_1.Vout.n13 And_Gate_1.Vout.t0 168.32
R26911 And_Gate_1.Vout.n4 And_Gate_1.Vout.t3 158.207
R26912 D_FlipFlop_7.CLK And_Gate_1.Vout.t5 158.202
R26913 And_Gate_1.Vout.n6 And_Gate_1.Vout.t4 150.293
R26914 And_Gate_1.Vout.t5 And_Gate_1.Vout.n9 150.293
R26915 And_Gate_1.Vout.t3 And_Gate_1.Vout.n3 150.273
R26916 And_Gate_1.Vout.n13 And_Gate_1.Vout.n12 81.2012
R26917 And_Gate_1.Vout.n1 And_Gate_1.Vout.t6 73.6406
R26918 And_Gate_1.Vout.n8 And_Gate_1.Vout.t2 73.6304
R26919 And_Gate_1.Vout.n7 And_Gate_1.Vout.t7 73.6304
R26920 And_Gate_1.Inverter_0.Vout And_Gate_1.Vout.t1 60.3943
R26921 And_Gate_1.Vout.n8 And_Gate_1.Vout.n7 16.332
R26922 And_Gate_1.Vout.n14 And_Gate_1.Vout.n0 1.62007
R26923 And_Gate_1.Inverter_0.Vout And_Gate_1.Vout.n14 1.25441
R26924 And_Gate_1.Vout.n2 And_Gate_1.Vout.n1 1.19615
R26925 And_Gate_1.Vout.n7 And_Gate_1.Vout.n6 1.1717
R26926 And_Gate_1.Vout.n9 And_Gate_1.Vout.n8 1.1717
R26927 And_Gate_1.Vout.n9 D_FlipFlop_7.3-input-nand_1.C 0.447191
R26928 And_Gate_1.Vout.n6 D_FlipFlop_7.Inverter_1.Vin 0.436162
R26929 And_Gate_1.Vout.n4 D_FlipFlop_7.CLK 0.321667
R26930 And_Gate_1.Vout.n5 D_FlipFlop_7.CLK 0.250383
R26931 And_Gate_1.Vout.n1 D_FlipFlop_7.3-input-nand_0.C 0.217464
R26932 And_Gate_1.Vout.n11 And_Gate_1.Vout.n10 0.186933
R26933 And_Gate_1.Vout.n11 D_FlipFlop_7.CLK 0.150776
R26934 And_Gate_1.Vout.n8 D_FlipFlop_7.3-input-nand_1.C 0.149957
R26935 And_Gate_1.Vout.n2 D_FlipFlop_7.3-input-nand_0.C 0.1255
R26936 And_Gate_1.Vout.n0 And_Gate_1.Inverter_0.Vout 0.1255
R26937 And_Gate_1.Vout.n7 D_FlipFlop_7.Inverter_1.Vin 0.117348
R26938 And_Gate_1.Vout.n5 And_Gate_1.Vout.n4 0.1039
R26939 And_Gate_1.Vout.n0 And_Gate_1.Inverter_0.Vout 0.063
R26940 And_Gate_1.Vout.n14 And_Gate_1.Vout.n13 0.063
R26941 And_Gate_1.Vout.n7 D_FlipFlop_7.Inverter_1.Vin 0.0454219
R26942 And_Gate_1.Vout.n8 D_FlipFlop_7.3-input-nand_1.C 0.0454219
R26943 And_Gate_1.Vout.n12 And_Gate_1.Vout.n5 0.024
R26944 And_Gate_1.Vout.n12 And_Gate_1.Vout.n11 0.024
R26945 And_Gate_1.Vout.n3 And_Gate_1.Vout.n2 0.0216397
R26946 And_Gate_1.Vout.n3 D_FlipFlop_7.3-input-nand_0.C 0.0216397
R26947 And_Gate_1.Vout.n10 D_FlipFlop_7.CLK 0.00441667
R26948 And_Gate_1.Vout.n10 D_FlipFlop_7.CLK 0.00406061
R26949 Nand_Gate_2.B.n6 Nand_Gate_2.B.t2 169.46
R26950 Nand_Gate_2.B.n6 Nand_Gate_2.B.t3 167.809
R26951 Nand_Gate_2.B.n5 Nand_Gate_2.B.t1 167.809
R26952 Nand_Gate_2.B Nand_Gate_2.B.t5 158.585
R26953 Nand_Gate_2.B.t5 Nand_Gate_2.B.n2 150.293
R26954 Nand_Gate_2.B.n28 Nand_Gate_2.B.t11 150.273
R26955 Nand_Gate_2.B.n18 Nand_Gate_2.B.t8 150.273
R26956 Nand_Gate_2.B.n12 Nand_Gate_2.B.t4 150.273
R26957 Nand_Gate_2.B.n16 Nand_Gate_2.B.t6 73.6406
R26958 Nand_Gate_2.B.n10 Nand_Gate_2.B.t7 73.6406
R26959 Nand_Gate_2.B.n25 Nand_Gate_2.B.t9 73.6304
R26960 Nand_Gate_2.B.n0 Nand_Gate_2.B.t10 73.6304
R26961 Nand_Gate_2.B.n34 Nand_Gate_2.B.t0 60.3809
R26962 Nand_Gate_2.B.n29 Nand_Gate_2.B.n28 40.8363
R26963 Nand_Gate_2.B.n7 Nand_Gate_2.B.n6 11.4489
R26964 Nand_Gate_2.B.n5 Nand_Gate_2.B.n4 8.21389
R26965 Nand_Gate_2.B.n22 Nand_Gate_2.B.n15 8.1418
R26966 Nand_Gate_2.B.n24 Nand_Gate_2.B.n23 6.47604
R26967 Nand_Gate_2.B.n23 Nand_Gate_2.B 5.35402
R26968 Nand_Gate_2.B.n32 Nand_Gate_2.B 4.55128
R26969 Nand_Gate_2.B.n22 Nand_Gate_2.B.n21 4.5005
R26970 Nand_Gate_2.B.n2 Nand_Gate_2.B.n1 1.19615
R26971 Nand_Gate_2.B.n27 Nand_Gate_2.B.n26 1.1717
R26972 Nand_Gate_2.B.n33 Nand_Gate_2.B 1.08746
R26973 Nand_Gate_2.B.n24 Nand_Gate_2.B 0.973326
R26974 Nand_Gate_2.B.n27 Nand_Gate_2.B 0.932141
R26975 Nand_Gate_2.B.n17 Nand_Gate_2.B 0.851043
R26976 Nand_Gate_2.B.n11 Nand_Gate_2.B 0.851043
R26977 Nand_Gate_2.B Nand_Gate_2.B.n34 0.848156
R26978 Nand_Gate_2.B.n9 Nand_Gate_2.B.n8 0.788543
R26979 Nand_Gate_2.B.n31 Nand_Gate_2.B.n30 0.755935
R26980 Nand_Gate_2.B.n34 Nand_Gate_2.B.n33 0.682565
R26981 Nand_Gate_2.B.n9 Nand_Gate_2.B 0.65675
R26982 Nand_Gate_2.B.n20 Nand_Gate_2.B.n19 0.55213
R26983 Nand_Gate_2.B.n14 Nand_Gate_2.B.n13 0.55213
R26984 Nand_Gate_2.B.n20 Nand_Gate_2.B 0.486828
R26985 Nand_Gate_2.B.n14 Nand_Gate_2.B 0.486828
R26986 Nand_Gate_2.B.n30 Nand_Gate_2.B 0.48023
R26987 Nand_Gate_2.B.n17 Nand_Gate_2.B.n16 0.470609
R26988 Nand_Gate_2.B.n11 Nand_Gate_2.B.n10 0.470609
R26989 Nand_Gate_2.B.n2 Nand_Gate_2.B 0.447191
R26990 Nand_Gate_2.B.n4 Nand_Gate_2.B.n3 0.425067
R26991 Nand_Gate_2.B.n4 Nand_Gate_2.B 0.39003
R26992 Nand_Gate_2.B.n7 Nand_Gate_2.B.n5 0.280391
R26993 Nand_Gate_2.B.n16 Nand_Gate_2.B 0.217464
R26994 Nand_Gate_2.B.n10 Nand_Gate_2.B 0.217464
R26995 Nand_Gate_2.B Nand_Gate_2.B.n7 0.200143
R26996 Nand_Gate_2.B.n26 Nand_Gate_2.B 0.1255
R26997 Nand_Gate_2.B.n19 Nand_Gate_2.B 0.1255
R26998 Nand_Gate_2.B.n13 Nand_Gate_2.B 0.1255
R26999 Nand_Gate_2.B.n1 Nand_Gate_2.B 0.1255
R27000 Nand_Gate_2.B.n8 Nand_Gate_2.B 0.1255
R27001 Nand_Gate_2.B.n28 Nand_Gate_2.B.n27 0.063
R27002 Nand_Gate_2.B.n21 Nand_Gate_2.B.n17 0.063
R27003 Nand_Gate_2.B.n21 Nand_Gate_2.B.n20 0.063
R27004 Nand_Gate_2.B.n15 Nand_Gate_2.B.n11 0.063
R27005 Nand_Gate_2.B.n15 Nand_Gate_2.B.n14 0.063
R27006 Nand_Gate_2.B.n23 Nand_Gate_2.B.n22 0.063
R27007 Nand_Gate_2.B.n29 Nand_Gate_2.B.n24 0.063
R27008 Nand_Gate_2.B.n30 Nand_Gate_2.B.n29 0.063
R27009 Nand_Gate_2.B.n8 Nand_Gate_2.B 0.063
R27010 Nand_Gate_2.B.n33 Nand_Gate_2.B.n32 0.063
R27011 Nand_Gate_2.B.n32 Nand_Gate_2.B.n9 0.063
R27012 Nand_Gate_2.B.n19 Nand_Gate_2.B.n18 0.0216397
R27013 Nand_Gate_2.B.n18 Nand_Gate_2.B 0.0216397
R27014 Nand_Gate_2.B.n13 Nand_Gate_2.B.n12 0.0216397
R27015 Nand_Gate_2.B.n12 Nand_Gate_2.B 0.0216397
R27016 Nand_Gate_2.B.n31 Nand_Gate_2.B 0.0168043
R27017 Nand_Gate_2.B Nand_Gate_2.B.n31 0.0122188
R27018 Nand_Gate_2.B.n26 Nand_Gate_2.B.n25 0.0107679
R27019 Nand_Gate_2.B.n25 Nand_Gate_2.B 0.0107679
R27020 Nand_Gate_2.B.n1 Nand_Gate_2.B.n0 0.0107679
R27021 Nand_Gate_2.B.n0 Nand_Gate_2.B 0.0107679
R27022 Nand_Gate_2.B.n3 Nand_Gate_2.B 0.00441667
R27023 Nand_Gate_2.B.n3 Nand_Gate_2.B 0.00406061
R27024 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 316.762
R27025 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 168.108
R27026 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 150.293
R27027 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 150.273
R27028 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 73.6406
R27029 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 73.6304
R27030 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 60.4568
R27031 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 12.0358
R27032 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 1.19615
R27033 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.981478
R27034 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 0.788543
R27035 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.769522
R27036 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 0.682565
R27037 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.580578
R27038 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 0.55213
R27039 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 0.484875
R27040 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 0.470609
R27041 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.447191
R27042 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.428234
R27043 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.217464
R27044 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R27045 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R27046 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R27047 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 0.063
R27048 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 0.063
R27049 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.063
R27050 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 0.063
R27051 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 0.063
R27052 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 0.0216397
R27053 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.0216397
R27054 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 0.0107679
R27055 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.0107679
R27056 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 179.256
R27057 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 168.089
R27058 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 150.293
R27059 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 73.6304
R27060 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 60.4568
R27061 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 12.0358
R27062 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.981478
R27063 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 0.788543
R27064 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.769522
R27065 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 0.720633
R27066 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 0.682565
R27067 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.580578
R27068 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 0.55213
R27069 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 0.470609
R27070 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.447191
R27071 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.428234
R27072 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1255
R27073 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1255
R27074 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 0.063
R27075 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 0.063
R27076 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.063
R27077 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 0.063
R27078 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 0.063
R27079 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 0.0435206
R27080 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 0.0107679
R27081 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.0107679
R27082 And_Gate_4.Vout.n14 And_Gate_4.Vout.t0 168.108
R27083 And_Gate_4.Vout.n5 And_Gate_4.Vout.t6 158.207
R27084 D_FlipFlop_2.CLK And_Gate_4.Vout.t2 158.202
R27085 And_Gate_4.Vout.n7 And_Gate_4.Vout.t7 150.293
R27086 And_Gate_4.Vout.t2 And_Gate_4.Vout.n10 150.293
R27087 And_Gate_4.Vout.t6 And_Gate_4.Vout.n4 150.273
R27088 And_Gate_4.Vout.n2 And_Gate_4.Vout.t5 73.6406
R27089 And_Gate_4.Vout.n9 And_Gate_4.Vout.t4 73.6304
R27090 And_Gate_4.Vout.n8 And_Gate_4.Vout.t3 73.6304
R27091 And_Gate_4.Vout.n12 And_Gate_4.Vout.n11 62.4488
R27092 And_Gate_4.Inverter_0.Vout And_Gate_4.Vout.t1 60.3943
R27093 And_Gate_4.Vout.n9 And_Gate_4.Vout.n8 16.332
R27094 And_Gate_4.Vout.n3 And_Gate_4.Vout.n2 1.19615
R27095 And_Gate_4.Vout.n8 And_Gate_4.Vout.n7 1.1717
R27096 And_Gate_4.Vout.n10 And_Gate_4.Vout.n9 1.1717
R27097 And_Gate_4.Vout.n13 And_Gate_4.Inverter_0.Vout 0.981478
R27098 And_Gate_4.Vout.n14 And_Gate_4.Vout.n13 0.788543
R27099 And_Gate_4.Vout.n1 And_Gate_4.Vout.n0 0.682565
R27100 And_Gate_4.Vout.n1 And_Gate_4.Inverter_0.Vout 0.580578
R27101 And_Gate_4.Inverter_0.Vout And_Gate_4.Vout.n14 0.484875
R27102 And_Gate_4.Vout.n10 D_FlipFlop_2.3-input-nand_1.C 0.447191
R27103 And_Gate_4.Vout.n7 D_FlipFlop_2.Inverter_1.Vin 0.436162
R27104 And_Gate_4.Vout.n5 D_FlipFlop_2.CLK 0.321667
R27105 And_Gate_4.Vout.n6 And_Gate_4.Vout.n5 0.295033
R27106 And_Gate_4.Vout.n2 D_FlipFlop_2.3-input-nand_0.C 0.217464
R27107 And_Gate_4.Vout.n9 D_FlipFlop_2.3-input-nand_1.C 0.149957
R27108 And_Gate_4.Vout.n3 D_FlipFlop_2.3-input-nand_0.C 0.1255
R27109 And_Gate_4.Vout.n0 And_Gate_4.Inverter_0.Vout 0.1255
R27110 And_Gate_4.Vout.n8 D_FlipFlop_2.Inverter_1.Vin 0.117348
R27111 And_Gate_4.Vout.n0 And_Gate_4.Inverter_0.Vout 0.063
R27112 And_Gate_4.Vout.n13 And_Gate_4.Vout.n12 0.063
R27113 And_Gate_4.Vout.n12 And_Gate_4.Vout.n1 0.063
R27114 And_Gate_4.Vout.n6 D_FlipFlop_2.CLK 0.05925
R27115 And_Gate_4.Vout.n8 D_FlipFlop_2.Inverter_1.Vin 0.0454219
R27116 And_Gate_4.Vout.n9 D_FlipFlop_2.3-input-nand_1.C 0.0454219
R27117 And_Gate_4.Vout.n11 And_Gate_4.Vout.n6 0.024
R27118 And_Gate_4.Vout.n11 D_FlipFlop_2.CLK 0.0233816
R27119 And_Gate_4.Vout.n4 And_Gate_4.Vout.n3 0.0216397
R27120 And_Gate_4.Vout.n4 D_FlipFlop_2.3-input-nand_0.C 0.0216397
R27121 D_FlipFlop_0.CLK.n15 D_FlipFlop_0.CLK.t0 168.108
R27122 D_FlipFlop_0.CLK.n3 D_FlipFlop_0.CLK.t6 158.207
R27123 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.t2 158.202
R27124 D_FlipFlop_0.CLK.n5 D_FlipFlop_0.CLK.t7 150.293
R27125 D_FlipFlop_0.CLK.t2 D_FlipFlop_0.CLK.n8 150.293
R27126 D_FlipFlop_0.CLK.t6 D_FlipFlop_0.CLK.n2 150.273
R27127 D_FlipFlop_0.CLK.n0 D_FlipFlop_0.CLK.t3 73.6406
R27128 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK.t5 73.6304
R27129 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK.t4 73.6304
R27130 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.t1 60.3072
R27131 D_FlipFlop_0.CLK.n12 D_FlipFlop_0.CLK.n11 21.9583
R27132 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK.n6 16.332
R27133 D_FlipFlop_0.CLK.n15 D_FlipFlop_0.CLK.n14 1.62007
R27134 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK.n0 1.19615
R27135 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK.n5 1.1717
R27136 D_FlipFlop_0.CLK.n8 D_FlipFlop_0.CLK.n7 1.1717
R27137 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.n15 0.484875
R27138 D_FlipFlop_0.CLK.n8 D_FlipFlop_0.CLK 0.447191
R27139 D_FlipFlop_0.CLK.n5 D_FlipFlop_0.CLK 0.436162
R27140 D_FlipFlop_0.CLK.n3 D_FlipFlop_0.CLK 0.321667
R27141 D_FlipFlop_0.CLK.n4 D_FlipFlop_0.CLK.n3 0.219833
R27142 D_FlipFlop_0.CLK.n0 D_FlipFlop_0.CLK 0.217464
R27143 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK 0.149957
R27144 D_FlipFlop_0.CLK.n14 D_FlipFlop_0.CLK 0.149957
R27145 D_FlipFlop_0.CLK.n4 D_FlipFlop_0.CLK 0.13445
R27146 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK 0.1255
R27147 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK 0.117348
R27148 D_FlipFlop_0.CLK.n13 D_FlipFlop_0.CLK 0.0903438
R27149 D_FlipFlop_0.CLK.n10 D_FlipFlop_0.CLK.n9 0.071
R27150 D_FlipFlop_0.CLK.n10 D_FlipFlop_0.CLK 0.05925
R27151 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK 0.0454219
R27152 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK 0.0454219
R27153 D_FlipFlop_0.CLK.n13 D_FlipFlop_0.CLK.n12 0.027881
R27154 D_FlipFlop_0.CLK.n12 D_FlipFlop_0.CLK 0.027881
R27155 D_FlipFlop_0.CLK.n11 D_FlipFlop_0.CLK.n4 0.024
R27156 D_FlipFlop_0.CLK.n11 D_FlipFlop_0.CLK.n10 0.024
R27157 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK.n1 0.0216397
R27158 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK 0.0216397
R27159 D_FlipFlop_0.CLK.n14 D_FlipFlop_0.CLK.n13 0.0180781
R27160 D_FlipFlop_0.CLK.n9 D_FlipFlop_0.CLK 0.00441667
R27161 D_FlipFlop_0.CLK.n9 D_FlipFlop_0.CLK 0.00406061
R27162 And_Gate_3.Vout.n12 And_Gate_3.Vout.t0 168.32
R27163 And_Gate_3.Vout.n4 And_Gate_3.Vout.t3 158.226
R27164 D_FlipFlop_4.CLK And_Gate_3.Vout.t6 158.202
R27165 And_Gate_3.Vout.n5 And_Gate_3.Vout.t4 150.293
R27166 And_Gate_3.Vout.t6 And_Gate_3.Vout.n8 150.293
R27167 And_Gate_3.Vout.t3 And_Gate_3.Vout.n3 150.273
R27168 And_Gate_3.Vout.n1 And_Gate_3.Vout.t5 73.6406
R27169 And_Gate_3.Vout.n7 And_Gate_3.Vout.t2 73.6304
R27170 And_Gate_3.Vout.n6 And_Gate_3.Vout.t7 73.6304
R27171 And_Gate_3.Inverter_0.Vout And_Gate_3.Vout.t1 60.3943
R27172 And_Gate_3.Vout.n12 And_Gate_3.Vout.n11 37.7699
R27173 And_Gate_3.Vout.n7 And_Gate_3.Vout.n6 16.332
R27174 And_Gate_3.Vout.n13 And_Gate_3.Vout.n0 1.62007
R27175 And_Gate_3.Inverter_0.Vout And_Gate_3.Vout.n13 1.25441
R27176 And_Gate_3.Vout.n2 And_Gate_3.Vout.n1 1.19615
R27177 And_Gate_3.Vout.n6 And_Gate_3.Vout.n5 1.1717
R27178 And_Gate_3.Vout.n8 And_Gate_3.Vout.n7 1.1717
R27179 And_Gate_3.Vout.n8 D_FlipFlop_4.3-input-nand_1.C 0.447191
R27180 And_Gate_3.Vout.n5 D_FlipFlop_4.Inverter_1.Vin 0.436162
R27181 And_Gate_3.Vout.n4 D_FlipFlop_4.CLK 0.302439
R27182 And_Gate_3.Vout.n10 And_Gate_3.Vout.n9 0.269183
R27183 And_Gate_3.Vout.n1 D_FlipFlop_4.3-input-nand_0.C 0.217464
R27184 And_Gate_3.Vout.n10 D_FlipFlop_4.CLK 0.215711
R27185 And_Gate_3.Vout.n7 D_FlipFlop_4.3-input-nand_1.C 0.149957
R27186 And_Gate_3.Vout.n2 D_FlipFlop_4.3-input-nand_0.C 0.1255
R27187 And_Gate_3.Vout.n0 And_Gate_3.Inverter_0.Vout 0.1255
R27188 And_Gate_3.Vout.n6 D_FlipFlop_4.Inverter_1.Vin 0.117348
R27189 And_Gate_3.Vout.n0 And_Gate_3.Inverter_0.Vout 0.063
R27190 And_Gate_3.Vout.n13 And_Gate_3.Vout.n12 0.063
R27191 And_Gate_3.Vout.n6 D_FlipFlop_4.Inverter_1.Vin 0.0454219
R27192 And_Gate_3.Vout.n7 D_FlipFlop_4.3-input-nand_1.C 0.0454219
R27193 And_Gate_3.Vout.n11 And_Gate_3.Vout.n4 0.024
R27194 And_Gate_3.Vout.n11 And_Gate_3.Vout.n10 0.024
R27195 And_Gate_3.Vout.n3 And_Gate_3.Vout.n2 0.0216397
R27196 And_Gate_3.Vout.n3 D_FlipFlop_4.3-input-nand_0.C 0.0216397
R27197 And_Gate_3.Vout.n9 D_FlipFlop_4.CLK 0.00441667
R27198 And_Gate_3.Vout.n9 D_FlipFlop_4.CLK 0.00406061
R27199 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 316.762
R27200 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 168.108
R27201 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 150.293
R27202 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 150.273
R27203 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 73.6406
R27204 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 73.6304
R27205 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 60.4568
R27206 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 12.0358
R27207 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 1.19615
R27208 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.981478
R27209 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 0.788543
R27210 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.769522
R27211 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 0.682565
R27212 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.580578
R27213 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 0.55213
R27214 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 0.484875
R27215 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 0.470609
R27216 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.447191
R27217 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.428234
R27218 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.217464
R27219 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R27220 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R27221 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R27222 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 0.063
R27223 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 0.063
R27224 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.063
R27225 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 0.063
R27226 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 0.063
R27227 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 0.0216397
R27228 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.0216397
R27229 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 0.0107679
R27230 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.0107679
R27231 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.t3 169.46
R27232 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R27233 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t0 167.809
R27234 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t6 167.226
R27235 D_FlipFlop_2.3-input-nand_2.C.t6 D_FlipFlop_2.3-input-nand_2.C.n10 150.273
R27236 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C.t4 150.273
R27237 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C.t7 73.6406
R27238 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C.t5 73.6304
R27239 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C.t1 60.4568
R27240 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C.n5 12.3891
R27241 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.n12 11.4489
R27242 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C 1.68257
R27243 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C.n0 1.38365
R27244 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C.n8 1.19615
R27245 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C.n3 1.1717
R27246 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C 1.08448
R27247 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C 0.932141
R27248 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.C.n14 0.720633
R27249 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.n11 0.280391
R27250 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C 0.217464
R27251 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27252 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27253 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27254 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.n7 0.0874565
R27255 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C.n4 0.063
R27256 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C 0.063
R27257 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C.n6 0.063
R27258 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C.n1 0.063
R27259 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.n13 0.0435206
R27260 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C.n9 0.0216397
R27261 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C 0.0216397
R27262 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C.n2 0.0107679
R27263 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C 0.0107679
R27264 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.t0 168.553
R27265 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.t2 168.542
R27266 CDAC8_0.switch_9.Z.n0 CDAC8_0.switch_9.Z.t3 60.321
R27267 CDAC8_0.switch_9.Z.n0 CDAC8_0.switch_9.Z.t1 60.321
R27268 CDAC8_0.switch_9.Z.n23 CDAC8_0.switch_9.Z.n22 14.237
R27269 CDAC8_0.switch_9.Z.n36 CDAC8_0.switch_9.Z.n35 11.3711
R27270 CDAC8_0.switch_9.Z.n35 CDAC8_0.switch_9.Z.n5 7.35843
R27271 CDAC8_0.switch_9.Z.n35 CDAC8_0.switch_9.Z.n34 6.87433
R27272 CDAC8_0.switch_9.Z.n2 CDAC8_0.switch_9.Z.n1 1.58202
R27273 CDAC8_0.switch_9.Z.n3 CDAC8_0.switch_9.Z.t25 0.77316
R27274 CDAC8_0.switch_9.Z.n6 CDAC8_0.switch_9.Z.t28 0.77316
R27275 CDAC8_0.switch_9.Z.n8 CDAC8_0.switch_9.Z.t31 0.77316
R27276 CDAC8_0.switch_9.Z.n20 CDAC8_0.switch_9.Z.t29 0.77316
R27277 CDAC8_0.switch_9.Z.n3 CDAC8_0.switch_9.Z.t23 0.611304
R27278 CDAC8_0.switch_9.Z.n4 CDAC8_0.switch_9.Z.t32 0.611304
R27279 CDAC8_0.switch_9.Z.n10 CDAC8_0.switch_9.Z.t30 0.611304
R27280 CDAC8_0.switch_9.Z.n11 CDAC8_0.switch_9.Z.t10 0.611304
R27281 CDAC8_0.switch_9.Z.n12 CDAC8_0.switch_9.Z.t14 0.611304
R27282 CDAC8_0.switch_9.Z.n13 CDAC8_0.switch_9.Z.t13 0.611304
R27283 CDAC8_0.switch_9.Z.n14 CDAC8_0.switch_9.Z.t18 0.611304
R27284 CDAC8_0.switch_9.Z.n15 CDAC8_0.switch_9.Z.t17 0.611304
R27285 CDAC8_0.switch_9.Z.n16 CDAC8_0.switch_9.Z.t34 0.611304
R27286 CDAC8_0.switch_9.Z.n17 CDAC8_0.switch_9.Z.t6 0.611304
R27287 CDAC8_0.switch_9.Z.n18 CDAC8_0.switch_9.Z.t5 0.611304
R27288 CDAC8_0.switch_9.Z.n19 CDAC8_0.switch_9.Z.t9 0.611304
R27289 CDAC8_0.switch_9.Z.n6 CDAC8_0.switch_9.Z.t27 0.611304
R27290 CDAC8_0.switch_9.Z.n7 CDAC8_0.switch_9.Z.t35 0.611304
R27291 CDAC8_0.switch_9.Z.n33 CDAC8_0.switch_9.Z.t33 0.611304
R27292 CDAC8_0.switch_9.Z.n32 CDAC8_0.switch_9.Z.t12 0.611304
R27293 CDAC8_0.switch_9.Z.n31 CDAC8_0.switch_9.Z.t16 0.611304
R27294 CDAC8_0.switch_9.Z.n30 CDAC8_0.switch_9.Z.t15 0.611304
R27295 CDAC8_0.switch_9.Z.n29 CDAC8_0.switch_9.Z.t21 0.611304
R27296 CDAC8_0.switch_9.Z.n28 CDAC8_0.switch_9.Z.t19 0.611304
R27297 CDAC8_0.switch_9.Z.n27 CDAC8_0.switch_9.Z.t4 0.611304
R27298 CDAC8_0.switch_9.Z.n26 CDAC8_0.switch_9.Z.t8 0.611304
R27299 CDAC8_0.switch_9.Z.n25 CDAC8_0.switch_9.Z.t7 0.611304
R27300 CDAC8_0.switch_9.Z.n24 CDAC8_0.switch_9.Z.t11 0.611304
R27301 CDAC8_0.switch_9.Z.n9 CDAC8_0.switch_9.Z.t26 0.611304
R27302 CDAC8_0.switch_9.Z.n8 CDAC8_0.switch_9.Z.t24 0.611304
R27303 CDAC8_0.switch_9.Z.n21 CDAC8_0.switch_9.Z.t22 0.611304
R27304 CDAC8_0.switch_9.Z.n20 CDAC8_0.switch_9.Z.t20 0.611304
R27305 CDAC8_0.switch_9.Z.n1 CDAC8_0.switch_9.Z 0.259656
R27306 CDAC8_0.switch_9.Z.n2 CDAC8_0.switch_9.Z 0.188
R27307 CDAC8_0.switch_9.Z.n7 CDAC8_0.switch_9.Z.n6 0.162356
R27308 CDAC8_0.switch_9.Z.n33 CDAC8_0.switch_9.Z.n32 0.162356
R27309 CDAC8_0.switch_9.Z.n32 CDAC8_0.switch_9.Z.n31 0.162356
R27310 CDAC8_0.switch_9.Z.n31 CDAC8_0.switch_9.Z.n30 0.162356
R27311 CDAC8_0.switch_9.Z.n30 CDAC8_0.switch_9.Z.n29 0.162356
R27312 CDAC8_0.switch_9.Z.n29 CDAC8_0.switch_9.Z.n28 0.162356
R27313 CDAC8_0.switch_9.Z.n28 CDAC8_0.switch_9.Z.n27 0.162356
R27314 CDAC8_0.switch_9.Z.n27 CDAC8_0.switch_9.Z.n26 0.162356
R27315 CDAC8_0.switch_9.Z.n26 CDAC8_0.switch_9.Z.n25 0.162356
R27316 CDAC8_0.switch_9.Z.n25 CDAC8_0.switch_9.Z.n24 0.162356
R27317 CDAC8_0.switch_9.Z.n9 CDAC8_0.switch_9.Z.n8 0.162356
R27318 CDAC8_0.switch_9.Z.n4 CDAC8_0.switch_9.Z.n3 0.162356
R27319 CDAC8_0.switch_9.Z.n11 CDAC8_0.switch_9.Z.n10 0.162356
R27320 CDAC8_0.switch_9.Z.n12 CDAC8_0.switch_9.Z.n11 0.162356
R27321 CDAC8_0.switch_9.Z.n13 CDAC8_0.switch_9.Z.n12 0.162356
R27322 CDAC8_0.switch_9.Z.n14 CDAC8_0.switch_9.Z.n13 0.162356
R27323 CDAC8_0.switch_9.Z.n15 CDAC8_0.switch_9.Z.n14 0.162356
R27324 CDAC8_0.switch_9.Z.n16 CDAC8_0.switch_9.Z.n15 0.162356
R27325 CDAC8_0.switch_9.Z.n17 CDAC8_0.switch_9.Z.n16 0.162356
R27326 CDAC8_0.switch_9.Z.n18 CDAC8_0.switch_9.Z.n17 0.162356
R27327 CDAC8_0.switch_9.Z.n19 CDAC8_0.switch_9.Z.n18 0.162356
R27328 CDAC8_0.switch_9.Z.n21 CDAC8_0.switch_9.Z.n20 0.162356
R27329 CDAC8_0.switch_9.Z.n34 CDAC8_0.switch_9.Z.n33 0.115412
R27330 CDAC8_0.switch_9.Z.n10 CDAC8_0.switch_9.Z.n5 0.115412
R27331 CDAC8_0.switch_9.Z.n23 CDAC8_0.switch_9.Z.n9 0.0845094
R27332 CDAC8_0.switch_9.Z.n22 CDAC8_0.switch_9.Z.n21 0.0845094
R27333 CDAC8_0.switch_9.Z.n24 CDAC8_0.switch_9.Z.n23 0.0783469
R27334 CDAC8_0.switch_9.Z.n22 CDAC8_0.switch_9.Z.n19 0.0783469
R27335 CDAC8_0.switch_9.Z.n36 CDAC8_0.switch_9.Z.n2 0.063
R27336 CDAC8_0.switch_9.Z.n34 CDAC8_0.switch_9.Z.n7 0.0474438
R27337 CDAC8_0.switch_9.Z.n5 CDAC8_0.switch_9.Z.n4 0.0474438
R27338 CDAC8_0.switch_9.Z CDAC8_0.switch_9.Z.n37 0.0454219
R27339 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.n36 0.0278438
R27340 CDAC8_0.switch_9.Z.n1 CDAC8_0.switch_9.Z.n0 0.0188121
R27341 Nand_Gate_5.B.n24 Nand_Gate_5.B.t3 169.46
R27342 Nand_Gate_5.B.n26 Nand_Gate_5.B.t2 167.809
R27343 Nand_Gate_5.B.n24 Nand_Gate_5.B.t0 167.809
R27344 Nand_Gate_5.B Nand_Gate_5.B.t7 158.585
R27345 Nand_Gate_5.B.t7 Nand_Gate_5.B.n20 150.293
R27346 Nand_Gate_5.B.n16 Nand_Gate_5.B.t6 150.273
R27347 Nand_Gate_5.B.n5 Nand_Gate_5.B.t11 150.273
R27348 Nand_Gate_5.B.n0 Nand_Gate_5.B.t9 150.273
R27349 Nand_Gate_5.B.t5 Nand_Gate_5.B.n17 82.5626
R27350 Nand_Gate_5.B Nand_Gate_5.B.t10 81.5603
R27351 Nand_Gate_5.B.n3 Nand_Gate_5.B.t8 73.6406
R27352 Nand_Gate_5.B.t10 Nand_Gate_5.B.n11 73.6406
R27353 Nand_Gate_5.B.n13 Nand_Gate_5.B.t4 73.6304
R27354 Nand_Gate_5.B.n18 Nand_Gate_5.B.t5 73.6304
R27355 Nand_Gate_5.B.n22 Nand_Gate_5.B.t1 60.3809
R27356 Nand_Gate_5.B.n17 Nand_Gate_5.B.n16 32.9078
R27357 Nand_Gate_5.B.n17 Nand_Gate_5.B.n12 25.3147
R27358 Nand_Gate_5.B.n9 Nand_Gate_5.B.n8 12.6418
R27359 Nand_Gate_5.B.n25 Nand_Gate_5.B.n24 11.4489
R27360 Nand_Gate_5.B.n27 Nand_Gate_5.B.n26 8.21389
R27361 Nand_Gate_5.B.n23 Nand_Gate_5.B.n22 1.64452
R27362 Nand_Gate_5.B.n20 Nand_Gate_5.B.n19 1.19615
R27363 Nand_Gate_5.B.n15 Nand_Gate_5.B.n14 1.1717
R27364 Nand_Gate_5.B.n15 Nand_Gate_5.B 0.932141
R27365 Nand_Gate_5.B.n4 Nand_Gate_5.B 0.851043
R27366 Nand_Gate_5.B.n10 Nand_Gate_5.B 0.851043
R27367 Nand_Gate_5.B.n22 Nand_Gate_5.B 0.848156
R27368 Nand_Gate_5.B.n7 Nand_Gate_5.B.n6 0.55213
R27369 Nand_Gate_5.B.n2 Nand_Gate_5.B.n1 0.55213
R27370 Nand_Gate_5.B.n7 Nand_Gate_5.B 0.486828
R27371 Nand_Gate_5.B.n2 Nand_Gate_5.B 0.486828
R27372 Nand_Gate_5.B.n4 Nand_Gate_5.B.n3 0.470609
R27373 Nand_Gate_5.B.n11 Nand_Gate_5.B.n10 0.470609
R27374 Nand_Gate_5.B.n20 Nand_Gate_5.B 0.447191
R27375 Nand_Gate_5.B.n27 Nand_Gate_5.B.n21 0.425067
R27376 Nand_Gate_5.B Nand_Gate_5.B.n27 0.39003
R27377 Nand_Gate_5.B.n26 Nand_Gate_5.B.n25 0.280391
R27378 Nand_Gate_5.B.n3 Nand_Gate_5.B 0.217464
R27379 Nand_Gate_5.B.n11 Nand_Gate_5.B 0.217464
R27380 Nand_Gate_5.B.n25 Nand_Gate_5.B 0.200143
R27381 Nand_Gate_5.B.n23 Nand_Gate_5.B 0.1255
R27382 Nand_Gate_5.B.n14 Nand_Gate_5.B 0.1255
R27383 Nand_Gate_5.B.n6 Nand_Gate_5.B 0.1255
R27384 Nand_Gate_5.B.n1 Nand_Gate_5.B 0.1255
R27385 Nand_Gate_5.B.n19 Nand_Gate_5.B 0.1255
R27386 Nand_Gate_5.B Nand_Gate_5.B.n23 0.063
R27387 Nand_Gate_5.B.n16 Nand_Gate_5.B.n15 0.063
R27388 Nand_Gate_5.B.n8 Nand_Gate_5.B.n4 0.063
R27389 Nand_Gate_5.B.n8 Nand_Gate_5.B.n7 0.063
R27390 Nand_Gate_5.B.n10 Nand_Gate_5.B.n9 0.063
R27391 Nand_Gate_5.B.n9 Nand_Gate_5.B.n2 0.063
R27392 Nand_Gate_5.B.n6 Nand_Gate_5.B.n5 0.0216397
R27393 Nand_Gate_5.B.n5 Nand_Gate_5.B 0.0216397
R27394 Nand_Gate_5.B.n1 Nand_Gate_5.B.n0 0.0216397
R27395 Nand_Gate_5.B.n0 Nand_Gate_5.B 0.0216397
R27396 Nand_Gate_5.B.n14 Nand_Gate_5.B.n13 0.0107679
R27397 Nand_Gate_5.B.n13 Nand_Gate_5.B 0.0107679
R27398 Nand_Gate_5.B.n19 Nand_Gate_5.B.n18 0.0107679
R27399 Nand_Gate_5.B.n18 Nand_Gate_5.B 0.0107679
R27400 Nand_Gate_5.B.n12 Nand_Gate_5.B 0.00441667
R27401 Nand_Gate_5.B.n21 Nand_Gate_5.B 0.00441667
R27402 Nand_Gate_5.B.n12 Nand_Gate_5.B 0.00406061
R27403 Nand_Gate_5.B.n21 Nand_Gate_5.B 0.00406061
R27404 Nand_Gate_6.A.n33 Nand_Gate_6.A.t1 169.46
R27405 Nand_Gate_6.A.n35 Nand_Gate_6.A.t3 167.809
R27406 Nand_Gate_6.A.n33 Nand_Gate_6.A.t0 167.809
R27407 Nand_Gate_6.A Nand_Gate_6.A.t11 158.585
R27408 Nand_Gate_6.A.n21 Nand_Gate_6.A.t9 150.293
R27409 Nand_Gate_6.A.t11 Nand_Gate_6.A.n2 150.293
R27410 Nand_Gate_6.A.n14 Nand_Gate_6.A.t8 150.273
R27411 Nand_Gate_6.A.n8 Nand_Gate_6.A.t10 150.273
R27412 Nand_Gate_6.A.n12 Nand_Gate_6.A.t6 73.6406
R27413 Nand_Gate_6.A.n6 Nand_Gate_6.A.t4 73.6406
R27414 Nand_Gate_6.A.n23 Nand_Gate_6.A.t5 73.6304
R27415 Nand_Gate_6.A.n0 Nand_Gate_6.A.t7 73.6304
R27416 Nand_Gate_6.A.n4 Nand_Gate_6.A.t2 60.3809
R27417 Nand_Gate_6.A.n27 Nand_Gate_6.A.n26 14.3097
R27418 Nand_Gate_6.A.n34 Nand_Gate_6.A.n33 11.4489
R27419 Nand_Gate_6.A.n36 Nand_Gate_6.A.n35 8.21389
R27420 Nand_Gate_6.A.n18 Nand_Gate_6.A.n11 8.1418
R27421 Nand_Gate_6.A.n29 Nand_Gate_6.A.n28 5.61191
R27422 Nand_Gate_6.A.n29 Nand_Gate_6.A 5.35402
R27423 Nand_Gate_6.A.n30 Nand_Gate_6.A.n29 4.563
R27424 Nand_Gate_6.A.n18 Nand_Gate_6.A.n17 4.5005
R27425 Nand_Gate_6.A.n28 Nand_Gate_6.A 1.83746
R27426 Nand_Gate_6.A.n20 Nand_Gate_6.A.n19 1.62007
R27427 Nand_Gate_6.A.n2 Nand_Gate_6.A.n1 1.19615
R27428 Nand_Gate_6.A.n5 Nand_Gate_6.A 1.08746
R27429 Nand_Gate_6.A.n20 Nand_Gate_6.A 1.01739
R27430 Nand_Gate_6.A.n13 Nand_Gate_6.A 0.851043
R27431 Nand_Gate_6.A.n7 Nand_Gate_6.A 0.851043
R27432 Nand_Gate_6.A.n4 Nand_Gate_6.A 0.848156
R27433 Nand_Gate_6.A.n32 Nand_Gate_6.A.n31 0.788543
R27434 Nand_Gate_6.A.n22 Nand_Gate_6.A 0.769522
R27435 Nand_Gate_6.A.n5 Nand_Gate_6.A.n4 0.682565
R27436 Nand_Gate_6.A.n31 Nand_Gate_6.A 0.65675
R27437 Nand_Gate_6.A.n22 Nand_Gate_6.A.n21 0.55213
R27438 Nand_Gate_6.A.n16 Nand_Gate_6.A.n15 0.55213
R27439 Nand_Gate_6.A.n10 Nand_Gate_6.A.n9 0.55213
R27440 Nand_Gate_6.A.n16 Nand_Gate_6.A 0.486828
R27441 Nand_Gate_6.A.n10 Nand_Gate_6.A 0.486828
R27442 Nand_Gate_6.A.n25 Nand_Gate_6.A.n24 0.470609
R27443 Nand_Gate_6.A.n13 Nand_Gate_6.A.n12 0.470609
R27444 Nand_Gate_6.A.n7 Nand_Gate_6.A.n6 0.470609
R27445 Nand_Gate_6.A.n21 Nand_Gate_6.A 0.447191
R27446 Nand_Gate_6.A.n2 Nand_Gate_6.A 0.447191
R27447 Nand_Gate_6.A.n25 Nand_Gate_6.A 0.428234
R27448 Nand_Gate_6.A.n36 Nand_Gate_6.A.n3 0.425067
R27449 Nand_Gate_6.A Nand_Gate_6.A.n36 0.39003
R27450 Nand_Gate_6.A.n35 Nand_Gate_6.A.n34 0.280391
R27451 Nand_Gate_6.A.n34 Nand_Gate_6.A.n32 0.262643
R27452 Nand_Gate_6.A.n12 Nand_Gate_6.A 0.217464
R27453 Nand_Gate_6.A.n6 Nand_Gate_6.A 0.217464
R27454 Nand_Gate_6.A.n24 Nand_Gate_6.A 0.1255
R27455 Nand_Gate_6.A.n15 Nand_Gate_6.A 0.1255
R27456 Nand_Gate_6.A.n9 Nand_Gate_6.A 0.1255
R27457 Nand_Gate_6.A.n32 Nand_Gate_6.A 0.1255
R27458 Nand_Gate_6.A.n1 Nand_Gate_6.A 0.1255
R27459 Nand_Gate_6.A.n26 Nand_Gate_6.A.n22 0.063
R27460 Nand_Gate_6.A.n26 Nand_Gate_6.A.n25 0.063
R27461 Nand_Gate_6.A.n17 Nand_Gate_6.A.n13 0.063
R27462 Nand_Gate_6.A.n17 Nand_Gate_6.A.n16 0.063
R27463 Nand_Gate_6.A.n11 Nand_Gate_6.A.n7 0.063
R27464 Nand_Gate_6.A.n11 Nand_Gate_6.A.n10 0.063
R27465 Nand_Gate_6.A.n28 Nand_Gate_6.A.n27 0.063
R27466 Nand_Gate_6.A.n27 Nand_Gate_6.A.n20 0.063
R27467 Nand_Gate_6.A.n30 Nand_Gate_6.A.n5 0.063
R27468 Nand_Gate_6.A.n31 Nand_Gate_6.A.n30 0.063
R27469 Nand_Gate_6.A.n32 Nand_Gate_6.A 0.063
R27470 Nand_Gate_6.A Nand_Gate_6.A.n18 0.0512812
R27471 Nand_Gate_6.A.n15 Nand_Gate_6.A.n14 0.0216397
R27472 Nand_Gate_6.A.n14 Nand_Gate_6.A 0.0216397
R27473 Nand_Gate_6.A.n9 Nand_Gate_6.A.n8 0.0216397
R27474 Nand_Gate_6.A.n8 Nand_Gate_6.A 0.0216397
R27475 Nand_Gate_6.A.n19 Nand_Gate_6.A 0.0168043
R27476 Nand_Gate_6.A.n19 Nand_Gate_6.A 0.0122188
R27477 Nand_Gate_6.A.n24 Nand_Gate_6.A.n23 0.0107679
R27478 Nand_Gate_6.A.n23 Nand_Gate_6.A 0.0107679
R27479 Nand_Gate_6.A.n1 Nand_Gate_6.A.n0 0.0107679
R27480 Nand_Gate_6.A.n0 Nand_Gate_6.A 0.0107679
R27481 Nand_Gate_6.A.n3 Nand_Gate_6.A 0.00441667
R27482 Nand_Gate_6.A.n3 Nand_Gate_6.A 0.00406061
R27483 FFCLR.n205 FFCLR.t1 169.46
R27484 FFCLR.n207 FFCLR.t3 167.809
R27485 FFCLR.n205 FFCLR.t0 167.809
R27486 FFCLR.n45 FFCLR.t27 158.988
R27487 FFCLR.n84 FFCLR.t7 158.965
R27488 FFCLR.n64 FFCLR.t45 158.965
R27489 FFCLR.n187 FFCLR.t55 158.965
R27490 FFCLR.n165 FFCLR.t5 158.965
R27491 FFCLR.n143 FFCLR.t9 158.965
R27492 FFCLR.n121 FFCLR.t49 158.965
R27493 FFCLR FFCLR.t6 158.585
R27494 FFCLR FFCLR.t44 158.581
R27495 FFCLR.n192 FFCLR.t16 150.293
R27496 FFCLR.n93 FFCLR.t56 150.293
R27497 FFCLR.n87 FFCLR.t24 150.293
R27498 FFCLR.n73 FFCLR.t22 150.293
R27499 FFCLR.n67 FFCLR.t50 150.293
R27500 FFCLR.n53 FFCLR.t8 150.293
R27501 FFCLR.n47 FFCLR.t33 150.293
R27502 FFCLR.n174 FFCLR.t30 150.293
R27503 FFCLR.n168 FFCLR.t58 150.293
R27504 FFCLR.n152 FFCLR.t51 150.293
R27505 FFCLR.n146 FFCLR.t21 150.293
R27506 FFCLR.n130 FFCLR.t36 150.293
R27507 FFCLR.n124 FFCLR.t10 150.293
R27508 FFCLR.n108 FFCLR.t28 150.293
R27509 FFCLR.n102 FFCLR.t54 150.293
R27510 FFCLR.t44 FFCLR.n38 150.293
R27511 FFCLR.t6 FFCLR.n2 150.293
R27512 FFCLR.t7 FFCLR.n83 150.273
R27513 FFCLR.t45 FFCLR.n63 150.273
R27514 FFCLR.t27 FFCLR.n44 150.273
R27515 FFCLR.t55 FFCLR.n186 150.273
R27516 FFCLR.t5 FFCLR.n164 150.273
R27517 FFCLR.t9 FFCLR.n142 150.273
R27518 FFCLR.t49 FFCLR.n120 150.273
R27519 FFCLR.n29 FFCLR.t38 150.273
R27520 FFCLR.n23 FFCLR.t11 150.273
R27521 FFCLR.n14 FFCLR.t40 150.273
R27522 FFCLR.n8 FFCLR.t34 150.273
R27523 FFCLR.n198 FFCLR.n191 88.4503
R27524 FFCLR.n81 FFCLR.t14 73.6406
R27525 FFCLR.n61 FFCLR.t37 73.6406
R27526 FFCLR.n42 FFCLR.t19 73.6406
R27527 FFCLR.n184 FFCLR.t20 73.6406
R27528 FFCLR.n162 FFCLR.t52 73.6406
R27529 FFCLR.n140 FFCLR.t15 73.6406
R27530 FFCLR.n118 FFCLR.t43 73.6406
R27531 FFCLR.n27 FFCLR.t13 73.6406
R27532 FFCLR.n21 FFCLR.t39 73.6406
R27533 FFCLR.n12 FFCLR.t32 73.6406
R27534 FFCLR.n6 FFCLR.t41 73.6406
R27535 FFCLR.n194 FFCLR.t48 73.6304
R27536 FFCLR.n95 FFCLR.t4 73.6304
R27537 FFCLR.n89 FFCLR.t31 73.6304
R27538 FFCLR.n75 FFCLR.t42 73.6304
R27539 FFCLR.n69 FFCLR.t12 73.6304
R27540 FFCLR.n55 FFCLR.t23 73.6304
R27541 FFCLR.n49 FFCLR.t53 73.6304
R27542 FFCLR.n176 FFCLR.t47 73.6304
R27543 FFCLR.n170 FFCLR.t18 73.6304
R27544 FFCLR.n154 FFCLR.t57 73.6304
R27545 FFCLR.n148 FFCLR.t25 73.6304
R27546 FFCLR.n132 FFCLR.t59 73.6304
R27547 FFCLR.n126 FFCLR.t29 73.6304
R27548 FFCLR.n110 FFCLR.t46 73.6304
R27549 FFCLR.n104 FFCLR.t17 73.6304
R27550 FFCLR.n36 FFCLR.t26 73.6304
R27551 FFCLR.n0 FFCLR.t35 73.6304
R27552 FFCLR.n4 FFCLR.t2 60.3809
R27553 FFCLR.n99 FFCLR.n92 15.5222
R27554 FFCLR.n79 FFCLR.n72 15.5222
R27555 FFCLR.n59 FFCLR.n52 15.5222
R27556 FFCLR.n180 FFCLR.n173 15.5222
R27557 FFCLR.n158 FFCLR.n151 15.5222
R27558 FFCLR.n136 FFCLR.n129 15.5222
R27559 FFCLR.n114 FFCLR.n107 15.5222
R27560 FFCLR.n33 FFCLR.n26 15.5222
R27561 FFCLR.n206 FFCLR.n205 11.4489
R27562 FFCLR.n189 FFCLR 10.7094
R27563 FFCLR.n190 FFCLR.n100 9.59712
R27564 FFCLR.n198 FFCLR.n197 9.57083
R27565 FFCLR.n188 FFCLR 9.51957
R27566 FFCLR.n190 FFCLR.n189 9.43184
R27567 FFCLR.n34 FFCLR.n33 8.26552
R27568 FFCLR.n208 FFCLR.n207 8.21389
R27569 FFCLR.n18 FFCLR.n11 8.1418
R27570 FFCLR.n167 FFCLR 7.84808
R27571 FFCLR.n100 FFCLR.n99 7.83713
R27572 FFCLR.n80 FFCLR.n79 7.83713
R27573 FFCLR.n60 FFCLR.n59 7.83713
R27574 FFCLR.n181 FFCLR.n180 7.83713
R27575 FFCLR.n159 FFCLR.n158 7.83713
R27576 FFCLR.n137 FFCLR.n136 7.83713
R27577 FFCLR.n115 FFCLR.n114 7.83713
R27578 FFCLR.n166 FFCLR 6.72777
R27579 FFCLR.n199 FFCLR.n198 6.58222
R27580 FFCLR.n20 FFCLR.n19 6.47604
R27581 FFCLR.n19 FFCLR 5.35402
R27582 FFCLR.n145 FFCLR 5.31008
R27583 FFCLR.n202 FFCLR 4.55128
R27584 FFCLR.n99 FFCLR.n98 4.5005
R27585 FFCLR.n79 FFCLR.n78 4.5005
R27586 FFCLR.n59 FFCLR.n58 4.5005
R27587 FFCLR.n180 FFCLR.n179 4.5005
R27588 FFCLR.n158 FFCLR.n157 4.5005
R27589 FFCLR.n136 FFCLR.n135 4.5005
R27590 FFCLR.n114 FFCLR.n113 4.5005
R27591 FFCLR.n33 FFCLR.n32 4.5005
R27592 FFCLR.n18 FFCLR.n17 4.5005
R27593 FFCLR.n144 FFCLR 3.93597
R27594 FFCLR.n191 FFCLR.n41 3.73088
R27595 FFCLR.n191 FFCLR.n190 3.4105
R27596 FFCLR.n123 FFCLR 2.77208
R27597 FFCLR.n189 FFCLR.n188 2.2612
R27598 FFCLR.n64 FFCLR.n60 1.95257
R27599 FFCLR.n84 FFCLR.n80 1.95257
R27600 FFCLR.n123 FFCLR.n122 1.90557
R27601 FFCLR.n145 FFCLR.n144 1.90557
R27602 FFCLR.n167 FFCLR.n166 1.90557
R27603 FFCLR.n82 FFCLR.n81 1.19615
R27604 FFCLR.n62 FFCLR.n61 1.19615
R27605 FFCLR.n43 FFCLR.n42 1.19615
R27606 FFCLR.n185 FFCLR.n184 1.19615
R27607 FFCLR.n163 FFCLR.n162 1.19615
R27608 FFCLR.n141 FFCLR.n140 1.19615
R27609 FFCLR.n119 FFCLR.n118 1.19615
R27610 FFCLR.n38 FFCLR.n37 1.19615
R27611 FFCLR.n2 FFCLR.n1 1.19615
R27612 FFCLR.n122 FFCLR 1.14417
R27613 FFCLR.n94 FFCLR 1.09561
R27614 FFCLR.n88 FFCLR 1.09561
R27615 FFCLR.n74 FFCLR 1.09561
R27616 FFCLR.n68 FFCLR 1.09561
R27617 FFCLR.n54 FFCLR 1.09561
R27618 FFCLR.n48 FFCLR 1.09561
R27619 FFCLR.n175 FFCLR 1.09561
R27620 FFCLR.n169 FFCLR 1.09561
R27621 FFCLR.n153 FFCLR 1.09561
R27622 FFCLR.n147 FFCLR 1.09561
R27623 FFCLR.n131 FFCLR 1.09561
R27624 FFCLR.n125 FFCLR 1.09561
R27625 FFCLR.n109 FFCLR 1.09561
R27626 FFCLR.n103 FFCLR 1.09561
R27627 FFCLR.n5 FFCLR 1.08746
R27628 FFCLR.n20 FFCLR 0.973326
R27629 FFCLR.n13 FFCLR 0.851043
R27630 FFCLR.n7 FFCLR 0.851043
R27631 FFCLR.n4 FFCLR 0.848156
R27632 FFCLR.n97 FFCLR.n96 0.796696
R27633 FFCLR.n91 FFCLR.n90 0.796696
R27634 FFCLR.n77 FFCLR.n76 0.796696
R27635 FFCLR.n71 FFCLR.n70 0.796696
R27636 FFCLR.n57 FFCLR.n56 0.796696
R27637 FFCLR.n51 FFCLR.n50 0.796696
R27638 FFCLR.n178 FFCLR.n177 0.796696
R27639 FFCLR.n172 FFCLR.n171 0.796696
R27640 FFCLR.n156 FFCLR.n155 0.796696
R27641 FFCLR.n150 FFCLR.n149 0.796696
R27642 FFCLR.n134 FFCLR.n133 0.796696
R27643 FFCLR.n128 FFCLR.n127 0.796696
R27644 FFCLR.n112 FFCLR.n111 0.796696
R27645 FFCLR.n106 FFCLR.n105 0.796696
R27646 FFCLR.n28 FFCLR.n27 0.796696
R27647 FFCLR.n22 FFCLR.n21 0.796696
R27648 FFCLR.n204 FFCLR.n203 0.788543
R27649 FFCLR.n46 FFCLR.n45 0.783833
R27650 FFCLR.n66 FFCLR.n65 0.783833
R27651 FFCLR.n86 FFCLR.n85 0.783833
R27652 FFCLR.n117 FFCLR.n116 0.783833
R27653 FFCLR.n139 FFCLR.n138 0.783833
R27654 FFCLR.n161 FFCLR.n160 0.783833
R27655 FFCLR.n183 FFCLR.n182 0.783833
R27656 FFCLR.n193 FFCLR 0.769522
R27657 FFCLR.n201 FFCLR.n200 0.755935
R27658 FFCLR.n45 FFCLR 0.716182
R27659 FFCLR.n65 FFCLR 0.716182
R27660 FFCLR.n85 FFCLR 0.716182
R27661 FFCLR.n117 FFCLR 0.716182
R27662 FFCLR.n139 FFCLR 0.716182
R27663 FFCLR.n161 FFCLR 0.716182
R27664 FFCLR.n183 FFCLR 0.716182
R27665 FFCLR.n34 FFCLR 0.716182
R27666 FFCLR.n5 FFCLR.n4 0.682565
R27667 FFCLR.n97 FFCLR 0.662609
R27668 FFCLR.n91 FFCLR 0.662609
R27669 FFCLR.n77 FFCLR 0.662609
R27670 FFCLR.n71 FFCLR 0.662609
R27671 FFCLR.n57 FFCLR 0.662609
R27672 FFCLR.n51 FFCLR 0.662609
R27673 FFCLR.n178 FFCLR 0.662609
R27674 FFCLR.n172 FFCLR 0.662609
R27675 FFCLR.n156 FFCLR 0.662609
R27676 FFCLR.n150 FFCLR 0.662609
R27677 FFCLR.n134 FFCLR 0.662609
R27678 FFCLR.n128 FFCLR 0.662609
R27679 FFCLR.n112 FFCLR 0.662609
R27680 FFCLR.n106 FFCLR 0.662609
R27681 FFCLR.n203 FFCLR 0.65675
R27682 FFCLR.n35 FFCLR.n34 0.565283
R27683 FFCLR.n193 FFCLR.n192 0.55213
R27684 FFCLR.n16 FFCLR.n15 0.55213
R27685 FFCLR.n10 FFCLR.n9 0.55213
R27686 FFCLR.n28 FFCLR 0.524957
R27687 FFCLR.n22 FFCLR 0.524957
R27688 FFCLR.n16 FFCLR 0.486828
R27689 FFCLR.n10 FFCLR 0.486828
R27690 FFCLR.n200 FFCLR 0.48023
R27691 FFCLR.n196 FFCLR.n195 0.470609
R27692 FFCLR.n13 FFCLR.n12 0.470609
R27693 FFCLR.n7 FFCLR.n6 0.470609
R27694 FFCLR.n192 FFCLR 0.447191
R27695 FFCLR.n93 FFCLR 0.447191
R27696 FFCLR.n87 FFCLR 0.447191
R27697 FFCLR.n73 FFCLR 0.447191
R27698 FFCLR.n67 FFCLR 0.447191
R27699 FFCLR.n53 FFCLR 0.447191
R27700 FFCLR.n47 FFCLR 0.447191
R27701 FFCLR.n174 FFCLR 0.447191
R27702 FFCLR.n168 FFCLR 0.447191
R27703 FFCLR.n152 FFCLR 0.447191
R27704 FFCLR.n146 FFCLR 0.447191
R27705 FFCLR.n130 FFCLR 0.447191
R27706 FFCLR.n124 FFCLR 0.447191
R27707 FFCLR.n108 FFCLR 0.447191
R27708 FFCLR.n102 FFCLR 0.447191
R27709 FFCLR.n38 FFCLR 0.447191
R27710 FFCLR.n2 FFCLR 0.447191
R27711 FFCLR.n196 FFCLR 0.428234
R27712 FFCLR.n208 FFCLR.n3 0.425067
R27713 FFCLR FFCLR.n208 0.39003
R27714 FFCLR.n207 FFCLR.n206 0.280391
R27715 FFCLR.n101 FFCLR 0.257433
R27716 FFCLR.n31 FFCLR 0.252453
R27717 FFCLR.n25 FFCLR 0.252453
R27718 FFCLR.n101 FFCLR 0.234076
R27719 FFCLR.n94 FFCLR.n93 0.226043
R27720 FFCLR.n88 FFCLR.n87 0.226043
R27721 FFCLR.n74 FFCLR.n73 0.226043
R27722 FFCLR.n68 FFCLR.n67 0.226043
R27723 FFCLR.n54 FFCLR.n53 0.226043
R27724 FFCLR.n48 FFCLR.n47 0.226043
R27725 FFCLR.n175 FFCLR.n174 0.226043
R27726 FFCLR.n169 FFCLR.n168 0.226043
R27727 FFCLR.n153 FFCLR.n152 0.226043
R27728 FFCLR.n147 FFCLR.n146 0.226043
R27729 FFCLR.n131 FFCLR.n130 0.226043
R27730 FFCLR.n125 FFCLR.n124 0.226043
R27731 FFCLR.n109 FFCLR.n108 0.226043
R27732 FFCLR.n103 FFCLR.n102 0.226043
R27733 FFCLR.n31 FFCLR.n30 0.226043
R27734 FFCLR.n25 FFCLR.n24 0.226043
R27735 FFCLR.n35 FFCLR 0.222967
R27736 FFCLR.n81 FFCLR 0.217464
R27737 FFCLR.n61 FFCLR 0.217464
R27738 FFCLR.n42 FFCLR 0.217464
R27739 FFCLR.n184 FFCLR 0.217464
R27740 FFCLR.n162 FFCLR 0.217464
R27741 FFCLR.n140 FFCLR 0.217464
R27742 FFCLR.n118 FFCLR 0.217464
R27743 FFCLR.n27 FFCLR 0.217464
R27744 FFCLR.n21 FFCLR 0.217464
R27745 FFCLR.n12 FFCLR 0.217464
R27746 FFCLR.n6 FFCLR 0.217464
R27747 FFCLR.n206 FFCLR 0.200143
R27748 FFCLR.n40 FFCLR.n39 0.159517
R27749 FFCLR.n40 FFCLR 0.129132
R27750 FFCLR.n195 FFCLR 0.1255
R27751 FFCLR.n96 FFCLR 0.1255
R27752 FFCLR.n90 FFCLR 0.1255
R27753 FFCLR.n82 FFCLR 0.1255
R27754 FFCLR.n76 FFCLR 0.1255
R27755 FFCLR.n70 FFCLR 0.1255
R27756 FFCLR.n62 FFCLR 0.1255
R27757 FFCLR.n56 FFCLR 0.1255
R27758 FFCLR.n50 FFCLR 0.1255
R27759 FFCLR.n43 FFCLR 0.1255
R27760 FFCLR.n185 FFCLR 0.1255
R27761 FFCLR.n177 FFCLR 0.1255
R27762 FFCLR.n171 FFCLR 0.1255
R27763 FFCLR.n163 FFCLR 0.1255
R27764 FFCLR.n155 FFCLR 0.1255
R27765 FFCLR.n149 FFCLR 0.1255
R27766 FFCLR.n141 FFCLR 0.1255
R27767 FFCLR.n133 FFCLR 0.1255
R27768 FFCLR.n127 FFCLR 0.1255
R27769 FFCLR.n119 FFCLR 0.1255
R27770 FFCLR.n111 FFCLR 0.1255
R27771 FFCLR.n105 FFCLR 0.1255
R27772 FFCLR.n30 FFCLR 0.1255
R27773 FFCLR.n24 FFCLR 0.1255
R27774 FFCLR.n37 FFCLR 0.1255
R27775 FFCLR.n15 FFCLR 0.1255
R27776 FFCLR.n9 FFCLR 0.1255
R27777 FFCLR.n204 FFCLR 0.1255
R27778 FFCLR.n1 FFCLR 0.1255
R27779 FFCLR.n197 FFCLR.n193 0.063
R27780 FFCLR.n197 FFCLR.n196 0.063
R27781 FFCLR.n98 FFCLR.n94 0.063
R27782 FFCLR.n98 FFCLR.n97 0.063
R27783 FFCLR.n92 FFCLR.n88 0.063
R27784 FFCLR.n92 FFCLR.n91 0.063
R27785 FFCLR.n78 FFCLR.n74 0.063
R27786 FFCLR.n78 FFCLR.n77 0.063
R27787 FFCLR.n72 FFCLR.n68 0.063
R27788 FFCLR.n72 FFCLR.n71 0.063
R27789 FFCLR.n58 FFCLR.n54 0.063
R27790 FFCLR.n58 FFCLR.n57 0.063
R27791 FFCLR.n52 FFCLR.n48 0.063
R27792 FFCLR.n52 FFCLR.n51 0.063
R27793 FFCLR.n179 FFCLR.n175 0.063
R27794 FFCLR.n179 FFCLR.n178 0.063
R27795 FFCLR.n173 FFCLR.n169 0.063
R27796 FFCLR.n173 FFCLR.n172 0.063
R27797 FFCLR.n157 FFCLR.n153 0.063
R27798 FFCLR.n157 FFCLR.n156 0.063
R27799 FFCLR.n151 FFCLR.n147 0.063
R27800 FFCLR.n151 FFCLR.n150 0.063
R27801 FFCLR.n135 FFCLR.n131 0.063
R27802 FFCLR.n135 FFCLR.n134 0.063
R27803 FFCLR.n129 FFCLR.n125 0.063
R27804 FFCLR.n129 FFCLR.n128 0.063
R27805 FFCLR.n113 FFCLR.n109 0.063
R27806 FFCLR.n113 FFCLR.n112 0.063
R27807 FFCLR.n107 FFCLR.n103 0.063
R27808 FFCLR.n107 FFCLR.n106 0.063
R27809 FFCLR.n32 FFCLR.n28 0.063
R27810 FFCLR.n32 FFCLR.n31 0.063
R27811 FFCLR.n26 FFCLR.n22 0.063
R27812 FFCLR.n26 FFCLR.n25 0.063
R27813 FFCLR.n17 FFCLR.n13 0.063
R27814 FFCLR.n17 FFCLR.n16 0.063
R27815 FFCLR.n11 FFCLR.n7 0.063
R27816 FFCLR.n11 FFCLR.n10 0.063
R27817 FFCLR.n19 FFCLR.n18 0.063
R27818 FFCLR.n199 FFCLR.n20 0.063
R27819 FFCLR.n200 FFCLR.n199 0.063
R27820 FFCLR.n202 FFCLR.n5 0.063
R27821 FFCLR.n203 FFCLR.n202 0.063
R27822 FFCLR FFCLR.n204 0.063
R27823 FFCLR.n65 FFCLR.n64 0.024
R27824 FFCLR.n85 FFCLR.n84 0.024
R27825 FFCLR.n115 FFCLR.n101 0.024
R27826 FFCLR.n122 FFCLR.n121 0.024
R27827 FFCLR.n121 FFCLR.n117 0.024
R27828 FFCLR.n137 FFCLR.n123 0.024
R27829 FFCLR.n144 FFCLR.n143 0.024
R27830 FFCLR.n143 FFCLR.n139 0.024
R27831 FFCLR.n159 FFCLR.n145 0.024
R27832 FFCLR.n166 FFCLR.n165 0.024
R27833 FFCLR.n165 FFCLR.n161 0.024
R27834 FFCLR.n181 FFCLR.n167 0.024
R27835 FFCLR.n188 FFCLR.n187 0.024
R27836 FFCLR.n187 FFCLR.n183 0.024
R27837 FFCLR.n41 FFCLR.n35 0.024
R27838 FFCLR.n41 FFCLR.n40 0.024
R27839 FFCLR.n83 FFCLR.n82 0.0216397
R27840 FFCLR.n83 FFCLR 0.0216397
R27841 FFCLR.n63 FFCLR.n62 0.0216397
R27842 FFCLR.n63 FFCLR 0.0216397
R27843 FFCLR.n44 FFCLR.n43 0.0216397
R27844 FFCLR.n44 FFCLR 0.0216397
R27845 FFCLR.n186 FFCLR.n185 0.0216397
R27846 FFCLR.n186 FFCLR 0.0216397
R27847 FFCLR.n164 FFCLR.n163 0.0216397
R27848 FFCLR.n164 FFCLR 0.0216397
R27849 FFCLR.n142 FFCLR.n141 0.0216397
R27850 FFCLR.n142 FFCLR 0.0216397
R27851 FFCLR.n120 FFCLR.n119 0.0216397
R27852 FFCLR.n120 FFCLR 0.0216397
R27853 FFCLR.n30 FFCLR.n29 0.0216397
R27854 FFCLR.n29 FFCLR 0.0216397
R27855 FFCLR.n24 FFCLR.n23 0.0216397
R27856 FFCLR.n23 FFCLR 0.0216397
R27857 FFCLR.n15 FFCLR.n14 0.0216397
R27858 FFCLR.n14 FFCLR 0.0216397
R27859 FFCLR.n9 FFCLR.n8 0.0216397
R27860 FFCLR.n8 FFCLR 0.0216397
R27861 FFCLR.n60 FFCLR 0.0204394
R27862 FFCLR.n80 FFCLR 0.0204394
R27863 FFCLR.n100 FFCLR 0.0204394
R27864 FFCLR FFCLR.n115 0.0204394
R27865 FFCLR FFCLR.n137 0.0204394
R27866 FFCLR FFCLR.n159 0.0204394
R27867 FFCLR FFCLR.n181 0.0204394
R27868 FFCLR.n201 FFCLR 0.0168043
R27869 FFCLR FFCLR.n201 0.0122188
R27870 FFCLR.n195 FFCLR.n194 0.0107679
R27871 FFCLR.n194 FFCLR 0.0107679
R27872 FFCLR.n96 FFCLR.n95 0.0107679
R27873 FFCLR.n95 FFCLR 0.0107679
R27874 FFCLR.n90 FFCLR.n89 0.0107679
R27875 FFCLR.n89 FFCLR 0.0107679
R27876 FFCLR.n76 FFCLR.n75 0.0107679
R27877 FFCLR.n75 FFCLR 0.0107679
R27878 FFCLR.n70 FFCLR.n69 0.0107679
R27879 FFCLR.n69 FFCLR 0.0107679
R27880 FFCLR.n56 FFCLR.n55 0.0107679
R27881 FFCLR.n55 FFCLR 0.0107679
R27882 FFCLR.n50 FFCLR.n49 0.0107679
R27883 FFCLR.n49 FFCLR 0.0107679
R27884 FFCLR.n177 FFCLR.n176 0.0107679
R27885 FFCLR.n176 FFCLR 0.0107679
R27886 FFCLR.n171 FFCLR.n170 0.0107679
R27887 FFCLR.n170 FFCLR 0.0107679
R27888 FFCLR.n155 FFCLR.n154 0.0107679
R27889 FFCLR.n154 FFCLR 0.0107679
R27890 FFCLR.n149 FFCLR.n148 0.0107679
R27891 FFCLR.n148 FFCLR 0.0107679
R27892 FFCLR.n133 FFCLR.n132 0.0107679
R27893 FFCLR.n132 FFCLR 0.0107679
R27894 FFCLR.n127 FFCLR.n126 0.0107679
R27895 FFCLR.n126 FFCLR 0.0107679
R27896 FFCLR.n111 FFCLR.n110 0.0107679
R27897 FFCLR.n110 FFCLR 0.0107679
R27898 FFCLR.n105 FFCLR.n104 0.0107679
R27899 FFCLR.n104 FFCLR 0.0107679
R27900 FFCLR.n37 FFCLR.n36 0.0107679
R27901 FFCLR.n36 FFCLR 0.0107679
R27902 FFCLR.n1 FFCLR.n0 0.0107679
R27903 FFCLR.n0 FFCLR 0.0107679
R27904 FFCLR.n46 FFCLR 0.00441667
R27905 FFCLR.n66 FFCLR 0.00441667
R27906 FFCLR.n86 FFCLR 0.00441667
R27907 FFCLR.n116 FFCLR 0.00441667
R27908 FFCLR.n138 FFCLR 0.00441667
R27909 FFCLR.n160 FFCLR 0.00441667
R27910 FFCLR.n182 FFCLR 0.00441667
R27911 FFCLR.n39 FFCLR 0.00441667
R27912 FFCLR.n3 FFCLR 0.00441667
R27913 FFCLR FFCLR.n46 0.00406061
R27914 FFCLR FFCLR.n66 0.00406061
R27915 FFCLR FFCLR.n86 0.00406061
R27916 FFCLR.n116 FFCLR 0.00406061
R27917 FFCLR.n138 FFCLR 0.00406061
R27918 FFCLR.n160 FFCLR 0.00406061
R27919 FFCLR.n182 FFCLR 0.00406061
R27920 FFCLR.n39 FFCLR 0.00406061
R27921 FFCLR.n3 FFCLR 0.00406061
R27922 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 316.762
R27923 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 168.108
R27924 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 150.293
R27925 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 150.273
R27926 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 73.6406
R27927 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 73.6304
R27928 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 60.3943
R27929 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 12.0358
R27930 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 1.19615
R27931 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.981478
R27932 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 0.788543
R27933 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.769522
R27934 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 0.682565
R27935 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.580578
R27936 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 0.55213
R27937 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 0.484875
R27938 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 0.470609
R27939 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.447191
R27940 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.428234
R27941 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.217464
R27942 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R27943 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R27944 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R27945 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 0.063
R27946 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 0.063
R27947 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.063
R27948 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 0.063
R27949 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 0.063
R27950 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 0.0216397
R27951 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.0216397
R27952 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 0.0107679
R27953 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.0107679
R27954 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 179.256
R27955 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 168.089
R27956 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 150.293
R27957 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 73.6304
R27958 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 60.3943
R27959 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 12.0358
R27960 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.981478
R27961 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 0.788543
R27962 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.769522
R27963 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 0.720633
R27964 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 0.682565
R27965 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.580578
R27966 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 0.55213
R27967 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 0.470609
R27968 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.447191
R27969 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.428234
R27970 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1255
R27971 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1255
R27972 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 0.063
R27973 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 0.063
R27974 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.063
R27975 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 0.063
R27976 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 0.063
R27977 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 0.0435206
R27978 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 0.0107679
R27979 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.0107679
R27980 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 316.762
R27981 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 168.108
R27982 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 150.293
R27983 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 150.273
R27984 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 73.6406
R27985 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 73.6304
R27986 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 60.4568
R27987 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 12.0358
R27988 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 1.19615
R27989 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.981478
R27990 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 0.788543
R27991 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.769522
R27992 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 0.682565
R27993 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.580578
R27994 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 0.55213
R27995 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 0.484875
R27996 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 0.470609
R27997 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.447191
R27998 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.428234
R27999 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.217464
R28000 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R28001 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R28002 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R28003 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 0.063
R28004 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 0.063
R28005 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.063
R28006 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 0.063
R28007 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 0.063
R28008 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 0.0216397
R28009 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.0216397
R28010 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 0.0107679
R28011 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.0107679
R28012 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 179.256
R28013 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 168.089
R28014 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 150.293
R28015 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 73.6304
R28016 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 60.4568
R28017 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 12.0358
R28018 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.981478
R28019 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 0.788543
R28020 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.769522
R28021 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.720633
R28022 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 0.682565
R28023 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.580578
R28024 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 0.55213
R28025 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 0.470609
R28026 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.447191
R28027 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.428234
R28028 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1255
R28029 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1255
R28030 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 0.063
R28031 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 0.063
R28032 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 0.063
R28033 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 0.063
R28034 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 0.063
R28035 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 0.0435206
R28036 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 0.0107679
R28037 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.0107679
R28038 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 169.46
R28039 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 167.809
R28040 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 167.809
R28041 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 167.226
R28042 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 150.273
R28043 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 150.273
R28044 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 73.6406
R28045 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 73.6304
R28046 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 60.3943
R28047 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 12.3891
R28048 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 11.4489
R28049 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 1.68257
R28050 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 1.38365
R28051 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 1.19615
R28052 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 1.1717
R28053 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 1.08448
R28054 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.932141
R28055 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.720633
R28056 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 0.280391
R28057 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.217464
R28058 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R28059 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R28060 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R28061 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 0.0874565
R28062 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 0.063
R28063 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 0.063
R28064 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 0.063
R28065 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 0.063
R28066 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 0.0435206
R28067 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 0.0216397
R28068 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.0216397
R28069 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 0.0107679
R28070 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.0107679
R28071 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 316.762
R28072 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 168.108
R28073 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 150.293
R28074 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 150.273
R28075 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 73.6406
R28076 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 73.6304
R28077 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 60.4568
R28078 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 12.0358
R28079 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 1.19615
R28080 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.981478
R28081 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 0.788543
R28082 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.769522
R28083 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 0.682565
R28084 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.580578
R28085 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 0.55213
R28086 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 0.484875
R28087 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 0.470609
R28088 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.447191
R28089 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.428234
R28090 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.217464
R28091 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R28092 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R28093 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R28094 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 0.063
R28095 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 0.063
R28096 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.063
R28097 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 0.063
R28098 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 0.063
R28099 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 0.0216397
R28100 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.0216397
R28101 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 0.0107679
R28102 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.0107679
R28103 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 169.46
R28104 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 168.089
R28105 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 167.809
R28106 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 150.293
R28107 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 73.6304
R28108 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 60.4568
R28109 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 12.0358
R28110 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 11.4489
R28111 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.981478
R28112 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 0.788543
R28113 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.769522
R28114 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 0.720633
R28115 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 0.682565
R28116 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.580578
R28117 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 0.55213
R28118 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 0.470609
R28119 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.447191
R28120 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.428234
R28121 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.1255
R28122 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.1255
R28123 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 0.063
R28124 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 0.063
R28125 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.063
R28126 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 0.063
R28127 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 0.063
R28128 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 0.0435206
R28129 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 0.0107679
R28130 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.0107679
R28131 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 169.46
R28132 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 167.809
R28133 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 167.809
R28134 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 167.226
R28135 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 150.273
R28136 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 150.273
R28137 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 73.6406
R28138 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 73.6304
R28139 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 60.3943
R28140 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 12.3891
R28141 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 11.4489
R28142 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 1.68257
R28143 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 1.38365
R28144 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 1.19615
R28145 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 1.1717
R28146 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 1.08448
R28147 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.932141
R28148 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 0.720633
R28149 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 0.280391
R28150 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.217464
R28151 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R28152 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R28153 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R28154 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 0.0874565
R28155 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 0.063
R28156 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.063
R28157 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 0.063
R28158 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 0.063
R28159 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 0.0435206
R28160 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 0.0216397
R28161 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.0216397
R28162 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 0.0107679
R28163 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.0107679
R28164 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 169.46
R28165 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 167.809
R28166 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 167.809
R28167 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 167.227
R28168 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 150.293
R28169 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 150.273
R28170 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 73.6406
R28171 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 73.6304
R28172 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 60.3809
R28173 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 12.3891
R28174 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 11.4489
R28175 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 1.38365
R28176 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 1.19615
R28177 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 1.1717
R28178 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.848156
R28179 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 0.447191
R28180 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R28181 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 0.280391
R28182 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.217464
R28183 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.200143
R28184 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R28185 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R28186 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R28187 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R28188 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 0.0874565
R28189 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 0.063
R28190 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 0.063
R28191 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 0.063
R28192 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R28193 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 0.0107679
R28194 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0107679
R28195 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 169.46
R28196 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 167.809
R28197 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 167.809
R28198 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 167.226
R28199 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 150.273
R28200 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 150.273
R28201 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 73.6406
R28202 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 73.6304
R28203 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 60.3943
R28204 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 12.3891
R28205 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 11.4489
R28206 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 1.68257
R28207 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 1.38365
R28208 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 1.19615
R28209 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 1.1717
R28210 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 1.08448
R28211 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.932141
R28212 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 0.720633
R28213 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 0.280391
R28214 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.217464
R28215 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R28216 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R28217 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R28218 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 0.0874565
R28219 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 0.063
R28220 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.063
R28221 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 0.063
R28222 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 0.063
R28223 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 0.0435206
R28224 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 0.0216397
R28225 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.0216397
R28226 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 0.0107679
R28227 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.0107679
R28228 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 169.46
R28229 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 167.809
R28230 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 167.809
R28231 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 167.226
R28232 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 150.273
R28233 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 150.273
R28234 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 73.6406
R28235 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 73.6304
R28236 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 60.3943
R28237 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 12.3891
R28238 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 11.4489
R28239 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 1.68257
R28240 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 1.38365
R28241 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 1.19615
R28242 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 1.1717
R28243 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 1.08448
R28244 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.932141
R28245 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.720633
R28246 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 0.280391
R28247 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.217464
R28248 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R28249 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R28250 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R28251 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 0.0874565
R28252 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 0.063
R28253 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.063
R28254 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 0.063
R28255 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 0.063
R28256 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 0.0435206
R28257 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 0.0216397
R28258 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 0.0216397
R28259 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 0.0107679
R28260 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.0107679
R28261 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 169.46
R28262 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 167.809
R28263 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 167.809
R28264 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 167.227
R28265 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 150.293
R28266 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 150.273
R28267 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 73.6406
R28268 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 73.6304
R28269 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 60.3809
R28270 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 12.3891
R28271 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 11.4489
R28272 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 1.38365
R28273 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 1.19615
R28274 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 1.1717
R28275 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 0.848156
R28276 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.447191
R28277 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R28278 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 0.280391
R28279 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.217464
R28280 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 0.200143
R28281 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R28282 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R28283 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R28284 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R28285 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 0.0874565
R28286 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.063
R28287 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 0.063
R28288 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 0.063
R28289 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R28290 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 0.0107679
R28291 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0107679
R28292 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 169.46
R28293 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 167.809
R28294 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 167.809
R28295 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 167.226
R28296 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 150.273
R28297 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 150.273
R28298 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 73.6406
R28299 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 73.6304
R28300 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 60.4568
R28301 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 12.3891
R28302 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 11.4489
R28303 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.68257
R28304 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 1.38365
R28305 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 1.19615
R28306 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 1.1717
R28307 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.08448
R28308 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.932141
R28309 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.720633
R28310 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 0.280391
R28311 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.217464
R28312 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R28313 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R28314 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R28315 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 0.0874565
R28316 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 0.063
R28317 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 0.063
R28318 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 0.063
R28319 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 0.063
R28320 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 0.0435206
R28321 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 0.0216397
R28322 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.0216397
R28323 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 0.0107679
R28324 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.0107679
R28325 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 169.46
R28326 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 167.809
R28327 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 167.809
R28328 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 167.227
R28329 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 150.293
R28330 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 150.273
R28331 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 73.6406
R28332 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 73.6304
R28333 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 60.3809
R28334 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 12.3891
R28335 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 11.4489
R28336 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 1.38365
R28337 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 1.19615
R28338 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 1.1717
R28339 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.848156
R28340 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 0.447191
R28341 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.38637
R28342 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 0.280391
R28343 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 0.262643
R28344 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.217464
R28345 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.152844
R28346 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.149957
R28347 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.1255
R28348 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.1255
R28349 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 0.0874565
R28350 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 0.063
R28351 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 0.063
R28352 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.063
R28353 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.0454219
R28354 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 0.0107679
R28355 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.0107679
R28356 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t1 169.46
R28357 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.t3 167.809
R28358 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t0 167.809
R28359 D_FlipFlop_0.3-input-nand_2.Vout.t4 D_FlipFlop_0.3-input-nand_2.Vout.n11 167.227
R28360 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.t4 150.293
R28361 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.t7 150.273
R28362 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout.t5 73.6406
R28363 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout.t6 73.6304
R28364 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout.t2 60.3809
R28365 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n5 12.3891
R28366 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout.n9 11.4489
R28367 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout.n2 1.38365
R28368 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.n1 1.19615
R28369 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.n4 1.1717
R28370 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout 0.848156
R28371 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.Vout.n12 0.447191
R28372 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout 0.38637
R28373 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.n10 0.280391
R28374 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout.n8 0.262643
R28375 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout 0.217464
R28376 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout 0.152844
R28377 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.149957
R28378 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R28379 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R28380 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout.n7 0.0874565
R28381 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n3 0.063
R28382 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout.n6 0.063
R28383 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout 0.063
R28384 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.0454219
R28385 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout.n0 0.0107679
R28386 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout 0.0107679
R28387 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 169.46
R28388 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 167.809
R28389 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 167.809
R28390 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 167.227
R28391 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 150.293
R28392 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 150.273
R28393 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 73.6406
R28394 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 73.6304
R28395 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 60.3809
R28396 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 12.3891
R28397 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 11.4489
R28398 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 1.38365
R28399 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 1.19615
R28400 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 1.1717
R28401 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.848156
R28402 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 0.447191
R28403 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.38637
R28404 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 0.280391
R28405 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 0.262643
R28406 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.217464
R28407 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.152844
R28408 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.149957
R28409 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.1255
R28410 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.1255
R28411 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 0.0874565
R28412 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 0.063
R28413 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 0.063
R28414 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.063
R28415 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.0454219
R28416 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 0.0107679
R28417 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.0107679
R28418 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 169.46
R28419 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 167.809
R28420 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 167.809
R28421 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 167.226
R28422 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 150.273
R28423 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 150.273
R28424 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 73.6406
R28425 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 73.6304
R28426 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 60.4568
R28427 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 12.3891
R28428 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 11.4489
R28429 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.68257
R28430 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 1.38365
R28431 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 1.19615
R28432 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 1.1717
R28433 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.08448
R28434 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.932141
R28435 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 0.720633
R28436 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 0.280391
R28437 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.217464
R28438 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R28439 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R28440 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R28441 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 0.0874565
R28442 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 0.063
R28443 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.063
R28444 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 0.063
R28445 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 0.063
R28446 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 0.0435206
R28447 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 0.0216397
R28448 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.0216397
R28449 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 0.0107679
R28450 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.0107679
R28451 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 169.46
R28452 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 167.809
R28453 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 167.809
R28454 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 167.227
R28455 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 150.293
R28456 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 150.273
R28457 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 73.6406
R28458 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 73.6304
R28459 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 60.3809
R28460 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 12.3891
R28461 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 11.4489
R28462 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 1.38365
R28463 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 1.19615
R28464 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 1.1717
R28465 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 0.848156
R28466 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.447191
R28467 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.38637
R28468 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 0.280391
R28469 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 0.262643
R28470 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.217464
R28471 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.152844
R28472 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.149957
R28473 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.1255
R28474 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.1255
R28475 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 0.0874565
R28476 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.063
R28477 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 0.063
R28478 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 0.063
R28479 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.0454219
R28480 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 0.0107679
R28481 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.0107679
R28482 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 169.46
R28483 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 167.809
R28484 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 167.809
R28485 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 167.226
R28486 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 150.273
R28487 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 150.273
R28488 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 73.6406
R28489 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 73.6304
R28490 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 60.4568
R28491 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 12.3891
R28492 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 11.4489
R28493 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.68257
R28494 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 1.38365
R28495 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 1.19615
R28496 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 1.1717
R28497 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.08448
R28498 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.932141
R28499 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.720633
R28500 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 0.280391
R28501 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.217464
R28502 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R28503 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R28504 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R28505 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 0.0874565
R28506 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 0.063
R28507 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.063
R28508 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 0.063
R28509 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 0.063
R28510 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 0.0435206
R28511 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 0.0216397
R28512 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 0.0216397
R28513 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 0.0107679
R28514 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.0107679
R28515 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 316.762
R28516 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 168.108
R28517 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 150.293
R28518 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 150.273
R28519 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 73.6406
R28520 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 73.6304
R28521 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 60.3943
R28522 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 12.0358
R28523 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 1.19615
R28524 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.981478
R28525 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 0.788543
R28526 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.769522
R28527 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 0.682565
R28528 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.580578
R28529 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 0.55213
R28530 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 0.484875
R28531 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 0.470609
R28532 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.447191
R28533 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.428234
R28534 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.217464
R28535 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R28536 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R28537 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R28538 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 0.063
R28539 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 0.063
R28540 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.063
R28541 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 0.063
R28542 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 0.063
R28543 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 0.0216397
R28544 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.0216397
R28545 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 0.0107679
R28546 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.0107679
R28547 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 169.46
R28548 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 167.809
R28549 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 167.809
R28550 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 167.227
R28551 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 150.293
R28552 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 150.273
R28553 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 73.6406
R28554 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 73.6304
R28555 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 60.3809
R28556 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 12.3891
R28557 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 11.4489
R28558 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 1.38365
R28559 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 1.19615
R28560 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 1.1717
R28561 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 0.848156
R28562 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.447191
R28563 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R28564 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 0.280391
R28565 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.217464
R28566 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 0.200143
R28567 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R28568 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R28569 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R28570 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R28571 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 0.0874565
R28572 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.063
R28573 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 0.063
R28574 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 0.063
R28575 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R28576 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 0.0107679
R28577 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0107679
R28578 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C.t1 169.46
R28579 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C.t3 167.809
R28580 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C.t2 167.809
R28581 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C.t6 167.226
R28582 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.t7 150.273
R28583 D_FlipFlop_5.3-input-nand_2.C.t6 D_FlipFlop_5.3-input-nand_2.C.n2 150.273
R28584 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C.t5 73.6406
R28585 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C.t4 73.6304
R28586 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.t0 60.4568
R28587 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n11 12.3891
R28588 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C.n4 11.4489
R28589 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C 1.68257
R28590 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.n13 1.38365
R28591 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C.n0 1.19615
R28592 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C.n9 1.1717
R28593 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C 1.08448
R28594 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C 0.932141
R28595 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C 0.720633
R28596 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C.n3 0.280391
R28597 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C 0.217464
R28598 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C 0.1255
R28599 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C 0.1255
R28600 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C 0.1255
R28601 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C.n6 0.0874565
R28602 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.n10 0.063
R28603 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n7 0.063
R28604 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C.n12 0.063
R28605 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.C.n14 0.063
R28606 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C.n5 0.0435206
R28607 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C.n1 0.0216397
R28608 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C 0.0216397
R28609 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C.n8 0.0107679
R28610 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C 0.0107679
R28611 Q6.n2 Q6.t0 169.46
R28612 Q6.n4 Q6.t2 167.809
R28613 Q6.n2 Q6.t1 167.809
R28614 Q6 Q6.t6 158.585
R28615 Q6 Q6.t7 154.823
R28616 Q6.n14 Q6.t9 150.869
R28617 Q6.t7 Q6.n15 150.869
R28618 Q6.t6 Q6.n9 150.293
R28619 Q6.n16 Q6.n13 137.644
R28620 Q6.n13 Q6 85.5731
R28621 Q6.n15 Q6.t4 74.1352
R28622 Q6.n14 Q6.t5 74.1352
R28623 Q6.n7 Q6.t8 73.6304
R28624 Q6.n0 Q6.t3 60.3809
R28625 Q6.n3 Q6.n2 11.4489
R28626 Q6.n5 Q6.n4 8.21389
R28627 Q6.n13 Q6.n12 3.473
R28628 Q6.n15 Q6.n14 1.66898
R28629 Q6.n1 Q6.n0 1.64452
R28630 Q6.n9 Q6.n8 1.19615
R28631 Q6.n0 Q6 0.848156
R28632 Q6.n9 Q6 0.447191
R28633 Q6.n5 Q6 0.39003
R28634 Q6.n4 Q6.n3 0.280391
R28635 Q6.n3 Q6.n1 0.262643
R28636 Q6.n6 Q6 0.2167
R28637 Q6.n6 Q6.n5 0.212783
R28638 Q6.n11 Q6.n10 0.161083
R28639 Q6.n11 Q6 0.150045
R28640 Q6.n1 Q6 0.1255
R28641 Q6.n8 Q6 0.1255
R28642 Q6.n14 Q6 0.063
R28643 Q6.n1 Q6 0.063
R28644 Q6.n12 Q6.n6 0.024
R28645 Q6.n12 Q6.n11 0.024
R28646 Q6 Q6.n16 0.0168043
R28647 Q6.n16 Q6 0.0122188
R28648 Q6.n8 Q6.n7 0.0107679
R28649 Q6.n7 Q6 0.0107679
R28650 Q6.n10 Q6 0.00441667
R28651 Q6.n10 Q6 0.00406061
R28652 CDAC8_0.switch_2.Z.n5 CDAC8_0.switch_2.Z.t3 168.548
R28653 CDAC8_0.switch_2.Z.n5 CDAC8_0.switch_2.Z.t0 168.548
R28654 CDAC8_0.switch_2.Z.n0 CDAC8_0.switch_2.Z.t1 60.321
R28655 CDAC8_0.switch_2.Z.n0 CDAC8_0.switch_2.Z.t2 60.321
R28656 CDAC8_0.switch_2.Z.n4 CDAC8_0.switch_2.Z.n3 11.3205
R28657 CDAC8_0.switch_2.Z.n3 CDAC8_0.switch_2.Z.t5 3.64361
R28658 CDAC8_0.switch_2.Z.n3 CDAC8_0.switch_2.Z.t4 3.16265
R28659 CDAC8_0.switch_2.Z.n2 CDAC8_0.switch_2.Z.n1 1.59289
R28660 CDAC8_0.switch_2.Z.n1 CDAC8_0.switch_2.Z 0.259656
R28661 CDAC8_0.switch_2.Z.n2 CDAC8_0.switch_2.Z 0.17713
R28662 CDAC8_0.switch_2.Z.n4 CDAC8_0.switch_2.Z.n2 0.063
R28663 CDAC8_0.switch_2.Z CDAC8_0.switch_2.Z.n5 0.0454219
R28664 CDAC8_0.switch_2.Z.n5 CDAC8_0.switch_2.Z.n4 0.0200312
R28665 CDAC8_0.switch_2.Z.n1 CDAC8_0.switch_2.Z.n0 0.0188121
R28666 Q3.n5 Q3.t1 169.46
R28667 Q3.n7 Q3.t3 167.809
R28668 Q3.n5 Q3.t0 167.809
R28669 Q3.n11 Q3.t5 155.12
R28670 Q3.n14 Q3.t6 150.869
R28671 Q3.n13 Q3.t7 150.869
R28672 Q3.t5 Q3.n2 150.293
R28673 Q3.n15 Q3.n12 137.644
R28674 Q3 Q3.t9 78.1811
R28675 Q3.n13 Q3.t4 74.1352
R28676 Q3.t9 Q3.n14 74.1352
R28677 Q3.n0 Q3.t8 73.6304
R28678 Q3.n3 Q3.t2 60.3809
R28679 Q3.n12 Q3 36.8166
R28680 Q3.n6 Q3.n5 11.4489
R28681 Q3.n8 Q3.n7 8.21389
R28682 Q3.n11 Q3.n10 1.6986
R28683 Q3.n14 Q3.n13 1.66898
R28684 Q3.n4 Q3.n3 1.64452
R28685 Q3.n2 Q3.n1 1.19615
R28686 Q3.n3 Q3 0.848156
R28687 Q3.n2 Q3 0.447191
R28688 Q3.n8 Q3 0.39003
R28689 Q3.n9 Q3.n8 0.3483
R28690 Q3.n7 Q3.n6 0.280391
R28691 Q3.n6 Q3.n4 0.262643
R28692 Q3.n4 Q3 0.1255
R28693 Q3.n1 Q3 0.1255
R28694 Q3.n9 Q3 0.0811833
R28695 Q3.n13 Q3 0.063
R28696 Q3.n4 Q3 0.063
R28697 Q3.n10 Q3.n9 0.0491718
R28698 Q3.n12 Q3.n11 0.0273895
R28699 Q3.n10 Q3 0.025816
R28700 Q3 Q3.n15 0.0168043
R28701 Q3.n15 Q3 0.0122188
R28702 Q3.n1 Q3.n0 0.0107679
R28703 Q3.n0 Q3 0.0107679
R28704 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.t3 168.609
R28705 CDAC8_0.switch_5.Z CDAC8_0.switch_5.Z.t0 168.565
R28706 CDAC8_0.switch_5.Z.n0 CDAC8_0.switch_5.Z.t1 60.321
R28707 CDAC8_0.switch_5.Z.n0 CDAC8_0.switch_5.Z.t2 60.321
R28708 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.n10 11.3205
R28709 CDAC8_0.switch_5.Z.n6 CDAC8_0.switch_5.Z.n5 5.49497
R28710 CDAC8_0.switch_5.Z.n10 CDAC8_0.switch_5.Z.n2 2.98587
R28711 CDAC8_0.switch_5.Z.n10 CDAC8_0.switch_5.Z.n9 2.5049
R28712 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.n1 1.60376
R28713 CDAC8_0.switch_5.Z.n9 CDAC8_0.switch_5.Z.t10 0.726216
R28714 CDAC8_0.switch_5.Z.n2 CDAC8_0.switch_5.Z.t6 0.726216
R28715 CDAC8_0.switch_5.Z.n5 CDAC8_0.switch_5.Z.t9 0.658247
R28716 CDAC8_0.switch_5.Z.n6 CDAC8_0.switch_5.Z.t5 0.658247
R28717 CDAC8_0.switch_5.Z.n7 CDAC8_0.switch_5.Z.t8 0.611304
R28718 CDAC8_0.switch_5.Z.n8 CDAC8_0.switch_5.Z.t11 0.611304
R28719 CDAC8_0.switch_5.Z.n4 CDAC8_0.switch_5.Z.t4 0.611304
R28720 CDAC8_0.switch_5.Z.n3 CDAC8_0.switch_5.Z.t7 0.611304
R28721 CDAC8_0.switch_5.Z.n1 CDAC8_0.switch_5.Z 0.259656
R28722 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z 0.166261
R28723 CDAC8_0.switch_5.Z.n8 CDAC8_0.switch_5.Z.n7 0.162356
R28724 CDAC8_0.switch_5.Z.n4 CDAC8_0.switch_5.Z.n3 0.162356
R28725 CDAC8_0.switch_5.Z.n7 CDAC8_0.switch_5.Z.n6 0.115412
R28726 CDAC8_0.switch_5.Z.n5 CDAC8_0.switch_5.Z.n4 0.115412
R28727 CDAC8_0.switch_5.Z.n9 CDAC8_0.switch_5.Z.n8 0.0474438
R28728 CDAC8_0.switch_5.Z.n3 CDAC8_0.switch_5.Z.n2 0.0474438
R28729 CDAC8_0.switch_5.Z CDAC8_0.switch_5.Z.n11 0.0454219
R28730 CDAC8_0.switch_5.Z.n1 CDAC8_0.switch_5.Z.n0 0.0188121
R28731 Nand_Gate_5.Vout.n10 Nand_Gate_5.Vout.t0 179.256
R28732 Nand_Gate_5.Vout.n10 Nand_Gate_5.Vout.t2 168.089
R28733 Nand_Gate_5.Vout.n2 Nand_Gate_5.Vout.t3 150.293
R28734 Nand_Gate_5.Vout.n4 Nand_Gate_5.Vout.t4 73.6304
R28735 Nand_Gate_5.Vout Nand_Gate_5.Vout.t1 60.3943
R28736 Nand_Gate_5.Vout.n8 Nand_Gate_5.Vout.n7 35.6663
R28737 Nand_Gate_5.Vout.n9 Nand_Gate_5.Vout 0.981478
R28738 Nand_Gate_5.Vout.n11 Nand_Gate_5.Vout.n9 0.788543
R28739 Nand_Gate_5.Vout.n3 Nand_Gate_5.Vout 0.769522
R28740 Nand_Gate_5.Vout Nand_Gate_5.Vout.n11 0.720633
R28741 Nand_Gate_5.Vout.n1 Nand_Gate_5.Vout.n0 0.682565
R28742 Nand_Gate_5.Vout.n1 Nand_Gate_5.Vout 0.580578
R28743 Nand_Gate_5.Vout.n3 Nand_Gate_5.Vout.n2 0.55213
R28744 Nand_Gate_5.Vout.n6 Nand_Gate_5.Vout.n5 0.470609
R28745 Nand_Gate_5.Vout.n2 Nand_Gate_5.Vout 0.447191
R28746 Nand_Gate_5.Vout.n6 Nand_Gate_5.Vout 0.428234
R28747 Nand_Gate_5.Vout.n5 Nand_Gate_5.Vout 0.1255
R28748 Nand_Gate_5.Vout.n0 Nand_Gate_5.Vout 0.1255
R28749 Nand_Gate_5.Vout.n7 Nand_Gate_5.Vout.n3 0.063
R28750 Nand_Gate_5.Vout.n7 Nand_Gate_5.Vout.n6 0.063
R28751 Nand_Gate_5.Vout.n0 Nand_Gate_5.Vout 0.063
R28752 Nand_Gate_5.Vout.n9 Nand_Gate_5.Vout.n8 0.063
R28753 Nand_Gate_5.Vout.n8 Nand_Gate_5.Vout.n1 0.063
R28754 Nand_Gate_5.Vout.n11 Nand_Gate_5.Vout.n10 0.0435206
R28755 Nand_Gate_5.Vout.n5 Nand_Gate_5.Vout.n4 0.0107679
R28756 Nand_Gate_5.Vout.n4 Nand_Gate_5.Vout 0.0107679
R28757 Nand_Gate_6.B.n51 Nand_Gate_6.B.t0 169.46
R28758 Nand_Gate_6.B.n51 Nand_Gate_6.B.t1 167.809
R28759 Nand_Gate_6.B.n53 Nand_Gate_6.B.t3 167.809
R28760 Nand_Gate_6.B Nand_Gate_6.B.t5 158.585
R28761 Nand_Gate_6.B Nand_Gate_6.B.t9 158.581
R28762 Nand_Gate_6.B.n42 Nand_Gate_6.B.t8 150.293
R28763 Nand_Gate_6.B.t9 Nand_Gate_6.B.n38 150.293
R28764 Nand_Gate_6.B.t5 Nand_Gate_6.B.n2 150.293
R28765 Nand_Gate_6.B.n29 Nand_Gate_6.B.t7 150.273
R28766 Nand_Gate_6.B.n23 Nand_Gate_6.B.t12 150.273
R28767 Nand_Gate_6.B.n14 Nand_Gate_6.B.t11 150.273
R28768 Nand_Gate_6.B.n8 Nand_Gate_6.B.t17 150.273
R28769 Nand_Gate_6.B.n27 Nand_Gate_6.B.t13 73.6406
R28770 Nand_Gate_6.B.n21 Nand_Gate_6.B.t6 73.6406
R28771 Nand_Gate_6.B.n12 Nand_Gate_6.B.t15 73.6406
R28772 Nand_Gate_6.B.n6 Nand_Gate_6.B.t10 73.6406
R28773 Nand_Gate_6.B.n43 Nand_Gate_6.B.t14 73.6304
R28774 Nand_Gate_6.B.n36 Nand_Gate_6.B.t4 73.6304
R28775 Nand_Gate_6.B.n0 Nand_Gate_6.B.t16 73.6304
R28776 Nand_Gate_6.B.n4 Nand_Gate_6.B.t2 60.3809
R28777 Nand_Gate_6.B.n44 Nand_Gate_6.B.n41 47.1622
R28778 Nand_Gate_6.B.n44 Nand_Gate_6.B.n43 34.7148
R28779 Nand_Gate_6.B.n33 Nand_Gate_6.B.n26 15.5222
R28780 Nand_Gate_6.B.n52 Nand_Gate_6.B.n51 11.4489
R28781 Nand_Gate_6.B.n34 Nand_Gate_6.B.n33 8.26552
R28782 Nand_Gate_6.B.n54 Nand_Gate_6.B.n53 8.21389
R28783 Nand_Gate_6.B.n18 Nand_Gate_6.B.n11 8.1418
R28784 Nand_Gate_6.B.n47 Nand_Gate_6.B.n46 5.61191
R28785 Nand_Gate_6.B.n47 Nand_Gate_6.B 5.35402
R28786 Nand_Gate_6.B.n45 Nand_Gate_6.B.n44 4.81893
R28787 Nand_Gate_6.B.n48 Nand_Gate_6.B.n47 4.563
R28788 Nand_Gate_6.B.n33 Nand_Gate_6.B.n32 4.5005
R28789 Nand_Gate_6.B.n18 Nand_Gate_6.B.n17 4.5005
R28790 Nand_Gate_6.B.n46 Nand_Gate_6.B 1.83746
R28791 Nand_Gate_6.B.n20 Nand_Gate_6.B.n19 1.62007
R28792 Nand_Gate_6.B.n38 Nand_Gate_6.B.n37 1.19615
R28793 Nand_Gate_6.B.n2 Nand_Gate_6.B.n1 1.19615
R28794 Nand_Gate_6.B.n43 Nand_Gate_6.B.n42 1.1717
R28795 Nand_Gate_6.B.n5 Nand_Gate_6.B 1.08746
R28796 Nand_Gate_6.B.n20 Nand_Gate_6.B 1.01739
R28797 Nand_Gate_6.B.n13 Nand_Gate_6.B 0.851043
R28798 Nand_Gate_6.B.n7 Nand_Gate_6.B 0.851043
R28799 Nand_Gate_6.B.n4 Nand_Gate_6.B 0.848156
R28800 Nand_Gate_6.B.n28 Nand_Gate_6.B.n27 0.796696
R28801 Nand_Gate_6.B.n22 Nand_Gate_6.B.n21 0.796696
R28802 Nand_Gate_6.B.n50 Nand_Gate_6.B.n49 0.788543
R28803 Nand_Gate_6.B.n34 Nand_Gate_6.B 0.716182
R28804 Nand_Gate_6.B.n5 Nand_Gate_6.B.n4 0.682565
R28805 Nand_Gate_6.B.n49 Nand_Gate_6.B 0.65675
R28806 Nand_Gate_6.B.n16 Nand_Gate_6.B.n15 0.55213
R28807 Nand_Gate_6.B.n10 Nand_Gate_6.B.n9 0.55213
R28808 Nand_Gate_6.B.n28 Nand_Gate_6.B 0.524957
R28809 Nand_Gate_6.B.n22 Nand_Gate_6.B 0.524957
R28810 Nand_Gate_6.B.n16 Nand_Gate_6.B 0.486828
R28811 Nand_Gate_6.B.n10 Nand_Gate_6.B 0.486828
R28812 Nand_Gate_6.B.n35 Nand_Gate_6.B 0.4846
R28813 Nand_Gate_6.B.n13 Nand_Gate_6.B.n12 0.470609
R28814 Nand_Gate_6.B.n7 Nand_Gate_6.B.n6 0.470609
R28815 Nand_Gate_6.B.n42 Nand_Gate_6.B 0.447191
R28816 Nand_Gate_6.B.n38 Nand_Gate_6.B 0.447191
R28817 Nand_Gate_6.B.n2 Nand_Gate_6.B 0.447191
R28818 Nand_Gate_6.B.n54 Nand_Gate_6.B.n3 0.425067
R28819 Nand_Gate_6.B.n40 Nand_Gate_6.B.n39 0.42115
R28820 Nand_Gate_6.B Nand_Gate_6.B.n54 0.39003
R28821 Nand_Gate_6.B.n40 Nand_Gate_6.B 0.335684
R28822 Nand_Gate_6.B.n35 Nand_Gate_6.B.n34 0.30365
R28823 Nand_Gate_6.B.n53 Nand_Gate_6.B.n52 0.280391
R28824 Nand_Gate_6.B.n52 Nand_Gate_6.B.n50 0.262643
R28825 Nand_Gate_6.B.n31 Nand_Gate_6.B 0.252453
R28826 Nand_Gate_6.B.n25 Nand_Gate_6.B 0.252453
R28827 Nand_Gate_6.B.n31 Nand_Gate_6.B.n30 0.226043
R28828 Nand_Gate_6.B.n25 Nand_Gate_6.B.n24 0.226043
R28829 Nand_Gate_6.B.n27 Nand_Gate_6.B 0.217464
R28830 Nand_Gate_6.B.n21 Nand_Gate_6.B 0.217464
R28831 Nand_Gate_6.B.n12 Nand_Gate_6.B 0.217464
R28832 Nand_Gate_6.B.n6 Nand_Gate_6.B 0.217464
R28833 Nand_Gate_6.B.n43 Nand_Gate_6.B 0.149957
R28834 Nand_Gate_6.B.n30 Nand_Gate_6.B 0.1255
R28835 Nand_Gate_6.B.n24 Nand_Gate_6.B 0.1255
R28836 Nand_Gate_6.B.n37 Nand_Gate_6.B 0.1255
R28837 Nand_Gate_6.B.n15 Nand_Gate_6.B 0.1255
R28838 Nand_Gate_6.B.n9 Nand_Gate_6.B 0.1255
R28839 Nand_Gate_6.B.n50 Nand_Gate_6.B 0.1255
R28840 Nand_Gate_6.B.n1 Nand_Gate_6.B 0.1255
R28841 Nand_Gate_6.B.n32 Nand_Gate_6.B.n28 0.063
R28842 Nand_Gate_6.B.n32 Nand_Gate_6.B.n31 0.063
R28843 Nand_Gate_6.B.n26 Nand_Gate_6.B.n22 0.063
R28844 Nand_Gate_6.B.n26 Nand_Gate_6.B.n25 0.063
R28845 Nand_Gate_6.B.n17 Nand_Gate_6.B.n13 0.063
R28846 Nand_Gate_6.B.n17 Nand_Gate_6.B.n16 0.063
R28847 Nand_Gate_6.B.n11 Nand_Gate_6.B.n7 0.063
R28848 Nand_Gate_6.B.n11 Nand_Gate_6.B.n10 0.063
R28849 Nand_Gate_6.B.n46 Nand_Gate_6.B.n45 0.063
R28850 Nand_Gate_6.B.n45 Nand_Gate_6.B.n20 0.063
R28851 Nand_Gate_6.B.n48 Nand_Gate_6.B.n5 0.063
R28852 Nand_Gate_6.B.n49 Nand_Gate_6.B.n48 0.063
R28853 Nand_Gate_6.B.n50 Nand_Gate_6.B 0.063
R28854 Nand_Gate_6.B Nand_Gate_6.B.n18 0.0512812
R28855 Nand_Gate_6.B.n43 Nand_Gate_6.B 0.0454219
R28856 Nand_Gate_6.B.n41 Nand_Gate_6.B.n35 0.024
R28857 Nand_Gate_6.B.n41 Nand_Gate_6.B.n40 0.024
R28858 Nand_Gate_6.B.n30 Nand_Gate_6.B.n29 0.0216397
R28859 Nand_Gate_6.B.n29 Nand_Gate_6.B 0.0216397
R28860 Nand_Gate_6.B.n24 Nand_Gate_6.B.n23 0.0216397
R28861 Nand_Gate_6.B.n23 Nand_Gate_6.B 0.0216397
R28862 Nand_Gate_6.B.n15 Nand_Gate_6.B.n14 0.0216397
R28863 Nand_Gate_6.B.n14 Nand_Gate_6.B 0.0216397
R28864 Nand_Gate_6.B.n9 Nand_Gate_6.B.n8 0.0216397
R28865 Nand_Gate_6.B.n8 Nand_Gate_6.B 0.0216397
R28866 Nand_Gate_6.B.n19 Nand_Gate_6.B 0.0168043
R28867 Nand_Gate_6.B.n19 Nand_Gate_6.B 0.0122188
R28868 Nand_Gate_6.B.n37 Nand_Gate_6.B.n36 0.0107679
R28869 Nand_Gate_6.B.n36 Nand_Gate_6.B 0.0107679
R28870 Nand_Gate_6.B.n1 Nand_Gate_6.B.n0 0.0107679
R28871 Nand_Gate_6.B.n0 Nand_Gate_6.B 0.0107679
R28872 Nand_Gate_6.B.n39 Nand_Gate_6.B 0.00441667
R28873 Nand_Gate_6.B.n3 Nand_Gate_6.B 0.00441667
R28874 Nand_Gate_6.B.n39 Nand_Gate_6.B 0.00406061
R28875 Nand_Gate_6.B.n3 Nand_Gate_6.B 0.00406061
R28876 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 169.46
R28877 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 168.089
R28878 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 167.809
R28879 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 150.273
R28880 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 73.6406
R28881 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 60.3809
R28882 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 12.0358
R28883 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 11.4489
R28884 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 1.08746
R28885 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.851043
R28886 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.848156
R28887 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 0.788543
R28888 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 0.682565
R28889 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.65675
R28890 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 0.55213
R28891 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.486828
R28892 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 0.470609
R28893 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 0.262643
R28894 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.217464
R28895 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.1255
R28896 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.1255
R28897 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 0.063
R28898 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 0.063
R28899 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 0.063
R28900 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 0.063
R28901 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 0.063
R28902 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 0.0216397
R28903 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0216397
R28904 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 179.256
R28905 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 168.089
R28906 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 150.293
R28907 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 73.6304
R28908 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 60.3943
R28909 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 12.0358
R28910 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.981478
R28911 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 0.788543
R28912 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.769522
R28913 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 0.720633
R28914 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 0.682565
R28915 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.580578
R28916 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 0.55213
R28917 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 0.470609
R28918 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.447191
R28919 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.428234
R28920 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1255
R28921 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1255
R28922 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 0.063
R28923 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 0.063
R28924 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.063
R28925 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 0.063
R28926 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 0.063
R28927 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 0.0435206
R28928 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 0.0107679
R28929 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.0107679
R28930 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 316.762
R28931 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 168.108
R28932 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 150.293
R28933 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 150.273
R28934 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 73.6406
R28935 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 73.6304
R28936 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 60.3943
R28937 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 12.0358
R28938 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 1.19615
R28939 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.981478
R28940 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 0.788543
R28941 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.769522
R28942 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 0.682565
R28943 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.580578
R28944 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 0.55213
R28945 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 0.484875
R28946 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 0.470609
R28947 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.447191
R28948 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.428234
R28949 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.217464
R28950 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R28951 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R28952 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R28953 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 0.063
R28954 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 0.063
R28955 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.063
R28956 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 0.063
R28957 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 0.063
R28958 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 0.0216397
R28959 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.0216397
R28960 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 0.0107679
R28961 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.0107679
R28962 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 316.762
R28963 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 168.108
R28964 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 150.293
R28965 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 150.273
R28966 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 73.6406
R28967 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 73.6304
R28968 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 60.4568
R28969 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 12.0358
R28970 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 1.19615
R28971 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.981478
R28972 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 0.788543
R28973 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.769522
R28974 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 0.682565
R28975 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.580578
R28976 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 0.55213
R28977 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 0.484875
R28978 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 0.470609
R28979 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.447191
R28980 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.428234
R28981 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.217464
R28982 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R28983 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R28984 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R28985 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 0.063
R28986 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 0.063
R28987 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.063
R28988 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 0.063
R28989 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 0.063
R28990 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 0.0216397
R28991 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.0216397
R28992 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 0.0107679
R28993 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.0107679
R28994 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 179.256
R28995 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 168.089
R28996 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 150.293
R28997 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 73.6304
R28998 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 60.4568
R28999 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 12.0358
R29000 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.981478
R29001 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 0.788543
R29002 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.769522
R29003 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 0.720633
R29004 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 0.682565
R29005 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.580578
R29006 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 0.55213
R29007 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 0.470609
R29008 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.447191
R29009 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.428234
R29010 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1255
R29011 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1255
R29012 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 0.063
R29013 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 0.063
R29014 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.063
R29015 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 0.063
R29016 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 0.063
R29017 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 0.0435206
R29018 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 0.0107679
R29019 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.0107679
R29020 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 169.46
R29021 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 168.089
R29022 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 167.809
R29023 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 150.273
R29024 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 73.6406
R29025 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 60.3809
R29026 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 12.0358
R29027 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 11.4489
R29028 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 1.08746
R29029 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.851043
R29030 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.848156
R29031 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 0.788543
R29032 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 0.682565
R29033 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.65675
R29034 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 0.55213
R29035 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.486828
R29036 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 0.470609
R29037 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 0.262643
R29038 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.217464
R29039 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.1255
R29040 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.1255
R29041 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 0.063
R29042 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 0.063
R29043 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 0.063
R29044 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 0.063
R29045 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 0.063
R29046 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 0.0216397
R29047 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.0216397
R29048 Nand_Gate_5.A.n55 Nand_Gate_5.A.t1 169.46
R29049 Nand_Gate_5.A.n57 Nand_Gate_5.A.t3 167.809
R29050 Nand_Gate_5.A.n55 Nand_Gate_5.A.t0 167.809
R29051 Nand_Gate_5.A Nand_Gate_5.A.t7 158.585
R29052 Nand_Gate_5.A Nand_Gate_5.A.t17 158.581
R29053 Nand_Gate_5.A.n42 Nand_Gate_5.A.t9 150.293
R29054 Nand_Gate_5.A.t17 Nand_Gate_5.A.n38 150.293
R29055 Nand_Gate_5.A.t7 Nand_Gate_5.A.n2 150.293
R29056 Nand_Gate_5.A.n29 Nand_Gate_5.A.t14 150.273
R29057 Nand_Gate_5.A.n23 Nand_Gate_5.A.t5 150.273
R29058 Nand_Gate_5.A.n14 Nand_Gate_5.A.t11 150.273
R29059 Nand_Gate_5.A.n8 Nand_Gate_5.A.t12 150.273
R29060 Nand_Gate_5.A.n27 Nand_Gate_5.A.t6 73.6406
R29061 Nand_Gate_5.A.n21 Nand_Gate_5.A.t15 73.6406
R29062 Nand_Gate_5.A.n12 Nand_Gate_5.A.t13 73.6406
R29063 Nand_Gate_5.A.n6 Nand_Gate_5.A.t8 73.6406
R29064 Nand_Gate_5.A.n44 Nand_Gate_5.A.t4 73.6304
R29065 Nand_Gate_5.A.n36 Nand_Gate_5.A.t10 73.6304
R29066 Nand_Gate_5.A.n0 Nand_Gate_5.A.t16 73.6304
R29067 Nand_Gate_5.A.n4 Nand_Gate_5.A.t2 60.3809
R29068 Nand_Gate_5.A.n48 Nand_Gate_5.A.n41 25.1004
R29069 Nand_Gate_5.A.n33 Nand_Gate_5.A.n26 15.5222
R29070 Nand_Gate_5.A.n56 Nand_Gate_5.A.n55 11.4489
R29071 Nand_Gate_5.A.n48 Nand_Gate_5.A.n47 9.57083
R29072 Nand_Gate_5.A.n34 Nand_Gate_5.A.n33 8.26552
R29073 Nand_Gate_5.A.n58 Nand_Gate_5.A.n57 8.21389
R29074 Nand_Gate_5.A.n18 Nand_Gate_5.A.n11 8.1418
R29075 Nand_Gate_5.A.n49 Nand_Gate_5.A.n48 6.58222
R29076 Nand_Gate_5.A.n20 Nand_Gate_5.A.n19 6.47604
R29077 Nand_Gate_5.A.n19 Nand_Gate_5.A 5.35402
R29078 Nand_Gate_5.A.n52 Nand_Gate_5.A 4.55128
R29079 Nand_Gate_5.A.n33 Nand_Gate_5.A.n32 4.5005
R29080 Nand_Gate_5.A.n18 Nand_Gate_5.A.n17 4.5005
R29081 Nand_Gate_5.A.n38 Nand_Gate_5.A.n37 1.19615
R29082 Nand_Gate_5.A.n2 Nand_Gate_5.A.n1 1.19615
R29083 Nand_Gate_5.A.n5 Nand_Gate_5.A 1.08746
R29084 Nand_Gate_5.A.n20 Nand_Gate_5.A 0.973326
R29085 Nand_Gate_5.A.n13 Nand_Gate_5.A 0.851043
R29086 Nand_Gate_5.A.n7 Nand_Gate_5.A 0.851043
R29087 Nand_Gate_5.A.n4 Nand_Gate_5.A 0.848156
R29088 Nand_Gate_5.A.n28 Nand_Gate_5.A.n27 0.796696
R29089 Nand_Gate_5.A.n22 Nand_Gate_5.A.n21 0.796696
R29090 Nand_Gate_5.A.n54 Nand_Gate_5.A.n53 0.788543
R29091 Nand_Gate_5.A.n43 Nand_Gate_5.A 0.769522
R29092 Nand_Gate_5.A.n51 Nand_Gate_5.A.n50 0.755935
R29093 Nand_Gate_5.A.n34 Nand_Gate_5.A 0.716182
R29094 Nand_Gate_5.A.n5 Nand_Gate_5.A.n4 0.682565
R29095 Nand_Gate_5.A.n53 Nand_Gate_5.A 0.65675
R29096 Nand_Gate_5.A.n43 Nand_Gate_5.A.n42 0.55213
R29097 Nand_Gate_5.A.n16 Nand_Gate_5.A.n15 0.55213
R29098 Nand_Gate_5.A.n10 Nand_Gate_5.A.n9 0.55213
R29099 Nand_Gate_5.A.n35 Nand_Gate_5.A.n34 0.546483
R29100 Nand_Gate_5.A.n28 Nand_Gate_5.A 0.524957
R29101 Nand_Gate_5.A.n22 Nand_Gate_5.A 0.524957
R29102 Nand_Gate_5.A.n16 Nand_Gate_5.A 0.486828
R29103 Nand_Gate_5.A.n10 Nand_Gate_5.A 0.486828
R29104 Nand_Gate_5.A.n50 Nand_Gate_5.A 0.48023
R29105 Nand_Gate_5.A.n46 Nand_Gate_5.A.n45 0.470609
R29106 Nand_Gate_5.A.n13 Nand_Gate_5.A.n12 0.470609
R29107 Nand_Gate_5.A.n7 Nand_Gate_5.A.n6 0.470609
R29108 Nand_Gate_5.A.n42 Nand_Gate_5.A 0.447191
R29109 Nand_Gate_5.A.n38 Nand_Gate_5.A 0.447191
R29110 Nand_Gate_5.A.n2 Nand_Gate_5.A 0.447191
R29111 Nand_Gate_5.A.n46 Nand_Gate_5.A 0.428234
R29112 Nand_Gate_5.A.n58 Nand_Gate_5.A.n3 0.425067
R29113 Nand_Gate_5.A Nand_Gate_5.A.n58 0.39003
R29114 Nand_Gate_5.A.n57 Nand_Gate_5.A.n56 0.280391
R29115 Nand_Gate_5.A.n31 Nand_Gate_5.A 0.252453
R29116 Nand_Gate_5.A.n25 Nand_Gate_5.A 0.252453
R29117 Nand_Gate_5.A.n35 Nand_Gate_5.A 0.241767
R29118 Nand_Gate_5.A.n31 Nand_Gate_5.A.n30 0.226043
R29119 Nand_Gate_5.A.n25 Nand_Gate_5.A.n24 0.226043
R29120 Nand_Gate_5.A.n27 Nand_Gate_5.A 0.217464
R29121 Nand_Gate_5.A.n21 Nand_Gate_5.A 0.217464
R29122 Nand_Gate_5.A.n12 Nand_Gate_5.A 0.217464
R29123 Nand_Gate_5.A.n6 Nand_Gate_5.A 0.217464
R29124 Nand_Gate_5.A.n56 Nand_Gate_5.A 0.200143
R29125 Nand_Gate_5.A.n40 Nand_Gate_5.A.n39 0.178317
R29126 Nand_Gate_5.A.n40 Nand_Gate_5.A 0.143974
R29127 Nand_Gate_5.A.n45 Nand_Gate_5.A 0.1255
R29128 Nand_Gate_5.A.n30 Nand_Gate_5.A 0.1255
R29129 Nand_Gate_5.A.n24 Nand_Gate_5.A 0.1255
R29130 Nand_Gate_5.A.n37 Nand_Gate_5.A 0.1255
R29131 Nand_Gate_5.A.n15 Nand_Gate_5.A 0.1255
R29132 Nand_Gate_5.A.n9 Nand_Gate_5.A 0.1255
R29133 Nand_Gate_5.A.n54 Nand_Gate_5.A 0.1255
R29134 Nand_Gate_5.A.n1 Nand_Gate_5.A 0.1255
R29135 Nand_Gate_5.A.n47 Nand_Gate_5.A.n43 0.063
R29136 Nand_Gate_5.A.n47 Nand_Gate_5.A.n46 0.063
R29137 Nand_Gate_5.A.n32 Nand_Gate_5.A.n28 0.063
R29138 Nand_Gate_5.A.n32 Nand_Gate_5.A.n31 0.063
R29139 Nand_Gate_5.A.n26 Nand_Gate_5.A.n22 0.063
R29140 Nand_Gate_5.A.n26 Nand_Gate_5.A.n25 0.063
R29141 Nand_Gate_5.A.n17 Nand_Gate_5.A.n13 0.063
R29142 Nand_Gate_5.A.n17 Nand_Gate_5.A.n16 0.063
R29143 Nand_Gate_5.A.n11 Nand_Gate_5.A.n7 0.063
R29144 Nand_Gate_5.A.n11 Nand_Gate_5.A.n10 0.063
R29145 Nand_Gate_5.A.n19 Nand_Gate_5.A.n18 0.063
R29146 Nand_Gate_5.A.n49 Nand_Gate_5.A.n20 0.063
R29147 Nand_Gate_5.A.n50 Nand_Gate_5.A.n49 0.063
R29148 Nand_Gate_5.A.n52 Nand_Gate_5.A.n5 0.063
R29149 Nand_Gate_5.A.n53 Nand_Gate_5.A.n52 0.063
R29150 Nand_Gate_5.A Nand_Gate_5.A.n54 0.063
R29151 Nand_Gate_5.A.n41 Nand_Gate_5.A.n35 0.024
R29152 Nand_Gate_5.A.n41 Nand_Gate_5.A.n40 0.024
R29153 Nand_Gate_5.A.n30 Nand_Gate_5.A.n29 0.0216397
R29154 Nand_Gate_5.A.n29 Nand_Gate_5.A 0.0216397
R29155 Nand_Gate_5.A.n24 Nand_Gate_5.A.n23 0.0216397
R29156 Nand_Gate_5.A.n23 Nand_Gate_5.A 0.0216397
R29157 Nand_Gate_5.A.n15 Nand_Gate_5.A.n14 0.0216397
R29158 Nand_Gate_5.A.n14 Nand_Gate_5.A 0.0216397
R29159 Nand_Gate_5.A.n9 Nand_Gate_5.A.n8 0.0216397
R29160 Nand_Gate_5.A.n8 Nand_Gate_5.A 0.0216397
R29161 Nand_Gate_5.A.n51 Nand_Gate_5.A 0.0168043
R29162 Nand_Gate_5.A Nand_Gate_5.A.n51 0.0122188
R29163 Nand_Gate_5.A.n45 Nand_Gate_5.A.n44 0.0107679
R29164 Nand_Gate_5.A.n44 Nand_Gate_5.A 0.0107679
R29165 Nand_Gate_5.A.n37 Nand_Gate_5.A.n36 0.0107679
R29166 Nand_Gate_5.A.n36 Nand_Gate_5.A 0.0107679
R29167 Nand_Gate_5.A.n1 Nand_Gate_5.A.n0 0.0107679
R29168 Nand_Gate_5.A.n0 Nand_Gate_5.A 0.0107679
R29169 Nand_Gate_5.A.n39 Nand_Gate_5.A 0.00441667
R29170 Nand_Gate_5.A.n3 Nand_Gate_5.A 0.00441667
R29171 Nand_Gate_5.A.n39 Nand_Gate_5.A 0.00406061
R29172 Nand_Gate_5.A.n3 Nand_Gate_5.A 0.00406061
R29173 a_138533_35417.n0 a_138533_35417.t3 1546.57
R29174 a_138533_35417.n1 a_138533_35417.t1 27.7124
R29175 a_138533_35417.t0 a_138533_35417.n1 21.1744
R29176 a_138533_35417.n0 a_138533_35417.t2 11.1233
R29177 a_138533_35417.n1 a_138533_35417.n0 5.89691
R29178 Nand_Gate_4.B.n51 Nand_Gate_4.B.t2 169.46
R29179 Nand_Gate_4.B.n51 Nand_Gate_4.B.t3 167.809
R29180 Nand_Gate_4.B.n53 Nand_Gate_4.B.t0 167.809
R29181 Nand_Gate_4.B Nand_Gate_4.B.t17 158.585
R29182 Nand_Gate_4.B Nand_Gate_4.B.t7 158.581
R29183 Nand_Gate_4.B.n42 Nand_Gate_4.B.t10 150.293
R29184 Nand_Gate_4.B.t7 Nand_Gate_4.B.n38 150.293
R29185 Nand_Gate_4.B.t17 Nand_Gate_4.B.n2 150.293
R29186 Nand_Gate_4.B.n29 Nand_Gate_4.B.t4 150.273
R29187 Nand_Gate_4.B.n23 Nand_Gate_4.B.t11 150.273
R29188 Nand_Gate_4.B.n14 Nand_Gate_4.B.t6 150.273
R29189 Nand_Gate_4.B.n8 Nand_Gate_4.B.t16 150.273
R29190 Nand_Gate_4.B.n44 Nand_Gate_4.B.n41 76.0985
R29191 Nand_Gate_4.B.n27 Nand_Gate_4.B.t12 73.6406
R29192 Nand_Gate_4.B.n21 Nand_Gate_4.B.t5 73.6406
R29193 Nand_Gate_4.B.n12 Nand_Gate_4.B.t14 73.6406
R29194 Nand_Gate_4.B.n6 Nand_Gate_4.B.t13 73.6406
R29195 Nand_Gate_4.B.n43 Nand_Gate_4.B.t8 73.6304
R29196 Nand_Gate_4.B.n36 Nand_Gate_4.B.t15 73.6304
R29197 Nand_Gate_4.B.n0 Nand_Gate_4.B.t9 73.6304
R29198 Nand_Gate_4.B.n4 Nand_Gate_4.B.t1 60.3809
R29199 Nand_Gate_4.B.n44 Nand_Gate_4.B.n43 34.7148
R29200 Nand_Gate_4.B.n33 Nand_Gate_4.B.n26 15.5222
R29201 Nand_Gate_4.B.n52 Nand_Gate_4.B.n51 11.4489
R29202 Nand_Gate_4.B.n34 Nand_Gate_4.B.n33 8.26552
R29203 Nand_Gate_4.B.n54 Nand_Gate_4.B.n53 8.21389
R29204 Nand_Gate_4.B.n18 Nand_Gate_4.B.n11 8.1418
R29205 Nand_Gate_4.B.n47 Nand_Gate_4.B.n46 5.61191
R29206 Nand_Gate_4.B.n47 Nand_Gate_4.B 5.35402
R29207 Nand_Gate_4.B.n45 Nand_Gate_4.B.n44 4.81893
R29208 Nand_Gate_4.B.n48 Nand_Gate_4.B.n47 4.563
R29209 Nand_Gate_4.B.n33 Nand_Gate_4.B.n32 4.5005
R29210 Nand_Gate_4.B.n18 Nand_Gate_4.B.n17 4.5005
R29211 Nand_Gate_4.B.n46 Nand_Gate_4.B 1.83746
R29212 Nand_Gate_4.B.n20 Nand_Gate_4.B.n19 1.62007
R29213 Nand_Gate_4.B.n38 Nand_Gate_4.B.n37 1.19615
R29214 Nand_Gate_4.B.n2 Nand_Gate_4.B.n1 1.19615
R29215 Nand_Gate_4.B.n43 Nand_Gate_4.B.n42 1.1717
R29216 Nand_Gate_4.B.n5 Nand_Gate_4.B 1.08746
R29217 Nand_Gate_4.B.n20 Nand_Gate_4.B 1.01739
R29218 Nand_Gate_4.B.n13 Nand_Gate_4.B 0.851043
R29219 Nand_Gate_4.B.n7 Nand_Gate_4.B 0.851043
R29220 Nand_Gate_4.B.n4 Nand_Gate_4.B 0.848156
R29221 Nand_Gate_4.B.n28 Nand_Gate_4.B.n27 0.796696
R29222 Nand_Gate_4.B.n22 Nand_Gate_4.B.n21 0.796696
R29223 Nand_Gate_4.B.n50 Nand_Gate_4.B.n49 0.788543
R29224 Nand_Gate_4.B.n34 Nand_Gate_4.B 0.716182
R29225 Nand_Gate_4.B.n5 Nand_Gate_4.B.n4 0.682565
R29226 Nand_Gate_4.B.n49 Nand_Gate_4.B 0.65675
R29227 Nand_Gate_4.B.n16 Nand_Gate_4.B.n15 0.55213
R29228 Nand_Gate_4.B.n10 Nand_Gate_4.B.n9 0.55213
R29229 Nand_Gate_4.B.n28 Nand_Gate_4.B 0.524957
R29230 Nand_Gate_4.B.n22 Nand_Gate_4.B 0.524957
R29231 Nand_Gate_4.B.n16 Nand_Gate_4.B 0.486828
R29232 Nand_Gate_4.B.n10 Nand_Gate_4.B 0.486828
R29233 Nand_Gate_4.B.n13 Nand_Gate_4.B.n12 0.470609
R29234 Nand_Gate_4.B.n7 Nand_Gate_4.B.n6 0.470609
R29235 Nand_Gate_4.B.n42 Nand_Gate_4.B 0.447191
R29236 Nand_Gate_4.B.n38 Nand_Gate_4.B 0.447191
R29237 Nand_Gate_4.B.n2 Nand_Gate_4.B 0.447191
R29238 Nand_Gate_4.B.n54 Nand_Gate_4.B.n3 0.425067
R29239 Nand_Gate_4.B.n35 Nand_Gate_4.B 0.412533
R29240 Nand_Gate_4.B Nand_Gate_4.B.n54 0.39003
R29241 Nand_Gate_4.B.n35 Nand_Gate_4.B.n34 0.375717
R29242 Nand_Gate_4.B.n40 Nand_Gate_4.B.n39 0.349083
R29243 Nand_Gate_4.B.n53 Nand_Gate_4.B.n52 0.280391
R29244 Nand_Gate_4.B.n40 Nand_Gate_4.B 0.278789
R29245 Nand_Gate_4.B.n52 Nand_Gate_4.B.n50 0.262643
R29246 Nand_Gate_4.B.n31 Nand_Gate_4.B 0.252453
R29247 Nand_Gate_4.B.n25 Nand_Gate_4.B 0.252453
R29248 Nand_Gate_4.B.n31 Nand_Gate_4.B.n30 0.226043
R29249 Nand_Gate_4.B.n25 Nand_Gate_4.B.n24 0.226043
R29250 Nand_Gate_4.B.n27 Nand_Gate_4.B 0.217464
R29251 Nand_Gate_4.B.n21 Nand_Gate_4.B 0.217464
R29252 Nand_Gate_4.B.n12 Nand_Gate_4.B 0.217464
R29253 Nand_Gate_4.B.n6 Nand_Gate_4.B 0.217464
R29254 Nand_Gate_4.B.n43 Nand_Gate_4.B 0.149957
R29255 Nand_Gate_4.B.n30 Nand_Gate_4.B 0.1255
R29256 Nand_Gate_4.B.n24 Nand_Gate_4.B 0.1255
R29257 Nand_Gate_4.B.n37 Nand_Gate_4.B 0.1255
R29258 Nand_Gate_4.B.n15 Nand_Gate_4.B 0.1255
R29259 Nand_Gate_4.B.n9 Nand_Gate_4.B 0.1255
R29260 Nand_Gate_4.B.n50 Nand_Gate_4.B 0.1255
R29261 Nand_Gate_4.B.n1 Nand_Gate_4.B 0.1255
R29262 Nand_Gate_4.B.n32 Nand_Gate_4.B.n28 0.063
R29263 Nand_Gate_4.B.n32 Nand_Gate_4.B.n31 0.063
R29264 Nand_Gate_4.B.n26 Nand_Gate_4.B.n22 0.063
R29265 Nand_Gate_4.B.n26 Nand_Gate_4.B.n25 0.063
R29266 Nand_Gate_4.B.n17 Nand_Gate_4.B.n13 0.063
R29267 Nand_Gate_4.B.n17 Nand_Gate_4.B.n16 0.063
R29268 Nand_Gate_4.B.n11 Nand_Gate_4.B.n7 0.063
R29269 Nand_Gate_4.B.n11 Nand_Gate_4.B.n10 0.063
R29270 Nand_Gate_4.B.n46 Nand_Gate_4.B.n45 0.063
R29271 Nand_Gate_4.B.n45 Nand_Gate_4.B.n20 0.063
R29272 Nand_Gate_4.B.n48 Nand_Gate_4.B.n5 0.063
R29273 Nand_Gate_4.B.n49 Nand_Gate_4.B.n48 0.063
R29274 Nand_Gate_4.B.n50 Nand_Gate_4.B 0.063
R29275 Nand_Gate_4.B Nand_Gate_4.B.n18 0.0512812
R29276 Nand_Gate_4.B.n43 Nand_Gate_4.B 0.0454219
R29277 Nand_Gate_4.B.n41 Nand_Gate_4.B.n35 0.024
R29278 Nand_Gate_4.B.n41 Nand_Gate_4.B.n40 0.024
R29279 Nand_Gate_4.B.n30 Nand_Gate_4.B.n29 0.0216397
R29280 Nand_Gate_4.B.n29 Nand_Gate_4.B 0.0216397
R29281 Nand_Gate_4.B.n24 Nand_Gate_4.B.n23 0.0216397
R29282 Nand_Gate_4.B.n23 Nand_Gate_4.B 0.0216397
R29283 Nand_Gate_4.B.n15 Nand_Gate_4.B.n14 0.0216397
R29284 Nand_Gate_4.B.n14 Nand_Gate_4.B 0.0216397
R29285 Nand_Gate_4.B.n9 Nand_Gate_4.B.n8 0.0216397
R29286 Nand_Gate_4.B.n8 Nand_Gate_4.B 0.0216397
R29287 Nand_Gate_4.B.n19 Nand_Gate_4.B 0.0168043
R29288 Nand_Gate_4.B.n19 Nand_Gate_4.B 0.0122188
R29289 Nand_Gate_4.B.n37 Nand_Gate_4.B.n36 0.0107679
R29290 Nand_Gate_4.B.n36 Nand_Gate_4.B 0.0107679
R29291 Nand_Gate_4.B.n1 Nand_Gate_4.B.n0 0.0107679
R29292 Nand_Gate_4.B.n0 Nand_Gate_4.B 0.0107679
R29293 Nand_Gate_4.B.n39 Nand_Gate_4.B 0.00441667
R29294 Nand_Gate_4.B.n3 Nand_Gate_4.B 0.00441667
R29295 Nand_Gate_4.B.n39 Nand_Gate_4.B 0.00406061
R29296 Nand_Gate_4.B.n3 Nand_Gate_4.B 0.00406061
R29297 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t0 169.46
R29298 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t1 167.809
R29299 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.t2 167.809
R29300 D_FlipFlop_3.3-input-nand_2.Vout.t6 D_FlipFlop_3.3-input-nand_2.Vout.n11 167.227
R29301 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.t6 150.293
R29302 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.t5 150.273
R29303 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout.t7 73.6406
R29304 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout.t4 73.6304
R29305 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout.t3 60.3809
R29306 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n5 12.3891
R29307 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout.n9 11.4489
R29308 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout.n2 1.38365
R29309 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.n1 1.19615
R29310 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.n4 1.1717
R29311 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout 0.848156
R29312 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.Vout.n12 0.447191
R29313 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R29314 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.n10 0.280391
R29315 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout.n8 0.262643
R29316 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout 0.217464
R29317 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R29318 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R29319 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R29320 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R29321 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout.n7 0.0874565
R29322 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n3 0.063
R29323 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout.n6 0.063
R29324 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout 0.063
R29325 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R29326 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout.n0 0.0107679
R29327 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout 0.0107679
R29328 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t0 169.46
R29329 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t3 167.809
R29330 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.t1 167.809
R29331 D_FlipFlop_3.3-input-nand_2.C.t4 D_FlipFlop_3.3-input-nand_2.C.n13 167.226
R29332 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.t5 150.273
R29333 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.t4 150.273
R29334 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C.t7 73.6406
R29335 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C.t6 73.6304
R29336 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C.t2 60.4568
R29337 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n7 12.3891
R29338 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n11 11.4489
R29339 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C 1.68257
R29340 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C.n2 1.38365
R29341 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C.n0 1.19615
R29342 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C.n5 1.1717
R29343 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C 1.08448
R29344 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C 0.932141
R29345 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C 0.720633
R29346 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.n12 0.280391
R29347 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C 0.217464
R29348 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29349 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29350 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29351 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C.n9 0.0874565
R29352 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.n6 0.063
R29353 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.063
R29354 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C.n8 0.063
R29355 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n3 0.063
R29356 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n10 0.0435206
R29357 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.n1 0.0216397
R29358 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.C.n14 0.0216397
R29359 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C.n4 0.0107679
R29360 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C 0.0107679
R29361 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.t3 169.46
R29362 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C.t2 167.809
R29363 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.t0 167.809
R29364 D_FlipFlop_0.3-input-nand_2.C.t7 D_FlipFlop_0.3-input-nand_2.C.n13 167.226
R29365 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C.t4 150.273
R29366 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.t7 150.273
R29367 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C.t6 73.6406
R29368 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C.t5 73.6304
R29369 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C.t1 60.4568
R29370 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C.n7 12.3891
R29371 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n11 11.4489
R29372 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C 1.68257
R29373 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C.n2 1.38365
R29374 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C.n0 1.19615
R29375 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C.n5 1.1717
R29376 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C 1.08448
R29377 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C 0.932141
R29378 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C 0.720633
R29379 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C.n12 0.280391
R29380 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C 0.217464
R29381 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C 0.1255
R29382 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C 0.1255
R29383 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C 0.1255
R29384 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C.n9 0.0874565
R29385 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C.n6 0.063
R29386 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C 0.063
R29387 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C.n8 0.063
R29388 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C.n3 0.063
R29389 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n10 0.0435206
R29390 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.n1 0.0216397
R29391 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_2.C.n14 0.0216397
R29392 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C.n4 0.0107679
R29393 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C 0.0107679
R29394 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 169.46
R29395 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 168.089
R29396 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 167.809
R29397 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 150.293
R29398 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 73.6304
R29399 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 60.3943
R29400 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 12.0358
R29401 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 11.4489
R29402 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.981478
R29403 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 0.788543
R29404 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.769522
R29405 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 0.720633
R29406 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 0.682565
R29407 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.580578
R29408 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 0.55213
R29409 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 0.470609
R29410 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.447191
R29411 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.428234
R29412 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.1255
R29413 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.1255
R29414 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 0.063
R29415 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 0.063
R29416 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.063
R29417 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 0.063
R29418 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 0.063
R29419 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 0.0435206
R29420 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 0.0107679
R29421 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.0107679
R29422 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 169.46
R29423 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 168.089
R29424 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 167.809
R29425 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 150.293
R29426 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 73.6304
R29427 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 60.4568
R29428 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 12.0358
R29429 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 11.4489
R29430 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.981478
R29431 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 0.788543
R29432 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.769522
R29433 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 0.720633
R29434 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 0.682565
R29435 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.580578
R29436 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 0.55213
R29437 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 0.470609
R29438 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.447191
R29439 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.428234
R29440 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.1255
R29441 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.1255
R29442 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 0.063
R29443 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 0.063
R29444 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.063
R29445 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 0.063
R29446 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 0.063
R29447 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 0.0435206
R29448 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 0.0107679
R29449 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.0107679
R29450 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 169.46
R29451 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 168.089
R29452 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 167.809
R29453 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 150.273
R29454 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 73.6406
R29455 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 60.3809
R29456 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 12.0358
R29457 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 11.4489
R29458 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 1.08746
R29459 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.851043
R29460 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.848156
R29461 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 0.788543
R29462 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 0.682565
R29463 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.65675
R29464 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 0.55213
R29465 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.486828
R29466 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 0.470609
R29467 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.217464
R29468 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 0.200143
R29469 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.1255
R29470 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.1255
R29471 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 0.063
R29472 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 0.063
R29473 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 0.063
R29474 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 0.063
R29475 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 0.063
R29476 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 0.0216397
R29477 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.0216397
R29478 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 169.46
R29479 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 167.809
R29480 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 167.809
R29481 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 167.226
R29482 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 150.273
R29483 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 150.273
R29484 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 73.6406
R29485 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 73.6304
R29486 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 60.4568
R29487 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 12.3891
R29488 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 11.4489
R29489 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.68257
R29490 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 1.38365
R29491 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 1.19615
R29492 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 1.1717
R29493 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.08448
R29494 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.932141
R29495 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.720633
R29496 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 0.280391
R29497 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.217464
R29498 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R29499 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R29500 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R29501 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 0.0874565
R29502 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 0.063
R29503 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.063
R29504 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 0.063
R29505 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 0.063
R29506 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 0.0435206
R29507 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 0.0216397
R29508 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 0.0216397
R29509 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 0.0107679
R29510 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.0107679
R29511 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 169.46
R29512 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 167.809
R29513 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 167.809
R29514 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 167.227
R29515 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 150.293
R29516 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 150.273
R29517 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 73.6406
R29518 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 73.6304
R29519 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 60.3809
R29520 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 12.3891
R29521 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 11.4489
R29522 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 1.38365
R29523 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 1.19615
R29524 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 1.1717
R29525 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.848156
R29526 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 0.447191
R29527 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.38637
R29528 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 0.280391
R29529 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 0.262643
R29530 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.217464
R29531 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.152844
R29532 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.149957
R29533 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.1255
R29534 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.1255
R29535 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 0.0874565
R29536 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 0.063
R29537 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 0.063
R29538 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.063
R29539 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.0454219
R29540 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 0.0107679
R29541 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.0107679
R29542 Nand_Gate_7.B.n6 Nand_Gate_7.B.t2 169.46
R29543 Nand_Gate_7.B.n6 Nand_Gate_7.B.t3 167.809
R29544 Nand_Gate_7.B.n5 Nand_Gate_7.B.t1 167.809
R29545 Nand_Gate_7.B Nand_Gate_7.B.t15 158.585
R29546 Nand_Gate_7.B Nand_Gate_7.B.t8 158.581
R29547 Nand_Gate_7.B.n46 Nand_Gate_7.B.t16 150.293
R29548 Nand_Gate_7.B.t8 Nand_Gate_7.B.n42 150.293
R29549 Nand_Gate_7.B.t15 Nand_Gate_7.B.n2 150.293
R29550 Nand_Gate_7.B.n33 Nand_Gate_7.B.t7 150.273
R29551 Nand_Gate_7.B.n27 Nand_Gate_7.B.t17 150.273
R29552 Nand_Gate_7.B.n18 Nand_Gate_7.B.t11 150.273
R29553 Nand_Gate_7.B.n12 Nand_Gate_7.B.t14 150.273
R29554 Nand_Gate_7.B.n31 Nand_Gate_7.B.t6 73.6406
R29555 Nand_Gate_7.B.n25 Nand_Gate_7.B.t12 73.6406
R29556 Nand_Gate_7.B.n16 Nand_Gate_7.B.t13 73.6406
R29557 Nand_Gate_7.B.n10 Nand_Gate_7.B.t10 73.6406
R29558 Nand_Gate_7.B.n47 Nand_Gate_7.B.t9 73.6304
R29559 Nand_Gate_7.B.n40 Nand_Gate_7.B.t4 73.6304
R29560 Nand_Gate_7.B.n0 Nand_Gate_7.B.t5 73.6304
R29561 Nand_Gate_7.B.n48 Nand_Gate_7.B.n45 61.6632
R29562 Nand_Gate_7.B.n54 Nand_Gate_7.B.t0 60.3809
R29563 Nand_Gate_7.B.n48 Nand_Gate_7.B.n47 34.7148
R29564 Nand_Gate_7.B.n37 Nand_Gate_7.B.n30 15.5222
R29565 Nand_Gate_7.B.n7 Nand_Gate_7.B.n6 11.4489
R29566 Nand_Gate_7.B.n38 Nand_Gate_7.B.n37 8.26552
R29567 Nand_Gate_7.B.n5 Nand_Gate_7.B.n4 8.21389
R29568 Nand_Gate_7.B.n22 Nand_Gate_7.B.n15 8.1418
R29569 Nand_Gate_7.B.n51 Nand_Gate_7.B.n50 5.61191
R29570 Nand_Gate_7.B.n51 Nand_Gate_7.B 5.35402
R29571 Nand_Gate_7.B.n49 Nand_Gate_7.B.n48 4.81893
R29572 Nand_Gate_7.B.n52 Nand_Gate_7.B.n51 4.563
R29573 Nand_Gate_7.B.n37 Nand_Gate_7.B.n36 4.5005
R29574 Nand_Gate_7.B.n22 Nand_Gate_7.B.n21 4.5005
R29575 Nand_Gate_7.B.n50 Nand_Gate_7.B 1.83746
R29576 Nand_Gate_7.B.n24 Nand_Gate_7.B.n23 1.62007
R29577 Nand_Gate_7.B.n42 Nand_Gate_7.B.n41 1.19615
R29578 Nand_Gate_7.B.n2 Nand_Gate_7.B.n1 1.19615
R29579 Nand_Gate_7.B.n47 Nand_Gate_7.B.n46 1.1717
R29580 Nand_Gate_7.B.n53 Nand_Gate_7.B 1.08746
R29581 Nand_Gate_7.B.n24 Nand_Gate_7.B 1.01739
R29582 Nand_Gate_7.B.n17 Nand_Gate_7.B 0.851043
R29583 Nand_Gate_7.B.n11 Nand_Gate_7.B 0.851043
R29584 Nand_Gate_7.B Nand_Gate_7.B.n54 0.848156
R29585 Nand_Gate_7.B.n32 Nand_Gate_7.B.n31 0.796696
R29586 Nand_Gate_7.B.n26 Nand_Gate_7.B.n25 0.796696
R29587 Nand_Gate_7.B.n9 Nand_Gate_7.B.n8 0.788543
R29588 Nand_Gate_7.B.n38 Nand_Gate_7.B 0.716182
R29589 Nand_Gate_7.B.n54 Nand_Gate_7.B.n53 0.682565
R29590 Nand_Gate_7.B.n9 Nand_Gate_7.B 0.65675
R29591 Nand_Gate_7.B.n20 Nand_Gate_7.B.n19 0.55213
R29592 Nand_Gate_7.B.n14 Nand_Gate_7.B.n13 0.55213
R29593 Nand_Gate_7.B.n32 Nand_Gate_7.B 0.524957
R29594 Nand_Gate_7.B.n26 Nand_Gate_7.B 0.524957
R29595 Nand_Gate_7.B.n20 Nand_Gate_7.B 0.486828
R29596 Nand_Gate_7.B.n14 Nand_Gate_7.B 0.486828
R29597 Nand_Gate_7.B.n39 Nand_Gate_7.B 0.481467
R29598 Nand_Gate_7.B.n17 Nand_Gate_7.B.n16 0.470609
R29599 Nand_Gate_7.B.n11 Nand_Gate_7.B.n10 0.470609
R29600 Nand_Gate_7.B.n46 Nand_Gate_7.B 0.447191
R29601 Nand_Gate_7.B.n42 Nand_Gate_7.B 0.447191
R29602 Nand_Gate_7.B.n2 Nand_Gate_7.B 0.447191
R29603 Nand_Gate_7.B.n4 Nand_Gate_7.B.n3 0.425067
R29604 Nand_Gate_7.B.n44 Nand_Gate_7.B.n43 0.418017
R29605 Nand_Gate_7.B.n4 Nand_Gate_7.B 0.39003
R29606 Nand_Gate_7.B.n44 Nand_Gate_7.B 0.333211
R29607 Nand_Gate_7.B.n39 Nand_Gate_7.B.n38 0.306783
R29608 Nand_Gate_7.B.n7 Nand_Gate_7.B.n5 0.280391
R29609 Nand_Gate_7.B.n8 Nand_Gate_7.B.n7 0.262643
R29610 Nand_Gate_7.B.n35 Nand_Gate_7.B 0.252453
R29611 Nand_Gate_7.B.n29 Nand_Gate_7.B 0.252453
R29612 Nand_Gate_7.B.n35 Nand_Gate_7.B.n34 0.226043
R29613 Nand_Gate_7.B.n29 Nand_Gate_7.B.n28 0.226043
R29614 Nand_Gate_7.B.n31 Nand_Gate_7.B 0.217464
R29615 Nand_Gate_7.B.n25 Nand_Gate_7.B 0.217464
R29616 Nand_Gate_7.B.n16 Nand_Gate_7.B 0.217464
R29617 Nand_Gate_7.B.n10 Nand_Gate_7.B 0.217464
R29618 Nand_Gate_7.B.n47 Nand_Gate_7.B 0.149957
R29619 Nand_Gate_7.B.n34 Nand_Gate_7.B 0.1255
R29620 Nand_Gate_7.B.n28 Nand_Gate_7.B 0.1255
R29621 Nand_Gate_7.B.n41 Nand_Gate_7.B 0.1255
R29622 Nand_Gate_7.B.n19 Nand_Gate_7.B 0.1255
R29623 Nand_Gate_7.B.n13 Nand_Gate_7.B 0.1255
R29624 Nand_Gate_7.B.n1 Nand_Gate_7.B 0.1255
R29625 Nand_Gate_7.B.n8 Nand_Gate_7.B 0.1255
R29626 Nand_Gate_7.B.n36 Nand_Gate_7.B.n32 0.063
R29627 Nand_Gate_7.B.n36 Nand_Gate_7.B.n35 0.063
R29628 Nand_Gate_7.B.n30 Nand_Gate_7.B.n26 0.063
R29629 Nand_Gate_7.B.n30 Nand_Gate_7.B.n29 0.063
R29630 Nand_Gate_7.B.n21 Nand_Gate_7.B.n17 0.063
R29631 Nand_Gate_7.B.n21 Nand_Gate_7.B.n20 0.063
R29632 Nand_Gate_7.B.n15 Nand_Gate_7.B.n11 0.063
R29633 Nand_Gate_7.B.n15 Nand_Gate_7.B.n14 0.063
R29634 Nand_Gate_7.B.n50 Nand_Gate_7.B.n49 0.063
R29635 Nand_Gate_7.B.n49 Nand_Gate_7.B.n24 0.063
R29636 Nand_Gate_7.B.n8 Nand_Gate_7.B 0.063
R29637 Nand_Gate_7.B.n53 Nand_Gate_7.B.n52 0.063
R29638 Nand_Gate_7.B.n52 Nand_Gate_7.B.n9 0.063
R29639 Nand_Gate_7.B Nand_Gate_7.B.n22 0.0512812
R29640 Nand_Gate_7.B.n47 Nand_Gate_7.B 0.0454219
R29641 Nand_Gate_7.B.n45 Nand_Gate_7.B.n39 0.024
R29642 Nand_Gate_7.B.n45 Nand_Gate_7.B.n44 0.024
R29643 Nand_Gate_7.B.n34 Nand_Gate_7.B.n33 0.0216397
R29644 Nand_Gate_7.B.n33 Nand_Gate_7.B 0.0216397
R29645 Nand_Gate_7.B.n28 Nand_Gate_7.B.n27 0.0216397
R29646 Nand_Gate_7.B.n27 Nand_Gate_7.B 0.0216397
R29647 Nand_Gate_7.B.n19 Nand_Gate_7.B.n18 0.0216397
R29648 Nand_Gate_7.B.n18 Nand_Gate_7.B 0.0216397
R29649 Nand_Gate_7.B.n13 Nand_Gate_7.B.n12 0.0216397
R29650 Nand_Gate_7.B.n12 Nand_Gate_7.B 0.0216397
R29651 Nand_Gate_7.B.n23 Nand_Gate_7.B 0.0168043
R29652 Nand_Gate_7.B.n23 Nand_Gate_7.B 0.0122188
R29653 Nand_Gate_7.B.n41 Nand_Gate_7.B.n40 0.0107679
R29654 Nand_Gate_7.B.n40 Nand_Gate_7.B 0.0107679
R29655 Nand_Gate_7.B.n1 Nand_Gate_7.B.n0 0.0107679
R29656 Nand_Gate_7.B.n0 Nand_Gate_7.B 0.0107679
R29657 Nand_Gate_7.B.n43 Nand_Gate_7.B 0.00441667
R29658 Nand_Gate_7.B.n3 Nand_Gate_7.B 0.00441667
R29659 Nand_Gate_7.B.n43 Nand_Gate_7.B 0.00406061
R29660 Nand_Gate_7.B.n3 Nand_Gate_7.B 0.00406061
R29661 Q1.n5 Q1.t1 169.46
R29662 Q1.n7 Q1.t2 167.809
R29663 Q1.n5 Q1.t0 167.809
R29664 Q1.n11 Q1.t4 155.124
R29665 Q1.n14 Q1.t7 150.869
R29666 Q1.n13 Q1.t9 150.869
R29667 Q1.t4 Q1.n2 150.293
R29668 Q1.n15 Q1.n12 137.644
R29669 Q1 Q1.t5 78.1811
R29670 Q1.n13 Q1.t6 74.1352
R29671 Q1.t5 Q1.n14 74.1352
R29672 Q1.n0 Q1.t8 73.6304
R29673 Q1.n3 Q1.t3 60.3809
R29674 Q1.n12 Q1 41.1198
R29675 Q1.n6 Q1.n5 11.4489
R29676 Q1.n8 Q1.n7 8.21389
R29677 Q1.n11 Q1.n10 1.70176
R29678 Q1.n14 Q1.n13 1.66898
R29679 Q1.n4 Q1.n3 1.64452
R29680 Q1.n2 Q1.n1 1.19615
R29681 Q1.n3 Q1 0.848156
R29682 Q1.n2 Q1 0.447191
R29683 Q1.n8 Q1 0.39003
R29684 Q1.n9 Q1.n8 0.3624
R29685 Q1.n7 Q1.n6 0.280391
R29686 Q1.n6 Q1.n4 0.262643
R29687 Q1.n4 Q1 0.1255
R29688 Q1.n1 Q1 0.1255
R29689 Q1.n9 Q1 0.0670833
R29690 Q1.n13 Q1 0.063
R29691 Q1.n4 Q1 0.063
R29692 Q1.n10 Q1.n9 0.0428618
R29693 Q1.n12 Q1.n11 0.0305325
R29694 Q1.n10 Q1 0.0194691
R29695 Q1 Q1.n15 0.0168043
R29696 Q1.n15 Q1 0.0122188
R29697 Q1.n1 Q1.n0 0.0107679
R29698 Q1.n0 Q1 0.0107679
R29699 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 169.46
R29700 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 167.809
R29701 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 167.809
R29702 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 167.227
R29703 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 150.293
R29704 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 150.273
R29705 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 73.6406
R29706 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 73.6304
R29707 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 60.3809
R29708 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 12.3891
R29709 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 11.4489
R29710 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 1.38365
R29711 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 1.19615
R29712 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 1.1717
R29713 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 0.848156
R29714 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.447191
R29715 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.38637
R29716 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 0.280391
R29717 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 0.262643
R29718 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.217464
R29719 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.152844
R29720 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.149957
R29721 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.1255
R29722 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.1255
R29723 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 0.0874565
R29724 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.063
R29725 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 0.063
R29726 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 0.063
R29727 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.0454219
R29728 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 0.0107679
R29729 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.0107679
R29730 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 169.46
R29731 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 167.809
R29732 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 167.809
R29733 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 167.226
R29734 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 150.273
R29735 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 150.273
R29736 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 73.6406
R29737 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 73.6304
R29738 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 60.4568
R29739 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 12.3891
R29740 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 11.4489
R29741 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.68257
R29742 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 1.38365
R29743 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 1.19615
R29744 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 1.1717
R29745 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.08448
R29746 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.932141
R29747 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.720633
R29748 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 0.280391
R29749 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.217464
R29750 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R29751 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R29752 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R29753 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 0.0874565
R29754 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 0.063
R29755 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.063
R29756 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 0.063
R29757 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 0.063
R29758 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 0.0435206
R29759 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 0.0216397
R29760 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 0.0216397
R29761 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 0.0107679
R29762 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.0107679
R29763 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 169.46
R29764 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 167.809
R29765 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 167.809
R29766 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 167.227
R29767 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 150.293
R29768 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 150.273
R29769 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 73.6406
R29770 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 73.6304
R29771 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 60.3809
R29772 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 12.3891
R29773 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 11.4489
R29774 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 1.38365
R29775 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 1.19615
R29776 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 1.1717
R29777 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.848156
R29778 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 0.447191
R29779 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.38637
R29780 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 0.280391
R29781 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.217464
R29782 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.200143
R29783 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.152844
R29784 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.149957
R29785 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.1255
R29786 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.1255
R29787 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 0.0874565
R29788 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 0.063
R29789 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 0.063
R29790 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 0.063
R29791 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0454219
R29792 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 0.0107679
R29793 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0107679
R29794 CDAC8_0.switch_1.Z.n4 CDAC8_0.switch_1.Z.t2 168.075
R29795 CDAC8_0.switch_1.Z.n4 CDAC8_0.switch_1.Z.t0 168.075
R29796 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z.t3 60.6851
R29797 CDAC8_0.switch_1.Z CDAC8_0.switch_1.Z.t1 60.6226
R29798 CDAC8_0.switch_1.Z.n2 CDAC8_0.switch_1.Z.t4 14.5332
R29799 CDAC8_0.switch_1.Z.n5 CDAC8_0.switch_1.Z.n3 1.29126
R29800 CDAC8_0.switch_1.Z.n3 CDAC8_0.switch_1.Z 0.478761
R29801 CDAC8_0.switch_1.Z.n1 CDAC8_0.switch_1.Z 0.21925
R29802 CDAC8_0.switch_1.Z.n1 CDAC8_0.switch_1.Z.n0 0.179848
R29803 CDAC8_0.switch_1.Z CDAC8_0.switch_1.Z.n5 0.178175
R29804 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z 0.1255
R29805 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z 0.063
R29806 CDAC8_0.switch_1.Z.n3 CDAC8_0.switch_1.Z.n2 0.063
R29807 CDAC8_0.switch_1.Z.n2 CDAC8_0.switch_1.Z.n1 0.063
R29808 CDAC8_0.switch_1.Z.n5 CDAC8_0.switch_1.Z.n4 0.0130546
R29809 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 169.46
R29810 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 167.809
R29811 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 167.809
R29812 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 167.227
R29813 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 150.293
R29814 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 150.273
R29815 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 73.6406
R29816 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 73.6304
R29817 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 60.3809
R29818 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 12.3891
R29819 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 11.4489
R29820 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 1.38365
R29821 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 1.19615
R29822 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 1.1717
R29823 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 0.848156
R29824 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.447191
R29825 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R29826 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 0.280391
R29827 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.217464
R29828 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 0.200143
R29829 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R29830 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R29831 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R29832 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R29833 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 0.0874565
R29834 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.063
R29835 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 0.063
R29836 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 0.063
R29837 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R29838 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 0.0107679
R29839 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0107679
R29840 Nand_Gate_2.Vout.n10 Nand_Gate_2.Vout.t0 179.256
R29841 Nand_Gate_2.Vout.n10 Nand_Gate_2.Vout.t2 168.089
R29842 Nand_Gate_2.Vout.n2 Nand_Gate_2.Vout.t4 150.293
R29843 Nand_Gate_2.Vout.n4 Nand_Gate_2.Vout.t3 73.6304
R29844 Nand_Gate_2.Vout Nand_Gate_2.Vout.t1 60.3943
R29845 Nand_Gate_2.Vout.n8 Nand_Gate_2.Vout.n7 35.6663
R29846 Nand_Gate_2.Vout.n9 Nand_Gate_2.Vout 0.981478
R29847 Nand_Gate_2.Vout.n11 Nand_Gate_2.Vout.n9 0.788543
R29848 Nand_Gate_2.Vout.n3 Nand_Gate_2.Vout 0.769522
R29849 Nand_Gate_2.Vout Nand_Gate_2.Vout.n11 0.720633
R29850 Nand_Gate_2.Vout.n1 Nand_Gate_2.Vout.n0 0.682565
R29851 Nand_Gate_2.Vout.n1 Nand_Gate_2.Vout 0.580578
R29852 Nand_Gate_2.Vout.n3 Nand_Gate_2.Vout.n2 0.55213
R29853 Nand_Gate_2.Vout.n6 Nand_Gate_2.Vout.n5 0.470609
R29854 Nand_Gate_2.Vout.n2 Nand_Gate_2.Vout 0.447191
R29855 Nand_Gate_2.Vout.n6 Nand_Gate_2.Vout 0.428234
R29856 Nand_Gate_2.Vout.n5 Nand_Gate_2.Vout 0.1255
R29857 Nand_Gate_2.Vout.n0 Nand_Gate_2.Vout 0.1255
R29858 Nand_Gate_2.Vout.n7 Nand_Gate_2.Vout.n3 0.063
R29859 Nand_Gate_2.Vout.n7 Nand_Gate_2.Vout.n6 0.063
R29860 Nand_Gate_2.Vout.n0 Nand_Gate_2.Vout 0.063
R29861 Nand_Gate_2.Vout.n9 Nand_Gate_2.Vout.n8 0.063
R29862 Nand_Gate_2.Vout.n8 Nand_Gate_2.Vout.n1 0.063
R29863 Nand_Gate_2.Vout.n11 Nand_Gate_2.Vout.n10 0.0435206
R29864 Nand_Gate_2.Vout.n5 Nand_Gate_2.Vout.n4 0.0107679
R29865 Nand_Gate_2.Vout.n4 Nand_Gate_2.Vout 0.0107679
R29866 Nand_Gate_3.B.n6 Nand_Gate_3.B.t3 169.46
R29867 Nand_Gate_3.B.n6 Nand_Gate_3.B.t2 167.809
R29868 Nand_Gate_3.B.n5 Nand_Gate_3.B.t1 167.809
R29869 Nand_Gate_3.B Nand_Gate_3.B.t7 158.585
R29870 Nand_Gate_3.B.t7 Nand_Gate_3.B.n2 150.293
R29871 Nand_Gate_3.B.n28 Nand_Gate_3.B.t6 150.273
R29872 Nand_Gate_3.B.n18 Nand_Gate_3.B.t10 150.273
R29873 Nand_Gate_3.B.n12 Nand_Gate_3.B.t5 150.273
R29874 Nand_Gate_3.B.n16 Nand_Gate_3.B.t4 73.6406
R29875 Nand_Gate_3.B.n10 Nand_Gate_3.B.t11 73.6406
R29876 Nand_Gate_3.B.n25 Nand_Gate_3.B.t8 73.6304
R29877 Nand_Gate_3.B.n0 Nand_Gate_3.B.t9 73.6304
R29878 Nand_Gate_3.B.n34 Nand_Gate_3.B.t0 60.3809
R29879 Nand_Gate_3.B.n29 Nand_Gate_3.B.n28 40.8363
R29880 Nand_Gate_3.B.n7 Nand_Gate_3.B.n6 11.4489
R29881 Nand_Gate_3.B.n5 Nand_Gate_3.B.n4 8.21389
R29882 Nand_Gate_3.B.n22 Nand_Gate_3.B.n15 8.1418
R29883 Nand_Gate_3.B.n24 Nand_Gate_3.B.n23 6.47604
R29884 Nand_Gate_3.B.n23 Nand_Gate_3.B 5.35402
R29885 Nand_Gate_3.B.n32 Nand_Gate_3.B 4.55128
R29886 Nand_Gate_3.B.n22 Nand_Gate_3.B.n21 4.5005
R29887 Nand_Gate_3.B.n2 Nand_Gate_3.B.n1 1.19615
R29888 Nand_Gate_3.B.n27 Nand_Gate_3.B.n26 1.1717
R29889 Nand_Gate_3.B.n33 Nand_Gate_3.B 1.08746
R29890 Nand_Gate_3.B.n24 Nand_Gate_3.B 0.973326
R29891 Nand_Gate_3.B.n27 Nand_Gate_3.B 0.932141
R29892 Nand_Gate_3.B.n17 Nand_Gate_3.B 0.851043
R29893 Nand_Gate_3.B.n11 Nand_Gate_3.B 0.851043
R29894 Nand_Gate_3.B Nand_Gate_3.B.n34 0.848156
R29895 Nand_Gate_3.B.n9 Nand_Gate_3.B.n8 0.788543
R29896 Nand_Gate_3.B.n31 Nand_Gate_3.B.n30 0.755935
R29897 Nand_Gate_3.B.n34 Nand_Gate_3.B.n33 0.682565
R29898 Nand_Gate_3.B.n9 Nand_Gate_3.B 0.65675
R29899 Nand_Gate_3.B.n20 Nand_Gate_3.B.n19 0.55213
R29900 Nand_Gate_3.B.n14 Nand_Gate_3.B.n13 0.55213
R29901 Nand_Gate_3.B.n20 Nand_Gate_3.B 0.486828
R29902 Nand_Gate_3.B.n14 Nand_Gate_3.B 0.486828
R29903 Nand_Gate_3.B.n30 Nand_Gate_3.B 0.48023
R29904 Nand_Gate_3.B.n17 Nand_Gate_3.B.n16 0.470609
R29905 Nand_Gate_3.B.n11 Nand_Gate_3.B.n10 0.470609
R29906 Nand_Gate_3.B.n2 Nand_Gate_3.B 0.447191
R29907 Nand_Gate_3.B.n4 Nand_Gate_3.B.n3 0.425067
R29908 Nand_Gate_3.B.n4 Nand_Gate_3.B 0.39003
R29909 Nand_Gate_3.B.n7 Nand_Gate_3.B.n5 0.280391
R29910 Nand_Gate_3.B.n16 Nand_Gate_3.B 0.217464
R29911 Nand_Gate_3.B.n10 Nand_Gate_3.B 0.217464
R29912 Nand_Gate_3.B Nand_Gate_3.B.n7 0.200143
R29913 Nand_Gate_3.B.n26 Nand_Gate_3.B 0.1255
R29914 Nand_Gate_3.B.n19 Nand_Gate_3.B 0.1255
R29915 Nand_Gate_3.B.n13 Nand_Gate_3.B 0.1255
R29916 Nand_Gate_3.B.n1 Nand_Gate_3.B 0.1255
R29917 Nand_Gate_3.B.n8 Nand_Gate_3.B 0.1255
R29918 Nand_Gate_3.B.n28 Nand_Gate_3.B.n27 0.063
R29919 Nand_Gate_3.B.n21 Nand_Gate_3.B.n17 0.063
R29920 Nand_Gate_3.B.n21 Nand_Gate_3.B.n20 0.063
R29921 Nand_Gate_3.B.n15 Nand_Gate_3.B.n11 0.063
R29922 Nand_Gate_3.B.n15 Nand_Gate_3.B.n14 0.063
R29923 Nand_Gate_3.B.n23 Nand_Gate_3.B.n22 0.063
R29924 Nand_Gate_3.B.n29 Nand_Gate_3.B.n24 0.063
R29925 Nand_Gate_3.B.n30 Nand_Gate_3.B.n29 0.063
R29926 Nand_Gate_3.B.n8 Nand_Gate_3.B 0.063
R29927 Nand_Gate_3.B.n33 Nand_Gate_3.B.n32 0.063
R29928 Nand_Gate_3.B.n32 Nand_Gate_3.B.n9 0.063
R29929 Nand_Gate_3.B.n19 Nand_Gate_3.B.n18 0.0216397
R29930 Nand_Gate_3.B.n18 Nand_Gate_3.B 0.0216397
R29931 Nand_Gate_3.B.n13 Nand_Gate_3.B.n12 0.0216397
R29932 Nand_Gate_3.B.n12 Nand_Gate_3.B 0.0216397
R29933 Nand_Gate_3.B.n31 Nand_Gate_3.B 0.0168043
R29934 Nand_Gate_3.B Nand_Gate_3.B.n31 0.0122188
R29935 Nand_Gate_3.B.n26 Nand_Gate_3.B.n25 0.0107679
R29936 Nand_Gate_3.B.n25 Nand_Gate_3.B 0.0107679
R29937 Nand_Gate_3.B.n1 Nand_Gate_3.B.n0 0.0107679
R29938 Nand_Gate_3.B.n0 Nand_Gate_3.B 0.0107679
R29939 Nand_Gate_3.B.n3 Nand_Gate_3.B 0.00441667
R29940 Nand_Gate_3.B.n3 Nand_Gate_3.B 0.00406061
R29941 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 316.762
R29942 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 168.108
R29943 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 150.293
R29944 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 150.273
R29945 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 73.6406
R29946 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 73.6304
R29947 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 60.4568
R29948 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 12.0358
R29949 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 1.19615
R29950 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.981478
R29951 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 0.788543
R29952 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.769522
R29953 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 0.682565
R29954 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.580578
R29955 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 0.55213
R29956 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 0.484875
R29957 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 0.470609
R29958 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.447191
R29959 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.428234
R29960 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.217464
R29961 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R29962 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R29963 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R29964 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 0.063
R29965 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 0.063
R29966 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.063
R29967 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 0.063
R29968 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 0.063
R29969 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 0.0216397
R29970 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.0216397
R29971 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 0.0107679
R29972 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.0107679
R29973 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 169.46
R29974 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 167.809
R29975 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 167.809
R29976 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 167.227
R29977 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 150.293
R29978 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 150.273
R29979 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 73.6406
R29980 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 73.6304
R29981 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 60.3809
R29982 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 12.3891
R29983 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 11.4489
R29984 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 1.38365
R29985 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 1.19615
R29986 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 1.1717
R29987 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.848156
R29988 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 0.447191
R29989 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R29990 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 0.280391
R29991 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.217464
R29992 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.200143
R29993 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R29994 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R29995 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R29996 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R29997 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 0.0874565
R29998 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 0.063
R29999 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 0.063
R30000 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 0.063
R30001 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R30002 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 0.0107679
R30003 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0107679
R30004 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 316.762
R30005 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 168.108
R30006 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 150.293
R30007 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 150.273
R30008 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 73.6406
R30009 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 73.6304
R30010 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 60.3943
R30011 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 12.0358
R30012 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 1.19615
R30013 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.981478
R30014 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 0.788543
R30015 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.769522
R30016 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 0.682565
R30017 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.580578
R30018 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 0.55213
R30019 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 0.484875
R30020 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 0.470609
R30021 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.447191
R30022 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.428234
R30023 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.217464
R30024 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R30025 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R30026 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R30027 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 0.063
R30028 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 0.063
R30029 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.063
R30030 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 0.063
R30031 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 0.063
R30032 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 0.0216397
R30033 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.0216397
R30034 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 0.0107679
R30035 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.0107679
R30036 Nand_Gate_1.B.n51 Nand_Gate_1.B.t1 169.46
R30037 Nand_Gate_1.B.n53 Nand_Gate_1.B.t3 167.809
R30038 Nand_Gate_1.B.n51 Nand_Gate_1.B.t0 167.809
R30039 Nand_Gate_1.B Nand_Gate_1.B.t16 158.585
R30040 Nand_Gate_1.B Nand_Gate_1.B.t9 158.581
R30041 Nand_Gate_1.B.n42 Nand_Gate_1.B.t4 150.293
R30042 Nand_Gate_1.B.t9 Nand_Gate_1.B.n38 150.293
R30043 Nand_Gate_1.B.t16 Nand_Gate_1.B.n2 150.293
R30044 Nand_Gate_1.B.n29 Nand_Gate_1.B.t7 150.273
R30045 Nand_Gate_1.B.n23 Nand_Gate_1.B.t14 150.273
R30046 Nand_Gate_1.B.n14 Nand_Gate_1.B.t11 150.273
R30047 Nand_Gate_1.B.n8 Nand_Gate_1.B.t6 150.273
R30048 Nand_Gate_1.B.n27 Nand_Gate_1.B.t8 73.6406
R30049 Nand_Gate_1.B.n21 Nand_Gate_1.B.t15 73.6406
R30050 Nand_Gate_1.B.n12 Nand_Gate_1.B.t5 73.6406
R30051 Nand_Gate_1.B.n6 Nand_Gate_1.B.t10 73.6406
R30052 Nand_Gate_1.B.n43 Nand_Gate_1.B.t12 73.6304
R30053 Nand_Gate_1.B.n36 Nand_Gate_1.B.t17 73.6304
R30054 Nand_Gate_1.B.n0 Nand_Gate_1.B.t13 73.6304
R30055 Nand_Gate_1.B.n4 Nand_Gate_1.B.t2 60.3809
R30056 Nand_Gate_1.B.n44 Nand_Gate_1.B.n43 34.7148
R30057 Nand_Gate_1.B.n44 Nand_Gate_1.B.n41 32.6611
R30058 Nand_Gate_1.B.n33 Nand_Gate_1.B.n26 15.5222
R30059 Nand_Gate_1.B.n52 Nand_Gate_1.B.n51 11.4489
R30060 Nand_Gate_1.B.n34 Nand_Gate_1.B.n33 8.26552
R30061 Nand_Gate_1.B.n54 Nand_Gate_1.B.n53 8.21389
R30062 Nand_Gate_1.B.n18 Nand_Gate_1.B.n11 8.1418
R30063 Nand_Gate_1.B.n47 Nand_Gate_1.B.n46 5.61191
R30064 Nand_Gate_1.B.n47 Nand_Gate_1.B 5.35402
R30065 Nand_Gate_1.B.n45 Nand_Gate_1.B.n44 4.81893
R30066 Nand_Gate_1.B.n48 Nand_Gate_1.B.n47 4.563
R30067 Nand_Gate_1.B.n33 Nand_Gate_1.B.n32 4.5005
R30068 Nand_Gate_1.B.n18 Nand_Gate_1.B.n17 4.5005
R30069 Nand_Gate_1.B.n46 Nand_Gate_1.B 1.83746
R30070 Nand_Gate_1.B.n20 Nand_Gate_1.B.n19 1.62007
R30071 Nand_Gate_1.B.n38 Nand_Gate_1.B.n37 1.19615
R30072 Nand_Gate_1.B.n2 Nand_Gate_1.B.n1 1.19615
R30073 Nand_Gate_1.B.n43 Nand_Gate_1.B.n42 1.1717
R30074 Nand_Gate_1.B.n5 Nand_Gate_1.B 1.08746
R30075 Nand_Gate_1.B.n20 Nand_Gate_1.B 1.01739
R30076 Nand_Gate_1.B.n13 Nand_Gate_1.B 0.851043
R30077 Nand_Gate_1.B.n7 Nand_Gate_1.B 0.851043
R30078 Nand_Gate_1.B.n4 Nand_Gate_1.B 0.848156
R30079 Nand_Gate_1.B.n28 Nand_Gate_1.B.n27 0.796696
R30080 Nand_Gate_1.B.n22 Nand_Gate_1.B.n21 0.796696
R30081 Nand_Gate_1.B.n50 Nand_Gate_1.B.n49 0.788543
R30082 Nand_Gate_1.B.n34 Nand_Gate_1.B 0.716182
R30083 Nand_Gate_1.B.n5 Nand_Gate_1.B.n4 0.682565
R30084 Nand_Gate_1.B.n49 Nand_Gate_1.B 0.65675
R30085 Nand_Gate_1.B.n16 Nand_Gate_1.B.n15 0.55213
R30086 Nand_Gate_1.B.n10 Nand_Gate_1.B.n9 0.55213
R30087 Nand_Gate_1.B.n28 Nand_Gate_1.B 0.524957
R30088 Nand_Gate_1.B.n22 Nand_Gate_1.B 0.524957
R30089 Nand_Gate_1.B.n35 Nand_Gate_1.B 0.487733
R30090 Nand_Gate_1.B.n16 Nand_Gate_1.B 0.486828
R30091 Nand_Gate_1.B.n10 Nand_Gate_1.B 0.486828
R30092 Nand_Gate_1.B.n13 Nand_Gate_1.B.n12 0.470609
R30093 Nand_Gate_1.B.n7 Nand_Gate_1.B.n6 0.470609
R30094 Nand_Gate_1.B.n42 Nand_Gate_1.B 0.447191
R30095 Nand_Gate_1.B.n38 Nand_Gate_1.B 0.447191
R30096 Nand_Gate_1.B.n2 Nand_Gate_1.B 0.447191
R30097 Nand_Gate_1.B.n54 Nand_Gate_1.B.n3 0.425067
R30098 Nand_Gate_1.B.n40 Nand_Gate_1.B.n39 0.424283
R30099 Nand_Gate_1.B Nand_Gate_1.B.n54 0.39003
R30100 Nand_Gate_1.B.n40 Nand_Gate_1.B 0.338158
R30101 Nand_Gate_1.B.n35 Nand_Gate_1.B.n34 0.300517
R30102 Nand_Gate_1.B.n53 Nand_Gate_1.B.n52 0.280391
R30103 Nand_Gate_1.B.n52 Nand_Gate_1.B.n50 0.262643
R30104 Nand_Gate_1.B.n31 Nand_Gate_1.B 0.252453
R30105 Nand_Gate_1.B.n25 Nand_Gate_1.B 0.252453
R30106 Nand_Gate_1.B.n31 Nand_Gate_1.B.n30 0.226043
R30107 Nand_Gate_1.B.n25 Nand_Gate_1.B.n24 0.226043
R30108 Nand_Gate_1.B.n27 Nand_Gate_1.B 0.217464
R30109 Nand_Gate_1.B.n21 Nand_Gate_1.B 0.217464
R30110 Nand_Gate_1.B.n12 Nand_Gate_1.B 0.217464
R30111 Nand_Gate_1.B.n6 Nand_Gate_1.B 0.217464
R30112 Nand_Gate_1.B.n43 Nand_Gate_1.B 0.149957
R30113 Nand_Gate_1.B.n30 Nand_Gate_1.B 0.1255
R30114 Nand_Gate_1.B.n24 Nand_Gate_1.B 0.1255
R30115 Nand_Gate_1.B.n37 Nand_Gate_1.B 0.1255
R30116 Nand_Gate_1.B.n15 Nand_Gate_1.B 0.1255
R30117 Nand_Gate_1.B.n9 Nand_Gate_1.B 0.1255
R30118 Nand_Gate_1.B.n50 Nand_Gate_1.B 0.1255
R30119 Nand_Gate_1.B.n1 Nand_Gate_1.B 0.1255
R30120 Nand_Gate_1.B.n32 Nand_Gate_1.B.n28 0.063
R30121 Nand_Gate_1.B.n32 Nand_Gate_1.B.n31 0.063
R30122 Nand_Gate_1.B.n26 Nand_Gate_1.B.n22 0.063
R30123 Nand_Gate_1.B.n26 Nand_Gate_1.B.n25 0.063
R30124 Nand_Gate_1.B.n17 Nand_Gate_1.B.n13 0.063
R30125 Nand_Gate_1.B.n17 Nand_Gate_1.B.n16 0.063
R30126 Nand_Gate_1.B.n11 Nand_Gate_1.B.n7 0.063
R30127 Nand_Gate_1.B.n11 Nand_Gate_1.B.n10 0.063
R30128 Nand_Gate_1.B.n46 Nand_Gate_1.B.n45 0.063
R30129 Nand_Gate_1.B.n45 Nand_Gate_1.B.n20 0.063
R30130 Nand_Gate_1.B.n48 Nand_Gate_1.B.n5 0.063
R30131 Nand_Gate_1.B.n49 Nand_Gate_1.B.n48 0.063
R30132 Nand_Gate_1.B.n50 Nand_Gate_1.B 0.063
R30133 Nand_Gate_1.B Nand_Gate_1.B.n18 0.0512812
R30134 Nand_Gate_1.B.n43 Nand_Gate_1.B 0.0454219
R30135 Nand_Gate_1.B.n41 Nand_Gate_1.B.n35 0.024
R30136 Nand_Gate_1.B.n41 Nand_Gate_1.B.n40 0.024
R30137 Nand_Gate_1.B.n30 Nand_Gate_1.B.n29 0.0216397
R30138 Nand_Gate_1.B.n29 Nand_Gate_1.B 0.0216397
R30139 Nand_Gate_1.B.n24 Nand_Gate_1.B.n23 0.0216397
R30140 Nand_Gate_1.B.n23 Nand_Gate_1.B 0.0216397
R30141 Nand_Gate_1.B.n15 Nand_Gate_1.B.n14 0.0216397
R30142 Nand_Gate_1.B.n14 Nand_Gate_1.B 0.0216397
R30143 Nand_Gate_1.B.n9 Nand_Gate_1.B.n8 0.0216397
R30144 Nand_Gate_1.B.n8 Nand_Gate_1.B 0.0216397
R30145 Nand_Gate_1.B.n19 Nand_Gate_1.B 0.0168043
R30146 Nand_Gate_1.B.n19 Nand_Gate_1.B 0.0122188
R30147 Nand_Gate_1.B.n37 Nand_Gate_1.B.n36 0.0107679
R30148 Nand_Gate_1.B.n36 Nand_Gate_1.B 0.0107679
R30149 Nand_Gate_1.B.n1 Nand_Gate_1.B.n0 0.0107679
R30150 Nand_Gate_1.B.n0 Nand_Gate_1.B 0.0107679
R30151 Nand_Gate_1.B.n39 Nand_Gate_1.B 0.00441667
R30152 Nand_Gate_1.B.n3 Nand_Gate_1.B 0.00441667
R30153 Nand_Gate_1.B.n39 Nand_Gate_1.B 0.00406061
R30154 Nand_Gate_1.B.n3 Nand_Gate_1.B 0.00406061
R30155 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 169.46
R30156 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 168.089
R30157 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 167.809
R30158 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 150.293
R30159 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 73.6304
R30160 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 60.3943
R30161 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 12.0358
R30162 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 11.4489
R30163 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.981478
R30164 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 0.788543
R30165 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.769522
R30166 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 0.720633
R30167 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 0.682565
R30168 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.580578
R30169 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 0.55213
R30170 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 0.470609
R30171 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.447191
R30172 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.428234
R30173 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.1255
R30174 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.1255
R30175 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 0.063
R30176 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 0.063
R30177 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.063
R30178 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 0.063
R30179 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 0.063
R30180 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 0.0435206
R30181 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 0.0107679
R30182 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.0107679
R30183 Q7.n2 Q7.t2 169.46
R30184 Q7.n4 Q7.t0 167.809
R30185 Q7.n2 Q7.t3 167.809
R30186 Q7 Q7.t6 158.585
R30187 Q7 Q7.t9 154.823
R30188 Q7.n14 Q7.t4 150.869
R30189 Q7.t9 Q7.n15 150.869
R30190 Q7.t6 Q7.n9 150.293
R30191 Q7.n16 Q7.n13 137.644
R30192 Q7.n13 Q7 85.5731
R30193 Q7.n15 Q7.t7 74.1352
R30194 Q7.n14 Q7.t8 74.1352
R30195 Q7.n7 Q7.t5 73.6304
R30196 Q7.n0 Q7.t1 60.3809
R30197 Q7.n3 Q7.n2 11.4489
R30198 Q7.n5 Q7.n4 8.21389
R30199 Q7.n13 Q7.n12 3.473
R30200 Q7.n15 Q7.n14 1.66898
R30201 Q7.n1 Q7.n0 1.64452
R30202 Q7.n9 Q7.n8 1.19615
R30203 Q7.n0 Q7 0.848156
R30204 Q7.n9 Q7 0.447191
R30205 Q7.n5 Q7 0.39003
R30206 Q7.n4 Q7.n3 0.280391
R30207 Q7.n3 Q7.n1 0.262643
R30208 Q7.n6 Q7.n5 0.224533
R30209 Q7.n6 Q7 0.20495
R30210 Q7.n11 Q7.n10 0.149333
R30211 Q7.n11 Q7 0.139364
R30212 Q7.n1 Q7 0.1255
R30213 Q7.n8 Q7 0.1255
R30214 Q7.n14 Q7 0.063
R30215 Q7.n1 Q7 0.063
R30216 Q7.n12 Q7.n6 0.024
R30217 Q7.n12 Q7.n11 0.024
R30218 Q7 Q7.n16 0.0168043
R30219 Q7.n16 Q7 0.0122188
R30220 Q7.n8 Q7.n7 0.0107679
R30221 Q7.n7 Q7 0.0107679
R30222 Q7.n10 Q7 0.00441667
R30223 Q7.n10 Q7 0.00406061
R30224 And_Gate_5.Vout.n15 And_Gate_5.Vout.t0 168.108
R30225 And_Gate_5.Vout.n5 And_Gate_5.Vout.t6 158.207
R30226 D_FlipFlop_1.CLK And_Gate_5.Vout.t2 158.202
R30227 And_Gate_5.Vout.n7 And_Gate_5.Vout.t7 150.293
R30228 And_Gate_5.Vout.t2 And_Gate_5.Vout.n10 150.293
R30229 And_Gate_5.Vout.t6 And_Gate_5.Vout.n4 150.273
R30230 And_Gate_5.Vout.n13 And_Gate_5.Vout.n12 89.3276
R30231 And_Gate_5.Vout.n2 And_Gate_5.Vout.t3 73.6406
R30232 And_Gate_5.Vout.n9 And_Gate_5.Vout.t5 73.6304
R30233 And_Gate_5.Vout.n8 And_Gate_5.Vout.t4 73.6304
R30234 And_Gate_5.Inverter_0.Vout And_Gate_5.Vout.t1 60.3943
R30235 And_Gate_5.Vout.n9 And_Gate_5.Vout.n8 16.332
R30236 And_Gate_5.Vout.n3 And_Gate_5.Vout.n2 1.19615
R30237 And_Gate_5.Vout.n8 And_Gate_5.Vout.n7 1.1717
R30238 And_Gate_5.Vout.n10 And_Gate_5.Vout.n9 1.1717
R30239 And_Gate_5.Vout.n14 And_Gate_5.Inverter_0.Vout 0.981478
R30240 And_Gate_5.Vout.n15 And_Gate_5.Vout.n14 0.788543
R30241 And_Gate_5.Vout.n1 And_Gate_5.Vout.n0 0.682565
R30242 And_Gate_5.Vout.n1 And_Gate_5.Inverter_0.Vout 0.580578
R30243 And_Gate_5.Inverter_0.Vout And_Gate_5.Vout.n15 0.484875
R30244 And_Gate_5.Vout.n10 D_FlipFlop_1.3-input-nand_1.C 0.447191
R30245 And_Gate_5.Vout.n7 D_FlipFlop_1.Inverter_1.Vin 0.436162
R30246 And_Gate_5.Vout.n5 D_FlipFlop_1.CLK 0.321667
R30247 And_Gate_5.Vout.n6 And_Gate_5.Vout.n5 0.283283
R30248 And_Gate_5.Vout.n2 D_FlipFlop_1.3-input-nand_0.C 0.217464
R30249 And_Gate_5.Vout.n9 D_FlipFlop_1.3-input-nand_1.C 0.149957
R30250 And_Gate_5.Vout.n3 D_FlipFlop_1.3-input-nand_0.C 0.1255
R30251 And_Gate_5.Vout.n0 And_Gate_5.Inverter_0.Vout 0.1255
R30252 And_Gate_5.Vout.n8 D_FlipFlop_1.Inverter_1.Vin 0.117348
R30253 And_Gate_5.Vout.n6 D_FlipFlop_1.CLK 0.071
R30254 And_Gate_5.Vout.n0 And_Gate_5.Inverter_0.Vout 0.063
R30255 And_Gate_5.Vout.n14 And_Gate_5.Vout.n13 0.063
R30256 And_Gate_5.Vout.n13 And_Gate_5.Vout.n1 0.063
R30257 And_Gate_5.Vout.n8 D_FlipFlop_1.Inverter_1.Vin 0.0454219
R30258 And_Gate_5.Vout.n9 D_FlipFlop_1.3-input-nand_1.C 0.0454219
R30259 And_Gate_5.Vout.n12 And_Gate_5.Vout.n6 0.024
R30260 And_Gate_5.Vout.n12 And_Gate_5.Vout.n11 0.024
R30261 And_Gate_5.Vout.n4 And_Gate_5.Vout.n3 0.0216397
R30262 And_Gate_5.Vout.n4 D_FlipFlop_1.3-input-nand_0.C 0.0216397
R30263 And_Gate_5.Vout.n11 D_FlipFlop_1.CLK 0.0104697
R30264 And_Gate_5.Vout.n11 D_FlipFlop_1.CLK 0.0091579
R30265 Q5.n2 Q5.t1 169.46
R30266 Q5.n4 Q5.t3 167.809
R30267 Q5.n2 Q5.t0 167.809
R30268 Q5 Q5.t9 158.585
R30269 Q5 Q5.t4 154.823
R30270 Q5.n14 Q5.t5 150.869
R30271 Q5.t4 Q5.n15 150.869
R30272 Q5.t9 Q5.n9 150.293
R30273 Q5.n16 Q5.n13 137.644
R30274 Q5.n13 Q5 85.5731
R30275 Q5.n15 Q5.t6 74.1352
R30276 Q5.n14 Q5.t7 74.1352
R30277 Q5.n7 Q5.t8 73.6304
R30278 Q5.n0 Q5.t2 60.3809
R30279 Q5.n3 Q5.n2 11.4489
R30280 Q5.n5 Q5.n4 8.21389
R30281 Q5.n13 Q5.n12 3.473
R30282 Q5.n15 Q5.n14 1.66898
R30283 Q5.n1 Q5.n0 1.64452
R30284 Q5.n9 Q5.n8 1.19615
R30285 Q5.n0 Q5 0.848156
R30286 Q5.n9 Q5 0.447191
R30287 Q5.n5 Q5 0.39003
R30288 Q5.n4 Q5.n3 0.280391
R30289 Q5.n3 Q5.n1 0.262643
R30290 Q5.n6 Q5 0.222967
R30291 Q5.n6 Q5.n5 0.206517
R30292 Q5.n11 Q5.n10 0.16735
R30293 Q5.n11 Q5 0.155742
R30294 Q5.n1 Q5 0.1255
R30295 Q5.n8 Q5 0.1255
R30296 Q5.n14 Q5 0.063
R30297 Q5.n1 Q5 0.063
R30298 Q5.n12 Q5.n6 0.024
R30299 Q5.n12 Q5.n11 0.024
R30300 Q5 Q5.n16 0.0168043
R30301 Q5.n16 Q5 0.0122188
R30302 Q5.n8 Q5.n7 0.0107679
R30303 Q5.n7 Q5 0.0107679
R30304 Q5.n10 Q5 0.00441667
R30305 Q5.n10 Q5 0.00406061
R30306 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t1 169.46
R30307 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.t3 167.809
R30308 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t0 167.809
R30309 D_FlipFlop_7.3-input-nand_2.C.t4 D_FlipFlop_7.3-input-nand_2.C.n13 167.226
R30310 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C.t5 150.273
R30311 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.t4 150.273
R30312 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C.t7 73.6406
R30313 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C.t6 73.6304
R30314 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C.t2 60.4568
R30315 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C.n7 12.3891
R30316 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.n11 11.4489
R30317 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C 1.68257
R30318 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C.n2 1.38365
R30319 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C.n0 1.19615
R30320 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C.n5 1.1717
R30321 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C 1.08448
R30322 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C 0.932141
R30323 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C 0.720633
R30324 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.n12 0.280391
R30325 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C 0.217464
R30326 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30327 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30328 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30329 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C.n9 0.0874565
R30330 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C.n6 0.063
R30331 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C 0.063
R30332 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C.n8 0.063
R30333 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C.n3 0.063
R30334 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.n10 0.0435206
R30335 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.n1 0.0216397
R30336 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.C.n14 0.0216397
R30337 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C.n4 0.0107679
R30338 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C 0.0107679
R30339 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t3 169.46
R30340 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.t2 167.809
R30341 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t0 167.809
R30342 D_FlipFlop_7.3-input-nand_2.Vout.t6 D_FlipFlop_7.3-input-nand_2.Vout.n11 167.227
R30343 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.t6 150.293
R30344 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.t5 150.273
R30345 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout.t7 73.6406
R30346 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout.t4 73.6304
R30347 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout.t1 60.3809
R30348 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n5 12.3891
R30349 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout.n9 11.4489
R30350 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout.n2 1.38365
R30351 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.n1 1.19615
R30352 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.n4 1.1717
R30353 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout 0.848156
R30354 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.Vout.n12 0.447191
R30355 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R30356 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.n10 0.280391
R30357 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout.n8 0.262643
R30358 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout 0.217464
R30359 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R30360 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R30361 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R30362 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R30363 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout.n7 0.0874565
R30364 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n3 0.063
R30365 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout.n6 0.063
R30366 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout 0.063
R30367 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R30368 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout.n0 0.0107679
R30369 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout 0.0107679
R30370 Nand_Gate_1.Vout.n10 Nand_Gate_1.Vout.t2 179.256
R30371 Nand_Gate_1.Vout.n10 Nand_Gate_1.Vout.t0 168.089
R30372 Nand_Gate_1.Vout.n2 Nand_Gate_1.Vout.t4 150.293
R30373 Nand_Gate_1.Vout.n4 Nand_Gate_1.Vout.t3 73.6304
R30374 Nand_Gate_1.Vout Nand_Gate_1.Vout.t1 60.3943
R30375 Nand_Gate_1.Vout.n8 Nand_Gate_1.Vout.n7 37.3347
R30376 Nand_Gate_1.Vout.n9 Nand_Gate_1.Vout 0.981478
R30377 Nand_Gate_1.Vout.n11 Nand_Gate_1.Vout.n9 0.788543
R30378 Nand_Gate_1.Vout.n3 Nand_Gate_1.Vout 0.769522
R30379 Nand_Gate_1.Vout Nand_Gate_1.Vout.n11 0.720633
R30380 Nand_Gate_1.Vout.n1 Nand_Gate_1.Vout.n0 0.682565
R30381 Nand_Gate_1.Vout.n1 Nand_Gate_1.Vout 0.580578
R30382 Nand_Gate_1.Vout.n3 Nand_Gate_1.Vout.n2 0.55213
R30383 Nand_Gate_1.Vout.n6 Nand_Gate_1.Vout.n5 0.470609
R30384 Nand_Gate_1.Vout.n2 Nand_Gate_1.Vout 0.447191
R30385 Nand_Gate_1.Vout.n6 Nand_Gate_1.Vout 0.428234
R30386 Nand_Gate_1.Vout.n5 Nand_Gate_1.Vout 0.1255
R30387 Nand_Gate_1.Vout.n0 Nand_Gate_1.Vout 0.1255
R30388 Nand_Gate_1.Vout.n7 Nand_Gate_1.Vout.n3 0.063
R30389 Nand_Gate_1.Vout.n7 Nand_Gate_1.Vout.n6 0.063
R30390 Nand_Gate_1.Vout.n0 Nand_Gate_1.Vout 0.063
R30391 Nand_Gate_1.Vout.n9 Nand_Gate_1.Vout.n8 0.063
R30392 Nand_Gate_1.Vout.n8 Nand_Gate_1.Vout.n1 0.063
R30393 Nand_Gate_1.Vout.n11 Nand_Gate_1.Vout.n10 0.0435206
R30394 Nand_Gate_1.Vout.n5 Nand_Gate_1.Vout.n4 0.0107679
R30395 Nand_Gate_1.Vout.n4 Nand_Gate_1.Vout 0.0107679
R30396 Nand_Gate_7.A.n32 Nand_Gate_7.A.t0 169.46
R30397 Nand_Gate_7.A.n32 Nand_Gate_7.A.t3 167.809
R30398 Nand_Gate_7.A.n34 Nand_Gate_7.A.t2 167.809
R30399 Nand_Gate_7.A Nand_Gate_7.A.t6 158.585
R30400 Nand_Gate_7.A.n20 Nand_Gate_7.A.t9 150.293
R30401 Nand_Gate_7.A.t6 Nand_Gate_7.A.n2 150.293
R30402 Nand_Gate_7.A.n14 Nand_Gate_7.A.t8 150.273
R30403 Nand_Gate_7.A.n8 Nand_Gate_7.A.t5 150.273
R30404 Nand_Gate_7.A.n12 Nand_Gate_7.A.t4 73.6406
R30405 Nand_Gate_7.A.n6 Nand_Gate_7.A.t7 73.6406
R30406 Nand_Gate_7.A.n22 Nand_Gate_7.A.t11 73.6304
R30407 Nand_Gate_7.A.n0 Nand_Gate_7.A.t10 73.6304
R30408 Nand_Gate_7.A.n4 Nand_Gate_7.A.t1 60.3809
R30409 Nand_Gate_7.A.n26 Nand_Gate_7.A.n25 14.3097
R30410 Nand_Gate_7.A.n33 Nand_Gate_7.A.n32 11.4489
R30411 Nand_Gate_7.A.n35 Nand_Gate_7.A.n34 8.21389
R30412 Nand_Gate_7.A.n18 Nand_Gate_7.A.n11 8.1418
R30413 Nand_Gate_7.A.n28 Nand_Gate_7.A.n27 5.61191
R30414 Nand_Gate_7.A.n28 Nand_Gate_7.A 5.3423
R30415 Nand_Gate_7.A.n29 Nand_Gate_7.A.n28 4.563
R30416 Nand_Gate_7.A.n18 Nand_Gate_7.A.n17 4.5005
R30417 Nand_Gate_7.A.n27 Nand_Gate_7.A 1.82115
R30418 Nand_Gate_7.A.n19 Nand_Gate_7.A 1.62007
R30419 Nand_Gate_7.A.n2 Nand_Gate_7.A.n1 1.19615
R30420 Nand_Gate_7.A.n5 Nand_Gate_7.A 1.08746
R30421 Nand_Gate_7.A.n19 Nand_Gate_7.A 1.00726
R30422 Nand_Gate_7.A.n13 Nand_Gate_7.A 0.851043
R30423 Nand_Gate_7.A.n7 Nand_Gate_7.A 0.851043
R30424 Nand_Gate_7.A.n4 Nand_Gate_7.A 0.848156
R30425 Nand_Gate_7.A.n31 Nand_Gate_7.A.n30 0.788543
R30426 Nand_Gate_7.A.n21 Nand_Gate_7.A 0.769522
R30427 Nand_Gate_7.A.n5 Nand_Gate_7.A.n4 0.682565
R30428 Nand_Gate_7.A.n30 Nand_Gate_7.A 0.65675
R30429 Nand_Gate_7.A.n21 Nand_Gate_7.A.n20 0.55213
R30430 Nand_Gate_7.A.n16 Nand_Gate_7.A.n15 0.55213
R30431 Nand_Gate_7.A.n10 Nand_Gate_7.A.n9 0.55213
R30432 Nand_Gate_7.A.n16 Nand_Gate_7.A 0.486828
R30433 Nand_Gate_7.A.n10 Nand_Gate_7.A 0.486828
R30434 Nand_Gate_7.A.n24 Nand_Gate_7.A.n23 0.470609
R30435 Nand_Gate_7.A.n13 Nand_Gate_7.A.n12 0.470609
R30436 Nand_Gate_7.A.n7 Nand_Gate_7.A.n6 0.470609
R30437 Nand_Gate_7.A.n20 Nand_Gate_7.A 0.447191
R30438 Nand_Gate_7.A.n2 Nand_Gate_7.A 0.447191
R30439 Nand_Gate_7.A.n24 Nand_Gate_7.A 0.428234
R30440 Nand_Gate_7.A.n35 Nand_Gate_7.A.n3 0.425067
R30441 Nand_Gate_7.A Nand_Gate_7.A.n35 0.39003
R30442 Nand_Gate_7.A.n34 Nand_Gate_7.A.n33 0.280391
R30443 Nand_Gate_7.A.n33 Nand_Gate_7.A.n31 0.262643
R30444 Nand_Gate_7.A.n12 Nand_Gate_7.A 0.217464
R30445 Nand_Gate_7.A.n6 Nand_Gate_7.A 0.217464
R30446 Nand_Gate_7.A.n23 Nand_Gate_7.A 0.1255
R30447 Nand_Gate_7.A.n15 Nand_Gate_7.A 0.1255
R30448 Nand_Gate_7.A.n9 Nand_Gate_7.A 0.1255
R30449 Nand_Gate_7.A.n31 Nand_Gate_7.A 0.1255
R30450 Nand_Gate_7.A.n1 Nand_Gate_7.A 0.1255
R30451 Nand_Gate_7.A.n25 Nand_Gate_7.A.n21 0.063
R30452 Nand_Gate_7.A.n25 Nand_Gate_7.A.n24 0.063
R30453 Nand_Gate_7.A.n17 Nand_Gate_7.A.n13 0.063
R30454 Nand_Gate_7.A.n17 Nand_Gate_7.A.n16 0.063
R30455 Nand_Gate_7.A.n11 Nand_Gate_7.A.n7 0.063
R30456 Nand_Gate_7.A.n11 Nand_Gate_7.A.n10 0.063
R30457 Nand_Gate_7.A Nand_Gate_7.A.n18 0.063
R30458 Nand_Gate_7.A.n27 Nand_Gate_7.A.n26 0.063
R30459 Nand_Gate_7.A.n26 Nand_Gate_7.A.n19 0.063
R30460 Nand_Gate_7.A.n29 Nand_Gate_7.A.n5 0.063
R30461 Nand_Gate_7.A.n30 Nand_Gate_7.A.n29 0.063
R30462 Nand_Gate_7.A.n31 Nand_Gate_7.A 0.063
R30463 Nand_Gate_7.A.n15 Nand_Gate_7.A.n14 0.0216397
R30464 Nand_Gate_7.A.n14 Nand_Gate_7.A 0.0216397
R30465 Nand_Gate_7.A.n9 Nand_Gate_7.A.n8 0.0216397
R30466 Nand_Gate_7.A.n8 Nand_Gate_7.A 0.0216397
R30467 Nand_Gate_7.A.n23 Nand_Gate_7.A.n22 0.0107679
R30468 Nand_Gate_7.A.n22 Nand_Gate_7.A 0.0107679
R30469 Nand_Gate_7.A.n1 Nand_Gate_7.A.n0 0.0107679
R30470 Nand_Gate_7.A.n0 Nand_Gate_7.A 0.0107679
R30471 Nand_Gate_7.A.n3 Nand_Gate_7.A 0.00441667
R30472 Nand_Gate_7.A.n3 Nand_Gate_7.A 0.00406061
R30473 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout.t3 169.46
R30474 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout.t2 167.809
R30475 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout.t1 167.809
R30476 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout.t6 167.227
R30477 D_FlipFlop_5.3-input-nand_2.Vout.t6 D_FlipFlop_5.3-input-nand_2.Vout.n2 150.293
R30478 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.t5 150.273
R30479 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout.t7 73.6406
R30480 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout.t4 73.6304
R30481 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.t0 60.3809
R30482 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n9 12.3891
R30483 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.n4 11.4489
R30484 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.n11 1.38365
R30485 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout.n1 1.19615
R30486 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.n8 1.1717
R30487 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.Vout.n12 0.848156
R30488 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout 0.447191
R30489 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R30490 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.n3 0.280391
R30491 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout.n5 0.262643
R30492 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout 0.217464
R30493 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R30494 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R30495 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R30496 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R30497 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout.n6 0.0874565
R30498 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout 0.063
R30499 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout.n10 0.063
R30500 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n7 0.063
R30501 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R30502 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout.n0 0.0107679
R30503 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout 0.0107679
R30504 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 169.46
R30505 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 168.089
R30506 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 167.809
R30507 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 150.293
R30508 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 73.6304
R30509 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 60.4568
R30510 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 12.0358
R30511 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 11.4489
R30512 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.981478
R30513 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 0.788543
R30514 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.769522
R30515 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 0.720633
R30516 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 0.682565
R30517 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.580578
R30518 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 0.55213
R30519 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 0.470609
R30520 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.447191
R30521 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.428234
R30522 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.1255
R30523 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.1255
R30524 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 0.063
R30525 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 0.063
R30526 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.063
R30527 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 0.063
R30528 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 0.063
R30529 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 0.0435206
R30530 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 0.0107679
R30531 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.0107679
R30532 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 169.46
R30533 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 167.809
R30534 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 167.809
R30535 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 167.227
R30536 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 150.293
R30537 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 150.273
R30538 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 73.6406
R30539 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 73.6304
R30540 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 60.3809
R30541 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 12.3891
R30542 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 11.4489
R30543 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 1.38365
R30544 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 1.19615
R30545 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 1.1717
R30546 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.848156
R30547 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 0.447191
R30548 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.38637
R30549 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 0.280391
R30550 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 0.262643
R30551 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.217464
R30552 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.152844
R30553 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.149957
R30554 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.1255
R30555 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.1255
R30556 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 0.0874565
R30557 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 0.063
R30558 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 0.063
R30559 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.063
R30560 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.0454219
R30561 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 0.0107679
R30562 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.0107679
R30563 And_Gate_2.Vout.n12 And_Gate_2.Vout.t0 168.32
R30564 And_Gate_2.Vout.n4 And_Gate_2.Vout.t4 158.23
R30565 D_FlipFlop_5.CLK And_Gate_2.Vout.t6 158.202
R30566 And_Gate_2.Vout.n5 And_Gate_2.Vout.t5 150.293
R30567 And_Gate_2.Vout.t6 And_Gate_2.Vout.n8 150.293
R30568 And_Gate_2.Vout.t4 And_Gate_2.Vout.n3 150.273
R30569 And_Gate_2.Vout.n1 And_Gate_2.Vout.t7 73.6406
R30570 And_Gate_2.Vout.n7 And_Gate_2.Vout.t3 73.6304
R30571 And_Gate_2.Vout.n6 And_Gate_2.Vout.t2 73.6304
R30572 And_Gate_2.Inverter_0.Vout And_Gate_2.Vout.t1 60.3943
R30573 And_Gate_2.Vout.n12 And_Gate_2.Vout.n11 52.2702
R30574 And_Gate_2.Vout.n7 And_Gate_2.Vout.n6 16.332
R30575 And_Gate_2.Vout.n13 And_Gate_2.Vout.n0 1.62007
R30576 And_Gate_2.Inverter_0.Vout And_Gate_2.Vout.n13 1.25441
R30577 And_Gate_2.Vout.n2 And_Gate_2.Vout.n1 1.19615
R30578 And_Gate_2.Vout.n6 And_Gate_2.Vout.n5 1.1717
R30579 And_Gate_2.Vout.n8 And_Gate_2.Vout.n7 1.1717
R30580 And_Gate_2.Vout.n8 D_FlipFlop_5.3-input-nand_1.C 0.447191
R30581 And_Gate_2.Vout.n5 D_FlipFlop_5.Inverter_1.Vin 0.436162
R30582 And_Gate_2.Vout.n4 D_FlipFlop_5.CLK 0.298879
R30583 And_Gate_2.Vout.n10 And_Gate_2.Vout.n9 0.265267
R30584 And_Gate_2.Vout.n1 D_FlipFlop_5.3-input-nand_0.C 0.217464
R30585 And_Gate_2.Vout.n10 D_FlipFlop_5.CLK 0.212618
R30586 And_Gate_2.Vout.n7 D_FlipFlop_5.3-input-nand_1.C 0.149957
R30587 And_Gate_2.Vout.n2 D_FlipFlop_5.3-input-nand_0.C 0.1255
R30588 And_Gate_2.Vout.n0 And_Gate_2.Inverter_0.Vout 0.1255
R30589 And_Gate_2.Vout.n6 D_FlipFlop_5.Inverter_1.Vin 0.117348
R30590 And_Gate_2.Vout.n0 And_Gate_2.Inverter_0.Vout 0.063
R30591 And_Gate_2.Vout.n13 And_Gate_2.Vout.n12 0.063
R30592 And_Gate_2.Vout.n6 D_FlipFlop_5.Inverter_1.Vin 0.0454219
R30593 And_Gate_2.Vout.n7 D_FlipFlop_5.3-input-nand_1.C 0.0454219
R30594 And_Gate_2.Vout.n11 And_Gate_2.Vout.n4 0.024
R30595 And_Gate_2.Vout.n11 And_Gate_2.Vout.n10 0.024
R30596 And_Gate_2.Vout.n3 And_Gate_2.Vout.n2 0.0216397
R30597 And_Gate_2.Vout.n3 D_FlipFlop_5.3-input-nand_0.C 0.0216397
R30598 And_Gate_2.Vout.n9 D_FlipFlop_5.CLK 0.00441667
R30599 And_Gate_2.Vout.n9 D_FlipFlop_5.CLK 0.00406061
R30600 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 169.46
R30601 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 168.089
R30602 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 167.809
R30603 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 150.293
R30604 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 73.6304
R30605 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 60.3943
R30606 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 12.0358
R30607 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 11.4489
R30608 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.981478
R30609 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 0.788543
R30610 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.769522
R30611 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 0.720633
R30612 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 0.682565
R30613 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.580578
R30614 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 0.55213
R30615 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 0.470609
R30616 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.447191
R30617 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.428234
R30618 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.1255
R30619 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.1255
R30620 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 0.063
R30621 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 0.063
R30622 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.063
R30623 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 0.063
R30624 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 0.063
R30625 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 0.0435206
R30626 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 0.0107679
R30627 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.0107679
R30628 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 169.46
R30629 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 168.089
R30630 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 167.809
R30631 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 150.293
R30632 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 73.6304
R30633 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 60.4568
R30634 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 12.0358
R30635 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 11.4489
R30636 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.981478
R30637 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 0.788543
R30638 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.769522
R30639 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 0.720633
R30640 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 0.682565
R30641 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.580578
R30642 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 0.55213
R30643 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 0.470609
R30644 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.447191
R30645 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.428234
R30646 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.1255
R30647 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.1255
R30648 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 0.063
R30649 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 0.063
R30650 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.063
R30651 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 0.063
R30652 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 0.063
R30653 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 0.0435206
R30654 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 0.0107679
R30655 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.0107679
R30656 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 169.46
R30657 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 167.809
R30658 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 167.809
R30659 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 167.226
R30660 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 150.273
R30661 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 150.273
R30662 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 73.6406
R30663 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 73.6304
R30664 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 60.3943
R30665 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 12.3891
R30666 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 11.4489
R30667 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 1.68257
R30668 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 1.38365
R30669 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 1.19615
R30670 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 1.1717
R30671 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 1.08448
R30672 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.932141
R30673 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 0.720633
R30674 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 0.280391
R30675 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.217464
R30676 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R30677 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R30678 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R30679 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 0.0874565
R30680 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 0.063
R30681 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.063
R30682 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 0.063
R30683 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 0.063
R30684 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 0.0435206
R30685 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 0.0216397
R30686 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.0216397
R30687 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 0.0107679
R30688 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.0107679
R30689 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 179.256
R30690 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 168.089
R30691 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 150.293
R30692 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 73.6304
R30693 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 60.3943
R30694 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 12.0358
R30695 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.981478
R30696 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 0.788543
R30697 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.769522
R30698 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 0.720633
R30699 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 0.682565
R30700 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.580578
R30701 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 0.55213
R30702 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 0.470609
R30703 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.447191
R30704 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.428234
R30705 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1255
R30706 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1255
R30707 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 0.063
R30708 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 0.063
R30709 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.063
R30710 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 0.063
R30711 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 0.063
R30712 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 0.0435206
R30713 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 0.0107679
R30714 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.0107679
R30715 And_Gate_4.A.n0 And_Gate_4.A.t2 179.256
R30716 And_Gate_4.A.n0 And_Gate_4.A.t1 168.089
R30717 And_Gate_4.A.n3 And_Gate_4.A.t3 150.293
R30718 And_Gate_4.A.n5 And_Gate_4.A.t4 73.6304
R30719 Nand_Gate_0.Vout And_Gate_4.A.t0 60.3943
R30720 And_Gate_4.A.n9 And_Gate_4.A.n8 35.6663
R30721 And_Gate_4.A.n2 Nand_Gate_0.Vout 0.981478
R30722 And_Gate_4.A.n2 And_Gate_4.A.n1 0.788543
R30723 And_Gate_4.A.n4 And_Gate_4.Nand_Gate_0.A 0.769522
R30724 And_Gate_4.A.n1 Nand_Gate_0.Vout 0.720633
R30725 And_Gate_4.A.n11 And_Gate_4.A.n10 0.682565
R30726 And_Gate_4.A.n10 Nand_Gate_0.Vout 0.580578
R30727 And_Gate_4.A.n4 And_Gate_4.A.n3 0.55213
R30728 And_Gate_4.A.n7 And_Gate_4.A.n6 0.470609
R30729 And_Gate_4.A.n3 And_Gate_4.Nand_Gate_0.A 0.447191
R30730 And_Gate_4.A.n7 And_Gate_4.Nand_Gate_0.A 0.428234
R30731 And_Gate_4.A.n6 And_Gate_4.Nand_Gate_0.A 0.1255
R30732 And_Gate_4.A.n11 Nand_Gate_0.Vout 0.1255
R30733 And_Gate_4.A.n8 And_Gate_4.A.n4 0.063
R30734 And_Gate_4.A.n8 And_Gate_4.A.n7 0.063
R30735 And_Gate_4.A.n9 And_Gate_4.A.n2 0.063
R30736 And_Gate_4.A.n10 And_Gate_4.A.n9 0.063
R30737 Nand_Gate_0.Vout And_Gate_4.A.n11 0.063
R30738 And_Gate_4.A.n1 And_Gate_4.A.n0 0.0435206
R30739 And_Gate_4.A.n6 And_Gate_4.A.n5 0.0107679
R30740 And_Gate_4.A.n5 And_Gate_4.Nand_Gate_0.A 0.0107679
R30741 Q2.n5 Q2.t3 169.46
R30742 Q2.n7 Q2.t0 167.809
R30743 Q2.n5 Q2.t2 167.809
R30744 Q2.n11 Q2.t8 155.121
R30745 Q2.n14 Q2.t4 150.869
R30746 Q2.n13 Q2.t5 150.869
R30747 Q2.t8 Q2.n2 150.293
R30748 Q2.n15 Q2.n12 137.644
R30749 Q2 Q2.t6 78.1811
R30750 Q2.n13 Q2.t7 74.1352
R30751 Q2.t6 Q2.n14 74.1352
R30752 Q2.n0 Q2.t9 73.6304
R30753 Q2.n3 Q2.t1 60.3809
R30754 Q2.n12 Q2 38.8494
R30755 Q2.n6 Q2.n5 11.4489
R30756 Q2.n8 Q2.n7 8.21389
R30757 Q2.n11 Q2.n10 1.70018
R30758 Q2.n14 Q2.n13 1.66898
R30759 Q2.n4 Q2.n3 1.64452
R30760 Q2.n2 Q2.n1 1.19615
R30761 Q2.n3 Q2 0.848156
R30762 Q2.n2 Q2 0.447191
R30763 Q2.n8 Q2 0.39003
R30764 Q2.n9 Q2.n8 0.35535
R30765 Q2.n7 Q2.n6 0.280391
R30766 Q2.n6 Q2.n4 0.262643
R30767 Q2.n4 Q2 0.1255
R30768 Q2.n1 Q2 0.1255
R30769 Q2.n9 Q2 0.0741333
R30770 Q2.n13 Q2 0.063
R30771 Q2.n4 Q2 0.063
R30772 Q2.n10 Q2.n9 0.0460197
R30773 Q2.n12 Q2.n11 0.0288742
R30774 Q2.n10 Q2 0.0226455
R30775 Q2 Q2.n15 0.0168043
R30776 Q2.n15 Q2 0.0122188
R30777 Q2.n1 Q2.n0 0.0107679
R30778 Q2.n0 Q2 0.0107679
R30779 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 179.256
R30780 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 168.089
R30781 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 150.293
R30782 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 73.6304
R30783 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 60.4568
R30784 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 12.0358
R30785 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.981478
R30786 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 0.788543
R30787 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.769522
R30788 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 0.720633
R30789 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 0.682565
R30790 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.580578
R30791 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 0.55213
R30792 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 0.470609
R30793 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.447191
R30794 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.428234
R30795 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1255
R30796 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1255
R30797 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 0.063
R30798 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 0.063
R30799 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.063
R30800 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 0.063
R30801 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 0.063
R30802 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 0.0435206
R30803 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 0.0107679
R30804 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.0107679
R30805 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 179.256
R30806 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 168.089
R30807 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 150.293
R30808 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 73.6304
R30809 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 60.4568
R30810 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 12.0358
R30811 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.981478
R30812 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 0.788543
R30813 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.769522
R30814 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 0.720633
R30815 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 0.682565
R30816 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.580578
R30817 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 0.55213
R30818 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 0.470609
R30819 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.447191
R30820 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.428234
R30821 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1255
R30822 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1255
R30823 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 0.063
R30824 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 0.063
R30825 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.063
R30826 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 0.063
R30827 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 0.063
R30828 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 0.0435206
R30829 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 0.0107679
R30830 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.0107679
R30831 Nand_Gate_1.A.n33 Nand_Gate_1.A.t0 169.46
R30832 Nand_Gate_1.A.n33 Nand_Gate_1.A.t3 167.809
R30833 Nand_Gate_1.A.n35 Nand_Gate_1.A.t2 167.809
R30834 Nand_Gate_1.A Nand_Gate_1.A.t6 158.585
R30835 Nand_Gate_1.A.n21 Nand_Gate_1.A.t5 150.293
R30836 Nand_Gate_1.A.t6 Nand_Gate_1.A.n2 150.293
R30837 Nand_Gate_1.A.n14 Nand_Gate_1.A.t4 150.273
R30838 Nand_Gate_1.A.n8 Nand_Gate_1.A.t11 150.273
R30839 Nand_Gate_1.A.n12 Nand_Gate_1.A.t9 73.6406
R30840 Nand_Gate_1.A.n6 Nand_Gate_1.A.t7 73.6406
R30841 Nand_Gate_1.A.n23 Nand_Gate_1.A.t8 73.6304
R30842 Nand_Gate_1.A.n0 Nand_Gate_1.A.t10 73.6304
R30843 Nand_Gate_1.A.n4 Nand_Gate_1.A.t1 60.3809
R30844 Nand_Gate_1.A.n27 Nand_Gate_1.A.n26 14.3097
R30845 Nand_Gate_1.A.n34 Nand_Gate_1.A.n33 11.4489
R30846 Nand_Gate_1.A.n36 Nand_Gate_1.A.n35 8.21389
R30847 Nand_Gate_1.A.n18 Nand_Gate_1.A.n11 8.1418
R30848 Nand_Gate_1.A.n29 Nand_Gate_1.A.n28 5.61191
R30849 Nand_Gate_1.A.n29 Nand_Gate_1.A 5.35402
R30850 Nand_Gate_1.A.n30 Nand_Gate_1.A.n29 4.563
R30851 Nand_Gate_1.A.n18 Nand_Gate_1.A.n17 4.5005
R30852 Nand_Gate_1.A.n28 Nand_Gate_1.A 1.83746
R30853 Nand_Gate_1.A.n20 Nand_Gate_1.A.n19 1.62007
R30854 Nand_Gate_1.A.n2 Nand_Gate_1.A.n1 1.19615
R30855 Nand_Gate_1.A.n5 Nand_Gate_1.A 1.08746
R30856 Nand_Gate_1.A.n20 Nand_Gate_1.A 1.01739
R30857 Nand_Gate_1.A.n13 Nand_Gate_1.A 0.851043
R30858 Nand_Gate_1.A.n7 Nand_Gate_1.A 0.851043
R30859 Nand_Gate_1.A.n4 Nand_Gate_1.A 0.848156
R30860 Nand_Gate_1.A.n32 Nand_Gate_1.A.n31 0.788543
R30861 Nand_Gate_1.A.n22 Nand_Gate_1.A 0.769522
R30862 Nand_Gate_1.A.n5 Nand_Gate_1.A.n4 0.682565
R30863 Nand_Gate_1.A.n31 Nand_Gate_1.A 0.65675
R30864 Nand_Gate_1.A.n22 Nand_Gate_1.A.n21 0.55213
R30865 Nand_Gate_1.A.n16 Nand_Gate_1.A.n15 0.55213
R30866 Nand_Gate_1.A.n10 Nand_Gate_1.A.n9 0.55213
R30867 Nand_Gate_1.A.n16 Nand_Gate_1.A 0.486828
R30868 Nand_Gate_1.A.n10 Nand_Gate_1.A 0.486828
R30869 Nand_Gate_1.A.n25 Nand_Gate_1.A.n24 0.470609
R30870 Nand_Gate_1.A.n13 Nand_Gate_1.A.n12 0.470609
R30871 Nand_Gate_1.A.n7 Nand_Gate_1.A.n6 0.470609
R30872 Nand_Gate_1.A.n21 Nand_Gate_1.A 0.447191
R30873 Nand_Gate_1.A.n2 Nand_Gate_1.A 0.447191
R30874 Nand_Gate_1.A.n25 Nand_Gate_1.A 0.428234
R30875 Nand_Gate_1.A.n36 Nand_Gate_1.A.n3 0.425067
R30876 Nand_Gate_1.A Nand_Gate_1.A.n36 0.39003
R30877 Nand_Gate_1.A.n35 Nand_Gate_1.A.n34 0.280391
R30878 Nand_Gate_1.A.n34 Nand_Gate_1.A.n32 0.262643
R30879 Nand_Gate_1.A.n12 Nand_Gate_1.A 0.217464
R30880 Nand_Gate_1.A.n6 Nand_Gate_1.A 0.217464
R30881 Nand_Gate_1.A.n24 Nand_Gate_1.A 0.1255
R30882 Nand_Gate_1.A.n15 Nand_Gate_1.A 0.1255
R30883 Nand_Gate_1.A.n9 Nand_Gate_1.A 0.1255
R30884 Nand_Gate_1.A.n32 Nand_Gate_1.A 0.1255
R30885 Nand_Gate_1.A.n1 Nand_Gate_1.A 0.1255
R30886 Nand_Gate_1.A.n26 Nand_Gate_1.A.n22 0.063
R30887 Nand_Gate_1.A.n26 Nand_Gate_1.A.n25 0.063
R30888 Nand_Gate_1.A.n17 Nand_Gate_1.A.n13 0.063
R30889 Nand_Gate_1.A.n17 Nand_Gate_1.A.n16 0.063
R30890 Nand_Gate_1.A.n11 Nand_Gate_1.A.n7 0.063
R30891 Nand_Gate_1.A.n11 Nand_Gate_1.A.n10 0.063
R30892 Nand_Gate_1.A.n28 Nand_Gate_1.A.n27 0.063
R30893 Nand_Gate_1.A.n27 Nand_Gate_1.A.n20 0.063
R30894 Nand_Gate_1.A.n30 Nand_Gate_1.A.n5 0.063
R30895 Nand_Gate_1.A.n31 Nand_Gate_1.A.n30 0.063
R30896 Nand_Gate_1.A.n32 Nand_Gate_1.A 0.063
R30897 Nand_Gate_1.A Nand_Gate_1.A.n18 0.0512812
R30898 Nand_Gate_1.A.n15 Nand_Gate_1.A.n14 0.0216397
R30899 Nand_Gate_1.A.n14 Nand_Gate_1.A 0.0216397
R30900 Nand_Gate_1.A.n9 Nand_Gate_1.A.n8 0.0216397
R30901 Nand_Gate_1.A.n8 Nand_Gate_1.A 0.0216397
R30902 Nand_Gate_1.A.n19 Nand_Gate_1.A 0.0168043
R30903 Nand_Gate_1.A.n19 Nand_Gate_1.A 0.0122188
R30904 Nand_Gate_1.A.n24 Nand_Gate_1.A.n23 0.0107679
R30905 Nand_Gate_1.A.n23 Nand_Gate_1.A 0.0107679
R30906 Nand_Gate_1.A.n1 Nand_Gate_1.A.n0 0.0107679
R30907 Nand_Gate_1.A.n0 Nand_Gate_1.A 0.0107679
R30908 Nand_Gate_1.A.n3 Nand_Gate_1.A 0.00441667
R30909 Nand_Gate_1.A.n3 Nand_Gate_1.A 0.00406061
R30910 Q4.n2 Q4.t3 169.46
R30911 Q4.n4 Q4.t1 167.809
R30912 Q4.n2 Q4.t2 167.809
R30913 Q4 Q4.t9 158.585
R30914 Q4.n15 Q4.t8 150.869
R30915 Q4.t9 Q4.n9 150.293
R30916 Q4.n17 Q4.t7 150.273
R30917 Q4.n14 Q4.n13 137.644
R30918 Q4.n13 Q4 85.5731
R30919 Q4.n16 Q4.t4 74.1352
R30920 Q4.n15 Q4.t6 74.1352
R30921 Q4.n7 Q4.t5 73.6304
R30922 Q4.n0 Q4.t0 60.3809
R30923 Q4.n3 Q4.n2 11.4489
R30924 Q4.n5 Q4.n4 8.21389
R30925 Q4 Q4.n17 4.54933
R30926 Q4.n13 Q4.n12 3.473
R30927 Q4.n16 Q4.n15 1.66898
R30928 Q4.n1 Q4.n0 1.64452
R30929 Q4.n9 Q4.n8 1.19615
R30930 Q4.n0 Q4 0.848156
R30931 Q4.n17 Q4.n16 0.55213
R30932 Q4.n9 Q4 0.447191
R30933 Q4.n5 Q4 0.39003
R30934 Q4.n4 Q4.n3 0.280391
R30935 Q4.n3 Q4.n1 0.262643
R30936 Q4.n6 Q4.n5 0.219833
R30937 Q4.n6 Q4 0.20965
R30938 Q4.n11 Q4.n10 0.154033
R30939 Q4.n11 Q4 0.143636
R30940 Q4.n1 Q4 0.1255
R30941 Q4.n8 Q4 0.1255
R30942 Q4.n15 Q4 0.063
R30943 Q4.n1 Q4 0.063
R30944 Q4.n12 Q4.n6 0.024
R30945 Q4.n12 Q4.n11 0.024
R30946 Q4.n14 Q4 0.0168043
R30947 Q4 Q4.n14 0.0122188
R30948 Q4.n8 Q4.n7 0.0107679
R30949 Q4.n7 Q4 0.0107679
R30950 Q4.n10 Q4 0.00441667
R30951 Q4.n10 Q4 0.00406061
R30952 And_Gate_6.Vout.n14 And_Gate_6.Vout.t0 168.108
R30953 And_Gate_6.Vout.n5 And_Gate_6.Vout.t2 158.207
R30954 D_FlipFlop_3.CLK And_Gate_6.Vout.t4 158.202
R30955 And_Gate_6.Vout.n7 And_Gate_6.Vout.t3 150.293
R30956 And_Gate_6.Vout.t4 And_Gate_6.Vout.n10 150.293
R30957 And_Gate_6.Vout.t2 And_Gate_6.Vout.n4 150.273
R30958 And_Gate_6.Vout.n2 And_Gate_6.Vout.t5 73.6406
R30959 And_Gate_6.Vout.n9 And_Gate_6.Vout.t7 73.6304
R30960 And_Gate_6.Vout.n8 And_Gate_6.Vout.t6 73.6304
R30961 And_Gate_6.Inverter_0.Vout And_Gate_6.Vout.t1 60.3943
R30962 And_Gate_6.Vout.n12 And_Gate_6.Vout.n11 42.3602
R30963 And_Gate_6.Vout.n9 And_Gate_6.Vout.n8 16.332
R30964 And_Gate_6.Vout.n3 And_Gate_6.Vout.n2 1.19615
R30965 And_Gate_6.Vout.n8 And_Gate_6.Vout.n7 1.1717
R30966 And_Gate_6.Vout.n10 And_Gate_6.Vout.n9 1.1717
R30967 And_Gate_6.Vout.n13 And_Gate_6.Inverter_0.Vout 0.981478
R30968 And_Gate_6.Vout.n14 And_Gate_6.Vout.n13 0.788543
R30969 And_Gate_6.Vout.n1 And_Gate_6.Vout.n0 0.682565
R30970 And_Gate_6.Vout.n1 And_Gate_6.Inverter_0.Vout 0.580578
R30971 And_Gate_6.Inverter_0.Vout And_Gate_6.Vout.n14 0.484875
R30972 And_Gate_6.Vout.n10 D_FlipFlop_3.3-input-nand_1.C 0.447191
R30973 And_Gate_6.Vout.n7 D_FlipFlop_3.Inverter_1.Vin 0.436162
R30974 And_Gate_6.Vout.n5 D_FlipFlop_3.CLK 0.321667
R30975 And_Gate_6.Vout.n6 And_Gate_6.Vout.n5 0.29425
R30976 And_Gate_6.Vout.n2 D_FlipFlop_3.3-input-nand_0.C 0.217464
R30977 And_Gate_6.Vout.n9 D_FlipFlop_3.3-input-nand_1.C 0.149957
R30978 And_Gate_6.Vout.n3 D_FlipFlop_3.3-input-nand_0.C 0.1255
R30979 And_Gate_6.Vout.n0 And_Gate_6.Inverter_0.Vout 0.1255
R30980 And_Gate_6.Vout.n8 D_FlipFlop_3.Inverter_1.Vin 0.117348
R30981 And_Gate_6.Vout.n0 And_Gate_6.Inverter_0.Vout 0.063
R30982 And_Gate_6.Vout.n13 And_Gate_6.Vout.n12 0.063
R30983 And_Gate_6.Vout.n12 And_Gate_6.Vout.n1 0.063
R30984 And_Gate_6.Vout.n6 D_FlipFlop_3.CLK 0.0600333
R30985 And_Gate_6.Vout.n8 D_FlipFlop_3.Inverter_1.Vin 0.0454219
R30986 And_Gate_6.Vout.n9 D_FlipFlop_3.3-input-nand_1.C 0.0454219
R30987 And_Gate_6.Vout.n11 And_Gate_6.Vout.n6 0.024
R30988 And_Gate_6.Vout.n11 D_FlipFlop_3.CLK 0.024
R30989 And_Gate_6.Vout.n4 And_Gate_6.Vout.n3 0.0216397
R30990 And_Gate_6.Vout.n4 D_FlipFlop_3.3-input-nand_0.C 0.0216397
R30991 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 169.46
R30992 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 168.089
R30993 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 167.809
R30994 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 150.273
R30995 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 73.6406
R30996 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 60.3809
R30997 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 12.0358
R30998 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 11.4489
R30999 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 1.08746
R31000 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.851043
R31001 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.848156
R31002 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 0.788543
R31003 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 0.682565
R31004 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.65675
R31005 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 0.55213
R31006 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.486828
R31007 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 0.470609
R31008 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 0.262643
R31009 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.217464
R31010 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.1255
R31011 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.1255
R31012 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 0.063
R31013 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 0.063
R31014 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 0.063
R31015 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 0.063
R31016 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 0.063
R31017 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 0.0216397
R31018 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0216397
R31019 And_Gate_0.Vout.n12 And_Gate_0.Vout.t0 168.32
R31020 And_Gate_0.Vout.n4 And_Gate_0.Vout.t5 158.246
R31021 D_FlipFlop_6.CLK And_Gate_0.Vout.t7 158.202
R31022 And_Gate_0.Vout.n5 And_Gate_0.Vout.t6 150.293
R31023 And_Gate_0.Vout.t7 And_Gate_0.Vout.n8 150.293
R31024 And_Gate_0.Vout.t5 And_Gate_0.Vout.n3 150.273
R31025 And_Gate_0.Vout.n1 And_Gate_0.Vout.t4 73.6406
R31026 And_Gate_0.Vout.n7 And_Gate_0.Vout.t3 73.6304
R31027 And_Gate_0.Vout.n6 And_Gate_0.Vout.t2 73.6304
R31028 And_Gate_0.Vout.n12 And_Gate_0.Vout.n11 66.7548
R31029 And_Gate_0.Inverter_0.Vout And_Gate_0.Vout.t1 60.3943
R31030 And_Gate_0.Vout.n7 And_Gate_0.Vout.n6 16.332
R31031 And_Gate_0.Vout.n13 And_Gate_0.Vout.n0 1.62007
R31032 And_Gate_0.Inverter_0.Vout And_Gate_0.Vout.n13 1.25441
R31033 And_Gate_0.Vout.n2 And_Gate_0.Vout.n1 1.19615
R31034 And_Gate_0.Vout.n6 And_Gate_0.Vout.n5 1.1717
R31035 And_Gate_0.Vout.n8 And_Gate_0.Vout.n7 1.1717
R31036 And_Gate_0.Vout.n8 D_FlipFlop_6.3-input-nand_1.C 0.447191
R31037 And_Gate_0.Vout.n5 D_FlipFlop_6.Inverter_1.Vin 0.436162
R31038 And_Gate_0.Vout.n4 D_FlipFlop_6.CLK 0.281076
R31039 And_Gate_0.Vout.n10 And_Gate_0.Vout.n9 0.245683
R31040 And_Gate_0.Vout.n1 D_FlipFlop_6.3-input-nand_0.C 0.217464
R31041 And_Gate_0.Vout.n10 D_FlipFlop_6.CLK 0.197158
R31042 And_Gate_0.Vout.n7 D_FlipFlop_6.3-input-nand_1.C 0.149957
R31043 And_Gate_0.Vout.n2 D_FlipFlop_6.3-input-nand_0.C 0.1255
R31044 And_Gate_0.Vout.n0 And_Gate_0.Inverter_0.Vout 0.1255
R31045 And_Gate_0.Vout.n6 D_FlipFlop_6.Inverter_1.Vin 0.117348
R31046 And_Gate_0.Vout.n0 And_Gate_0.Inverter_0.Vout 0.063
R31047 And_Gate_0.Vout.n13 And_Gate_0.Vout.n12 0.063
R31048 And_Gate_0.Vout.n6 D_FlipFlop_6.Inverter_1.Vin 0.0454219
R31049 And_Gate_0.Vout.n7 D_FlipFlop_6.3-input-nand_1.C 0.0454219
R31050 And_Gate_0.Vout.n11 And_Gate_0.Vout.n4 0.024
R31051 And_Gate_0.Vout.n11 And_Gate_0.Vout.n10 0.024
R31052 And_Gate_0.Vout.n3 And_Gate_0.Vout.n2 0.0216397
R31053 And_Gate_0.Vout.n3 D_FlipFlop_6.3-input-nand_0.C 0.0216397
R31054 And_Gate_0.Vout.n9 D_FlipFlop_6.CLK 0.00441667
R31055 And_Gate_0.Vout.n9 D_FlipFlop_6.CLK 0.00406061
R31056 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 169.46
R31057 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 167.809
R31058 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 167.809
R31059 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 167.226
R31060 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 150.273
R31061 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 150.273
R31062 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 73.6406
R31063 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 73.6304
R31064 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 60.4568
R31065 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 12.3891
R31066 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 11.4489
R31067 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.68257
R31068 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 1.38365
R31069 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 1.19615
R31070 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 1.1717
R31071 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.08448
R31072 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.932141
R31073 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 0.720633
R31074 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 0.280391
R31075 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.217464
R31076 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R31077 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R31078 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R31079 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 0.0874565
R31080 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 0.063
R31081 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.063
R31082 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 0.063
R31083 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 0.063
R31084 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 0.0435206
R31085 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 0.0216397
R31086 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.0216397
R31087 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 0.0107679
R31088 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.0107679
R31089 And_Gate_5.A.n10 And_Gate_5.A.t0 179.256
R31090 And_Gate_5.A.n10 And_Gate_5.A.t2 168.089
R31091 And_Gate_5.A.n2 And_Gate_5.A.t4 150.293
R31092 And_Gate_5.A.n4 And_Gate_5.A.t3 73.6304
R31093 Nand_Gate_3.Vout And_Gate_5.A.t1 60.3943
R31094 And_Gate_5.A.n8 And_Gate_5.A.n7 35.6663
R31095 And_Gate_5.A.n9 Nand_Gate_3.Vout 0.981478
R31096 And_Gate_5.A.n11 And_Gate_5.A.n9 0.788543
R31097 And_Gate_5.A.n3 And_Gate_5.Nand_Gate_0.A 0.769522
R31098 Nand_Gate_3.Vout And_Gate_5.A.n11 0.720633
R31099 And_Gate_5.A.n1 And_Gate_5.A.n0 0.682565
R31100 And_Gate_5.A.n1 Nand_Gate_3.Vout 0.580578
R31101 And_Gate_5.A.n3 And_Gate_5.A.n2 0.55213
R31102 And_Gate_5.A.n6 And_Gate_5.A.n5 0.470609
R31103 And_Gate_5.A.n2 And_Gate_5.Nand_Gate_0.A 0.447191
R31104 And_Gate_5.A.n6 And_Gate_5.Nand_Gate_0.A 0.428234
R31105 And_Gate_5.A.n5 And_Gate_5.Nand_Gate_0.A 0.1255
R31106 And_Gate_5.A.n0 Nand_Gate_3.Vout 0.1255
R31107 And_Gate_5.A.n7 And_Gate_5.A.n3 0.063
R31108 And_Gate_5.A.n7 And_Gate_5.A.n6 0.063
R31109 And_Gate_5.A.n0 Nand_Gate_3.Vout 0.063
R31110 And_Gate_5.A.n9 And_Gate_5.A.n8 0.063
R31111 And_Gate_5.A.n8 And_Gate_5.A.n1 0.063
R31112 And_Gate_5.A.n11 And_Gate_5.A.n10 0.0435206
R31113 And_Gate_5.A.n5 And_Gate_5.A.n4 0.0107679
R31114 And_Gate_5.A.n4 And_Gate_5.Nand_Gate_0.A 0.0107679
R31115 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 169.46
R31116 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 168.089
R31117 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 167.809
R31118 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 150.273
R31119 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 73.6406
R31120 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 60.3809
R31121 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 12.0358
R31122 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 11.4489
R31123 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 1.08746
R31124 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.851043
R31125 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.848156
R31126 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 0.788543
R31127 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 0.682565
R31128 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.65675
R31129 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 0.55213
R31130 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.486828
R31131 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 0.470609
R31132 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 0.262643
R31133 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.217464
R31134 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.1255
R31135 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.1255
R31136 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 0.063
R31137 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 0.063
R31138 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 0.063
R31139 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 0.063
R31140 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 0.063
R31141 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 0.0216397
R31142 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0216397
R31143 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 169.46
R31144 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 168.089
R31145 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 167.809
R31146 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 150.273
R31147 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 73.6406
R31148 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 60.3809
R31149 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 12.0358
R31150 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 11.4489
R31151 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 1.08746
R31152 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.851043
R31153 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.848156
R31154 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 0.788543
R31155 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 0.682565
R31156 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.65675
R31157 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 0.55213
R31158 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.486828
R31159 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 0.470609
R31160 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 0.262643
R31161 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.217464
R31162 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.1255
R31163 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.1255
R31164 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 0.063
R31165 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 0.063
R31166 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 0.063
R31167 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 0.063
R31168 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 0.063
R31169 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 0.0216397
R31170 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.0216397
R31171 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 169.46
R31172 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 168.089
R31173 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 167.809
R31174 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 150.293
R31175 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 73.6304
R31176 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 60.3943
R31177 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 12.0358
R31178 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 11.4489
R31179 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.981478
R31180 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 0.788543
R31181 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.769522
R31182 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 0.720633
R31183 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 0.682565
R31184 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.580578
R31185 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 0.55213
R31186 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 0.470609
R31187 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.447191
R31188 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.428234
R31189 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.1255
R31190 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.1255
R31191 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 0.063
R31192 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 0.063
R31193 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.063
R31194 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 0.063
R31195 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 0.063
R31196 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 0.0435206
R31197 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 0.0107679
R31198 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.0107679
R31199 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t1 169.46
R31200 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.t2 167.809
R31201 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t0 167.809
R31202 D_FlipFlop_4.3-input-nand_2.Vout.t7 D_FlipFlop_4.3-input-nand_2.Vout.n11 167.227
R31203 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.t7 150.293
R31204 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.t5 150.273
R31205 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6406
R31206 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout.t4 73.6304
R31207 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout.t3 60.3809
R31208 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n5 12.3891
R31209 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout.n9 11.4489
R31210 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout.n2 1.38365
R31211 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.n1 1.19615
R31212 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.n4 1.1717
R31213 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout 0.848156
R31214 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.Vout.n12 0.447191
R31215 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout 0.38637
R31216 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.n10 0.280391
R31217 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout.n8 0.262643
R31218 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout 0.217464
R31219 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R31220 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R31221 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R31222 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R31223 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout.n7 0.0874565
R31224 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n3 0.063
R31225 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout.n6 0.063
R31226 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout 0.063
R31227 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R31228 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout.n0 0.0107679
R31229 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout 0.0107679
R31230 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.t1 169.46
R31231 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C.t3 167.809
R31232 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.t0 167.809
R31233 D_FlipFlop_4.3-input-nand_2.C.t4 D_FlipFlop_4.3-input-nand_2.C.n13 167.226
R31234 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C.t6 150.273
R31235 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.t4 150.273
R31236 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C.t5 73.6406
R31237 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C.t7 73.6304
R31238 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C.t2 60.4568
R31239 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C.n7 12.3891
R31240 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.n11 11.4489
R31241 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C 1.68257
R31242 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C.n2 1.38365
R31243 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C.n0 1.19615
R31244 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C.n5 1.1717
R31245 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C 1.08448
R31246 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C 0.932141
R31247 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C 0.720633
R31248 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C.n12 0.280391
R31249 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C 0.217464
R31250 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C 0.1255
R31251 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C 0.1255
R31252 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C 0.1255
R31253 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C.n9 0.0874565
R31254 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C.n6 0.063
R31255 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C 0.063
R31256 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C.n8 0.063
R31257 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C.n3 0.063
R31258 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.n10 0.0435206
R31259 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.n1 0.0216397
R31260 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_2.C.n14 0.0216397
R31261 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C.n4 0.0107679
R31262 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C 0.0107679
R31263 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 179.256
R31264 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 168.089
R31265 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 150.293
R31266 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 73.6304
R31267 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 60.4568
R31268 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 12.0358
R31269 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.981478
R31270 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 0.788543
R31271 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.769522
R31272 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.720633
R31273 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 0.682565
R31274 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.580578
R31275 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 0.55213
R31276 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 0.470609
R31277 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.447191
R31278 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.428234
R31279 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1255
R31280 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1255
R31281 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 0.063
R31282 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 0.063
R31283 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 0.063
R31284 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 0.063
R31285 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 0.063
R31286 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 0.0435206
R31287 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 0.0107679
R31288 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.0107679
R31289 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z.t3 168.609
R31290 CDAC8_0.switch_0.Z CDAC8_0.switch_0.Z.t0 168.565
R31291 CDAC8_0.switch_0.Z.n0 CDAC8_0.switch_0.Z.t1 60.321
R31292 CDAC8_0.switch_0.Z.n0 CDAC8_0.switch_0.Z.t2 60.321
R31293 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z.n6 11.3205
R31294 CDAC8_0.switch_0.Z.n4 CDAC8_0.switch_0.Z.n3 5.58885
R31295 CDAC8_0.switch_0.Z.n6 CDAC8_0.switch_0.Z.n2 2.98587
R31296 CDAC8_0.switch_0.Z.n6 CDAC8_0.switch_0.Z.n5 2.5049
R31297 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z.n1 1.60376
R31298 CDAC8_0.switch_0.Z.n2 CDAC8_0.switch_0.Z.t5 0.658247
R31299 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z.t7 0.658247
R31300 CDAC8_0.switch_0.Z.n3 CDAC8_0.switch_0.Z.t6 0.611304
R31301 CDAC8_0.switch_0.Z.n4 CDAC8_0.switch_0.Z.t4 0.611304
R31302 CDAC8_0.switch_0.Z.n1 CDAC8_0.switch_0.Z 0.259656
R31303 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z 0.166261
R31304 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z.n4 0.115412
R31305 CDAC8_0.switch_0.Z.n3 CDAC8_0.switch_0.Z.n2 0.115412
R31306 CDAC8_0.switch_0.Z CDAC8_0.switch_0.Z.n7 0.0454219
R31307 CDAC8_0.switch_0.Z.n1 CDAC8_0.switch_0.Z.n0 0.0188121
R31308 RingCounter_0.D_FlipFlop_16.Q.n20 RingCounter_0.D_FlipFlop_16.Q.t3 169.46
R31309 RingCounter_0.D_FlipFlop_16.Q.n20 RingCounter_0.D_FlipFlop_16.Q.t2 167.809
R31310 RingCounter_0.D_FlipFlop_16.Q.n19 RingCounter_0.D_FlipFlop_16.Q.t1 167.809
R31311 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Q.t8 158.585
R31312 RingCounter_0.D_FlipFlop_16.Q.t8 RingCounter_0.D_FlipFlop_16.Q.n15 150.293
R31313 RingCounter_0.D_FlipFlop_16.Q.n8 RingCounter_0.D_FlipFlop_16.Q.t7 150.273
R31314 RingCounter_0.D_FlipFlop_16.Q.n2 RingCounter_0.D_FlipFlop_16.Q.t6 150.273
R31315 RingCounter_0.D_FlipFlop_16.Q.n6 RingCounter_0.D_FlipFlop_16.Q.t9 73.6406
R31316 RingCounter_0.D_FlipFlop_16.Q.n0 RingCounter_0.D_FlipFlop_16.Q.t4 73.6406
R31317 RingCounter_0.D_FlipFlop_16.Q.n13 RingCounter_0.D_FlipFlop_16.Q.t5 73.6304
R31318 RingCounter_0.D_FlipFlop_16.Q.n18 RingCounter_0.D_FlipFlop_16.Q.n12 62.8776
R31319 RingCounter_0.D_FlipFlop_16.Q.n23 RingCounter_0.D_FlipFlop_16.Q.t0 60.3809
R31320 RingCounter_0.D_FlipFlop_16.Q.n21 RingCounter_0.D_FlipFlop_16.Q.n20 11.4489
R31321 RingCounter_0.D_FlipFlop_16.Q.n19 RingCounter_0.D_FlipFlop_16.Q.n18 8.19039
R31322 RingCounter_0.D_FlipFlop_16.Q.n12 RingCounter_0.D_FlipFlop_16.Q.n5 8.1418
R31323 RingCounter_0.D_FlipFlop_16.Q.n12 RingCounter_0.D_FlipFlop_16.Q.n11 4.5005
R31324 RingCounter_0.D_FlipFlop_16.Q.n23 RingCounter_0.D_FlipFlop_16.Q.n22 1.64452
R31325 RingCounter_0.D_FlipFlop_16.Q.n15 RingCounter_0.D_FlipFlop_16.Q.n14 1.19615
R31326 RingCounter_0.D_FlipFlop_16.Q.n7 RingCounter_0.D_FlipFlop_16.Q 0.851043
R31327 RingCounter_0.D_FlipFlop_16.Q.n1 RingCounter_0.D_FlipFlop_16.Q 0.851043
R31328 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Q.n23 0.848156
R31329 RingCounter_0.D_FlipFlop_16.Q.n10 RingCounter_0.D_FlipFlop_16.Q.n9 0.55213
R31330 RingCounter_0.D_FlipFlop_16.Q.n4 RingCounter_0.D_FlipFlop_16.Q.n3 0.55213
R31331 RingCounter_0.D_FlipFlop_16.Q.n10 RingCounter_0.D_FlipFlop_16.Q 0.486828
R31332 RingCounter_0.D_FlipFlop_16.Q.n4 RingCounter_0.D_FlipFlop_16.Q 0.486828
R31333 RingCounter_0.D_FlipFlop_16.Q.n7 RingCounter_0.D_FlipFlop_16.Q.n6 0.470609
R31334 RingCounter_0.D_FlipFlop_16.Q.n1 RingCounter_0.D_FlipFlop_16.Q.n0 0.470609
R31335 RingCounter_0.D_FlipFlop_16.Q.n15 RingCounter_0.D_FlipFlop_16.Q 0.447191
R31336 RingCounter_0.D_FlipFlop_16.Q.n17 RingCounter_0.D_FlipFlop_16.Q.n16 0.425067
R31337 RingCounter_0.D_FlipFlop_16.Q.n17 RingCounter_0.D_FlipFlop_16.Q 0.39003
R31338 RingCounter_0.D_FlipFlop_16.Q.n21 RingCounter_0.D_FlipFlop_16.Q.n19 0.280391
R31339 RingCounter_0.D_FlipFlop_16.Q.n22 RingCounter_0.D_FlipFlop_16.Q.n21 0.262643
R31340 RingCounter_0.D_FlipFlop_16.Q.n6 RingCounter_0.D_FlipFlop_16.Q 0.217464
R31341 RingCounter_0.D_FlipFlop_16.Q.n0 RingCounter_0.D_FlipFlop_16.Q 0.217464
R31342 RingCounter_0.D_FlipFlop_16.Q.n9 RingCounter_0.D_FlipFlop_16.Q 0.1255
R31343 RingCounter_0.D_FlipFlop_16.Q.n3 RingCounter_0.D_FlipFlop_16.Q 0.1255
R31344 RingCounter_0.D_FlipFlop_16.Q.n14 RingCounter_0.D_FlipFlop_16.Q 0.1255
R31345 RingCounter_0.D_FlipFlop_16.Q.n22 RingCounter_0.D_FlipFlop_16.Q 0.1255
R31346 RingCounter_0.D_FlipFlop_16.Q.n11 RingCounter_0.D_FlipFlop_16.Q.n7 0.063
R31347 RingCounter_0.D_FlipFlop_16.Q.n11 RingCounter_0.D_FlipFlop_16.Q.n10 0.063
R31348 RingCounter_0.D_FlipFlop_16.Q.n5 RingCounter_0.D_FlipFlop_16.Q.n1 0.063
R31349 RingCounter_0.D_FlipFlop_16.Q.n5 RingCounter_0.D_FlipFlop_16.Q.n4 0.063
R31350 RingCounter_0.D_FlipFlop_16.Q.n22 RingCounter_0.D_FlipFlop_16.Q 0.063
R31351 RingCounter_0.D_FlipFlop_16.Q.n18 RingCounter_0.D_FlipFlop_16.Q.n17 0.024
R31352 RingCounter_0.D_FlipFlop_16.Q.n9 RingCounter_0.D_FlipFlop_16.Q.n8 0.0216397
R31353 RingCounter_0.D_FlipFlop_16.Q.n8 RingCounter_0.D_FlipFlop_16.Q 0.0216397
R31354 RingCounter_0.D_FlipFlop_16.Q.n3 RingCounter_0.D_FlipFlop_16.Q.n2 0.0216397
R31355 RingCounter_0.D_FlipFlop_16.Q.n2 RingCounter_0.D_FlipFlop_16.Q 0.0216397
R31356 RingCounter_0.D_FlipFlop_16.Q.n14 RingCounter_0.D_FlipFlop_16.Q.n13 0.0107679
R31357 RingCounter_0.D_FlipFlop_16.Q.n13 RingCounter_0.D_FlipFlop_16.Q 0.0107679
R31358 RingCounter_0.D_FlipFlop_16.Q.n16 RingCounter_0.D_FlipFlop_16.Q 0.00441667
R31359 RingCounter_0.D_FlipFlop_16.Q.n16 RingCounter_0.D_FlipFlop_16.Q 0.00406061
R31360 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 316.762
R31361 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 168.108
R31362 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 150.293
R31363 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 150.273
R31364 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 73.6406
R31365 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 73.6304
R31366 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 60.3943
R31367 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 12.0358
R31368 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 1.19615
R31369 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.981478
R31370 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 0.788543
R31371 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.769522
R31372 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 0.682565
R31373 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.580578
R31374 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 0.55213
R31375 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 0.484875
R31376 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 0.470609
R31377 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.447191
R31378 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.428234
R31379 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.217464
R31380 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R31381 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R31382 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R31383 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 0.063
R31384 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 0.063
R31385 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.063
R31386 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 0.063
R31387 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 0.063
R31388 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 0.0216397
R31389 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.0216397
R31390 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 0.0107679
R31391 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.0107679
R31392 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 179.256
R31393 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 168.089
R31394 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 150.273
R31395 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 73.6406
R31396 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 60.3809
R31397 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 12.0358
R31398 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 1.08746
R31399 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.851043
R31400 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.848156
R31401 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 0.788543
R31402 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 0.682565
R31403 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.65675
R31404 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 0.55213
R31405 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.486828
R31406 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 0.470609
R31407 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.217464
R31408 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 0.200143
R31409 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.1255
R31410 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.1255
R31411 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 0.063
R31412 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 0.063
R31413 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 0.063
R31414 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 0.063
R31415 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 0.063
R31416 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 0.0216397
R31417 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.0216397
R31418 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 316.762
R31419 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 168.108
R31420 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 150.293
R31421 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 150.273
R31422 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 73.6406
R31423 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 73.6304
R31424 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 60.3943
R31425 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 12.0358
R31426 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 1.19615
R31427 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.981478
R31428 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 0.788543
R31429 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.769522
R31430 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 0.682565
R31431 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.580578
R31432 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 0.55213
R31433 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 0.484875
R31434 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 0.470609
R31435 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.447191
R31436 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.428234
R31437 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.217464
R31438 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R31439 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R31440 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R31441 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 0.063
R31442 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 0.063
R31443 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.063
R31444 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 0.063
R31445 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 0.063
R31446 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 0.0216397
R31447 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.0216397
R31448 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 0.0107679
R31449 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.0107679
R31450 a_138485_16882.n0 a_138485_16882.t4 575.905
R31451 a_138485_16882.n1 a_138485_16882.t1 575.905
R31452 a_138485_16882.n0 a_138485_16882.t3 338.675
R31453 a_138485_16882.t0 a_138485_16882.n2 13.268
R31454 a_138485_16882.n2 a_138485_16882.t2 9.51806
R31455 a_138485_16882.n1 a_138485_16882.n0 1.7505
R31456 a_138485_16882.n2 a_138485_16882.n1 0.484196
R31457 Vbias.n26 Vbias.n18 93853.1
R31458 Vbias.n26 Vbias.n19 93853.1
R31459 Vbias.n22 Vbias.n18 93853.1
R31460 Vbias.n18 Vbias.n17 41816.1
R31461 Vbias.n64 Vbias.n9 7992.36
R31462 Vbias.n65 Vbias.n9 7992.36
R31463 Vbias.n65 Vbias.n8 7992.36
R31464 Vbias.n64 Vbias.n8 7992.36
R31465 Vbias.n33 Vbias.n14 7992.36
R31466 Vbias.n33 Vbias.n15 7992.36
R31467 Vbias.n29 Vbias.n15 7992.36
R31468 Vbias.n29 Vbias.n14 7992.36
R31469 Vbias.n57 Vbias.n43 6345.81
R31470 Vbias.n57 Vbias.n44 6345.81
R31471 Vbias.n61 Vbias.n44 6345.81
R31472 Vbias.n61 Vbias.n43 6345.81
R31473 Vbias.n40 Vbias.n11 6345.81
R31474 Vbias.n40 Vbias.n12 6345.81
R31475 Vbias.n36 Vbias.n12 6345.81
R31476 Vbias.n36 Vbias.n11 6345.81
R31477 Vbias.n25 Vbias.n20 6098.07
R31478 Vbias.n23 Vbias.n20 6098.07
R31479 Vbias.n25 Vbias.n24 5912.48
R31480 Vbias.n24 Vbias.n23 5912.48
R31481 Vbias.n54 Vbias.n46 4699.26
R31482 Vbias.n54 Vbias.n47 4699.26
R31483 Vbias.n50 Vbias.n47 4699.26
R31484 Vbias.n32 Vbias.n31 918.212
R31485 Vbias.n63 Vbias.n7 918.212
R31486 Vbias.n63 Vbias.n6 918.212
R31487 Vbias.n31 Vbias.n30 918.212
R31488 Vbias.n66 Vbias.n7 861.144
R31489 Vbias.n30 Vbias.n16 861.144
R31490 Vbias.n32 Vbias.n5 819.201
R31491 Vbias.n67 Vbias.n6 819.201
R31492 Vbias.n58 Vbias.n45 729.976
R31493 Vbias.n59 Vbias.n58 729.976
R31494 Vbias.n60 Vbias.n59 729.976
R31495 Vbias.n60 Vbias.n45 729.976
R31496 Vbias.n39 Vbias.n13 729.976
R31497 Vbias.n39 Vbias.n38 729.976
R31498 Vbias.n38 Vbias.n37 729.976
R31499 Vbias.n37 Vbias.n13 729.976
R31500 Vbias.n51 Vbias.n48 541.741
R31501 Vbias.n53 Vbias.n48 541.741
R31502 Vbias.n52 Vbias.n51 484.675
R31503 Vbias.n53 Vbias.n52 484.675
R31504 Vbias.n28 Vbias.n27 296.86
R31505 Vbias.n22 Vbias.n21 190.803
R31506 Vbias.n27 Vbias.n17 186.645
R31507 Vbias.n56 Vbias.n55 164.214
R31508 Vbias.n31 Vbias.n14 117.001
R31509 Vbias.n14 Vbias.t5 117.001
R31510 Vbias.n16 Vbias.n15 117.001
R31511 Vbias.n15 Vbias.t5 117.001
R31512 Vbias.n64 Vbias.n63 117.001
R31513 Vbias.t3 Vbias.n64 117.001
R31514 Vbias.n66 Vbias.n65 117.001
R31515 Vbias.n65 Vbias.t3 117.001
R31516 Vbias.n13 Vbias.n11 117.001
R31517 Vbias.t9 Vbias.n11 117.001
R31518 Vbias.n38 Vbias.n12 117.001
R31519 Vbias.t9 Vbias.n12 117.001
R31520 Vbias.n45 Vbias.n43 117.001
R31521 Vbias.t1 Vbias.n43 117.001
R31522 Vbias.n59 Vbias.n44 117.001
R31523 Vbias.t1 Vbias.n44 117.001
R31524 Vbias.n48 Vbias.n46 117.001
R31525 Vbias.n52 Vbias.n47 117.001
R31526 Vbias.n47 Vbias.t7 117.001
R31527 Vbias.n49 Vbias.n46 112.052
R31528 Vbias.n50 Vbias.n49 86.728
R31529 Vbias.n28 Vbias.t5 72.8308
R31530 Vbias.n56 Vbias.t1 72.8308
R31531 Vbias.n55 Vbias.t7 72.8308
R31532 Vbias.n35 Vbias.n34 71.4462
R31533 Vbias.n62 Vbias.n42 71.4462
R31534 Vbias.n41 Vbias.n10 41.5387
R31535 Vbias.n20 Vbias.n18 32.5005
R31536 Vbias.n24 Vbias.n19 32.5005
R31537 Vbias.n21 Vbias.n19 32.4237
R31538 Vbias.t9 Vbias.n10 31.2926
R31539 Vbias.t3 Vbias.n41 31.2926
R31540 Vbias.n51 Vbias.n50 17.7278
R31541 Vbias.n54 Vbias.n53 17.7278
R31542 Vbias.n55 Vbias.n54 17.7278
R31543 Vbias.n16 Vbias.n5 17.443
R31544 Vbias.n67 Vbias.n66 17.443
R31545 Vbias.n2 Vbias.t8 16.8637
R31546 Vbias.n0 Vbias.t6 14.4765
R31547 Vbias.n1 Vbias.t4 14.02
R31548 Vbias.n37 Vbias.n36 12.4473
R31549 Vbias.n36 Vbias.n35 12.4473
R31550 Vbias.n40 Vbias.n39 12.4473
R31551 Vbias.n41 Vbias.n40 12.4473
R31552 Vbias.n61 Vbias.n60 12.4473
R31553 Vbias.n62 Vbias.n61 12.4473
R31554 Vbias.n58 Vbias.n57 12.4473
R31555 Vbias.n57 Vbias.n56 12.4473
R31556 Vbias.n69 Vbias.n0 11.6088
R31557 Vbias.n3 Vbias.t0 9.73694
R31558 Vbias.n30 Vbias.n29 9.43598
R31559 Vbias.n29 Vbias.n28 9.43598
R31560 Vbias.n33 Vbias.n32 9.43598
R31561 Vbias.n34 Vbias.n33 9.43598
R31562 Vbias.n8 Vbias.n6 9.43598
R31563 Vbias.n10 Vbias.n8 9.43598
R31564 Vbias.n9 Vbias.n7 9.43598
R31565 Vbias.n42 Vbias.n9 9.43598
R31566 Vbias.n4 Vbias.n3 8.19877
R31567 Vbias.n24 Vbias 6.10462
R31568 Vbias.n68 Vbias.n5 3.91345
R31569 Vbias.n68 Vbias.n67 3.91345
R31570 Vbias.n52 Vbias.n4 3.61865
R31571 Vbias.n3 Vbias.n2 3.4105
R31572 Vbias.t2 Vbias.n17 3.30535
R31573 Vbias.n69 Vbias.n4 2.813
R31574 Vbias.n49 Vbias.t7 2.16029
R31575 Vbias.n2 Vbias.n1 1.57387
R31576 Vbias.n35 Vbias.t5 1.38511
R31577 Vbias.n34 Vbias.t9 1.38511
R31578 Vbias.t3 Vbias.n62 1.38511
R31579 Vbias.t1 Vbias.n42 1.38511
R31580 Vbias.n26 Vbias.n25 1.28905
R31581 Vbias.n27 Vbias.n26 1.28905
R31582 Vbias.n23 Vbias.n22 1.28905
R31583 Vbias.n1 Vbias.n0 1.16354
R31584 Vbias.n69 Vbias.n68 0.664786
R31585 Vbias.n21 Vbias.t2 0.0670719
R31586 Vbias Vbias.n69 0.0512812
R31587 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 169.46
R31588 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 167.809
R31589 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 167.809
R31590 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 167.226
R31591 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 150.273
R31592 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 150.273
R31593 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 73.6406
R31594 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 73.6304
R31595 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 60.4568
R31596 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 12.3891
R31597 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 11.4489
R31598 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.68257
R31599 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 1.38365
R31600 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 1.19615
R31601 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 1.1717
R31602 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.08448
R31603 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.932141
R31604 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.720633
R31605 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 0.280391
R31606 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.217464
R31607 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R31608 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R31609 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R31610 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 0.0874565
R31611 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 0.063
R31612 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.063
R31613 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 0.063
R31614 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 0.063
R31615 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 0.0435206
R31616 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 0.0216397
R31617 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 0.0216397
R31618 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 0.0107679
R31619 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.0107679
R31620 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 169.46
R31621 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 168.089
R31622 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 167.809
R31623 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 150.293
R31624 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 73.6304
R31625 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 60.3943
R31626 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 12.0358
R31627 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 11.4489
R31628 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.981478
R31629 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 0.788543
R31630 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.769522
R31631 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 0.720633
R31632 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 0.682565
R31633 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.580578
R31634 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 0.55213
R31635 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 0.470609
R31636 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.447191
R31637 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.428234
R31638 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.1255
R31639 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.1255
R31640 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 0.063
R31641 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 0.063
R31642 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.063
R31643 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 0.063
R31644 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 0.063
R31645 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 0.0435206
R31646 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 0.0107679
R31647 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.0107679
R31648 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 169.46
R31649 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 168.089
R31650 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 167.809
R31651 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 150.293
R31652 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 73.6304
R31653 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 60.4568
R31654 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 12.0358
R31655 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 11.4489
R31656 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.981478
R31657 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 0.788543
R31658 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.769522
R31659 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 0.720633
R31660 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 0.682565
R31661 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.580578
R31662 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 0.55213
R31663 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 0.470609
R31664 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.447191
R31665 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.428234
R31666 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.1255
R31667 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.1255
R31668 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 0.063
R31669 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 0.063
R31670 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.063
R31671 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 0.063
R31672 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 0.063
R31673 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 0.0435206
R31674 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 0.0107679
R31675 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.0107679
R31676 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 169.46
R31677 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 167.809
R31678 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 167.809
R31679 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 167.226
R31680 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 150.273
R31681 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 150.273
R31682 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 73.6406
R31683 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 73.6304
R31684 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 60.4568
R31685 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 12.3891
R31686 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 11.4489
R31687 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.68257
R31688 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 1.38365
R31689 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 1.19615
R31690 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 1.1717
R31691 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.08448
R31692 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.932141
R31693 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 0.720633
R31694 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 0.280391
R31695 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.217464
R31696 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R31697 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R31698 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R31699 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 0.0874565
R31700 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 0.063
R31701 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.063
R31702 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 0.063
R31703 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 0.063
R31704 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 0.0435206
R31705 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 0.0216397
R31706 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.0216397
R31707 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 0.0107679
R31708 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.0107679
R31709 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 179.256
R31710 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 168.089
R31711 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 150.293
R31712 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 73.6304
R31713 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 60.4568
R31714 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 12.0358
R31715 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.981478
R31716 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 0.788543
R31717 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.769522
R31718 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.720633
R31719 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 0.682565
R31720 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.580578
R31721 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 0.55213
R31722 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 0.470609
R31723 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.447191
R31724 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.428234
R31725 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1255
R31726 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1255
R31727 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 0.063
R31728 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 0.063
R31729 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 0.063
R31730 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 0.063
R31731 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 0.063
R31732 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 0.0435206
R31733 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 0.0107679
R31734 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.0107679
R31735 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 316.762
R31736 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 168.108
R31737 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 150.293
R31738 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 150.273
R31739 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 73.6406
R31740 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 73.6304
R31741 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 60.4568
R31742 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 12.0358
R31743 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 1.19615
R31744 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.981478
R31745 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 0.788543
R31746 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.769522
R31747 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 0.682565
R31748 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.580578
R31749 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 0.55213
R31750 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 0.484875
R31751 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 0.470609
R31752 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.447191
R31753 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.428234
R31754 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.217464
R31755 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R31756 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R31757 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R31758 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 0.063
R31759 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 0.063
R31760 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.063
R31761 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 0.063
R31762 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 0.063
R31763 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 0.0216397
R31764 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.0216397
R31765 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 0.0107679
R31766 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.0107679
R31767 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 169.46
R31768 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 167.809
R31769 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 167.809
R31770 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 167.227
R31771 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 150.293
R31772 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 150.273
R31773 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 73.6406
R31774 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6304
R31775 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 60.3809
R31776 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 12.3891
R31777 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 11.4489
R31778 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 1.38365
R31779 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 1.19615
R31780 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 1.1717
R31781 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.848156
R31782 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 0.447191
R31783 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.38637
R31784 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 0.280391
R31785 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.217464
R31786 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.200143
R31787 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R31788 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R31789 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R31790 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R31791 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 0.0874565
R31792 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 0.063
R31793 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 0.063
R31794 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 0.063
R31795 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R31796 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 0.0107679
R31797 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0107679
R31798 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 169.46
R31799 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 167.809
R31800 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 167.809
R31801 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 167.226
R31802 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 150.273
R31803 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 150.273
R31804 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 73.6406
R31805 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 73.6304
R31806 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 60.4568
R31807 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 12.3891
R31808 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 11.4489
R31809 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.68257
R31810 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 1.38365
R31811 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 1.19615
R31812 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 1.1717
R31813 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.08448
R31814 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.932141
R31815 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 0.720633
R31816 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 0.280391
R31817 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.217464
R31818 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R31819 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R31820 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R31821 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 0.0874565
R31822 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 0.063
R31823 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.063
R31824 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 0.063
R31825 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 0.063
R31826 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 0.0435206
R31827 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 0.0216397
R31828 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.0216397
R31829 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 0.0107679
R31830 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.0107679
R31831 And_Gate_1.B.n0 And_Gate_1.B.t2 179.256
R31832 And_Gate_1.B.n0 And_Gate_1.B.t1 168.089
R31833 And_Gate_1.B.n3 And_Gate_1.B.t3 150.293
R31834 And_Gate_1.B.n5 And_Gate_1.B.t4 73.6304
R31835 Nand_Gate_4.Vout And_Gate_1.B.t0 60.3943
R31836 And_Gate_1.B.n9 And_Gate_1.B.n8 37.3347
R31837 And_Gate_1.B.n2 Nand_Gate_4.Vout 0.981478
R31838 And_Gate_1.B.n2 And_Gate_1.B.n1 0.788543
R31839 And_Gate_1.B.n4 And_Gate_1.Nand_Gate_0.B 0.769522
R31840 And_Gate_1.B.n1 Nand_Gate_4.Vout 0.720633
R31841 And_Gate_1.B.n11 And_Gate_1.B.n10 0.682565
R31842 And_Gate_1.B.n10 Nand_Gate_4.Vout 0.580578
R31843 And_Gate_1.B.n4 And_Gate_1.B.n3 0.55213
R31844 And_Gate_1.B.n7 And_Gate_1.B.n6 0.470609
R31845 And_Gate_1.B.n3 And_Gate_1.Nand_Gate_0.B 0.447191
R31846 And_Gate_1.B.n7 And_Gate_1.Nand_Gate_0.B 0.428234
R31847 And_Gate_1.B.n6 And_Gate_1.Nand_Gate_0.B 0.1255
R31848 And_Gate_1.B.n11 Nand_Gate_4.Vout 0.1255
R31849 And_Gate_1.B.n8 And_Gate_1.B.n4 0.063
R31850 And_Gate_1.B.n8 And_Gate_1.B.n7 0.063
R31851 And_Gate_1.B.n9 And_Gate_1.B.n2 0.063
R31852 And_Gate_1.B.n10 And_Gate_1.B.n9 0.063
R31853 Nand_Gate_4.Vout And_Gate_1.B.n11 0.063
R31854 And_Gate_1.B.n1 And_Gate_1.B.n0 0.0435206
R31855 And_Gate_1.B.n6 And_Gate_1.B.n5 0.0107679
R31856 And_Gate_1.B.n5 And_Gate_1.Nand_Gate_0.B 0.0107679
R31857 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 179.256
R31858 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 168.089
R31859 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 150.293
R31860 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 73.6304
R31861 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 60.3943
R31862 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 12.0358
R31863 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.981478
R31864 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 0.788543
R31865 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.769522
R31866 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 0.720633
R31867 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 0.682565
R31868 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.580578
R31869 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 0.55213
R31870 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 0.470609
R31871 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.447191
R31872 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.428234
R31873 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1255
R31874 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1255
R31875 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 0.063
R31876 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 0.063
R31877 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.063
R31878 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 0.063
R31879 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 0.063
R31880 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 0.0435206
R31881 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 0.0107679
R31882 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.0107679
R31883 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout.t2 169.46
R31884 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout.t3 167.809
R31885 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout.t1 167.809
R31886 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout.t7 167.227
R31887 D_FlipFlop_2.3-input-nand_2.Vout.t7 D_FlipFlop_2.3-input-nand_2.Vout.n2 150.293
R31888 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.t6 150.273
R31889 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout.t4 73.6406
R31890 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout.t5 73.6304
R31891 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.t0 60.3809
R31892 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout.n9 12.3891
R31893 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.n4 11.4489
R31894 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.n11 1.38365
R31895 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout.n1 1.19615
R31896 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.n8 1.1717
R31897 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.Vout.n12 0.848156
R31898 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout 0.447191
R31899 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R31900 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.n3 0.280391
R31901 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout.n5 0.262643
R31902 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout 0.217464
R31903 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R31904 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R31905 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R31906 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R31907 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout.n6 0.0874565
R31908 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout 0.063
R31909 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout.n10 0.063
R31910 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout.n7 0.063
R31911 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R31912 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout.n0 0.0107679
R31913 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout 0.0107679
R31914 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 179.256
R31915 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 168.089
R31916 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 150.293
R31917 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 73.6304
R31918 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 60.3943
R31919 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 12.0358
R31920 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.981478
R31921 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 0.788543
R31922 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.769522
R31923 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 0.720633
R31924 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 0.682565
R31925 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.580578
R31926 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 0.55213
R31927 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 0.470609
R31928 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.447191
R31929 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.428234
R31930 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1255
R31931 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1255
R31932 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 0.063
R31933 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 0.063
R31934 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.063
R31935 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 0.063
R31936 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 0.063
R31937 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 0.0435206
R31938 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 0.0107679
R31939 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.0107679
R31940 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout.t3 169.46
R31941 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout.t2 167.809
R31942 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout.t1 167.809
R31943 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout.t7 167.227
R31944 D_FlipFlop_6.3-input-nand_2.Vout.t7 D_FlipFlop_6.3-input-nand_2.Vout.n2 150.293
R31945 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.t6 150.273
R31946 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout.t4 73.6406
R31947 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout.t5 73.6304
R31948 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.t0 60.3809
R31949 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout.n9 12.3891
R31950 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.n4 11.4489
R31951 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.n11 1.38365
R31952 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout.n1 1.19615
R31953 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.n8 1.1717
R31954 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.Vout.n12 0.848156
R31955 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout 0.447191
R31956 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R31957 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.n3 0.280391
R31958 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout.n5 0.262643
R31959 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout 0.217464
R31960 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R31961 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R31962 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R31963 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R31964 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout.n6 0.0874565
R31965 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout 0.063
R31966 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout.n10 0.063
R31967 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout.n7 0.063
R31968 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R31969 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout.n0 0.0107679
R31970 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout 0.0107679
R31971 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 316.762
R31972 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 168.108
R31973 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 150.293
R31974 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 150.273
R31975 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 73.6406
R31976 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 73.6304
R31977 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 60.4568
R31978 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 12.0358
R31979 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 1.19615
R31980 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.981478
R31981 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 0.788543
R31982 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.769522
R31983 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 0.682565
R31984 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.580578
R31985 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 0.55213
R31986 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 0.484875
R31987 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 0.470609
R31988 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.447191
R31989 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.428234
R31990 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.217464
R31991 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R31992 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R31993 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R31994 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 0.063
R31995 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 0.063
R31996 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.063
R31997 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 0.063
R31998 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 0.063
R31999 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 0.0216397
R32000 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.0216397
R32001 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 0.0107679
R32002 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.0107679
R32003 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 169.46
R32004 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 167.809
R32005 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 167.809
R32006 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 167.227
R32007 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 150.293
R32008 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 150.273
R32009 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 73.6406
R32010 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 73.6304
R32011 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 60.3809
R32012 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 12.3891
R32013 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 11.4489
R32014 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 1.38365
R32015 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 1.19615
R32016 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 1.1717
R32017 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.848156
R32018 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 0.447191
R32019 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.38637
R32020 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 0.280391
R32021 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 0.262643
R32022 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.217464
R32023 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.152844
R32024 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.149957
R32025 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.1255
R32026 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.1255
R32027 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 0.0874565
R32028 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 0.063
R32029 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 0.063
R32030 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.063
R32031 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.0454219
R32032 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 0.0107679
R32033 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.0107679
R32034 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 169.46
R32035 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 167.809
R32036 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 167.809
R32037 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 167.227
R32038 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 150.293
R32039 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 150.273
R32040 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 73.6406
R32041 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 73.6304
R32042 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 60.3809
R32043 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 12.3891
R32044 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 11.4489
R32045 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 1.38365
R32046 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 1.19615
R32047 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 1.1717
R32048 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.848156
R32049 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 0.447191
R32050 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.38637
R32051 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 0.280391
R32052 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 0.262643
R32053 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.217464
R32054 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.152844
R32055 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.149957
R32056 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.1255
R32057 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.1255
R32058 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 0.0874565
R32059 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 0.063
R32060 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 0.063
R32061 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.063
R32062 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.0454219
R32063 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 0.0107679
R32064 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.0107679
R32065 Nand_Gate_6.Vout.n10 Nand_Gate_6.Vout.t0 179.256
R32066 Nand_Gate_6.Vout.n10 Nand_Gate_6.Vout.t2 168.089
R32067 Nand_Gate_6.Vout.n2 Nand_Gate_6.Vout.t3 150.293
R32068 Nand_Gate_6.Vout.n4 Nand_Gate_6.Vout.t4 73.6304
R32069 Nand_Gate_6.Vout Nand_Gate_6.Vout.t1 60.3943
R32070 Nand_Gate_6.Vout.n8 Nand_Gate_6.Vout.n7 37.3347
R32071 Nand_Gate_6.Vout.n9 Nand_Gate_6.Vout 0.981478
R32072 Nand_Gate_6.Vout.n11 Nand_Gate_6.Vout.n9 0.788543
R32073 Nand_Gate_6.Vout.n3 Nand_Gate_6.Vout 0.769522
R32074 Nand_Gate_6.Vout Nand_Gate_6.Vout.n11 0.720633
R32075 Nand_Gate_6.Vout.n1 Nand_Gate_6.Vout.n0 0.682565
R32076 Nand_Gate_6.Vout.n1 Nand_Gate_6.Vout 0.580578
R32077 Nand_Gate_6.Vout.n3 Nand_Gate_6.Vout.n2 0.55213
R32078 Nand_Gate_6.Vout.n6 Nand_Gate_6.Vout.n5 0.470609
R32079 Nand_Gate_6.Vout.n2 Nand_Gate_6.Vout 0.447191
R32080 Nand_Gate_6.Vout.n6 Nand_Gate_6.Vout 0.428234
R32081 Nand_Gate_6.Vout.n5 Nand_Gate_6.Vout 0.1255
R32082 Nand_Gate_6.Vout.n0 Nand_Gate_6.Vout 0.1255
R32083 Nand_Gate_6.Vout.n7 Nand_Gate_6.Vout.n3 0.063
R32084 Nand_Gate_6.Vout.n7 Nand_Gate_6.Vout.n6 0.063
R32085 Nand_Gate_6.Vout.n0 Nand_Gate_6.Vout 0.063
R32086 Nand_Gate_6.Vout.n9 Nand_Gate_6.Vout.n8 0.063
R32087 Nand_Gate_6.Vout.n8 Nand_Gate_6.Vout.n1 0.063
R32088 Nand_Gate_6.Vout.n11 Nand_Gate_6.Vout.n10 0.0435206
R32089 Nand_Gate_6.Vout.n5 Nand_Gate_6.Vout.n4 0.0107679
R32090 Nand_Gate_6.Vout.n4 Nand_Gate_6.Vout 0.0107679
R32091 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 169.46
R32092 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 167.809
R32093 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 167.809
R32094 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 167.227
R32095 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 150.293
R32096 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 150.273
R32097 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 73.6406
R32098 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 73.6304
R32099 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 60.3809
R32100 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 12.3891
R32101 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 11.4489
R32102 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 1.38365
R32103 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 1.19615
R32104 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 1.1717
R32105 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.848156
R32106 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 0.447191
R32107 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.38637
R32108 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 0.280391
R32109 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 0.262643
R32110 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.217464
R32111 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.152844
R32112 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.149957
R32113 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.1255
R32114 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.1255
R32115 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 0.0874565
R32116 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 0.063
R32117 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 0.063
R32118 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.063
R32119 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.0454219
R32120 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 0.0107679
R32121 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.0107679
R32122 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 169.46
R32123 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 167.809
R32124 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 167.809
R32125 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 167.227
R32126 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 150.293
R32127 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 150.273
R32128 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 73.6406
R32129 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 73.6304
R32130 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 60.3809
R32131 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 12.3891
R32132 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 11.4489
R32133 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 1.38365
R32134 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 1.19615
R32135 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 1.1717
R32136 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.848156
R32137 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 0.447191
R32138 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R32139 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 0.280391
R32140 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.217464
R32141 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.200143
R32142 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R32143 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R32144 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R32145 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R32146 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 0.0874565
R32147 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 0.063
R32148 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 0.063
R32149 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 0.063
R32150 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R32151 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 0.0107679
R32152 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0107679
R32153 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 316.762
R32154 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 168.108
R32155 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 150.293
R32156 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 150.273
R32157 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 73.6406
R32158 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 73.6304
R32159 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 60.3943
R32160 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 12.0358
R32161 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 1.19615
R32162 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.981478
R32163 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 0.788543
R32164 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.769522
R32165 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 0.682565
R32166 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.580578
R32167 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 0.55213
R32168 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 0.484875
R32169 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 0.470609
R32170 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.447191
R32171 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.428234
R32172 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.217464
R32173 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R32174 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R32175 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R32176 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 0.063
R32177 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 0.063
R32178 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.063
R32179 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 0.063
R32180 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 0.063
R32181 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 0.0216397
R32182 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.0216397
R32183 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 0.0107679
R32184 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.0107679
R32185 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 316.762
R32186 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 168.108
R32187 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 150.293
R32188 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 150.273
R32189 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 73.6406
R32190 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 73.6304
R32191 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 60.4568
R32192 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 12.0358
R32193 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 1.19615
R32194 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.981478
R32195 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 0.788543
R32196 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.769522
R32197 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 0.682565
R32198 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.580578
R32199 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 0.55213
R32200 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 0.484875
R32201 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 0.470609
R32202 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.447191
R32203 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.428234
R32204 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.217464
R32205 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R32206 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R32207 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R32208 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 0.063
R32209 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 0.063
R32210 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.063
R32211 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 0.063
R32212 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 0.063
R32213 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 0.0216397
R32214 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.0216397
R32215 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 0.0107679
R32216 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.0107679
R32217 Q0.n7 Q0.t1 169.46
R32218 Q0.n9 Q0.t3 167.809
R32219 Q0.n7 Q0.t0 167.809
R32220 Q0 Q0.t9 158.585
R32221 Q0.n13 Q0.t7 150.869
R32222 Q0.n12 Q0.t8 150.869
R32223 Q0.t9 Q0.n2 150.293
R32224 Q0.n14 Q0.n11 137.644
R32225 Q0 Q0.t4 78.1811
R32226 Q0.n12 Q0.t5 74.1352
R32227 Q0.t4 Q0.n13 74.1352
R32228 Q0.n0 Q0.t6 73.6304
R32229 Q0.n5 Q0.t2 60.3809
R32230 Q0.n11 Q0 41.1198
R32231 Q0.n8 Q0.n7 11.4489
R32232 Q0.n10 Q0.n9 4.78039
R32233 Q0.n10 Q0.n4 1.74412
R32234 Q0.n13 Q0.n12 1.66898
R32235 Q0.n6 Q0.n5 1.64452
R32236 Q0.n2 Q0.n1 1.19615
R32237 Q0.n5 Q0 0.848156
R32238 Q0.n2 Q0 0.447191
R32239 Q0.n4 Q0.n3 0.3624
R32240 Q0.n4 Q0 0.333061
R32241 Q0.n9 Q0.n8 0.280391
R32242 Q0.n8 Q0.n6 0.262643
R32243 Q0.n6 Q0 0.1255
R32244 Q0.n1 Q0 0.1255
R32245 Q0.n12 Q0 0.063
R32246 Q0.n6 Q0 0.063
R32247 Q0.n11 Q0.n10 0.0305325
R32248 Q0 Q0.n14 0.0168043
R32249 Q0.n14 Q0 0.0122188
R32250 Q0.n1 Q0.n0 0.0107679
R32251 Q0.n0 Q0 0.0107679
R32252 Q0.n3 Q0 0.00441667
R32253 Q0.n3 Q0 0.00406061
R32254 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 179.256
R32255 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 168.089
R32256 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 150.293
R32257 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 73.6304
R32258 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 60.4568
R32259 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 12.0358
R32260 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.981478
R32261 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 0.788543
R32262 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.769522
R32263 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 0.720633
R32264 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 0.682565
R32265 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.580578
R32266 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 0.55213
R32267 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 0.470609
R32268 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.447191
R32269 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.428234
R32270 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1255
R32271 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1255
R32272 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 0.063
R32273 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 0.063
R32274 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.063
R32275 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 0.063
R32276 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 0.063
R32277 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 0.0435206
R32278 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 0.0107679
R32279 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.0107679
R32280 Vin Vin.t0 467.404
R32281 a_139804_27676.t0 a_139804_27676.n0 25.9955
R32282 a_139804_27676.n0 a_139804_27676.t1 14.4333
R32283 a_139804_27676.n0 a_139804_27676.t2 14.4333
R32284 Nand_Gate_0.B.n6 Nand_Gate_0.B.t3 169.46
R32285 Nand_Gate_0.B.n6 Nand_Gate_0.B.t2 167.809
R32286 Nand_Gate_0.B.n5 Nand_Gate_0.B.t1 167.809
R32287 Nand_Gate_0.B Nand_Gate_0.B.t5 158.585
R32288 Nand_Gate_0.B.t5 Nand_Gate_0.B.n2 150.293
R32289 Nand_Gate_0.B.n28 Nand_Gate_0.B.t4 150.273
R32290 Nand_Gate_0.B.n18 Nand_Gate_0.B.t7 150.273
R32291 Nand_Gate_0.B.n12 Nand_Gate_0.B.t10 150.273
R32292 Nand_Gate_0.B.n16 Nand_Gate_0.B.t6 73.6406
R32293 Nand_Gate_0.B.n10 Nand_Gate_0.B.t9 73.6406
R32294 Nand_Gate_0.B.n25 Nand_Gate_0.B.t8 73.6304
R32295 Nand_Gate_0.B.n0 Nand_Gate_0.B.t11 73.6304
R32296 Nand_Gate_0.B.n34 Nand_Gate_0.B.t0 60.3809
R32297 Nand_Gate_0.B.n29 Nand_Gate_0.B.n28 40.8363
R32298 Nand_Gate_0.B.n7 Nand_Gate_0.B.n6 11.4489
R32299 Nand_Gate_0.B.n5 Nand_Gate_0.B.n4 8.21389
R32300 Nand_Gate_0.B.n22 Nand_Gate_0.B.n15 8.1418
R32301 Nand_Gate_0.B.n24 Nand_Gate_0.B.n23 6.47604
R32302 Nand_Gate_0.B.n23 Nand_Gate_0.B 5.35402
R32303 Nand_Gate_0.B.n32 Nand_Gate_0.B 4.55128
R32304 Nand_Gate_0.B.n22 Nand_Gate_0.B.n21 4.5005
R32305 Nand_Gate_0.B.n2 Nand_Gate_0.B.n1 1.19615
R32306 Nand_Gate_0.B.n27 Nand_Gate_0.B.n26 1.1717
R32307 Nand_Gate_0.B.n33 Nand_Gate_0.B 1.08746
R32308 Nand_Gate_0.B.n24 Nand_Gate_0.B 0.973326
R32309 Nand_Gate_0.B.n27 Nand_Gate_0.B 0.932141
R32310 Nand_Gate_0.B.n17 Nand_Gate_0.B 0.851043
R32311 Nand_Gate_0.B.n11 Nand_Gate_0.B 0.851043
R32312 Nand_Gate_0.B Nand_Gate_0.B.n34 0.848156
R32313 Nand_Gate_0.B.n9 Nand_Gate_0.B.n8 0.788543
R32314 Nand_Gate_0.B.n31 Nand_Gate_0.B.n30 0.755935
R32315 Nand_Gate_0.B.n34 Nand_Gate_0.B.n33 0.682565
R32316 Nand_Gate_0.B.n9 Nand_Gate_0.B 0.65675
R32317 Nand_Gate_0.B.n20 Nand_Gate_0.B.n19 0.55213
R32318 Nand_Gate_0.B.n14 Nand_Gate_0.B.n13 0.55213
R32319 Nand_Gate_0.B.n20 Nand_Gate_0.B 0.486828
R32320 Nand_Gate_0.B.n14 Nand_Gate_0.B 0.486828
R32321 Nand_Gate_0.B.n30 Nand_Gate_0.B 0.48023
R32322 Nand_Gate_0.B.n17 Nand_Gate_0.B.n16 0.470609
R32323 Nand_Gate_0.B.n11 Nand_Gate_0.B.n10 0.470609
R32324 Nand_Gate_0.B.n2 Nand_Gate_0.B 0.447191
R32325 Nand_Gate_0.B.n4 Nand_Gate_0.B.n3 0.425067
R32326 Nand_Gate_0.B.n4 Nand_Gate_0.B 0.39003
R32327 Nand_Gate_0.B.n7 Nand_Gate_0.B.n5 0.280391
R32328 Nand_Gate_0.B.n16 Nand_Gate_0.B 0.217464
R32329 Nand_Gate_0.B.n10 Nand_Gate_0.B 0.217464
R32330 Nand_Gate_0.B Nand_Gate_0.B.n7 0.200143
R32331 Nand_Gate_0.B.n26 Nand_Gate_0.B 0.1255
R32332 Nand_Gate_0.B.n19 Nand_Gate_0.B 0.1255
R32333 Nand_Gate_0.B.n13 Nand_Gate_0.B 0.1255
R32334 Nand_Gate_0.B.n1 Nand_Gate_0.B 0.1255
R32335 Nand_Gate_0.B.n8 Nand_Gate_0.B 0.1255
R32336 Nand_Gate_0.B.n28 Nand_Gate_0.B.n27 0.063
R32337 Nand_Gate_0.B.n21 Nand_Gate_0.B.n17 0.063
R32338 Nand_Gate_0.B.n21 Nand_Gate_0.B.n20 0.063
R32339 Nand_Gate_0.B.n15 Nand_Gate_0.B.n11 0.063
R32340 Nand_Gate_0.B.n15 Nand_Gate_0.B.n14 0.063
R32341 Nand_Gate_0.B.n23 Nand_Gate_0.B.n22 0.063
R32342 Nand_Gate_0.B.n29 Nand_Gate_0.B.n24 0.063
R32343 Nand_Gate_0.B.n30 Nand_Gate_0.B.n29 0.063
R32344 Nand_Gate_0.B.n8 Nand_Gate_0.B 0.063
R32345 Nand_Gate_0.B.n33 Nand_Gate_0.B.n32 0.063
R32346 Nand_Gate_0.B.n32 Nand_Gate_0.B.n9 0.063
R32347 Nand_Gate_0.B.n19 Nand_Gate_0.B.n18 0.0216397
R32348 Nand_Gate_0.B.n18 Nand_Gate_0.B 0.0216397
R32349 Nand_Gate_0.B.n13 Nand_Gate_0.B.n12 0.0216397
R32350 Nand_Gate_0.B.n12 Nand_Gate_0.B 0.0216397
R32351 Nand_Gate_0.B.n31 Nand_Gate_0.B 0.0168043
R32352 Nand_Gate_0.B Nand_Gate_0.B.n31 0.0122188
R32353 Nand_Gate_0.B.n26 Nand_Gate_0.B.n25 0.0107679
R32354 Nand_Gate_0.B.n25 Nand_Gate_0.B 0.0107679
R32355 Nand_Gate_0.B.n1 Nand_Gate_0.B.n0 0.0107679
R32356 Nand_Gate_0.B.n0 Nand_Gate_0.B 0.0107679
R32357 Nand_Gate_0.B.n3 Nand_Gate_0.B 0.00441667
R32358 Nand_Gate_0.B.n3 Nand_Gate_0.B 0.00406061
R32359 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 169.46
R32360 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 168.089
R32361 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 167.809
R32362 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 150.293
R32363 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 73.6304
R32364 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 60.3943
R32365 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 12.0358
R32366 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 11.4489
R32367 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.981478
R32368 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 0.788543
R32369 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.769522
R32370 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 0.720633
R32371 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 0.682565
R32372 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.580578
R32373 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 0.55213
R32374 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 0.470609
R32375 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.447191
R32376 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.428234
R32377 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.1255
R32378 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.1255
R32379 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 0.063
R32380 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 0.063
R32381 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.063
R32382 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 0.063
R32383 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 0.063
R32384 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 0.0435206
R32385 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 0.0107679
R32386 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.0107679
R32387 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 169.46
R32388 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 168.089
R32389 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 167.809
R32390 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 150.293
R32391 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 73.6304
R32392 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 60.4568
R32393 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 12.0358
R32394 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 11.4489
R32395 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.981478
R32396 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 0.788543
R32397 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.769522
R32398 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 0.720633
R32399 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 0.682565
R32400 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.580578
R32401 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 0.55213
R32402 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 0.470609
R32403 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.447191
R32404 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.428234
R32405 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.1255
R32406 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.1255
R32407 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 0.063
R32408 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 0.063
R32409 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.063
R32410 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 0.063
R32411 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 0.063
R32412 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 0.0435206
R32413 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 0.0107679
R32414 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.0107679
R32415 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 169.46
R32416 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 168.089
R32417 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 167.809
R32418 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 150.273
R32419 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 73.6406
R32420 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 60.3809
R32421 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 12.0358
R32422 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 11.4489
R32423 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 1.08746
R32424 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.851043
R32425 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.848156
R32426 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 0.788543
R32427 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 0.682565
R32428 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.65675
R32429 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 0.55213
R32430 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.486828
R32431 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 0.470609
R32432 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 0.262643
R32433 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.217464
R32434 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.1255
R32435 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.1255
R32436 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 0.063
R32437 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 0.063
R32438 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 0.063
R32439 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 0.063
R32440 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 0.063
R32441 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 0.0216397
R32442 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.0216397
R32443 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 169.46
R32444 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 168.089
R32445 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 167.809
R32446 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 150.293
R32447 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 73.6304
R32448 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 60.4568
R32449 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 12.0358
R32450 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 11.4489
R32451 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.981478
R32452 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 0.788543
R32453 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.769522
R32454 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 0.720633
R32455 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 0.682565
R32456 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.580578
R32457 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 0.55213
R32458 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 0.470609
R32459 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.447191
R32460 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.428234
R32461 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.1255
R32462 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.1255
R32463 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 0.063
R32464 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 0.063
R32465 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.063
R32466 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 0.063
R32467 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 0.063
R32468 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 0.0435206
R32469 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 0.0107679
R32470 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.0107679
R32471 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 169.46
R32472 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 168.089
R32473 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 167.809
R32474 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 150.273
R32475 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 73.6406
R32476 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 60.3809
R32477 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 12.0358
R32478 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 11.4489
R32479 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 1.08746
R32480 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.851043
R32481 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.848156
R32482 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 0.788543
R32483 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 0.682565
R32484 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.65675
R32485 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 0.55213
R32486 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.486828
R32487 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 0.470609
R32488 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 0.262643
R32489 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.217464
R32490 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.1255
R32491 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.1255
R32492 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 0.063
R32493 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 0.063
R32494 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 0.063
R32495 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 0.063
R32496 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 0.063
R32497 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 0.0216397
R32498 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0216397
R32499 And_Gate_0.B.n10 And_Gate_0.B.t0 179.256
R32500 And_Gate_0.B.n10 And_Gate_0.B.t1 168.089
R32501 And_Gate_0.B.n2 And_Gate_0.B.t3 150.293
R32502 And_Gate_0.B.n4 And_Gate_0.B.t4 73.6304
R32503 Nand_Gate_7.Vout And_Gate_0.B.t2 60.3943
R32504 And_Gate_0.B.n8 And_Gate_0.B.n7 37.3347
R32505 And_Gate_0.B.n9 Nand_Gate_7.Vout 0.981478
R32506 And_Gate_0.B.n11 And_Gate_0.B.n9 0.788543
R32507 And_Gate_0.B.n3 And_Gate_0.Nand_Gate_0.B 0.769522
R32508 Nand_Gate_7.Vout And_Gate_0.B.n11 0.720633
R32509 And_Gate_0.B.n1 And_Gate_0.B.n0 0.682565
R32510 And_Gate_0.B.n1 Nand_Gate_7.Vout 0.580578
R32511 And_Gate_0.B.n3 And_Gate_0.B.n2 0.55213
R32512 And_Gate_0.B.n6 And_Gate_0.B.n5 0.470609
R32513 And_Gate_0.B.n2 And_Gate_0.Nand_Gate_0.B 0.447191
R32514 And_Gate_0.B.n6 And_Gate_0.Nand_Gate_0.B 0.428234
R32515 And_Gate_0.B.n5 And_Gate_0.Nand_Gate_0.B 0.1255
R32516 And_Gate_0.B.n0 Nand_Gate_7.Vout 0.1255
R32517 And_Gate_0.B.n7 And_Gate_0.B.n3 0.063
R32518 And_Gate_0.B.n7 And_Gate_0.B.n6 0.063
R32519 And_Gate_0.B.n0 Nand_Gate_7.Vout 0.063
R32520 And_Gate_0.B.n9 And_Gate_0.B.n8 0.063
R32521 And_Gate_0.B.n8 And_Gate_0.B.n1 0.063
R32522 And_Gate_0.B.n11 And_Gate_0.B.n10 0.0435206
R32523 And_Gate_0.B.n5 And_Gate_0.B.n4 0.0107679
R32524 And_Gate_0.B.n4 And_Gate_0.Nand_Gate_0.B 0.0107679
R32525 a_139663_37417.n0 a_139663_37417.t3 1302.5
R32526 a_139663_37417.n0 a_139663_37417.t0 1301.07
R32527 a_139663_37417.n1 a_139663_37417.t2 30.7707
R32528 a_139663_37417.t1 a_139663_37417.n1 18.2748
R32529 a_139663_37417.n1 a_139663_37417.n0 0.340816
R32530 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 169.46
R32531 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 167.809
R32532 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 167.809
R32533 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 167.226
R32534 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 150.273
R32535 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 150.273
R32536 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 73.6406
R32537 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 73.6304
R32538 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 60.3943
R32539 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 12.3891
R32540 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 11.4489
R32541 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 1.68257
R32542 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 1.38365
R32543 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 1.19615
R32544 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 1.1717
R32545 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 1.08448
R32546 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.932141
R32547 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.720633
R32548 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 0.280391
R32549 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.217464
R32550 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R32551 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R32552 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R32553 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 0.0874565
R32554 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 0.063
R32555 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.063
R32556 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 0.063
R32557 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 0.063
R32558 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 0.0435206
R32559 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 0.0216397
R32560 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 0.0216397
R32561 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 0.0107679
R32562 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.0107679
R32563 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 179.256
R32564 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 168.089
R32565 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 150.293
R32566 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 73.6304
R32567 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 60.3943
R32568 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 12.0358
R32569 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.981478
R32570 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 0.788543
R32571 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.769522
R32572 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 0.720633
R32573 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 0.682565
R32574 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.580578
R32575 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 0.55213
R32576 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 0.470609
R32577 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.447191
R32578 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.428234
R32579 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1255
R32580 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1255
R32581 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 0.063
R32582 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 0.063
R32583 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.063
R32584 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 0.063
R32585 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 0.063
R32586 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 0.0435206
R32587 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 0.0107679
R32588 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.0107679
R32589 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 169.46
R32590 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R32591 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 167.809
R32592 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 167.226
R32593 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 150.273
R32594 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 150.273
R32595 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 73.6406
R32596 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 73.6304
R32597 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 60.3943
R32598 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 12.3891
R32599 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 11.4489
R32600 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 1.68257
R32601 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 1.38365
R32602 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 1.19615
R32603 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 1.1717
R32604 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 1.08448
R32605 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.932141
R32606 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.720633
R32607 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 0.280391
R32608 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.217464
R32609 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R32610 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R32611 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R32612 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 0.0874565
R32613 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 0.063
R32614 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.063
R32615 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 0.063
R32616 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 0.063
R32617 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 0.0435206
R32618 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 0.0216397
R32619 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 0.0216397
R32620 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 0.0107679
R32621 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.0107679
C0 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_119711_49858# 0.04543f
C1 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout VDD 2.07863f
C2 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.1182f
C3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_66483_15797# 0.01335f
C4 D_FlipFlop_3.3-input-nand_2.Vout a_132311_40571# 0.04443f
C5 D_FlipFlop_1.Qbar Q6 0.01194f
C6 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.04107f
C7 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.06935f
C8 D_FlipFlop_6.Inverter_1.Vout VDD 1.73058f
C9 FFCLR D_FlipFlop_7.Nand_Gate_1.Vout 0.61318f
C10 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_76165_49858# 0.04444f
C11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout VDD 2.88547f
C12 Nand_Gate_2.Vout EN 0.11847f
C13 a_101705_49858# VDD 0.06015f
C14 a_134897_24200# VDD 0.01186f
C15 D_FlipFlop_3.Qbar a_128237_43285# 0.04443f
C16 D_FlipFlop_0.3-input-nand_1.B VDD 1.32602f
C17 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout CLK 0.03574f
C18 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.0846f
C19 D_FlipFlop_0.Nand_Gate_1.Vout a_130209_44135# 0.05964f
C20 Nand_Gate_2.A a_134897_40571# 0.0468f
C21 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_118967_15797# 0.04443f
C22 Nand_Gate_5.B RingCounter_0.D_FlipFlop_10.3-input-nand_1.B 0.29683f
C23 Nand_Gate_5.B RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.08377f
C24 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_45147_49858# 0.04443f
C25 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1541f
C26 a_52113_49858# EN 0.01149f
C27 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B EN 0.26843f
C28 a_134283_37007# a_134897_37007# 0.05935f
C29 FFCLR RingCounter_0.D_FlipFlop_1.3-input-nand_1.B 0.29683f
C30 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout EN 1.0224f
C31 D_FlipFlop_4.Inverter_1.Vout VDD 1.73058f
C32 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.30154f
C33 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C VDD 3.61245f
C34 a_128237_46849# a_128851_46849# 0.05935f
C35 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_2.Vout 0.92942f
C36 D_FlipFlop_0.Qbar D_FlipFlop_0.Nand_Gate_0.Vout 0.07122f
C37 CDAC8_0.switch_2.Z Q1 0.50863f
C38 D_FlipFlop_1.Qbar Comparator_0.Vinm 0.01573f
C39 a_45761_15797# CLK 0.04619f
C40 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 1.09975f
C41 Nand_Gate_0.B a_80239_49858# 0.04741f
C42 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout EN 0.78685f
C43 a_44403_15797# VDD 0.03339f
C44 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B a_78881_13083# 0.04443f
C45 a_128237_20636# a_128851_20636# 0.05935f
C46 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.3-input-nand_2.C 0.26069f
C47 a_59605_47663# CLK 0.04443f
C48 a_48937_47663# VDD 0.02521f
C49 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C VDD 3.56545f
C50 D_FlipFlop_4.Nand_Gate_0.Vout a_130209_30478# 0.05964f
C51 Nand_Gate_6.B Q0 0.06521f
C52 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.25963f
C53 D_FlipFlop_7.Nand_Gate_1.Vout a_128851_17072# 0.04995f
C54 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_2.Vout 0.92857f
C55 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B CLK 0.16166f
C56 a_84619_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.01335f
C57 Nand_Gate_5.A Comparator_0.Vinm 1.94937f
C58 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout EN 0.13192f
C59 D_FlipFlop_1.3-input-nand_1.Vout a_132311_33443# 0.04444f
C60 RingCounter_0.D_FlipFlop_3.Qbar a_80239_52572# 0.04443f
C61 D_FlipFlop_0.3-input-nand_1.Vout VDD 1.78032f
C62 a_128237_24200# a_128851_24200# 0.05935f
C63 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_74807_15797# 0.04443f
C64 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B a_45761_13083# 0.04443f
C65 a_132925_46849# VDD 0.01186f
C66 VDD Q2 3.59925f
C67 a_57545_49858# VDD 0.06015f
C68 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_123785_49858# 0.04995f
C69 D_FlipFlop_0.3-input-nand_2.C a_132925_44135# 0.01335f
C70 RingCounter_0.D_FlipFlop_8.Qbar a_39715_13083# 0.06113f
C71 EN Q5 0.2481f
C72 CDAC8_0.switch_8.Z Q4 0.5562f
C73 a_90535_13083# VDD 0.01327f
C74 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_110029_15797# 0.04444f
C75 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_80239_49858# 0.04444f
C76 Nand_Gate_0.B a_85233_52572# 0.04443f
C77 D_FlipFlop_3.3-input-nand_0.Vout VDD 1.77946f
C78 CDAC8_0.switch_0.Z CDAC8_0.switch_2.Z 0.1201f
C79 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout EN 0.08852f
C80 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B a_123655_13083# 0.04995f
C81 a_128237_27764# a_128851_27764# 0.05935f
C82 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B VDD 1.66713f
C83 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_43045_52572# 0.04443f
C84 a_123041_15797# a_123655_15797# 0.05935f
C85 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_121683_15797# 0.04995f
C86 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_7.Inverter_1.Vout 0.01422f
C87 a_75898_39392# CDAC8_0.switch_6.Z 0.29129f
C88 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C VDD 3.54707f
C89 a_130209_39721# VDD 0.02521f
C90 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_43789_15797# 0.04443f
C91 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout VDD 2.46653f
C92 CDAC8_0.switch_7.Z Q3 1.50848f
C93 Nand_Gate_7.B a_72835_15797# 0.06113f
C94 CDAC8_0.switch_5.Z CDAC8_0.switch_0.Z 0.09134f
C95 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.Vout 0.01194f
C96 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.C 0.01194f
C97 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout VDD 1.60037f
C98 a_124399_49858# VDD 0.02521f
C99 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout EN 1.03583f
C100 Nand_Gate_6.B Nand_Gate_4.B 0.062f
C101 Nand_Gate_7.B VDD 8.03863f
C102 Nand_Gate_1.A VDD 4.17892f
C103 a_128237_43285# a_128851_43285# 0.05935f
C104 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B a_84619_49858# 0.04995f
C105 a_98989_15797# VDD 0.03178f
C106 D_FlipFlop_3.Qbar D_FlipFlop_3.Nand_Gate_0.Vout 0.07122f
C107 Nand_Gate_1.A a_100961_15797# 0.04443f
C108 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_30647_15797# 0.04443f
C109 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_118967_13083# 0.04443f
C110 Nand_Gate_5.A a_134897_44135# 0.0468f
C111 Nand_Gate_5.B Q5 0.06203f
C112 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout CLK 0.30735f
C113 RingCounter_0.D_FlipFlop_12.Qbar a_84489_13083# 0.01335f
C114 a_50755_15797# a_51369_15797# 0.05935f
C115 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_75551_49858# 0.01335f
C116 a_84489_15797# VDD 0.01571f
C117 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_109285_52572# 0.04443f
C118 a_75898_18814# VDD 1.34284f
C119 D_FlipFlop_7.3-input-nand_0.Vout a_134283_19786# 0.05964f
C120 a_57545_52572# EN 0.04443f
C121 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.3-input-nand_2.C 0.26069f
C122 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B CLK 0.16274f
C123 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout a_122427_52572# 0.04443f
C124 D_FlipFlop_0.Nand_Gate_0.Vout a_128851_46849# 0.04995f
C125 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout CLK 0.29759f
C126 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.3-input-nand_2.Vout 0.16429f
C127 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout VDD 2.31704f
C128 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_83875_15797# 0.04444f
C129 a_57415_15797# VDD 0.06072f
C130 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B EN 0.26843f
C131 D_FlipFlop_2.3-input-nand_0.Vout a_132311_39721# 0.04444f
C132 a_46375_13083# VDD 0.01327f
C133 a_78881_15797# a_79495_15797# 0.05935f
C134 D_FlipFlop_0.CLK D_FlipFlop_0.Qbar 0.10195f
C135 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout CLK 0.23566f
C136 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_77523_15797# 0.04995f
C137 a_105955_13083# a_106569_13083# 0.05935f
C138 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD 1.56255f
C139 a_109285_52572# VDD 0.02521f
C140 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B a_74193_49858# 0.04443f
C141 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout a_118967_15797# 0.04443f
C142 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_43789_13083# 0.04443f
C143 D_FlipFlop_5.Qbar VDD 1.89808f
C144 RingCounter_0.D_FlipFlop_16.Q CDAC8_0.switch_7.Z 0.08064f
C145 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_46375_15797# 0.01335f
C146 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_0.Vout 1.03544f
C147 Nand_Gate_0.B RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.08524f
C148 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.3-input-nand_2.C 0.26069f
C149 a_132925_17072# VDD 0.01186f
C150 Nand_Gate_4.B a_45761_15797# 0.04443f
C151 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.3-input-nand_2.Vout 0.16429f
C152 Nand_Gate_0.A D_FlipFlop_2.Nand_Gate_0.Vout 0.65009f
C153 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Qbar 0.07122f
C154 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_80239_52572# 0.04444f
C155 FFCLR a_134897_36157# 0.04581f
C156 CLK Q0 1.75855f
C157 a_80239_49858# VDD 0.02906f
C158 D_FlipFlop_0.Nand_Gate_1.Vout VDD 1.46545f
C159 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.16429f
C160 CDAC8_0.switch_6.Z CDAC8_0.switch_5.Z 3.08882f
C161 D_FlipFlop_0.3-input-nand_1.Vout a_132925_44135# 0.04543f
C162 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout a_76165_49858# 0.04443f
C163 a_116995_13083# VDD 0.02521f
C164 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.3-input-nand_2.C 0.26069f
C165 Nand_Gate_0.B a_71017_47663# 0.04443f
C166 Nand_Gate_0.A CDAC8_0.switch_7.Z 7.14466f
C167 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C EN 0.07664f
C168 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C EN 0.07732f
C169 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout VDD 2.74107f
C170 FFCLR RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.08377f
C171 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_67227_49858# 0.04443f
C172 a_128237_40571# VDD 0.02521f
C173 CDAC8_0.switch_1.Z Q0 0.17328f
C174 RingCounter_0.D_FlipFlop_3.Qbar CLK 0.09276f
C175 RingCounter_0.D_FlipFlop_9.Qbar CLK 0.09276f
C176 a_34721_15797# a_35335_15797# 0.05935f
C177 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_33363_15797# 0.04995f
C178 RingCounter_0.D_FlipFlop_15.Qbar CLK 0.09276f
C179 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_54829_15797# 0.04443f
C180 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout a_74807_15797# 0.04443f
C181 a_91279_52572# Nand_Gate_2.A 0.06113f
C182 a_128237_19786# VDD 0.02521f
C183 D_FlipFlop_1.Qbar EN 0.04711f
C184 a_132311_39721# VDD 0.02521f
C185 a_83875_13083# a_84489_13083# 0.05935f
C186 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.08641f
C187 D_FlipFlop_3.Nand_Gate_1.Vout a_128237_40571# 0.04444f
C188 Nand_Gate_5.A a_115177_47663# 0.04443f
C189 D_FlipFlop_3.3-input-nand_2.C a_132311_40571# 0.05964f
C190 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B a_41073_49858# 0.04443f
C191 D_FlipFlop_7.3-input-nand_1.Vout a_132311_17072# 0.04444f
C192 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK 0.29644f
C193 And_Gate_3.Nand_Gate_0.Vout CLK 0.49672f
C194 RingCounter_0.D_FlipFlop_4.Qbar a_91279_49858# 0.06113f
C195 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout a_63767_13083# 0.04995f
C196 a_85233_52572# VDD 0.02521f
C197 a_75898_46095# Comparator_0.Vinm 0.04537f
C198 a_119711_52572# a_120325_52572# 0.05935f
C199 D_FlipFlop_7.Qbar a_128237_19786# 0.04443f
C200 D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.48313f
C201 D_FlipFlop_3.Nand_Gate_0.Vout a_128851_43285# 0.04995f
C202 a_130209_44135# VDD 0.02521f
C203 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_98245_52572# 0.04444f
C204 Nand_Gate_3.B Comparator_0.Vinm 0.03473f
C205 RingCounter_0.D_FlipFlop_15.Qbar a_50755_13083# 0.06113f
C206 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD 2.04843f
C207 Nand_Gate_5.A EN 0.49283f
C208 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_2.3-input-nand_0.Vout 0.01418f
C209 Nand_Gate_4.B CLK 0.53838f
C210 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout EN 0.78734f
C211 CDAC8_0.switch_9.Z Q5 0.65512f
C212 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_87949_15797# 0.05964f
C213 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_85233_49858# 0.05964f
C214 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_2.C 0.11436f
C215 a_72835_13083# VDD 0.02521f
C216 a_134283_43285# VDD 0.02521f
C217 Nand_Gate_0.B VDD 4.34021f
C218 CDAC8_0.switch_1.Z Nand_Gate_4.B 1.47073f
C219 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.08671f
C220 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout a_30647_15797# 0.04443f
C221 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1541f
C222 Nand_Gate_6.A EN 0.42008f
C223 D_FlipFlop_1.Qbar a_128237_33443# 0.06113f
C224 D_FlipFlop_6.Nand_Gate_1.Vout a_128851_20636# 0.04995f
C225 a_53471_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.01335f
C226 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.26069f
C227 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_90665_52572# 0.04995f
C228 Nand_Gate_4.B a_50755_13083# 0.04443f
C229 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B a_35335_13083# 0.04995f
C230 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.08641f
C231 Nand_Gate_5.A RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.08514f
C232 a_128851_19786# Q0 0.01335f
C233 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout a_67227_52572# 0.04443f
C234 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.04107f
C235 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_2.C 0.1129f
C236 Nand_Gate_2.A D_FlipFlop_3.Nand_Gate_0.Vout 0.65077f
C237 a_117739_49858# a_118353_49858# 0.05935f
C238 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.30154f
C239 a_107313_49858# CLK 0.04619f
C240 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.06935f
C241 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.16429f
C242 a_61795_13083# a_62409_13083# 0.05935f
C243 a_106699_49858# VDD 0.01712f
C244 Nand_Gate_5.A Nand_Gate_5.B 0.13955f
C245 D_FlipFlop_1.3-input-nand_1.B a_134283_33443# 0.04443f
C246 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C EN 0.07664f
C247 And_Gate_3.Nand_Gate_0.Vout Q0 0.05258f
C248 And_Gate_2.Nand_Gate_0.Vout EN 0.01805f
C249 D_FlipFlop_5.Nand_Gate_1.Vout a_128851_24200# 0.04995f
C250 RingCounter_0.D_FlipFlop_16.Qbar RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.11654f
C251 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B EN 0.43162f
C252 CLK Q4 0.11898f
C253 Nand_Gate_7.A EN 0.42008f
C254 Nand_Gate_2.A CDAC8_0.switch_6.Z 3.68553f
C255 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout EN 0.06649f
C256 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout VDD 2.16852f
C257 Nand_Gate_4.B Q0 1.41286f
C258 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_30647_13083# 0.04443f
C259 D_FlipFlop_3.3-input-nand_1.Vout VDD 1.78032f
C260 D_FlipFlop_6.3-input-nand_2.Vout VDD 2.77266f
C261 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.04109f
C262 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout CLK 0.03479f
C263 a_78267_52572# VDD 0.02521f
C264 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B CLK 0.16274f
C265 Nand_Gate_7.A a_62409_15797# 0.01335f
C266 D_FlipFlop_4.Nand_Gate_1.Vout a_128851_27764# 0.04995f
C267 FFCLR Nand_Gate_0.A 0.92681f
C268 a_28675_13083# VDD 0.02521f
C269 a_46375_15797# VDD 0.06072f
C270 a_101705_52572# VDD 0.01186f
C271 a_81685_47663# CLK 0.07396f
C272 D_FlipFlop_2.3-input-nand_0.Vout VDD 1.77946f
C273 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout CLK 0.23566f
C274 a_71017_47663# VDD 0.02521f
C275 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_108671_52572# 0.04995f
C276 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_43789_15797# 0.05964f
C277 a_54085_52572# VDD 0.02521f
C278 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Qbar 1.05791f
C279 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B a_95659_49858# 0.04995f
C280 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_89307_49858# 0.05964f
C281 D_FlipFlop_4.3-input-nand_2.Vout VDD 2.77266f
C282 Nand_Gate_0.A D_FlipFlop_2.Inverter_1.Vout 0.16179f
C283 Nand_Gate_4.B a_128851_19786# 0.04685f
C284 D_FlipFlop_1.3-input-nand_1.Vout a_134283_33443# 0.05964f
C285 a_95659_49858# a_96273_49858# 0.05935f
C286 a_63153_49858# CLK 0.04619f
C287 a_130209_36157# VDD 0.02521f
C288 Nand_Gate_1.Vout EN 0.10633f
C289 a_39715_13083# a_40329_13083# 0.05935f
C290 a_62539_49858# VDD 0.01712f
C291 RingCounter_0.D_FlipFlop_16.Q a_40459_52572# 0.04995f
C292 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.C 1.09975f
C293 a_128237_43285# Q5 0.06113f
C294 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_76909_13083# 0.05964f
C295 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout CLK 0.23566f
C296 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout EN 0.06649f
C297 a_95529_13083# VDD 0.0563f
C298 FFCLR a_134897_23350# 0.08436f
C299 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_112001_15797# 0.05964f
C300 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.30154f
C301 Nand_Gate_7.B a_132925_23350# 0.0478f
C302 a_64511_52572# a_65125_52572# 0.05935f
C303 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.08641f
C304 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_87205_49858# 0.05964f
C305 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout a_78267_52572# 0.04443f
C306 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.08671f
C307 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout a_111387_49858# 0.04995f
C308 a_55443_15797# EN 0.045f
C309 a_95659_52572# a_96273_52572# 0.05935f
C310 And_Gate_6.Nand_Gate_0.Vout a_103765_47663# 0.05964f
C311 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C VDD 3.61245f
C312 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_123655_15797# 0.01335f
C313 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout EN 0.09127f
C314 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.04107f
C315 FFCLR a_134897_30478# 0.08435f
C316 a_65869_15797# a_66483_15797# 0.05935f
C317 a_72835_15797# VDD 0.02906f
C318 Nand_Gate_6.B a_132925_26914# 0.04784f
C319 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout EN 0.06649f
C320 And_Gate_5.Nand_Gate_0.Vout VDD 1.43186f
C321 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B EN 0.26843f
C322 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.08671f
C323 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout EN 0.97979f
C324 Comparator_0.Vinm Q2 1.64425f
C325 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Qbar 0.07122f
C326 a_100961_15797# VDD 0.03119f
C327 Nand_Gate_1.A RingCounter_0.D_FlipFlop_11.3-input-nand_1.B 0.2969f
C328 RingCounter_0.D_FlipFlop_7.Qbar a_112745_49858# 0.01335f
C329 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121683_13083# 0.01335f
C330 Nand_Gate_1.A RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.08377f
C331 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B CLK 0.16166f
C332 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_98989_15797# 0.04444f
C333 a_130209_26914# VDD 0.02521f
C334 FFCLR D_FlipFlop_7.3-input-nand_0.Vout 0.1263f
C335 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout CLK 0.03479f
C336 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_78267_49858# 0.04443f
C337 D_FlipFlop_0.3-input-nand_1.B a_134897_44135# 0.04995f
C338 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout VDD 2.07863f
C339 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout CLK 0.1215f
C340 a_73579_49858# a_74193_49858# 0.05935f
C341 D_FlipFlop_7.Qbar VDD 1.89473f
C342 Nand_Gate_4.A a_34721_15797# 0.04443f
C343 Nand_Gate_3.B EN 0.99738f
C344 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.06935f
C345 D_FlipFlop_7.Nand_Gate_0.Vout Q0 0.1147f
C346 D_FlipFlop_3.Nand_Gate_1.Vout VDD 1.46545f
C347 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout CLK 0.03342f
C348 CDAC8_0.switch_7.Z CDAC8_0.switch_5.Z 3.08191f
C349 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.25963f
C350 a_45147_52572# VDD 0.02865f
C351 a_51369_13083# VDD 0.0563f
C352 D_FlipFlop_2.3-input-nand_0.Vout a_134283_39721# 0.05964f
C353 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_79495_15797# 0.01335f
C354 a_128851_30478# Q3 0.01335f
C355 RingCounter_0.D_FlipFlop_13.Qbar RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.11654f
C356 Nand_Gate_2.A a_96273_52572# 0.04443f
C357 D_FlipFlop_6.3-input-nand_1.Vout a_132311_20636# 0.04444f
C358 RingCounter_0.D_FlipFlop_4.Qbar Nand_Gate_2.A 1.10693f
C359 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout EN 0.08852f
C360 a_128237_37007# VDD 0.02521f
C361 RingCounter_0.D_FlipFlop_5.Qbar a_102319_49858# 0.06113f
C362 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_118967_15797# 0.05964f
C363 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.1182f
C364 D_FlipFlop_3.3-input-nand_1.B D_FlipFlop_3.3-input-nand_1.Vout 0.08641f
C365 a_112001_15797# a_112615_15797# 0.05935f
C366 Nand_Gate_7.B Comparator_0.Vinm 2.56398f
C367 Nand_Gate_2.A D_FlipFlop_3.Inverter_1.Vout 0.16207f
C368 Nand_Gate_4.B RingCounter_0.D_FlipFlop_8.3-input-nand_1.B 0.2969f
C369 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.C 1.09975f
C370 a_134897_17072# VDD 0.01186f
C371 D_FlipFlop_7.Nand_Gate_0.Vout a_128851_19786# 0.04995f
C372 a_86591_49858# CLK 0.03129f
C373 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout VDD 2.46653f
C374 Nand_Gate_5.A a_113359_49858# 0.04741f
C375 a_85233_49858# VDD 0.0325f
C376 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.07084f
C377 a_132311_36157# VDD 0.02521f
C378 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C CLK 0.30966f
C379 D_FlipFlop_5.3-input-nand_1.Vout a_132311_24200# 0.04444f
C380 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout EN 1.03583f
C381 Nand_Gate_1.B Q3 0.25213f
C382 a_75898_18814# Comparator_0.Vinm 0.0277f
C383 D_FlipFlop_0.3-input-nand_1.Vout a_134897_44135# 0.01335f
C384 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout VDD 2.73822f
C385 a_41687_15797# VDD 0.02906f
C386 a_121069_13083# CLK 0.03129f
C387 D_FlipFlop_1.3-input-nand_2.Vout a_132925_36157# 0.01335f
C388 Nand_Gate_4.B a_37897_16975# 0.04443f
C389 D_FlipFlop_3.Nand_Gate_0.Vout Q5 0.11443f
C390 a_118967_13083# VDD 0.02578f
C391 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.C 1.09975f
C392 a_130209_40571# VDD 0.02521f
C393 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.30154f
C394 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C VDD 3.56545f
C395 a_51499_49858# a_52113_49858# 0.05935f
C396 D_FlipFlop_2.3-input-nand_2.Vout a_132311_37007# 0.04443f
C397 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_35335_15797# 0.01335f
C398 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.04107f
C399 D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_4.B 0.66906f
C400 D_FlipFlop_4.3-input-nand_1.Vout a_132311_27764# 0.04444f
C401 CDAC8_0.switch_6.Z Q5 0.58263f
C402 a_79625_52572# EN 0.04443f
C403 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout EN 0.62384f
C404 D_FlipFlop_2.Qbar a_128237_39721# 0.04443f
C405 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1541f
C406 D_FlipFlop_1.Qbar D_FlipFlop_1.Nand_Gate_1.Vout 0.11654f
C407 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_74807_15797# 0.05964f
C408 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_54085_52572# 0.04443f
C409 Nand_Gate_4.A a_39715_13083# 0.04443f
C410 D_FlipFlop_7.Inverter_1.Vout VDD 1.73058f
C411 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_3.Inverter_1.Vout 0.01422f
C412 a_134283_39721# VDD 0.02521f
C413 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.C 1.09975f
C414 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout CLK 0.71127f
C415 RingCounter_0.D_FlipFlop_11.Qbar RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.07122f
C416 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.30154f
C417 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout CLK 0.30735f
C418 D_FlipFlop_3.Nand_Gate_1.Vout a_130209_40571# 0.05964f
C419 Nand_Gate_5.A D_FlipFlop_0.Qbar 0.06453f
C420 Nand_Gate_5.Vout VDD 1.47723f
C421 D_FlipFlop_7.3-input-nand_1.Vout a_134283_17072# 0.05964f
C422 a_117609_15797# VDD 0.01571f
C423 a_132311_33443# a_132925_33443# 0.05935f
C424 a_120325_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.05964f
C425 FFCLR D_FlipFlop_3.Qbar 0.03748f
C426 a_132925_44135# VDD 0.01186f
C427 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.06955f
C428 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout EN 0.78734f
C429 D_FlipFlop_7.3-input-nand_2.C a_130209_17072# 0.04443f
C430 FFCLR D_FlipFlop_5.3-input-nand_1.B 0.44757f
C431 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_51499_49858# 0.01335f
C432 a_128237_23350# Q1 0.06113f
C433 a_132311_26914# VDD 0.02521f
C434 a_42431_49858# CLK 0.03129f
C435 FFCLR a_47119_49858# 0.04741f
C436 a_41073_49858# VDD 0.02521f
C437 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout VDD 2.88547f
C438 a_76909_13083# CLK 0.03129f
C439 Nand_Gate_6.B a_89921_15797# 0.04443f
C440 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_87205_49858# 0.04444f
C441 D_FlipFlop_3.3-input-nand_1.B VDD 1.32602f
C442 a_101705_52572# Nand_Gate_2.B 0.01335f
C443 a_74807_13083# VDD 0.02578f
C444 D_FlipFlop_6.3-input-nand_2.C VDD 2.74431f
C445 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.08671f
C446 Nand_Gate_2.A CDAC8_0.switch_7.Z 7.18772f
C447 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C EN 0.07732f
C448 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_30647_15797# 0.05964f
C449 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_108671_49858# 0.01335f
C450 RingCounter_0.D_FlipFlop_5.Qbar CLK 0.09276f
C451 D_FlipFlop_2.3-input-nand_1.Vout VDD 1.78032f
C452 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_2.A 0.12214f
C453 a_44403_15797# EN 0.045f
C454 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout CLK 0.20785f
C455 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout VDD 2.73822f
C456 a_29289_15797# VDD 0.01186f
C457 Nand_Gate_6.A a_78881_15797# 0.04443f
C458 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C VDD 3.61242f
C459 D_FlipFlop_6.3-input-nand_2.Vout a_132925_23350# 0.01335f
C460 D_FlipFlop_4.3-input-nand_2.C VDD 2.74431f
C461 a_109285_49858# CLK 0.03129f
C462 And_Gate_2.Nand_Gate_0.Vout a_92725_16975# 0.05964f
C463 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C EN 0.07601f
C464 a_46505_52572# a_47119_52572# 0.05935f
C465 a_108671_49858# VDD 0.06071f
C466 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout VDD 2.01342f
C467 RingCounter_0.D_FlipFlop_10.Qbar RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.11654f
C468 FFCLR D_FlipFlop_5.3-input-nand_1.Vout 0.95879f
C469 D_FlipFlop_1.3-input-nand_0.Vout VDD 1.77126f
C470 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK 0.29644f
C471 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout CLK 0.71245f
C472 D_FlipFlop_4.Nand_Gate_0.Vout Q3 0.11443f
C473 CDAC8_0.switch_8.Z a_75898_42964# 0.01003f
C474 a_107313_52572# VDD 0.02521f
C475 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B a_107313_49858# 0.04443f
C476 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_1.Vout 0.07411f
C477 EN Q2 0.2481f
C478 D_FlipFlop_5.3-input-nand_2.Vout a_132925_26914# 0.01335f
C479 a_134283_19786# a_134897_19786# 0.05935f
C480 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_98245_49858# 0.05964f
C481 FFCLR a_128851_20636# 0.04443f
C482 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B CLK 0.16166f
C483 a_75898_35820# CDAC8_0.switch_7.Z 0.27082f
C484 Nand_Gate_0.B Comparator_0.Vinm 0.03263f
C485 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_33363_13083# 0.01335f
C486 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout a_122427_49858# 0.04995f
C487 a_90535_13083# EN 0.0452f
C488 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout a_45147_52572# 0.04443f
C489 a_32749_13083# CLK 0.02953f
C490 Nand_Gate_6.A Nand_Gate_6.Vout 0.0689f
C491 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout a_109285_49858# 0.04443f
C492 a_30647_13083# VDD 0.02578f
C493 a_128237_39721# a_128851_39721# 0.05935f
C494 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.09975f
C495 D_FlipFlop_2.Qbar D_FlipFlop_2.Nand_Gate_0.Vout 0.07122f
C496 Nand_Gate_2.B VDD 4.34021f
C497 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B EN 0.497f
C498 a_103765_47663# CLK 0.07396f
C499 D_FlipFlop_4.3-input-nand_2.Vout a_132925_30478# 0.01335f
C500 FFCLR a_128851_27764# 0.04443f
C501 a_89307_52572# RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.05964f
C502 a_93097_47663# VDD 0.02521f
C503 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0846f
C504 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout CLK 0.03574f
C505 Nand_Gate_5.A a_128851_46849# 0.04628f
C506 RingCounter_0.D_FlipFlop_6.Qbar a_123785_49858# 0.01335f
C507 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_91279_49858# 0.04444f
C508 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C EN 0.09031f
C509 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout EN 0.08852f
C510 a_48565_16975# VDD 0.02521f
C511 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout EN 0.6138f
C512 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B a_89921_13083# 0.04443f
C513 Nand_Gate_6.Vout And_Gate_2.Nand_Gate_0.Vout 0.24808f
C514 a_65125_49858# CLK 0.03129f
C515 Nand_Gate_5.B Q2 0.06203f
C516 Nand_Gate_7.B EN 1.37686f
C517 D_FlipFlop_7.Nand_Gate_1.Vout Q0 0.06993f
C518 Nand_Gate_1.A EN 0.42008f
C519 D_FlipFlop_5.3-input-nand_0.Vout VDD 1.77946f
C520 a_64511_49858# VDD 0.06071f
C521 a_112745_52572# a_113359_52572# 0.05935f
C522 D_FlipFlop_1.3-input-nand_0.Vout a_132311_36157# 0.04444f
C523 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.08377f
C524 a_99603_13083# CLK 0.03129f
C525 a_84489_15797# EN 0.04443f
C526 a_98989_13083# VDD 0.02578f
C527 a_132925_23350# VDD 0.01186f
C528 a_65125_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.05964f
C529 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_2.Vout 0.88855f
C530 Nand_Gate_7.A a_61795_13083# 0.04443f
C531 a_89921_15797# CLK 0.04619f
C532 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout EN 0.09127f
C533 a_96273_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.05964f
C534 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout a_43045_52572# 0.04444f
C535 a_46375_13083# EN 0.0452f
C536 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout CLK 0.03479f
C537 a_88563_15797# VDD 0.03339f
C538 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout CLK 0.03479f
C539 D_FlipFlop_6.3-input-nand_1.B a_134283_20636# 0.04443f
C540 D_FlipFlop_2.Nand_Gate_1.Vout VDD 1.46545f
C541 a_100347_52572# VDD 0.02521f
C542 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout EN 0.62384f
C543 Nand_Gate_0.A CDAC8_0.switch_8.Z 2.01979f
C544 FFCLR D_FlipFlop_0.CLK 0.60023f
C545 D_FlipFlop_3.3-input-nand_1.Vout a_132925_40571# 0.04543f
C546 FFCLR Nand_Gate_2.A 0.93855f
C547 Nand_Gate_5.B a_124399_49858# 0.04484f
C548 a_132925_30478# VDD 0.01186f
C549 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout VDD 2.31704f
C550 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.1182f
C551 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD 1.84669f
C552 Nand_Gate_5.B Nand_Gate_7.B 0.06463f
C553 a_123785_52572# VDD 0.01186f
C554 D_FlipFlop_0.Nand_Gate_0.Vout a_130209_46849# 0.05964f
C555 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout CLK 0.23566f
C556 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B VDD 1.73782f
C557 FFCLR D_FlipFlop_5.Nand_Gate_1.Vout 0.61318f
C558 a_76165_52572# VDD 0.02521f
C559 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD 2.04843f
C560 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_100961_15797# 0.05964f
C561 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout CLK 0.23566f
C562 D_FlipFlop_5.3-input-nand_1.B a_134283_24200# 0.04443f
C563 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_51369_15797# 0.04995f
C564 VDD Q6 3.79776f
C565 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_53471_52572# 0.04995f
C566 Nand_Gate_4.A RingCounter_0.D_FlipFlop_16.3-input-nand_1.B 0.2969f
C567 Nand_Gate_4.A RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.08377f
C568 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout EN 0.13192f
C569 D_FlipFlop_2.Nand_Gate_1.Vout a_128237_37007# 0.04444f
C570 a_55443_13083# CLK 0.03129f
C571 RingCounter_0.D_FlipFlop_11.Qbar a_95529_13083# 0.01335f
C572 D_FlipFlop_2.3-input-nand_2.C a_132311_37007# 0.05964f
C573 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_105955_13083# 0.04444f
C574 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_98989_13083# 0.04444f
C575 a_54829_13083# VDD 0.02578f
C576 D_FlipFlop_4.3-input-nand_1.B a_134283_27764# 0.04443f
C577 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121069_13083# 0.04443f
C578 Nand_Gate_3.B RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.08524f
C579 D_FlipFlop_2.Nand_Gate_0.Vout a_128851_39721# 0.04995f
C580 D_FlipFlop_6.3-input-nand_1.Vout a_134283_20636# 0.05964f
C581 FFCLR D_FlipFlop_0.Inverter_1.Vout 0.56808f
C582 a_130209_37007# VDD 0.02521f
C583 And_Gate_5.Nand_Gate_0.Vout Comparator_0.Vinm 0.02725f
C584 D_FlipFlop_4.Qbar a_128237_27764# 0.06113f
C585 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_1.3-input-nand_0.Vout 0.01418f
C586 D_FlipFlop_6.3-input-nand_0.Vout a_132311_23350# 0.04444f
C587 Comparator_0.Vinm VDD 17.402f
C588 D_FlipFlop_0.Qbar a_128237_44135# 0.06113f
C589 CDAC8_0.switch_7.Z Q5 1.11487f
C590 a_128237_37007# Q6 0.04443f
C591 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C CLK 0.30966f
C592 RingCounter_0.D_FlipFlop_12.Qbar a_83875_15797# 0.04443f
C593 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 1.09975f
C594 a_134283_36157# VDD 0.02521f
C595 a_52727_15797# VDD 0.02906f
C596 a_87205_49858# VDD 0.0301f
C597 D_FlipFlop_5.3-input-nand_1.Vout a_134283_24200# 0.05964f
C598 RingCounter_0.D_FlipFlop_11.Qbar VDD 1.95446f
C599 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.26069f
C600 a_123041_13083# CLK 0.04443f
C601 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.08641f
C602 CDAC8_0.switch_9.Z Q2 0.38677f
C603 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.04107f
C604 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.06935f
C605 a_121683_13083# VDD 0.05686f
C606 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout EN 0.97979f
C607 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.25963f
C608 D_FlipFlop_5.3-input-nand_0.Vout a_132311_26914# 0.04444f
C609 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK 0.29644f
C610 FFCLR D_FlipFlop_2.Qbar 0.03748f
C611 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_2.Vout 0.8898f
C612 a_106699_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.01335f
C613 a_52113_52572# VDD 0.02521f
C614 a_132925_40571# VDD 0.01186f
C615 RingCounter_0.D_FlipFlop_5.Qbar a_102319_52572# 0.04443f
C616 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_119711_49858# 0.01335f
C617 RingCounter_0.D_FlipFlop_8.Qbar RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.11654f
C618 D_FlipFlop_3.Nand_Gate_0.Vout a_130209_43285# 0.05964f
C619 D_FlipFlop_4.3-input-nand_1.Vout a_134283_27764# 0.05964f
C620 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.07084f
C621 Nand_Gate_0.B EN 0.99738f
C622 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.08641f
C623 Nand_Gate_6.B a_82057_16975# 0.04443f
C624 D_FlipFlop_2.3-input-nand_1.B VDD 1.32602f
C625 D_FlipFlop_4.3-input-nand_0.Vout a_132311_30478# 0.04444f
C626 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.04109f
C627 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout CLK 0.03479f
C628 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_96273_49858# 0.05964f
C629 Nand_Gate_2.B a_107313_52572# 0.04443f
C630 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout CLK 0.23566f
C631 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.07084f
C632 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B a_118353_49858# 0.04443f
C633 CDAC8_0.switch_9.Z Nand_Gate_7.B 1.10291f
C634 a_134897_44135# VDD 0.01186f
C635 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_55443_15797# 0.01335f
C636 D_FlipFlop_7.3-input-nand_2.C a_132925_17072# 0.01335f
C637 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_53471_49858# 0.04543f
C638 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.04107f
C639 a_106699_49858# EN 0.07058f
C640 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_46505_49858# 0.04995f
C641 CLK Q3 0.1175f
C642 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_41073_49858# 0.05964f
C643 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.06935f
C644 D_FlipFlop_7.3-input-nand_2.Vout VDD 2.77266f
C645 a_43045_49858# VDD 0.02568f
C646 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Nand_Gate_1.Vout 0.04109f
C647 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout VDD 2.46653f
C648 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout a_74807_13083# 0.04995f
C649 a_78881_13083# CLK 0.04619f
C650 Nand_Gate_6.B RingCounter_0.D_FlipFlop_12.3-input-nand_1.B 0.2969f
C651 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0846f
C652 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout a_120325_49858# 0.04443f
C653 Nand_Gate_6.B RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0839f
C654 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110643_15797# 0.01335f
C655 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1541f
C656 a_77523_13083# VDD 0.05686f
C657 Nand_Gate_2.B a_93097_47663# 0.04443f
C658 RingCounter_0.D_FlipFlop_14.Qbar a_61795_13083# 0.06113f
C659 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1541f
C660 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_111387_49858# 0.04443f
C661 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout CLK 0.30735f
C662 Nand_Gate_2.A RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.08514f
C663 a_40329_15797# VDD 0.01571f
C664 Nand_Gate_5.Vout Comparator_0.Vinm 0.02011f
C665 RingCounter_0.D_FlipFlop_17.Qbar a_47119_49858# 0.06113f
C666 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout VDD 2.74107f
C667 Nand_Gate_6.A RingCounter_0.D_FlipFlop_13.3-input-nand_1.B 0.2969f
C668 a_101705_52572# EN 0.04443f
C669 a_119711_49858# a_120325_49858# 0.05935f
C670 a_75898_35820# Q7 0.5017f
C671 Nand_Gate_6.A RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.08377f
C672 Nand_Gate_1.B a_104137_16975# 0.04443f
C673 D_FlipFlop_0.Inverter_1.Vout a_130209_46849# 0.04443f
C674 a_47119_52572# FFCLR 0.06113f
C675 a_111387_49858# VDD 0.04111f
C676 RingCounter_0.D_FlipFlop_16.Q CLK 0.06841f
C677 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.06935f
C678 FFCLR a_134897_19786# 0.08436f
C679 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_107927_13083# 0.04443f
C680 a_62539_49858# EN 0.07058f
C681 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_100347_49858# 0.05964f
C682 Nand_Gate_0.B And_Gate_4.Nand_Gate_0.Vout 0.02391f
C683 Nand_Gate_1.B a_112001_15797# 0.04443f
C684 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.08671f
C685 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_63767_15797# 0.04443f
C686 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_2.C 0.14842f
C687 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 1.09975f
C688 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_102319_52572# 0.04444f
C689 a_34721_13083# CLK 0.04619f
C690 a_42431_52572# VDD 0.05686f
C691 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_57545_49858# 0.04995f
C692 Nand_Gate_0.A CLK 0.70685f
C693 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.16429f
C694 a_33363_13083# VDD 0.05686f
C695 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout VDD 2.73822f
C696 a_69199_52572# VDD 0.02521f
C697 a_132311_20636# a_132925_20636# 0.05935f
C698 a_125845_47663# CLK 0.07396f
C699 Nand_Gate_5.A CDAC8_0.switch_7.Z 3.15716f
C700 a_115177_47663# VDD 0.03918f
C701 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C EN 0.07732f
C702 And_Gate_7.Nand_Gate_0.Vout CLK 0.32457f
C703 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_116995_15797# 0.04444f
C704 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_32749_13083# 0.04443f
C705 Nand_Gate_1.Vout a_114805_16975# 0.04995f
C706 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.3-input-nand_2.Vout 0.06935f
C707 CDAC8_0.switch_8.Z CDAC8_0.switch_5.Z 0.09134f
C708 a_70645_16975# VDD 0.02521f
C709 RingCounter_0.D_FlipFlop_12.Qbar RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.11654f
C710 And_Gate_5.Nand_Gate_0.Vout EN 0.0623f
C711 a_97631_49858# a_98245_49858# 0.05935f
C712 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C VDD 3.61242f
C713 a_132311_24200# a_132925_24200# 0.05935f
C714 VDD EN 0.14517p
C715 a_113359_52572# Nand_Gate_5.A 0.06113f
C716 Nand_Gate_7.B Q1 0.35004f
C717 a_67227_49858# VDD 0.04111f
C718 D_FlipFlop_1.3-input-nand_0.Vout a_134283_36157# 0.05964f
C719 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.30154f
C720 a_94915_15797# a_95529_15797# 0.05935f
C721 CDAC8_0.switch_0.Z Q2 0.50733f
C722 a_76909_15797# VDD 0.03178f
C723 Nand_Gate_1.A a_105955_13083# 0.04443f
C724 a_100961_13083# VDD 0.02865f
C725 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_1.B 0.27887f
C726 a_134283_23350# VDD 0.02521f
C727 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout CLK 0.30735f
C728 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1541f
C729 D_FlipFlop_2.3-input-nand_1.B D_FlipFlop_2.3-input-nand_1.Vout 0.08641f
C730 a_62409_15797# VDD 0.01571f
C731 D_FlipFlop_3.Inverter_1.Vout a_130209_43285# 0.04443f
C732 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_120325_52572# 0.04444f
C733 a_132311_27764# a_132925_27764# 0.05935f
C734 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B CLK 0.16166f
C735 Nand_Gate_2.B Comparator_0.Vinm 0.03245f
C736 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_87949_13083# 0.05964f
C737 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B CLK 0.16274f
C738 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.04107f
C739 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout CLK 0.29759f
C740 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.C 0.01194f
C741 a_90535_15797# VDD 0.06072f
C742 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.Vout 0.01194f
C743 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_72835_15797# 0.04444f
C744 D_FlipFlop_3.3-input-nand_1.Vout a_134897_40571# 0.01335f
C745 D_FlipFlop_4.Qbar D_FlipFlop_4.Nand_Gate_1.Vout 0.11654f
C746 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout VDD 2.16852f
C747 a_67841_15797# a_68455_15797# 0.05935f
C748 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_66483_15797# 0.04995f
C749 a_128237_17072# a_128851_17072# 0.05935f
C750 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_1.B 0.27878f
C751 a_134283_30478# VDD 0.02521f
C752 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD 1.56255f
C753 D_FlipFlop_0.Qbar D_FlipFlop_0.Nand_Gate_1.Vout 0.11654f
C754 Nand_Gate_5.B VDD 4.31948f
C755 D_FlipFlop_2.Nand_Gate_1.Vout Q6 0.06993f
C756 FFCLR a_134283_33443# 0.01803f
C757 a_128237_33443# VDD 0.02521f
C758 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1541f
C759 CDAC8_0.switch_0.Z Nand_Gate_7.B 3.36457f
C760 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.26069f
C761 a_75551_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.01335f
C762 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout EN 0.08852f
C763 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_112745_52572# 0.04995f
C764 a_85233_49858# EN 0.01149f
C765 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0846f
C766 a_75551_49858# a_76165_49858# 0.05935f
C767 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout VDD 2.73822f
C768 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout EN 0.06649f
C769 D_FlipFlop_1.Qbar a_128237_36157# 0.04443f
C770 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout a_89307_52572# 0.04443f
C771 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_2.C 0.1486f
C772 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout 0.30154f
C773 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_1.Vout 0.07303f
C774 Nand_Gate_0.A a_132925_39721# 0.04682f
C775 D_FlipFlop_2.Nand_Gate_1.Vout a_130209_37007# 0.05964f
C776 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_107927_13083# 0.05964f
C777 D_FlipFlop_7.Nand_Gate_0.Vout a_130209_19786# 0.05964f
C778 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_100961_13083# 0.05964f
C779 a_56801_13083# VDD 0.02865f
C780 CDAC8_0.switch_6.Z Q2 0.74768f
C781 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_95529_13083# 0.04995f
C782 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C EN 0.07664f
C783 a_57545_52572# a_58159_52572# 0.05935f
C784 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_88563_13083# 0.04543f
C785 a_110029_13083# a_110643_13083# 0.05935f
C786 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_83875_13083# 0.04444f
C787 Nand_Gate_5.Vout a_115177_47663# 0.05964f
C788 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_98989_15797# 0.04443f
C789 FFCLR D_FlipFlop_1.Qbar 0.0683f
C790 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_76909_13083# 0.04444f
C791 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_28675_15797# 0.04444f
C792 RingCounter_0.D_FlipFlop_12.Qbar CLK 0.09276f
C793 a_132925_37007# VDD 0.01186f
C794 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121069_15797# 0.05964f
C795 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout 0.30154f
C796 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_1.Vout 0.07299f
C797 And_Gate_4.Nand_Gate_0.Vout VDD 1.43186f
C798 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout a_63767_15797# 0.04443f
C799 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0846f
C800 RingCounter_0.D_FlipFlop_16.Q a_28675_15797# 0.07417f
C801 Nand_Gate_5.Vout EN 0.10962f
C802 a_122427_52572# VDD 0.02521f
C803 a_117609_15797# EN 0.04443f
C804 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_0.Vout 0.25997f
C805 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B a_57415_13083# 0.04995f
C806 FFCLR a_132925_24200# 0.045f
C807 a_90665_49858# VDD 0.06015f
C808 D_FlipFlop_1.3-input-nand_1.B VDD 1.32602f
C809 FFCLR Nand_Gate_5.A 0.61687f
C810 Comparator_0.Vinm Q6 0.56023f
C811 D_FlipFlop_6.Nand_Gate_0.Vout Q1 0.11443f
C812 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout VDD 2.07863f
C813 D_FlipFlop_7.3-input-nand_2.C VDD 2.74431f
C814 FFCLR D_FlipFlop_0.3-input-nand_2.Vout 0.06105f
C815 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout CLK 0.23566f
C816 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout 0.30154f
C817 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.30154f
C818 a_123655_13083# VDD 0.01327f
C819 a_123041_15797# CLK 0.04443f
C820 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.16429f
C821 a_98245_52572# VDD 0.02521f
C822 D_FlipFlop_6.Inverter_1.Vout a_130209_20636# 0.04995f
C823 a_121683_15797# VDD 0.03339f
C824 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.09975f
C825 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_40329_13083# 0.04995f
C826 CDAC8_0.switch_6.Z Nand_Gate_7.B 3.32256f
C827 a_134897_40571# VDD 0.01186f
C828 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Qbar 1.05791f
C829 D_FlipFlop_6.Qbar a_128851_20636# 0.01335f
C830 a_41073_49858# EN 0.01767f
C831 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_33363_13083# 0.04543f
C832 a_53471_49858# a_54085_49858# 0.05935f
C833 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_28675_13083# 0.04444f
C834 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_122427_49858# 0.04443f
C835 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout EN 0.78734f
C836 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_62539_49858# 0.01335f
C837 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_52727_13083# 0.04443f
C838 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_76909_15797# 0.05964f
C839 D_FlipFlop_5.Inverter_1.Vout a_130209_24200# 0.04995f
C840 Nand_Gate_5.B Nand_Gate_5.Vout 2.12832f
C841 a_87949_13083# a_88563_13083# 0.05935f
C842 D_FlipFlop_5.Qbar a_128851_24200# 0.01335f
C843 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_98245_49858# 0.04444f
C844 a_86591_52572# a_87205_52572# 0.05935f
C845 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout EN 0.06649f
C846 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.06955f
C847 a_29289_15797# EN 0.04443f
C848 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_65125_52572# 0.04444f
C849 a_134283_33443# a_134897_33443# 0.05935f
C850 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C EN 0.07732f
C851 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout a_100347_52572# 0.04443f
C852 D_FlipFlop_1.3-input-nand_1.Vout VDD 1.7803f
C853 CDAC8_0.switch_9.Z VDD 12.5516f
C854 a_117739_52572# a_118353_52572# 0.05935f
C855 a_134897_26914# VDD 0.01186f
C856 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout CLK 0.30716f
C857 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout 0.01681f
C858 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_43045_49858# 0.04444f
C859 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout EN 0.58846f
C860 D_FlipFlop_4.Inverter_1.Vout a_130209_27764# 0.04995f
C861 a_34721_15797# CLK 0.04619f
C862 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.16429f
C863 D_FlipFlop_1.3-input-nand_0.Vout EN 0.08617f
C864 a_46505_49858# VDD 0.01571f
C865 a_33363_15797# VDD 0.02954f
C866 a_128237_36157# a_128851_36157# 0.05935f
C867 CDAC8_0.switch_2.Z CLK 0.08199f
C868 D_FlipFlop_1.Qbar D_FlipFlop_1.Nand_Gate_0.Vout 0.07122f
C869 Nand_Gate_2.A a_132925_43285# 0.04684f
C870 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout VDD 2.74107f
C871 a_75898_21528# VDD 1.33597f
C872 a_79495_13083# VDD 0.01327f
C873 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_39715_15797# 0.04444f
C874 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_0.Vout 1.02519f
C875 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Qbar 0.07122f
C876 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1541f
C877 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK 0.29644f
C878 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_32749_15797# 0.05964f
C879 a_74193_52572# VDD 0.02521f
C880 FFCLR a_128851_36157# 0.04623f
C881 RingCounter_0.D_FlipFlop_2.Qbar VDD 1.96503f
C882 CDAC8_0.switch_2.Z CDAC8_0.switch_1.Z 0.06088f
C883 Nand_Gate_2.Vout And_Gate_6.Nand_Gate_0.Vout 0.10129f
C884 CDAC8_0.switch_5.Z CLK 0.21166f
C885 a_51499_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.01335f
C886 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout VDD 2.07863f
C887 a_75898_28676# VDD 1.30969f
C888 Nand_Gate_2.B EN 0.99738f
C889 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.06935f
C890 D_FlipFlop_1.Qbar Q7 1.06172f
C891 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.3-input-nand_2.C 0.26069f
C892 a_65869_13083# a_66483_13083# 0.05935f
C893 a_113359_49858# VDD 0.02906f
C894 Nand_Gate_5.A a_118353_52572# 0.04443f
C895 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.16429f
C896 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout CLK 0.03574f
C897 RingCounter_0.D_FlipFlop_7.Qbar Nand_Gate_5.A 1.10693f
C898 a_132925_19786# VDD 0.01186f
C899 RingCounter_0.D_FlipFlop_6.Qbar RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.11654f
C900 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout CLK 0.71127f
C901 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110643_13083# 0.01335f
C902 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_102319_49858# 0.04444f
C903 a_128237_20636# VDD 0.02521f
C904 Nand_Gate_1.B RingCounter_0.D_FlipFlop_9.3-input-nand_1.B 0.2969f
C905 D_FlipFlop_0.3-input-nand_2.Vout a_130209_46849# 0.04443f
C906 D_FlipFlop_2.3-input-nand_1.Vout a_132925_37007# 0.04543f
C907 D_FlipFlop_3.Qbar a_128851_40571# 0.01335f
C908 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_110643_13083# 0.04543f
C909 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout VDD 2.41001f
C910 RingCounter_0.D_FlipFlop_17.Qbar a_47119_52572# 0.04443f
C911 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.07084f
C912 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout VDD 3.68398f
C913 a_35335_13083# VDD 0.01327f
C914 RingCounter_0.D_FlipFlop_8.Qbar VDD 1.95446f
C915 D_FlipFlop_0.Qbar VDD 1.89794f
C916 a_88563_15797# EN 0.045f
C917 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.25963f
C918 D_FlipFlop_3.3-input-nand_1.B a_134897_40571# 0.04995f
C919 a_128237_27764# VDD 0.02521f
C920 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.06955f
C921 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.26069f
C922 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.06993f
C923 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.06955f
C924 a_128237_23350# a_128851_23350# 0.05935f
C925 a_92725_16975# VDD 0.02521f
C926 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout EN 0.09127f
C927 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.15399f
C928 a_128237_46849# Q4 0.06113f
C929 a_128237_43285# VDD 0.02521f
C930 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout EN 0.97839f
C931 D_FlipFlop_1.Nand_Gate_1.Vout VDD 1.46545f
C932 a_123785_52572# EN 0.04443f
C933 a_54829_15797# a_55443_15797# 0.05935f
C934 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout a_45147_52572# 0.04443f
C935 a_50755_15797# VDD 0.02906f
C936 a_43789_13083# a_44403_13083# 0.05935f
C937 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_76165_52572# 0.04443f
C938 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B EN 0.26843f
C939 a_69199_49858# VDD 0.02906f
C940 VDD Q1 3.61075f
C941 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout EN 0.97979f
C942 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.06955f
C943 FFCLR Nand_Gate_3.B 0.0826f
C944 a_78881_15797# VDD 0.03119f
C945 D_FlipFlop_1.Nand_Gate_0.Vout a_128851_36157# 0.04995f
C946 a_134283_46849# a_134897_46849# 0.05935f
C947 a_105955_13083# VDD 0.02521f
C948 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_43789_13083# 0.04444f
C949 EN Q6 0.2481f
C950 CDAC8_0.switch_8.Z Q5 0.32925f
C951 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Nand_Gate_1.Vout 0.04109f
C952 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B a_100961_13083# 0.04443f
C953 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_87949_15797# 0.04444f
C954 a_112001_15797# CLK 0.04619f
C955 a_128237_26914# a_128851_26914# 0.05935f
C956 D_FlipFlop_6.3-input-nand_1.B VDD 1.32726f
C957 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout VDD 2.16852f
C958 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout CLK 0.03479f
C959 D_FlipFlop_7.Qbar Q1 0.01194f
C960 a_110643_15797# VDD 0.03339f
C961 a_62539_52572# a_63153_52572# 0.05935f
C962 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_107927_15797# 0.05964f
C963 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.48392f
C964 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.06955f
C965 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.25963f
C966 D_FlipFlop_0.CLK CLK 0.01464f
C967 Nand_Gate_2.A CLK 0.64539f
C968 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout a_107927_13083# 0.04995f
C969 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_68455_15797# 0.01335f
C970 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Nand_Gate_1.Vout 0.04109f
C971 a_128237_30478# a_128851_30478# 0.05935f
C972 a_128851_36157# Q7 0.01335f
C973 CDAC8_0.switch_7.Z Q2 1.5084f
C974 D_FlipFlop_4.3-input-nand_1.B VDD 1.32727f
C975 a_91279_52572# VDD 0.02521f
C976 a_123785_52572# Nand_Gate_5.B 0.01335f
C977 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_121683_13083# 0.04543f
C978 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.16429f
C979 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_116995_13083# 0.04444f
C980 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_107927_15797# 0.04443f
C981 FFCLR D_FlipFlop_4.Qbar 0.03748f
C982 Comparator_0.Vinm EN 15.5364f
C983 D_FlipFlop_3.3-input-nand_2.Vout a_130209_43285# 0.04443f
C984 a_130209_33443# VDD 0.02521f
C985 Nand_Gate_3.B a_62539_52572# 0.04995f
C986 Nand_Gate_6.Vout VDD 1.36733f
C987 CDAC8_0.switch_0.Z VDD 1.38999f
C988 D_FlipFlop_1.3-input-nand_2.Vout a_132311_33443# 0.04443f
C989 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.03449f
C990 D_FlipFlop_2.Nand_Gate_0.Vout a_130209_39721# 0.05964f
C991 Nand_Gate_5.B Q6 0.06203f
C992 a_40459_52572# a_41073_52572# 0.05935f
C993 FFCLR D_FlipFlop_0.3-input-nand_2.C 0.76213f
C994 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_5.A 0.12214f
C995 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.04109f
C996 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout CLK 0.03574f
C997 D_FlipFlop_3.Qbar Q4 0.01194f
C998 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C VDD 3.61242f
C999 D_FlipFlop_6.3-input-nand_1.Vout VDD 1.78032f
C1000 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Qbar 1.05791f
C1001 D_FlipFlop_0.3-input-nand_2.Vout a_132311_46849# 0.05964f
C1002 a_61795_13083# VDD 0.02521f
C1003 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout m3_125329_49141# 0.01611f
C1004 And_Gate_0.Nand_Gate_0.Vout CLK 0.63116f
C1005 a_58159_52572# Nand_Gate_3.B 0.06113f
C1006 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_90535_13083# 0.01335f
C1007 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C VDD 3.56545f
C1008 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_85847_13083# 0.05964f
C1009 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_78881_13083# 0.05964f
C1010 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.25963f
C1011 CDAC8_0.switch_7.Z Nand_Gate_7.B 7.65138f
C1012 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_73449_13083# 0.04995f
C1013 a_134897_37007# VDD 0.01186f
C1014 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_66483_13083# 0.04543f
C1015 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B a_112615_13083# 0.04995f
C1016 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_61795_13083# 0.04444f
C1017 a_128851_46849# VDD 0.01186f
C1018 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B CLK 0.16166f
C1019 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_54829_13083# 0.04444f
C1020 Nand_Gate_5.B Comparator_0.Vinm 0.14544f
C1021 D_FlipFlop_6.3-input-nand_0.Vout a_134897_23350# 0.01335f
C1022 D_FlipFlop_4.3-input-nand_1.Vout VDD 1.78032f
C1023 RingCounter_0.D_FlipFlop_9.Qbar a_106569_13083# 0.01335f
C1024 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_63767_15797# 0.05964f
C1025 FFCLR D_FlipFlop_6.Inverter_1.Vout 0.56927f
C1026 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.07084f
C1027 a_96273_49858# CLK 0.04619f
C1028 D_FlipFlop_0.Nand_Gate_0.Vout Q4 0.11443f
C1029 FFCLR a_134897_24200# 0.04023f
C1030 RingCounter_0.D_FlipFlop_12.Qbar RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.07122f
C1031 D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.48313f
C1032 And_Gate_1.Nand_Gate_0.Vout CLK 0.59514f
C1033 a_95659_49858# VDD 0.01712f
C1034 a_128851_24200# VDD 0.01186f
C1035 FFCLR D_FlipFlop_0.3-input-nand_1.B 0.44507f
C1036 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.04107f
C1037 a_64511_52572# VDD 0.01186f
C1038 a_111387_52572# RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.05964f
C1039 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B CLK 0.06986f
C1040 D_FlipFlop_5.3-input-nand_0.Vout a_134897_26914# 0.01335f
C1041 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout CLK 0.28375f
C1042 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_107313_49858# 0.05964f
C1043 a_123655_15797# VDD 0.05687f
C1044 CDAC8_0.switch_6.Z VDD 13.0122f
C1045 Nand_Gate_4.B a_51369_15797# 0.01335f
C1046 Nand_Gate_6.B a_94915_15797# 0.06113f
C1047 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_35335_13083# 0.01335f
C1048 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout EN 0.08852f
C1049 FFCLR D_FlipFlop_4.Inverter_1.Vout 0.56808f
C1050 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_30647_13083# 0.05964f
C1051 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Nand_Gate_1.Vout 0.04109f
C1052 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.08641f
C1053 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_64511_49858# 0.04543f
C1054 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.06935f
C1055 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_55443_13083# 0.01335f
C1056 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout VDD 2.88547f
C1057 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_57545_52572# 0.04995f
C1058 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.C 0.01194f
C1059 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.Vout 0.01194f
C1060 D_FlipFlop_4.3-input-nand_0.Vout a_134897_30478# 0.01335f
C1061 And_Gate_4.Nand_Gate_0.Vout Comparator_0.Vinm 0.02739f
C1062 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.08671f
C1063 FFCLR a_48937_47663# 0.04705f
C1064 Nand_Gate_6.A a_83875_15797# 0.06113f
C1065 Nand_Gate_2.Vout CLK 2.32679f
C1066 a_40329_15797# EN 0.04443f
C1067 a_87205_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.05964f
C1068 D_FlipFlop_0.CLK a_132311_44135# 0.0315f
C1069 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout EN 0.1313f
C1070 D_FlipFlop_1.3-input-nand_1.B Comparator_0.Vinm 0.03198f
C1071 Nand_Gate_1.B Nand_Gate_1.Vout 2.35665f
C1072 D_FlipFlop_3.3-input-nand_2.Vout a_132311_43285# 0.05964f
C1073 Nand_Gate_3.B RingCounter_0.D_FlipFlop_2.3-input-nand_1.B 0.29683f
C1074 a_118353_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.05964f
C1075 FFCLR D_FlipFlop_0.3-input-nand_1.Vout 0.95879f
C1076 a_52113_49858# CLK 0.04619f
C1077 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B CLK 0.16274f
C1078 a_51499_49858# VDD 0.01712f
C1079 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout CLK 0.27362f
C1080 a_35335_15797# VDD 0.06072f
C1081 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1541f
C1082 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_0.Vout 1.01929f
C1083 CDAC8_0.switch_9.Z Q6 0.24469f
C1084 a_68585_52572# Nand_Gate_0.A 0.01335f
C1085 D_FlipFlop_0.3-input-nand_0.Vout a_134283_46849# 0.05964f
C1086 RingCounter_0.D_FlipFlop_11.Qbar RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.11654f
C1087 RingCounter_0.D_FlipFlop_10.Qbar CLK 0.09298f
C1088 D_FlipFlop_6.Nand_Gate_1.Vout VDD 1.46545f
C1089 D_FlipFlop_4.Nand_Gate_0.Vout a_128237_30478# 0.04444f
C1090 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_0.Vout 0.0846f
C1091 a_84489_13083# VDD 0.0563f
C1092 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.25963f
C1093 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout CLK 0.1215f
C1094 FFCLR D_FlipFlop_3.3-input-nand_0.Vout 0.1263f
C1095 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout a_107927_15797# 0.04443f
C1096 a_120325_52572# VDD 0.02521f
C1097 Nand_Gate_0.A RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.08514f
C1098 Nand_Gate_7.A a_56801_15797# 0.04443f
C1099 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout a_85847_13083# 0.04995f
C1100 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_75551_52572# 0.04995f
C1101 Vbias Vin 0.78432f
C1102 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout EN 0.06649f
C1103 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_111387_49858# 0.05964f
C1104 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_1.Vout 0.08671f
C1105 D_FlipFlop_4.Nand_Gate_1.Vout VDD 1.46545f
C1106 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout CLK 0.71127f
C1107 RingCounter_0.D_FlipFlop_13.Qbar a_72835_13083# 0.06113f
C1108 FFCLR RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.08514f
C1109 a_128237_26914# Q2 0.06113f
C1110 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.06935f
C1111 a_119711_49858# CLK 0.02953f
C1112 D_FlipFlop_1.3-input-nand_1.Vout Comparator_0.Vinm 0.03205f
C1113 CDAC8_0.switch_9.Z Comparator_0.Vinm 0.22008p
C1114 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.09975f
C1115 a_118353_49858# VDD 0.0325f
C1116 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD 2.04843f
C1117 FFCLR Nand_Gate_7.B 0.93969f
C1118 a_46505_52572# VDD 0.0563f
C1119 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_68585_49858# 0.04995f
C1120 D_FlipFlop_0.CLK Q4 0.19645f
C1121 Nand_Gate_2.A Q4 0.06203f
C1122 D_FlipFlop_2.Inverter_1.Vout a_130209_39721# 0.04443f
C1123 a_134283_19786# VDD 0.02521f
C1124 CLK Q5 0.1175f
C1125 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C EN 0.07732f
C1126 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_1.Vout 0.08671f
C1127 a_75898_21528# Comparator_0.Vinm 0.04177f
C1128 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout CLK 0.30716f
C1129 a_128237_39721# VDD 0.02521f
C1130 a_130209_20636# VDD 0.02521f
C1131 Nand_Gate_4.B And_Gate_1.Nand_Gate_0.Vout 0.06473f
C1132 D_FlipFlop_2.3-input-nand_1.Vout a_134897_37007# 0.01335f
C1133 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1541f
C1134 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.C 1.09975f
C1135 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.06955f
C1136 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_112615_13083# 0.01335f
C1137 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.08641f
C1138 a_62409_15797# EN 0.04443f
C1139 a_40329_13083# VDD 0.0563f
C1140 a_134283_20636# a_134897_20636# 0.05935f
C1141 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout VDD 2.07863f
C1142 RingCounter_0.D_FlipFlop_10.Qbar a_117609_13083# 0.01335f
C1143 a_75898_28676# Comparator_0.Vinm 0.03583f
C1144 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_1.Vout 0.08671f
C1145 Nand_Gate_5.B a_115177_47663# 0.04443f
C1146 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK 0.29644f
C1147 FFCLR D_FlipFlop_5.Qbar 0.03748f
C1148 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.25963f
C1149 a_130209_27764# VDD 0.02521f
C1150 a_96273_52572# VDD 0.02521f
C1151 a_67841_15797# CLK 0.04619f
C1152 RingCounter_0.D_FlipFlop_4.Qbar VDD 1.96503f
C1153 FFCLR a_132925_17072# 0.045f
C1154 RingCounter_0.D_FlipFlop_6.Qbar a_124399_52572# 0.04443f
C1155 Nand_Gate_7.B a_68455_15797# 0.04995f
C1156 a_66483_15797# VDD 0.03339f
C1157 a_114805_16975# VDD 0.02521f
C1158 D_FlipFlop_4.Qbar Nand_Gate_1.B 0.03509f
C1159 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_0.Vout 0.0846f
C1160 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout EN 0.62384f
C1161 D_FlipFlop_6.Qbar a_128237_23350# 0.04443f
C1162 D_FlipFlop_3.Inverter_1.Vout VDD 1.73058f
C1163 a_105955_15797# a_106569_15797# 0.05935f
C1164 Nand_Gate_5.B EN 0.58357f
C1165 a_75551_49858# CLK 0.03129f
C1166 a_134283_24200# a_134897_24200# 0.05935f
C1167 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C VDD 2.99599f
C1168 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout VDD 2.31704f
C1169 D_FlipFlop_1.3-input-nand_2.C a_132311_33443# 0.05964f
C1170 FFCLR D_FlipFlop_0.Nand_Gate_1.Vout 0.61318f
C1171 a_74193_49858# VDD 0.0325f
C1172 a_110029_13083# CLK 0.03129f
C1173 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_95529_15797# 0.04995f
C1174 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1541f
C1175 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B VDD 1.73782f
C1176 Nand_Gate_6.B Nand_Gate_6.A 0.08001f
C1177 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD 2.04843f
C1178 RingCounter_0.D_FlipFlop_10.Qbar a_116995_15797# 0.04443f
C1179 a_107927_13083# VDD 0.02578f
C1180 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_45761_13083# 0.05964f
C1181 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B CLK 0.16279f
C1182 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout EN 0.06649f
C1183 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_89921_15797# 0.05964f
C1184 D_FlipFlop_0.3-input-nand_2.C a_132311_46849# 0.04443f
C1185 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout 0.30154f
C1186 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.04107f
C1187 a_112615_15797# VDD 0.06072f
C1188 D_FlipFlop_5.Qbar a_128237_26914# 0.04443f
C1189 a_63153_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.05964f
C1190 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_6.3-input-nand_0.Vout 0.01418f
C1191 a_134283_27764# a_134897_27764# 0.05935f
C1192 RingCounter_0.D_FlipFlop_1.Qbar Nand_Gate_3.B 1.10693f
C1193 Nand_Gate_6.B And_Gate_2.Nand_Gate_0.Vout 0.04751f
C1194 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.06993f
C1195 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.Nand_Gate_1.Vout 0.1541f
C1196 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_123655_13083# 0.01335f
C1197 D_FlipFlop_1.Nand_Gate_1.Vout Comparator_0.Vinm 0.0419f
C1198 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_118967_13083# 0.05964f
C1199 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_98989_13083# 0.05964f
C1200 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_5.3-input-nand_0.Vout 0.01418f
C1201 a_132925_33443# VDD 0.01186f
C1202 Nand_Gate_3.B RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.08377f
C1203 And_Gate_4.Nand_Gate_0.Vout EN 0.0623f
C1204 Comparator_0.Vinm Q1 1.64921f
C1205 a_128237_17072# Q0 0.04443f
C1206 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C CLK 0.30966f
C1207 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C CLK 0.30901f
C1208 a_41073_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.05964f
C1209 D_FlipFlop_1.3-input-nand_1.B EN 0.40481f
C1210 a_85847_15797# VDD 0.02906f
C1211 RingCounter_0.D_FlipFlop_13.Qbar a_72835_15797# 0.04443f
C1212 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.Nand_Gate_1.Vout 0.1541f
C1213 a_75898_46095# CDAC8_0.switch_8.Z 0.33809f
C1214 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout VDD 2.07863f
C1215 a_43789_15797# a_44403_15797# 0.05935f
C1216 D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.48313f
C1217 a_123655_13083# EN 0.0452f
C1218 Nand_Gate_1.B D_FlipFlop_4.Inverter_1.Vout 0.12092f
C1219 D_FlipFlop_7.3-input-nand_2.Vout a_132925_19786# 0.01335f
C1220 RingCounter_0.D_FlipFlop_13.Qbar VDD 1.95446f
C1221 D_FlipFlop_3.Inverter_1.Vout a_130209_40571# 0.04995f
C1222 a_65869_13083# CLK 0.03129f
C1223 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.26069f
C1224 a_121683_15797# EN 0.045f
C1225 a_63767_13083# VDD 0.02578f
C1226 a_112001_13083# a_112615_13083# 0.05935f
C1227 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.07084f
C1228 CDAC8_0.switch_7.Z VDD 26.5678f
C1229 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_68455_13083# 0.01335f
C1230 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.Nand_Gate_1.Vout 0.1541f
C1231 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.0846f
C1232 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_63767_13083# 0.05964f
C1233 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_56801_13083# 0.05964f
C1234 D_FlipFlop_6.3-input-nand_2.C a_130209_20636# 0.04443f
C1235 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout 0.01681f
C1236 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout a_43045_49858# 0.04443f
C1237 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_51369_13083# 0.04995f
C1238 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 1.09975f
C1239 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_124399_52572# 0.04444f
C1240 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.48392f
C1241 D_FlipFlop_3.3-input-nand_2.C a_132311_43285# 0.04443f
C1242 D_FlipFlop_4.Qbar D_FlipFlop_4.Nand_Gate_0.Vout 0.07122f
C1243 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.14519f
C1244 a_98245_49858# CLK 0.03129f
C1245 CDAC8_0.switch_0.Z Comparator_0.Vinm 25.94f
C1246 Nand_Gate_7.B a_128851_23350# 0.04723f
C1247 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_73579_49858# 0.01335f
C1248 Nand_Gate_5.A CLK 0.8887f
C1249 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.16429f
C1250 a_97631_49858# VDD 0.06071f
C1251 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_106569_15797# 0.04995f
C1252 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.30154f
C1253 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout CLK 0.23566f
C1254 a_132311_24200# VDD 0.02521f
C1255 a_113359_52572# VDD 0.02521f
C1256 Nand_Gate_1.B Q2 0.05915f
C1257 CDAC8_0.switch_9.Z EN 5.40382f
C1258 Nand_Gate_4.A VDD 4.19805f
C1259 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_99603_15797# 0.01335f
C1260 D_FlipFlop_1.3-input-nand_1.Vout EN 0.97934f
C1261 RingCounter_0.D_FlipFlop_16.Qbar a_28675_15797# 0.04443f
C1262 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout VDD 2.73822f
C1263 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout VDD 2.8604f
C1264 D_FlipFlop_5.3-input-nand_2.C a_130209_24200# 0.04443f
C1265 Nand_Gate_0.A a_73579_52572# 0.04995f
C1266 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_109285_49858# 0.04444f
C1267 RingCounter_0.D_FlipFlop_2.Qbar a_69199_52572# 0.04443f
C1268 a_46505_49858# EN 0.04443f
C1269 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B a_68455_13083# 0.04995f
C1270 a_132311_46849# a_132925_46849# 0.05935f
C1271 a_33363_15797# EN 0.04775f
C1272 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_0.Vout 0.07084f
C1273 FFCLR D_FlipFlop_3.3-input-nand_1.Vout 0.95879f
C1274 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.06935f
C1275 Nand_Gate_6.B a_128851_26914# 0.04727f
C1276 FFCLR D_FlipFlop_6.3-input-nand_2.Vout 0.06105f
C1277 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.04107f
C1278 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout EN 0.13192f
C1279 Nand_Gate_6.A CLK 0.39021f
C1280 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C VDD 3.59745f
C1281 a_79495_13083# EN 0.0452f
C1282 CDAC8_0.switch_6.Z Q6 0.84702f
C1283 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout Nand_Gate_3.B 0.12214f
C1284 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.0846f
C1285 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_6.Inverter_1.Vout 0.01422f
C1286 D_FlipFlop_4.3-input-nand_2.C a_130209_27764# 0.04443f
C1287 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.06955f
C1288 a_89921_13083# a_90535_13083# 0.05935f
C1289 FFCLR D_FlipFlop_2.3-input-nand_0.Vout 0.1263f
C1290 FFCLR D_FlipFlop_4.3-input-nand_2.Vout 0.06105f
C1291 D_FlipFlop_0.CLK a_134283_44135# 0.04443f
C1292 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_63767_13083# 0.04443f
C1293 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C CLK 0.30966f
C1294 RingCounter_0.D_FlipFlop_16.Qbar a_29289_13083# 0.01335f
C1295 Nand_Gate_1.B Nand_Gate_7.B 0.0543f
C1296 And_Gate_2.Nand_Gate_0.Vout CLK 0.63116f
C1297 a_107927_15797# VDD 0.02906f
C1298 Nand_Gate_1.B Nand_Gate_1.A 0.08001f
C1299 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B CLK 0.16166f
C1300 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout a_56187_49858# 0.04995f
C1301 Nand_Gate_7.A CLK 0.39021f
C1302 D_FlipFlop_2.Qbar a_128851_37007# 0.01335f
C1303 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_54829_13083# 0.04443f
C1304 a_42431_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.01335f
C1305 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.26069f
C1306 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_5.Inverter_1.Vout 0.01422f
C1307 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout CLK 0.71245f
C1308 a_54085_49858# CLK 0.03129f
C1309 a_128237_44135# a_128851_44135# 0.05935f
C1310 a_53471_49858# VDD 0.06071f
C1311 CDAC8_0.switch_6.Z Comparator_0.Vinm 0.45096p
C1312 a_88563_13083# CLK 0.03129f
C1313 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Inverter_1.Vout 0.25963f
C1314 a_87949_13083# VDD 0.02578f
C1315 D_FlipFlop_2.3-input-nand_1.B a_134897_37007# 0.04995f
C1316 a_86591_52572# VDD 0.01186f
C1317 RingCounter_0.D_FlipFlop_1.Qbar a_57545_49858# 0.01335f
C1318 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.26069f
C1319 a_97631_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.01335f
C1320 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.0846f
C1321 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout EN 0.0879f
C1322 And_Gate_7.Nand_Gate_0.Vout a_125845_47663# 0.05964f
C1323 Nand_Gate_7.A RingCounter_0.D_FlipFlop_15.3-input-nand_1.B 0.2969f
C1324 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_52727_15797# 0.04443f
C1325 a_56187_52572# RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.05964f
C1326 Nand_Gate_7.A RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.08377f
C1327 a_128237_36157# VDD 0.02521f
C1328 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0846f
C1329 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout EN 0.07459f
C1330 a_35335_13083# EN 0.0452f
C1331 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_113359_49858# 0.04444f
C1332 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout a_111387_52572# 0.04443f
C1333 a_123785_49858# a_124399_49858# 0.05935f
C1334 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.06955f
C1335 a_132311_43285# a_132925_43285# 0.05935f
C1336 a_120325_49858# VDD 0.0301f
C1337 a_67841_13083# a_68455_13083# 0.05935f
C1338 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_0.Vout 0.07084f
C1339 Nand_Gate_1.Vout CLK 2.75905f
C1340 D_FlipFlop_6.Nand_Gate_0.Vout a_128851_23350# 0.04995f
C1341 FFCLR VDD 28.0344f
C1342 a_79625_52572# a_80239_52572# 0.05935f
C1343 RingCounter_0.D_FlipFlop_5.Qbar RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.11654f
C1344 D_FlipFlop_1.3-input-nand_1.B D_FlipFlop_1.3-input-nand_1.Vout 0.08641f
C1345 D_FlipFlop_1.Nand_Gate_1.Vout EN 0.6447f
C1346 D_FlipFlop_7.3-input-nand_1.B VDD 1.40016f
C1347 And_Gate_2.Nand_Gate_0.Vout Q0 0.05118f
C1348 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout CLK 0.71245f
C1349 Nand_Gate_1.B a_116995_13083# 0.04443f
C1350 Nand_Gate_0.A RingCounter_0.D_FlipFlop_3.3-input-nand_1.B 0.29683f
C1351 EN Q1 0.2481f
C1352 FFCLR D_FlipFlop_7.Qbar 0.03748f
C1353 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.04107f
C1354 D_FlipFlop_0.3-input-nand_2.Vout a_132311_44135# 0.04443f
C1355 Nand_Gate_7.B a_134897_20636# 0.04548f
C1356 a_132925_20636# VDD 0.01186f
C1357 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_69199_52572# 0.04444f
C1358 D_FlipFlop_2.Inverter_1.Vout VDD 1.73058f
C1359 D_FlipFlop_7.3-input-nand_0.Vout a_132311_19786# 0.04444f
C1360 D_FlipFlop_0.3-input-nand_0.Vout a_132925_46849# 0.04995f
C1361 FFCLR D_FlipFlop_3.Nand_Gate_1.Vout 0.61318f
C1362 RingCounter_0.D_FlipFlop_17.Qbar RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.11654f
C1363 D_FlipFlop_5.Nand_Gate_0.Vout a_128851_26914# 0.04995f
C1364 Nand_Gate_3.B a_58159_49858# 0.04741f
C1365 a_83875_15797# a_84489_15797# 0.05935f
C1366 a_44403_13083# CLK 0.03129f
C1367 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout a_47119_52572# 0.04444f
C1368 Nand_Gate_1.A a_106569_15797# 0.01335f
C1369 a_54829_15797# VDD 0.03178f
C1370 a_128237_39721# Q6 0.06113f
C1371 a_110643_15797# EN 0.045f
C1372 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout CLK 0.30735f
C1373 a_43789_13083# VDD 0.02578f
C1374 D_FlipFlop_2.3-input-nand_2.Vout a_130209_39721# 0.04443f
C1375 a_95529_15797# VDD 0.01571f
C1376 a_63153_52572# CLK 0.04619f
C1377 a_128237_26914# VDD 0.02521f
C1378 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout CLK 0.71245f
C1379 a_62539_52572# VDD 0.0564f
C1380 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.06955f
C1381 Nand_Gate_6.B a_134897_24200# 0.04546f
C1382 D_FlipFlop_1.Nand_Gate_0.Vout a_130209_36157# 0.05964f
C1383 a_132925_27764# VDD 0.01186f
C1384 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout EN 0.61318f
C1385 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_43789_15797# 0.04444f
C1386 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout VDD 2.74107f
C1387 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B CLK 0.16274f
C1388 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout CLK 0.29759f
C1389 a_68455_15797# VDD 0.06072f
C1390 a_128851_17072# VDD 0.01186f
C1391 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_61795_15797# 0.04444f
C1392 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.08671f
C1393 a_101705_49858# a_102319_49858# 0.05935f
C1394 a_41073_52572# CLK 0.04443f
C1395 D_FlipFlop_7.3-input-nand_1.B a_134897_17072# 0.04995f
C1396 a_56801_15797# a_57415_15797# 0.05935f
C1397 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_55443_15797# 0.04995f
C1398 D_FlipFlop_1.Nand_Gate_1.Vout a_128237_33443# 0.04444f
C1399 Nand_Gate_5.B Q1 0.06203f
C1400 a_40459_52572# VDD 0.01606f
C1401 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD 1.56255f
C1402 a_45761_13083# a_46375_13083# 0.05935f
C1403 a_76165_49858# VDD 0.0301f
C1404 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout CLK 0.03574f
C1405 Nand_Gate_1.Vout Q0 0.05051f
C1406 Nand_Gate_6.Vout EN 0.10992f
C1407 CDAC8_0.switch_0.Z EN 0.56688f
C1408 D_FlipFlop_7.Qbar a_128851_17072# 0.01335f
C1409 Nand_Gate_3.B CLK 0.28415f
C1410 a_112001_13083# CLK 0.04619f
C1411 a_108671_52572# a_109285_52572# 0.05935f
C1412 a_58159_52572# VDD 0.02521f
C1413 a_110643_13083# VDD 0.05686f
C1414 Nand_Gate_5.A Q4 0.46277f
C1415 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_87205_52572# 0.04444f
C1416 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C EN 0.07732f
C1417 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout a_122427_52572# 0.04443f
C1418 D_FlipFlop_3.3-input-nand_2.Vout VDD 2.77266f
C1419 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout CLK 0.30716f
C1420 D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.48313f
C1421 FFCLR D_FlipFlop_7.Inverter_1.Vout 0.56927f
C1422 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C EN 0.07664f
C1423 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_41687_13083# 0.04443f
C1424 a_132311_17072# a_132925_17072# 0.05935f
C1425 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_87949_15797# 0.04443f
C1426 Nand_Gate_6.B Q2 0.34858f
C1427 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Qbar 0.07122f
C1428 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B a_62539_49858# 0.04995f
C1429 D_FlipFlop_3.3-input-nand_0.Vout a_132925_43285# 0.04995f
C1430 RingCounter_0.D_FlipFlop_14.Qbar CLK 0.09276f
C1431 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK 0.27229f
C1432 a_134897_33443# VDD 0.01186f
C1433 CDAC8_0.switch_5.Z Q3 0.59604f
C1434 Nand_Gate_0.A a_75898_39392# 0.01513f
C1435 Nand_Gate_1.Vout And_Gate_3.Nand_Gate_0.Vout 0.2638f
C1436 RingCounter_0.D_FlipFlop_9.Qbar a_105955_15797# 0.04443f
C1437 a_118353_52572# VDD 0.02521f
C1438 FFCLR a_132925_44135# 0.045f
C1439 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.04109f
C1440 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_53471_49858# 0.01335f
C1441 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Nand_Gate_1.Vout 0.04109f
C1442 RingCounter_0.D_FlipFlop_7.Qbar VDD 1.96539f
C1443 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.25963f
C1444 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout a_52727_15797# 0.04443f
C1445 a_95659_49858# EN 0.07058f
C1446 D_FlipFlop_6.Qbar Q2 0.01194f
C1447 RingCounter_0.D_FlipFlop_6.Qbar m3_125329_49141# 0.04886f
C1448 a_73579_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.01335f
C1449 a_79625_49858# a_80239_49858# 0.05935f
C1450 VDD Q7 3.79323f
C1451 a_130209_46849# VDD 0.02521f
C1452 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.06935f
C1453 a_64511_52572# EN 0.045f
C1454 a_67841_13083# CLK 0.04619f
C1455 FFCLR D_FlipFlop_6.3-input-nand_2.C 0.76213f
C1456 FFCLR D_FlipFlop_3.3-input-nand_1.B 0.44757f
C1457 CDAC8_0.switch_6.Z EN 11.3849f
C1458 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout CLK 0.03479f
C1459 a_66483_13083# VDD 0.05686f
C1460 D_FlipFlop_2.Nand_Gate_0.Vout Q6 0.11443f
C1461 D_FlipFlop_2.3-input-nand_2.Vout a_132311_39721# 0.05964f
C1462 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B a_52113_49858# 0.04443f
C1463 Nand_Gate_2.Vout a_103765_47663# 0.04443f
C1464 RingCounter_0.D_FlipFlop_9.Qbar RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.11654f
C1465 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout EN 0.78734f
C1466 FFCLR D_FlipFlop_2.3-input-nand_1.Vout 0.96009f
C1467 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_118353_49858# 0.05964f
C1468 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout CLK 0.03574f
C1469 Nand_Gate_6.B Nand_Gate_7.B 0.05683f
C1470 D_FlipFlop_6.3-input-nand_2.C a_132925_20636# 0.01335f
C1471 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B VDD 1.79521f
C1472 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout VDD 2.16852f
C1473 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_2.Vout 0.92808f
C1474 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_65869_15797# 0.05964f
C1475 FFCLR D_FlipFlop_4.3-input-nand_2.C 0.76213f
C1476 CDAC8_0.switch_7.Z Q6 1.11431f
C1477 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout CLK 0.23566f
C1478 a_128851_23350# VDD 0.01186f
C1479 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_75551_49858# 0.04543f
C1480 a_100347_49858# VDD 0.04111f
C1481 a_134283_24200# VDD 0.02521f
C1482 D_FlipFlop_6.Qbar Nand_Gate_7.B 0.03706f
C1483 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout a_54085_49858# 0.04443f
C1484 FFCLR D_FlipFlop_1.3-input-nand_0.Vout 1.1811f
C1485 a_134897_46849# VDD 0.01186f
C1486 D_FlipFlop_0.Nand_Gate_1.Vout a_128851_44135# 0.04995f
C1487 CDAC8_0.switch_9.Z Q1 0.36574f
C1488 D_FlipFlop_5.3-input-nand_2.C a_132925_24200# 0.01335f
C1489 Nand_Gate_0.A RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.08377f
C1490 Nand_Gate_5.B a_123655_15797# 0.04995f
C1491 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.08641f
C1492 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_43045_49858# 0.05964f
C1493 a_51499_49858# EN 0.07058f
C1494 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.1182f
C1495 a_57545_49858# a_58159_49858# 0.05935f
C1496 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C CLK 0.30901f
C1497 a_128851_30478# VDD 0.01186f
C1498 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.16429f
C1499 D_FlipFlop_5.Qbar Nand_Gate_6.B 0.03561f
C1500 a_75898_21528# Q1 0.50347f
C1501 CDAC8_0.switch_7.Z Comparator_0.Vinm 0.90922p
C1502 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_98245_52572# 0.04443f
C1503 a_43789_15797# VDD 0.03178f
C1504 D_FlipFlop_4.3-input-nand_2.C a_132925_27764# 0.01335f
C1505 D_FlipFlop_1.Inverter_1.Vout a_130209_36157# 0.04443f
C1506 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1541f
C1507 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C CLK 0.30966f
C1508 RingCounter_0.D_FlipFlop_2.Qbar a_69199_49858# 0.06113f
C1509 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.06955f
C1510 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.1182f
C1511 a_118967_15797# VDD 0.02906f
C1512 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout a_67227_52572# 0.04443f
C1513 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_1.Vout 0.08671f
C1514 D_FlipFlop_5.Nand_Gate_0.Vout Q2 0.11443f
C1515 D_FlipFlop_7.Nand_Gate_1.Vout a_128237_17072# 0.04444f
C1516 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_66483_13083# 0.01335f
C1517 a_84619_52572# a_85233_52572# 0.05935f
C1518 Nand_Gate_1.B VDD 7.72762f
C1519 RingCounter_0.D_FlipFlop_9.Qbar RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.07122f
C1520 a_118353_49858# EN 0.01149f
C1521 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout EN 0.97979f
C1522 CLK Q2 0.1175f
C1523 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.48392f
C1524 FFCLR D_FlipFlop_5.3-input-nand_0.Vout 0.1261f
C1525 CDAC8_0.switch_9.Z CDAC8_0.switch_0.Z 3.66237f
C1526 a_132311_46849# VDD 0.02521f
C1527 a_56187_49858# VDD 0.04111f
C1528 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_122427_49858# 0.05964f
C1529 D_FlipFlop_0.3-input-nand_2.C a_132311_44135# 0.05964f
C1530 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Qbar 0.07122f
C1531 a_75898_46095# Q4 0.57913f
C1532 a_89921_13083# VDD 0.02865f
C1533 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.08641f
C1534 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout VDD 2.8604f
C1535 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_79625_49858# 0.04995f
C1536 Nand_Gate_0.B a_84619_52572# 0.04995f
C1537 a_128237_20636# Q1 0.04443f
C1538 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B a_123041_13083# 0.04443f
C1539 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B CLK 0.06986f
C1540 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_0.Vout 0.0846f
C1541 D_FlipFlop_1.Inverter_1.Vout VDD 1.73058f
C1542 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_121069_15797# 0.04444f
C1543 FFCLR D_FlipFlop_2.Nand_Gate_1.Vout 0.61702f
C1544 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C CLK 0.19377f
C1545 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout CLK 0.30716f
C1546 a_30647_15797# VDD 0.02521f
C1547 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout CLK 0.03436f
C1548 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.3-input-nand_2.Vout 0.16429f
C1549 a_123785_49858# VDD 0.0563f
C1550 Nand_Gate_7.B CLK 0.58704f
C1551 Nand_Gate_1.A CLK 0.39021f
C1552 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout a_96887_13083# 0.04995f
C1553 a_80239_52572# Nand_Gate_0.B 0.06113f
C1554 a_66483_15797# EN 0.045f
C1555 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout 0.30154f
C1556 D_FlipFlop_6.Qbar D_FlipFlop_6.Nand_Gate_0.Vout 0.07122f
C1557 a_98989_15797# a_99603_15797# 0.05935f
C1558 RingCounter_0.D_FlipFlop_12.Qbar a_83875_13083# 0.06113f
C1559 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout EN 0.09127f
C1560 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C EN 0.76392f
C1561 a_74193_49858# EN 0.01149f
C1562 a_83875_15797# VDD 0.02906f
C1563 Nand_Gate_7.B CDAC8_0.switch_1.Z 0.33175f
C1564 a_134897_20636# VDD 0.01186f
C1565 RingCounter_0.D_FlipFlop_1.Qbar VDD 1.96503f
C1566 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.08641f
C1567 a_128237_44135# Q4 0.04443f
C1568 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B EN 0.26843f
C1569 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.07084f
C1570 CDAC8_0.switch_9.Z CDAC8_0.switch_6.Z 10.0827f
C1571 D_FlipFlop_6.Inverter_1.Vout a_130209_23350# 0.04443f
C1572 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout EN 0.97979f
C1573 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout CLK 0.30735f
C1574 D_FlipFlop_3.3-input-nand_2.C VDD 2.74431f
C1575 D_FlipFlop_0.Nand_Gate_0.Vout a_128237_46849# 0.04444f
C1576 a_106569_15797# VDD 0.01571f
C1577 D_FlipFlop_5.Qbar D_FlipFlop_5.Nand_Gate_0.Vout 0.07122f
C1578 RingCounter_0.D_FlipFlop_17.Qbar VDD 1.9286f
C1579 a_56801_15797# VDD 0.03119f
C1580 a_45761_13083# VDD 0.02865f
C1581 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout CLK 0.03479f
C1582 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_76909_15797# 0.04444f
C1583 a_75898_18814# CDAC8_0.switch_1.Z 0.28283f
C1584 a_108671_52572# VDD 0.01186f
C1585 And_Gate_7.Nand_Gate_0.Vout D_FlipFlop_0.CLK 0.25434f
C1586 D_FlipFlop_5.Inverter_1.Vout VDD 1.73058f
C1587 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD 1.86552f
C1588 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B a_73579_49858# 0.04995f
C1589 a_134897_27764# VDD 0.01186f
C1590 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_45761_15797# 0.05964f
C1591 D_FlipFlop_2.3-input-nand_2.Vout VDD 2.77266f
C1592 Nand_Gate_4.A a_40329_15797# 0.01335f
C1593 FFCLR Comparator_0.Vinm 7.22775f
C1594 Nand_Gate_1.B a_117609_15797# 0.01335f
C1595 And_Gate_6.Nand_Gate_0.Vout VDD 1.43186f
C1596 D_FlipFlop_5.Inverter_1.Vout a_130209_26914# 0.04443f
C1597 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.Nand_Gate_1.Vout 0.1541f
C1598 a_132311_17072# VDD 0.02521f
C1599 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.25963f
C1600 D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.48313f
C1601 Nand_Gate_6.Vout a_92725_16975# 0.04995f
C1602 D_FlipFlop_2.Inverter_1.Vout a_130209_37007# 0.04995f
C1603 D_FlipFlop_1.Nand_Gate_1.Vout a_130209_33443# 0.05964f
C1604 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_79625_52572# 0.04995f
C1605 FFCLR a_134283_36157# 0.01145f
C1606 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_57415_15797# 0.01335f
C1607 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout VDD 2.75863f
C1608 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1541f
C1609 a_79625_49858# VDD 0.06015f
C1610 a_132925_33443# EN 0.05084f
C1611 CDAC8_0.switch_8.Z VDD 1.45517f
C1612 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout a_56187_52572# 0.04443f
C1613 CDAC8_0.switch_6.Z a_75898_28676# 0.01232f
C1614 D_FlipFlop_0.3-input-nand_1.Vout a_132311_44135# 0.04444f
C1615 D_FlipFlop_0.3-input-nand_0.Vout VDD 1.77946f
C1616 CDAC8_0.switch_0.Z Q1 0.0732f
C1617 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.04107f
C1618 a_112615_13083# VDD 0.01327f
C1619 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout CLK 0.71127f
C1620 a_109285_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.05964f
C1621 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.08671f
C1622 D_FlipFlop_4.Inverter_1.Vout a_130209_30478# 0.04443f
C1623 RingCounter_0.D_FlipFlop_10.Qbar RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.07122f
C1624 FFCLR a_132925_40571# 0.045f
C1625 FFCLR a_52113_52572# 0.04443f
C1626 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout 0.01681f
C1627 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_65125_49858# 0.05964f
C1628 a_75898_18814# Q0 0.50347f
C1629 Nand_Gate_0.B RingCounter_0.D_FlipFlop_4.3-input-nand_1.B 0.29683f
C1630 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout a_89307_49858# 0.04995f
C1631 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_32749_15797# 0.04444f
C1632 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Qbar 1.05791f
C1633 D_FlipFlop_2.3-input-nand_2.C a_132311_39721# 0.04443f
C1634 a_90665_52572# Nand_Gate_2.A 0.01335f
C1635 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_44403_13083# 0.01335f
C1636 FFCLR D_FlipFlop_2.3-input-nand_1.B 0.44531f
C1637 D_FlipFlop_6.3-input-nand_1.B D_FlipFlop_6.3-input-nand_1.Vout 0.08641f
C1638 CDAC8_0.switch_7.Z EN 21.7044f
C1639 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C VDD 3.56545f
C1640 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_2.C 0.11237f
C1641 D_FlipFlop_3.3-input-nand_2.C a_130209_40571# 0.04443f
C1642 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B a_40459_49858# 0.04995f
C1643 D_FlipFlop_3.3-input-nand_0.Vout a_134897_43285# 0.01335f
C1644 a_85233_52572# CLK 0.04619f
C1645 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.08671f
C1646 RingCounter_0.D_FlipFlop_4.Qbar a_90665_49858# 0.01335f
C1647 a_84619_52572# VDD 0.0564f
C1648 Nand_Gate_0.A D_FlipFlop_2.Qbar 0.06938f
C1649 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout EN 0.61318f
C1650 FFCLR a_134897_44135# 0.04023f
C1651 D_FlipFlop_3.Nand_Gate_0.Vout a_128237_43285# 0.04444f
C1652 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_56187_49858# 0.04443f
C1653 a_128851_44135# VDD 0.01186f
C1654 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_97631_52572# 0.04995f
C1655 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout CLK 0.29759f
C1656 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_52727_15797# 0.05964f
C1657 FFCLR D_FlipFlop_7.3-input-nand_2.Vout 0.06105f
C1658 D_FlipFlop_5.3-input-nand_1.B D_FlipFlop_5.3-input-nand_1.Vout 0.08641f
C1659 RingCounter_0.D_FlipFlop_13.Qbar RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.07122f
C1660 Nand_Gate_4.A EN 0.42016f
C1661 a_45761_15797# a_46375_15797# 0.05935f
C1662 a_75898_42964# Q5 0.5017f
C1663 Nand_Gate_7.B Nand_Gate_4.B 0.0623f
C1664 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout EN 0.06649f
C1665 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout EN 0.78747f
C1666 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.48392f
C1667 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_84619_49858# 0.01335f
C1668 Nand_Gate_0.B CLK 0.41477f
C1669 a_132925_43285# VDD 0.01186f
C1670 a_68455_13083# VDD 0.01327f
C1671 a_80239_52572# VDD 0.02521f
C1672 CDAC8_0.switch_6.Z Q1 0.74949f
C1673 a_116995_13083# a_117609_13083# 0.05935f
C1674 a_75898_18814# Nand_Gate_4.B 0.0322f
C1675 Nand_Gate_5.B CDAC8_0.switch_7.Z 0.08438f
C1676 RingCounter_0.D_FlipFlop_3.Qbar a_80239_49858# 0.06113f
C1677 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C EN 0.07667f
C1678 D_FlipFlop_4.3-input-nand_1.B D_FlipFlop_4.3-input-nand_1.Vout 0.08641f
C1679 a_53471_52572# a_54085_52572# 0.05935f
C1680 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_120325_49858# 0.04444f
C1681 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout VDD 2.88547f
C1682 D_FlipFlop_6.Nand_Gate_1.Vout a_128237_20636# 0.04444f
C1683 Nand_Gate_6.B VDD 7.82571f
C1684 a_128237_40571# a_128851_40571# 0.05935f
C1685 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B a_34721_13083# 0.04443f
C1686 a_128237_19786# Q0 0.06113f
C1687 Nand_Gate_2.A a_91279_49858# 0.04741f
C1688 a_102319_49858# VDD 0.02906f
C1689 D_FlipFlop_6.Qbar VDD 1.89809f
C1690 Nand_Gate_7.A a_59977_16975# 0.0476f
C1691 Comparator_0.Vinm Q7 0.78864f
C1692 D_FlipFlop_5.Nand_Gate_1.Vout a_128237_24200# 0.04444f
C1693 RingCounter_0.D_FlipFlop_16.Qbar RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.07122f
C1694 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout VDD 2.07863f
C1695 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.09975f
C1696 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout a_41687_13083# 0.04995f
C1697 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.04107f
C1698 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout CLK 0.03574f
C1699 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Qbar 1.16087f
C1700 a_128237_19786# a_128851_19786# 0.05935f
C1701 D_FlipFlop_6.Nand_Gate_1.Vout Q1 0.06993f
C1702 a_132311_39721# a_132925_39721# 0.05935f
C1703 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.06955f
C1704 a_86591_52572# EN 0.045f
C1705 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_0.Vout 0.07084f
C1706 Nand_Gate_7.A a_61795_15797# 0.06113f
C1707 D_FlipFlop_4.Nand_Gate_1.Vout a_128237_27764# 0.04444f
C1708 a_45761_15797# VDD 0.03119f
C1709 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.06935f
C1710 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B a_79495_13083# 0.04995f
C1711 And_Gate_5.Nand_Gate_0.Vout a_59605_47663# 0.06113f
C1712 a_94915_13083# a_95529_13083# 0.05935f
C1713 a_71017_47663# CLK 0.02953f
C1714 a_59605_47663# VDD 0.02521f
C1715 Nand_Gate_1.B a_132925_30478# 0.04789f
C1716 a_53471_52572# VDD 0.01186f
C1717 Nand_Gate_2.A D_FlipFlop_3.Qbar 0.06962f
C1718 D_FlipFlop_7.Nand_Gate_1.Vout a_130209_17072# 0.05964f
C1719 a_85233_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.05964f
C1720 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1541f
C1721 Nand_Gate_0.A a_128851_39721# 0.04625f
C1722 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B VDD 1.79521f
C1723 RingCounter_0.D_FlipFlop_3.Qbar Nand_Gate_0.B 1.10693f
C1724 D_FlipFlop_1.3-input-nand_1.Vout a_132925_33443# 0.04543f
C1725 FFCLR EN 2.21589f
C1726 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.09975f
C1727 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B a_46375_13083# 0.04995f
C1728 a_58159_49858# VDD 0.02906f
C1729 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_124399_49858# 0.04444f
C1730 D_FlipFlop_1.3-input-nand_2.Vout a_130209_36157# 0.04443f
C1731 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_74807_13083# 0.04443f
C1732 RingCounter_0.D_FlipFlop_8.Qbar a_40329_13083# 0.01335f
C1733 a_94915_13083# VDD 0.02521f
C1734 D_FlipFlop_0.Nand_Gate_1.Vout Q4 0.06993f
C1735 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_110643_15797# 0.04995f
C1736 Nand_Gate_4.B RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0839f
C1737 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_65869_13083# 0.04443f
C1738 Nand_Gate_0.B RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.08377f
C1739 D_FlipFlop_6.Nand_Gate_0.Vout a_130209_23350# 0.05964f
C1740 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_86591_49858# 0.01335f
C1741 Nand_Gate_2.B And_Gate_6.Nand_Gate_0.Vout 0.02391f
C1742 D_FlipFlop_0.CLK D_FlipFlop_0.Nand_Gate_0.Vout 0.01448f
C1743 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C CLK 0.30901f
C1744 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 1.09946f
C1745 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_123041_15797# 0.05964f
C1746 CDAC8_0.switch_9.Z CDAC8_0.switch_7.Z 3.75058f
C1747 a_95529_15797# EN 0.04443f
C1748 D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.48313f
C1749 D_FlipFlop_2.3-input-nand_2.C VDD 2.74431f
C1750 Nand_Gate_1.B Comparator_0.Vinm 1.25742f
C1751 And_Gate_5.Nand_Gate_0.Vout CLK 0.4651f
C1752 Nand_Gate_7.B a_73449_15797# 0.01335f
C1753 RingCounter_0.D_FlipFlop_3.Qbar RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.11654f
C1754 a_134283_43285# a_134897_43285# 0.05935f
C1755 a_72835_13083# a_73449_13083# 0.05935f
C1756 D_FlipFlop_5.Nand_Gate_0.Vout a_130209_26914# 0.05964f
C1757 FFCLR Nand_Gate_5.B 0.06347f
C1758 VDD CLK 82.6031f
C1759 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout EN 0.13192f
C1760 a_100961_15797# CLK 0.04619f
C1761 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B a_85233_49858# 0.04443f
C1762 a_99603_15797# VDD 0.03339f
C1763 Nand_Gate_1.A a_101575_15797# 0.04995f
C1764 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.09975f
C1765 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121069_13083# 0.05964f
C1766 D_FlipFlop_1.3-input-nand_2.Vout VDD 2.77266f
C1767 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout CLK 0.03574f
C1768 a_40459_52572# EN 0.04454f
C1769 D_FlipFlop_0.3-input-nand_1.B a_134283_44135# 0.04443f
C1770 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_76165_49858# 0.05964f
C1771 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout EN 0.62384f
C1772 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout VDD 2.31704f
C1773 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout a_100347_49858# 0.04995f
C1774 CDAC8_0.switch_1.Z VDD 1.11469f
C1775 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 1.09975f
C1776 D_FlipFlop_7.3-input-nand_0.Vout a_134897_19786# 0.01335f
C1777 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.04109f
C1778 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.16429f
C1779 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Inverter_1.Vout 0.25963f
C1780 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout a_87205_49858# 0.04443f
C1781 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_84489_15797# 0.04995f
C1782 D_FlipFlop_1.Inverter_1.Vout Comparator_0.Vinm 0.0387f
C1783 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B VDD 1.73782f
C1784 D_FlipFlop_2.3-input-nand_0.Vout a_132925_39721# 0.04995f
C1785 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD 2.04843f
C1786 a_50755_13083# VDD 0.02521f
C1787 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.06955f
C1788 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_78881_15797# 0.05964f
C1789 a_128237_30478# Q3 0.06113f
C1790 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout VDD 2.8604f
C1791 FFCLR a_132925_37007# 0.045f
C1792 Nand_Gate_2.A a_95659_52572# 0.04995f
C1793 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.26069f
C1794 RingCounter_0.D_FlipFlop_4.Qbar a_91279_52572# 0.04443f
C1795 RingCounter_0.D_FlipFlop_5.Qbar a_101705_49858# 0.01335f
C1796 Nand_Gate_2.A a_128851_43285# 0.04627f
C1797 a_134283_17072# VDD 0.02521f
C1798 D_FlipFlop_6.3-input-nand_2.Vout a_130209_23350# 0.04443f
C1799 Nand_Gate_4.B a_46375_15797# 0.04995f
C1800 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.06955f
C1801 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.04107f
C1802 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout CLK 0.30716f
C1803 a_106699_49858# a_107313_49858# 0.05935f
C1804 D_FlipFlop_7.Nand_Gate_0.Vout a_128237_19786# 0.04444f
C1805 a_85233_49858# CLK 0.04619f
C1806 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout Nand_Gate_0.B 0.12214f
C1807 FFCLR D_FlipFlop_1.3-input-nand_1.B 0.46505f
C1808 a_50755_13083# a_51369_13083# 0.05935f
C1809 a_84619_49858# VDD 0.01712f
C1810 a_134897_33443# EN 0.04304f
C1811 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout CLK 0.71245f
C1812 VDD Q0 4.32049f
C1813 D_FlipFlop_0.3-input-nand_1.Vout a_134283_44135# 0.05964f
C1814 FFCLR D_FlipFlop_7.3-input-nand_2.C 0.76213f
C1815 D_FlipFlop_5.3-input-nand_2.Vout VDD 2.77266f
C1816 D_FlipFlop_1.3-input-nand_2.Vout a_132311_36157# 0.05964f
C1817 a_117609_13083# VDD 0.0563f
C1818 EN Q7 0.26571f
C1819 CDAC8_0.switch_8.Z Q6 0.24676f
C1820 D_FlipFlop_5.3-input-nand_2.Vout a_130209_26914# 0.04443f
C1821 FFCLR a_134897_40571# 0.04023f
C1822 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C CLK 0.30966f
C1823 a_128851_40571# VDD 0.01186f
C1824 D_FlipFlop_7.Qbar Q0 1.09842f
C1825 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_0.Vout 1.03458f
C1826 a_63767_15797# VDD 0.02906f
C1827 RingCounter_0.D_FlipFlop_14.Qbar a_61795_15797# 0.04443f
C1828 RingCounter_0.D_FlipFlop_3.Qbar VDD 1.96503f
C1829 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_34721_15797# 0.05964f
C1830 RingCounter_0.D_FlipFlop_9.Qbar VDD 1.95446f
C1831 RingCounter_0.D_FlipFlop_15.Qbar VDD 1.95446f
C1832 VDD Vbias 0.35746p
C1833 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.26069f
C1834 Nand_Gate_2.A D_FlipFlop_0.CLK 0.06055f
C1835 And_Gate_6.Nand_Gate_0.Vout Comparator_0.Vinm 0.02639f
C1836 Nand_Gate_2.B a_102319_49858# 0.04741f
C1837 a_128851_19786# VDD 0.01186f
C1838 a_134283_17072# a_134897_17072# 0.05935f
C1839 a_132925_39721# VDD 0.01186f
C1840 Nand_Gate_5.Vout CLK 2.38648f
C1841 D_FlipFlop_4.3-input-nand_2.Vout a_130209_30478# 0.04443f
C1842 CDAC8_0.switch_7.Z Q1 1.51854f
C1843 D_FlipFlop_3.Nand_Gate_1.Vout a_128851_40571# 0.04995f
C1844 D_FlipFlop_7.3-input-nand_1.Vout a_132925_17072# 0.04543f
C1845 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Qbar 1.05791f
C1846 D_FlipFlop_3.3-input-nand_2.C a_132925_40571# 0.01335f
C1847 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B EN 0.43216f
C1848 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_0.Vout 1.03511f
C1849 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.04109f
C1850 a_116995_15797# VDD 0.0299f
C1851 RingCounter_0.D_FlipFlop_7.Qbar RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.11654f
C1852 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.07084f
C1853 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD 1.86552f
C1854 CDAC8_0.switch_8.Z Comparator_0.Vinm 0.10659p
C1855 And_Gate_3.Nand_Gate_0.Vout VDD 1.53086f
C1856 a_119711_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.01335f
C1857 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.26069f
C1858 FFCLR D_FlipFlop_1.3-input-nand_1.Vout 0.15444f
C1859 FFCLR CDAC8_0.switch_9.Z 2.17565f
C1860 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Inverter_1.Vout 0.25963f
C1861 a_78267_52572# RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.05964f
C1862 a_132311_44135# VDD 0.02521f
C1863 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0846f
C1864 FFCLR a_134897_26914# 0.08436f
C1865 Nand_Gate_5.B Q7 0.06203f
C1866 RingCounter_0.D_FlipFlop_15.Qbar a_51369_13083# 0.01335f
C1867 a_84619_49858# a_85233_49858# 0.05935f
C1868 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.06955f
C1869 a_41073_49858# CLK 0.04443f
C1870 a_128237_33443# Q7 0.04443f
C1871 a_40459_49858# VDD 0.05707f
C1872 a_28675_13083# a_29289_13083# 0.05935f
C1873 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout CLK 0.23566f
C1874 Nand_Gate_4.B VDD 8.57999f
C1875 D_FlipFlop_3.Qbar Q5 1.06173f
C1876 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_88563_15797# 0.01335f
C1877 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_86591_49858# 0.04543f
C1878 a_130209_23350# VDD 0.02521f
C1879 a_134897_43285# VDD 0.01186f
C1880 a_101705_52572# a_102319_52572# 0.05935f
C1881 a_73449_13083# VDD 0.0563f
C1882 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.04109f
C1883 Nand_Gate_6.A a_82057_16975# 0.0476f
C1884 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_1.Vout 0.08671f
C1885 D_FlipFlop_0.CLK D_FlipFlop_0.Inverter_1.Vout 0.2871f
C1886 D_FlipFlop_7.Qbar Nand_Gate_4.B 0.06645f
C1887 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.26069f
C1888 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.06935f
C1889 D_FlipFlop_1.Qbar a_128851_33443# 0.01335f
C1890 a_54085_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.05964f
C1891 D_FlipFlop_6.Nand_Gate_1.Vout a_130209_20636# 0.05964f
C1892 Nand_Gate_2.A RingCounter_0.D_FlipFlop_5.3-input-nand_1.B 0.29683f
C1893 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout CLK 0.6891f
C1894 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_91279_52572# 0.04444f
C1895 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C CLK 0.30901f
C1896 a_28675_15797# VDD 0.02521f
C1897 D_FlipFlop_6.3-input-nand_2.Vout a_132311_23350# 0.05964f
C1898 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.16429f
C1899 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0846f
C1900 a_130209_30478# VDD 0.02521f
C1901 a_108671_49858# CLK 0.03129f
C1902 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout CLK 0.30606f
C1903 a_107313_49858# VDD 0.0325f
C1904 D_FlipFlop_1.3-input-nand_1.B a_134897_33443# 0.04995f
C1905 Nand_Gate_1.B EN 1.13628f
C1906 D_FlipFlop_7.3-input-nand_2.Vout a_132311_17072# 0.04443f
C1907 a_107313_52572# CLK 0.04619f
C1908 Nand_Gate_4.B a_134897_17072# 0.04583f
C1909 D_FlipFlop_5.Nand_Gate_1.Vout a_130209_24200# 0.05964f
C1910 a_106699_52572# VDD 0.0564f
C1911 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B a_106699_49858# 0.04995f
C1912 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_0.Vout 0.0846f
C1913 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout EN 0.61318f
C1914 VDD Q4 3.72299f
C1915 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.07084f
C1916 D_FlipFlop_5.3-input-nand_2.Vout a_132311_26914# 0.05964f
C1917 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_97631_49858# 0.01335f
C1918 a_62539_49858# a_63153_49858# 0.05935f
C1919 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_32749_13083# 0.05964f
C1920 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110029_15797# 0.04443f
C1921 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.48392f
C1922 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout EN 0.78747f
C1923 Nand_Gate_6.B Comparator_0.Vinm 1.96281f
C1924 D_FlipFlop_4.Nand_Gate_1.Vout a_130209_27764# 0.05964f
C1925 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.Vout 0.01194f
C1926 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.C 0.01194f
C1927 a_29289_13083# VDD 0.0563f
C1928 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B VDD 1.73782f
C1929 Nand_Gate_2.B CLK 0.41441f
C1930 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_96887_15797# 0.04443f
C1931 a_102319_52572# VDD 0.02521f
C1932 a_93097_47663# CLK 0.02953f
C1933 Nand_Gate_2.A Nand_Gate_2.Vout 0.11161f
C1934 FFCLR D_FlipFlop_0.Qbar 0.03748f
C1935 D_FlipFlop_1.Inverter_1.Vout EN 0.59727f
C1936 D_FlipFlop_4.3-input-nand_2.Vout a_132311_30478# 0.05964f
C1937 a_81685_47663# VDD 0.02521f
C1938 a_116995_15797# a_117609_15797# 0.05935f
C1939 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_109285_52572# 0.04444f
C1940 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_44403_15797# 0.01335f
C1941 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout VDD 2.8604f
C1942 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Qbar 1.05791f
C1943 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B a_96273_49858# 0.04443f
C1944 Nand_Gate_5.B Nand_Gate_1.B 0.06366f
C1945 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_90665_49858# 0.04995f
C1946 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.04109f
C1947 a_48565_16975# CLK 0.04479f
C1948 Nand_Gate_7.B a_59977_16975# 0.04443f
C1949 a_37897_16975# VDD 0.02521f
C1950 Nand_Gate_4.B D_FlipFlop_7.Inverter_1.Vout 0.16546f
C1951 D_FlipFlop_1.3-input-nand_1.Vout a_134897_33443# 0.01335f
C1952 CDAC8_0.switch_6.Z CDAC8_0.switch_7.Z 14.5275f
C1953 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.Vout 0.01194f
C1954 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.C 0.01194f
C1955 a_64511_49858# CLK 0.03129f
C1956 D_FlipFlop_1.3-input-nand_2.C VDD 2.74431f
C1957 a_132311_44135# a_132925_44135# 0.05935f
C1958 a_63153_49858# VDD 0.0325f
C1959 D_FlipFlop_4.Qbar Q3 1.06575f
C1960 RingCounter_0.D_FlipFlop_16.Q a_41073_52572# 0.04443f
C1961 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_77523_13083# 0.01335f
C1962 CDAC8_0.switch_9.Z Q7 0.29749f
C1963 a_128851_43285# Q5 0.01335f
C1964 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout VDD 2.0863f
C1965 D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.48313f
C1966 a_98989_13083# CLK 0.03129f
C1967 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout a_98245_49858# 0.04443f
C1968 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Qbar 1.05791f
C1969 a_96887_13083# VDD 0.02578f
C1970 FFCLR D_FlipFlop_6.3-input-nand_1.B 0.44757f
C1971 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout VDD 2.88547f
C1972 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_112615_15797# 0.01335f
C1973 a_64511_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.01335f
C1974 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.26069f
C1975 a_132311_23350# VDD 0.02521f
C1976 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_89307_49858# 0.04443f
C1977 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.Nand_Gate_1.Vout 0.1541f
C1978 a_40459_49858# a_41073_49858# 0.05935f
C1979 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.25963f
C1980 D_FlipFlop_7.Qbar D_FlipFlop_7.Nand_Gate_0.Vout 0.07122f
C1981 RingCounter_0.D_FlipFlop_17.Qbar EN 0.03751f
C1982 a_95659_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.01335f
C1983 a_106569_15797# EN 0.04443f
C1984 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout a_42431_52572# 0.04995f
C1985 a_87949_15797# VDD 0.03178f
C1986 a_72835_15797# a_73449_15797# 0.05935f
C1987 a_108671_52572# EN 0.045f
C1988 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout CLK 0.30735f
C1989 D_FlipFlop_3.3-input-nand_1.Vout a_132311_40571# 0.04444f
C1990 FFCLR D_FlipFlop_4.3-input-nand_1.B 0.44757f
C1991 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK 0.69908f
C1992 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout EN 1.03583f
C1993 a_73449_15797# VDD 0.01571f
C1994 a_132311_30478# VDD 0.02521f
C1995 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_0.Vout 0.0846f
C1996 And_Gate_6.Nand_Gate_0.Vout EN 0.0623f
C1997 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B CLK 0.16274f
C1998 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout CLK 0.29759f
C1999 a_101575_15797# VDD 0.06072f
C2000 a_75551_52572# VDD 0.01186f
C2001 RingCounter_0.D_FlipFlop_7.Qbar a_113359_49858# 0.06113f
C2002 Nand_Gate_2.A Q5 1.05014f
C2003 a_100961_15797# a_101575_15797# 0.05935f
C2004 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.08641f
C2005 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_99603_15797# 0.04995f
C2006 CLK Q6 0.1175f
C2007 D_FlipFlop_5.3-input-nand_2.C VDD 2.74431f
C2008 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121069_15797# 0.04443f
C2009 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_50755_15797# 0.04444f
C2010 D_FlipFlop_1.3-input-nand_2.C a_132311_36157# 0.04443f
C2011 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B VDD 1.79521f
C2012 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout EN 0.08653f
C2013 CDAC8_0.switch_8.Z EN 1.97671f
C2014 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD 1.56255f
C2015 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout VDD 2.86518f
C2016 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_0.Vout 0.0846f
C2017 FFCLR D_FlipFlop_6.3-input-nand_1.Vout 0.95879f
C2018 Nand_Gate_4.A a_35335_15797# 0.04995f
C2019 a_112615_13083# EN 0.0452f
C2020 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.30154f
C2021 a_54829_13083# CLK 0.03129f
C2022 D_FlipFlop_2.3-input-nand_2.C a_130209_37007# 0.04443f
C2023 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout VDD 2.14483f
C2024 RingCounter_0.D_FlipFlop_11.Qbar a_94915_13083# 0.06113f
C2025 D_FlipFlop_2.3-input-nand_0.Vout a_134897_39721# 0.01335f
C2026 a_52727_13083# VDD 0.02578f
C2027 a_28675_15797# a_29289_15797# 0.05935f
C2028 Nand_Gate_2.A RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.08377f
C2029 FFCLR a_134897_37007# 0.04073f
C2030 D_FlipFlop_2.Nand_Gate_0.Vout a_128237_39721# 0.04444f
C2031 D_FlipFlop_6.3-input-nand_1.Vout a_132925_20636# 0.04543f
C2032 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Nand_Gate_1.Vout 0.04109f
C2033 a_128851_37007# VDD 0.01186f
C2034 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_0.Vout 0.0846f
C2035 FFCLR D_FlipFlop_4.3-input-nand_1.Vout 0.95879f
C2036 Comparator_0.Vinm CLK 2.97464f
C2037 Nand_Gate_5.A D_FlipFlop_0.Nand_Gate_0.Vout 0.65107f
C2038 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C EN 0.07664f
C2039 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.3-input-nand_2.Vout 0.16429f
C2040 Nand_Gate_6.A a_83875_13083# 0.04443f
C2041 D_FlipFlop_1.3-input-nand_2.Vout Comparator_0.Vinm 0.01683f
C2042 D_FlipFlop_7.3-input-nand_1.Vout VDD 1.78032f
C2043 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_120325_52572# 0.04443f
C2044 a_87205_49858# CLK 0.03129f
C2045 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Inverter_1.Vout 0.25963f
C2046 a_45147_52572# RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.05964f
C2047 FFCLR a_128851_24200# 0.04443f
C2048 a_132925_36157# VDD 0.01186f
C2049 a_86591_49858# VDD 0.06071f
C2050 RingCounter_0.D_FlipFlop_11.Qbar CLK 0.09276f
C2051 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.08671f
C2052 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_76909_15797# 0.04443f
C2053 D_FlipFlop_5.3-input-nand_1.Vout a_132925_24200# 0.04543f
C2054 CDAC8_0.switch_1.Z Comparator_0.Vinm 6.31039f
C2055 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C VDD 3.56545f
C2056 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout a_96887_15797# 0.04443f
C2057 a_121683_13083# CLK 0.03129f
C2058 D_FlipFlop_1.Nand_Gate_1.Vout Q7 0.06993f
C2059 a_121069_13083# VDD 0.02578f
C2060 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout a_89307_52572# 0.04443f
C2061 a_52113_52572# CLK 0.04619f
C2062 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.30154f
C2063 FFCLR CDAC8_0.switch_6.Z 6.54715f
C2064 a_106699_52572# a_107313_52572# 0.05935f
C2065 a_132311_40571# VDD 0.02521f
C2066 a_51499_52572# VDD 0.0564f
C2067 D_FlipFlop_6.3-input-nand_0.Vout VDD 1.77946f
C2068 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout EN 0.61318f
C2069 a_128237_37007# a_128851_37007# 0.05935f
C2070 a_68455_13083# EN 0.0452f
C2071 D_FlipFlop_4.3-input-nand_1.Vout a_132925_27764# 0.04543f
C2072 D_FlipFlop_2.Qbar Q5 0.01194f
C2073 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 1.09975f
C2074 a_134897_39721# VDD 0.01186f
C2075 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Qbar 0.07122f
C2076 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout EN 0.78734f
C2077 D_FlipFlop_6.3-input-nand_2.C a_132311_23350# 0.04443f
C2078 D_FlipFlop_7.3-input-nand_1.Vout a_134897_17072# 0.01335f
C2079 Nand_Gate_6.B EN 1.25083f
C2080 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_95659_49858# 0.01335f
C2081 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout VDD 2.74107f
C2082 D_FlipFlop_4.3-input-nand_0.Vout VDD 1.77946f
C2083 Nand_Gate_2.B a_106699_52572# 0.04995f
C2084 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout VDD 2.31704f
C2085 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B a_117739_49858# 0.04995f
C2086 Comparator_0.Vinm Q0 0.13685f
C2087 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_32749_15797# 0.04443f
C2088 a_134283_44135# VDD 0.02521f
C2089 D_FlipFlop_7.3-input-nand_2.C a_132311_17072# 0.05964f
C2090 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_54829_15797# 0.05964f
C2091 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_52113_49858# 0.05964f
C2092 a_132925_26914# VDD 0.01186f
C2093 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_45147_49858# 0.05964f
C2094 a_128851_23350# Q1 0.01335f
C2095 a_132311_36157# a_132925_36157# 0.05935f
C2096 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_40459_49858# 0.01335f
C2097 a_43045_49858# CLK 0.03129f
C2098 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout CLK 0.30716f
C2099 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_0.Vout 0.07084f
C2100 a_42431_49858# VDD 0.01186f
C2101 D_FlipFlop_5.3-input-nand_2.C a_132311_26914# 0.04443f
C2102 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0846f
C2103 FFCLR D_FlipFlop_6.Nand_Gate_1.Vout 0.61318f
C2104 a_77523_13083# CLK 0.03129f
C2105 Nand_Gate_6.B a_90535_15797# 0.04995f
C2106 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110029_15797# 0.05964f
C2107 a_102319_52572# Nand_Gate_2.B 0.06113f
C2108 a_76909_13083# VDD 0.02578f
C2109 Comparator_0.Vinm Vbias 1.12875f
C2110 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.3-input-nand_2.Vout 0.16429f
C2111 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_109285_49858# 0.05964f
C2112 Nand_Gate_5.B Nand_Gate_6.B 0.06371f
C2113 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.16429f
C2114 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout CLK 0.68793f
C2115 a_39715_15797# VDD 0.02906f
C2116 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_17.3-input-nand_1.B 0.29683f
C2117 RingCounter_0.D_FlipFlop_17.Qbar a_46505_49858# 0.01335f
C2118 RingCounter_0.D_FlipFlop_5.Qbar VDD 1.96503f
C2119 D_FlipFlop_4.3-input-nand_2.C a_132311_30478# 0.04443f
C2120 FFCLR D_FlipFlop_4.Nand_Gate_1.Vout 0.61318f
C2121 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.07084f
C2122 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout VDD 2.29866f
C2123 Nand_Gate_6.A a_79495_15797# 0.04995f
C2124 Nand_Gate_5.A D_FlipFlop_0.CLK 3.64288f
C2125 D_FlipFlop_5.Qbar Q3 0.01194f
C2126 a_53471_52572# EN 0.045f
C2127 a_109285_49858# VDD 0.0301f
C2128 a_46505_52572# FFCLR 0.01335f
C2129 D_FlipFlop_7.Nand_Gate_1.Vout VDD 1.46545f
C2130 D_FlipFlop_0.CLK a_134283_46849# 0.04443f
C2131 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_2.Vout 0.18665f
C2132 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B EN 0.43216f
C2133 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.06955f
C2134 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.04107f
C2135 Nand_Gate_1.B Q1 0.05915f
C2136 Nand_Gate_4.B Comparator_0.Vinm 1.16732f
C2137 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout a_118967_13083# 0.04995f
C2138 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD 1.86552f
C2139 CDAC8_0.switch_8.Z CDAC8_0.switch_9.Z 7.4006f
C2140 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout VDD 2.73822f
C2141 D_FlipFlop_7.Qbar D_FlipFlop_7.Nand_Gate_1.Vout 0.11654f
C2142 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_100347_49858# 0.04443f
C2143 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B VDD 1.79521f
C2144 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_65125_52572# 0.04443f
C2145 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_101705_52572# 0.04995f
C2146 a_134283_39721# a_134897_39721# 0.05935f
C2147 CDAC8_0.switch_6.Z Q7 0.66797f
C2148 a_33363_13083# CLK 0.02953f
C2149 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.25963f
C2150 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_56187_49858# 0.05964f
C2151 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout CLK 0.69861f
C2152 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.1182f
C2153 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout a_78267_52572# 0.04443f
C2154 a_32749_13083# VDD 0.02578f
C2155 a_68585_52572# VDD 0.01186f
C2156 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout 0.30154f
C2157 a_115177_47663# CLK 0.06931f
C2158 a_103765_47663# VDD 0.02521f
C2159 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_1.B 0.27862f
C2160 Nand_Gate_5.A D_FlipFlop_0.Inverter_1.Vout 0.15693f
C2161 a_132311_23350# a_132925_23350# 0.05935f
C2162 RingCounter_0.D_FlipFlop_6.Qbar a_124399_49858# 0.06113f
C2163 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout VDD 2.16852f
C2164 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_0.Vout 0.07084f
C2165 a_70645_16975# CLK 0.04479f
C2166 Nand_Gate_2.B RingCounter_0.D_FlipFlop_7.3-input-nand_1.B 0.29683f
C2167 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.06993f
C2168 Nand_Gate_1.Vout a_104137_16975# 0.05964f
C2169 a_59977_16975# VDD 0.02521f
C2170 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.3-input-nand_2.Vout 0.06935f
C2171 FFCLR D_FlipFlop_3.Inverter_1.Vout 0.56927f
C2172 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C CLK 0.30901f
C2173 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B a_90535_13083# 0.04995f
C2174 EN CLK 8.56318f
C2175 Comparator_0.Vinm Q4 1.26254f
C2176 a_65125_49858# VDD 0.0301f
C2177 a_112745_52572# Nand_Gate_5.A 0.01335f
C2178 D_FlipFlop_1.3-input-nand_0.Vout a_132925_36157# 0.04995f
C2179 a_99603_15797# EN 0.045f
C2180 D_FlipFlop_1.3-input-nand_2.Vout EN 0.07759f
C2181 a_100961_13083# CLK 0.04619f
C2182 a_75898_25104# Q2 0.50364f
C2183 a_132311_26914# a_132925_26914# 0.05935f
C2184 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_0.Vout 0.07084f
C2185 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_2.Inverter_1.Vout 0.01422f
C2186 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout EN 0.09127f
C2187 a_87949_15797# a_88563_15797# 0.05935f
C2188 a_99603_13083# VDD 0.05686f
C2189 CDAC8_0.switch_1.Z EN 0.15062f
C2190 a_61795_15797# VDD 0.02906f
C2191 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_2.Vout 0.90723f
C2192 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_119711_52572# 0.04995f
C2193 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_85847_13083# 0.04443f
C2194 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B EN 0.26843f
C2195 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0846f
C2196 D_FlipFlop_1.Inverter_1.Vout a_130209_33443# 0.04995f
C2197 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout EN 0.97979f
C2198 a_89921_15797# VDD 0.03119f
C2199 RingCounter_0.D_FlipFlop_1.Qbar RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.11654f
C2200 D_FlipFlop_6.3-input-nand_1.B a_134897_20636# 0.04995f
C2201 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout 0.30154f
C2202 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD 1.56255f
C2203 a_132311_30478# a_132925_30478# 0.05935f
C2204 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout CLK 0.03574f
C2205 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.48392f
C2206 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout EN 0.78747f
C2207 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_0.Vout 0.07084f
C2208 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_76909_13083# 0.04443f
C2209 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_1.Vout 0.07295f
C2210 D_FlipFlop_3.3-input-nand_1.Vout a_134283_40571# 0.05964f
C2211 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout CLK 0.03479f
C2212 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_65869_15797# 0.04444f
C2213 Nand_Gate_5.B CLK 0.29423f
C2214 a_124399_52572# VDD 0.02521f
C2215 D_FlipFlop_1.3-input-nand_2.C Comparator_0.Vinm 0.03357f
C2216 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout VDD 2.8604f
C2217 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_101575_15797# 0.01335f
C2218 a_75551_52572# a_76165_52572# 0.05935f
C2219 D_FlipFlop_5.3-input-nand_1.B a_134897_24200# 0.04995f
C2220 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.25963f
C2221 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout VDD 2.88547f
C2222 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout CLK 0.71245f
C2223 a_84619_49858# EN 0.07058f
C2224 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_54085_52572# 0.04444f
C2225 a_128237_24200# Q2 0.04443f
C2226 EN Q0 0.24699f
C2227 a_56801_13083# CLK 0.04619f
C2228 D_FlipFlop_2.Nand_Gate_1.Vout a_128851_37007# 0.04995f
C2229 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_106569_13083# 0.04995f
C2230 D_FlipFlop_2.3-input-nand_2.C a_132925_37007# 0.01335f
C2231 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.3-input-nand_2.Vout 0.06935f
C2232 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_99603_13083# 0.04543f
C2233 a_55443_13083# VDD 0.05686f
C2234 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_94915_13083# 0.04444f
C2235 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.06955f
C2236 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_87949_13083# 0.04444f
C2237 D_FlipFlop_4.3-input-nand_1.B a_134897_27764# 0.04995f
C2238 FFCLR CDAC8_0.switch_7.Z 11.2108f
C2239 D_FlipFlop_6.3-input-nand_1.Vout a_134897_20636# 0.01335f
C2240 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Inverter_1.Vout 0.25963f
C2241 a_132311_37007# VDD 0.02521f
C2242 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.08641f
C2243 D_FlipFlop_4.Qbar a_128851_27764# 0.01335f
C2244 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.04107f
C2245 And_Gate_4.Nand_Gate_0.Vout CLK 0.50205f
C2246 D_FlipFlop_6.3-input-nand_0.Vout a_132925_23350# 0.04995f
C2247 D_FlipFlop_0.Qbar a_128851_44135# 0.01335f
C2248 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_41687_15797# 0.05964f
C2249 a_108671_49858# a_109285_49858# 0.05935f
C2250 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B a_56801_13083# 0.04443f
C2251 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C VDD 3.56545f
C2252 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout EN 1.03583f
C2253 Nand_Gate_5.B Q0 0.06203f
C2254 a_134897_36157# VDD 0.01186f
C2255 a_89307_49858# VDD 0.04111f
C2256 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.06935f
C2257 And_Gate_3.Nand_Gate_0.Vout EN 0.02316f
C2258 D_FlipFlop_5.3-input-nand_1.Vout a_134897_24200# 0.01335f
C2259 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout CLK 0.03574f
C2260 Nand_Gate_0.A Nand_Gate_0.B 0.08217f
C2261 a_130209_19786# VDD 0.02521f
C2262 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_96887_15797# 0.05964f
C2263 a_123041_13083# VDD 0.02865f
C2264 D_FlipFlop_5.3-input-nand_0.Vout a_132925_26914# 0.04995f
C2265 a_97631_52572# VDD 0.01186f
C2266 a_121069_15797# VDD 0.03178f
C2267 a_107313_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.05964f
C2268 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.04109f
C2269 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_39715_13083# 0.04444f
C2270 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_41687_15797# 0.04443f
C2271 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD 1.86552f
C2272 a_40459_49858# EN 0.02716f
C2273 D_FlipFlop_6.Qbar a_128237_20636# 0.06113f
C2274 a_134283_40571# VDD 0.02521f
C2275 Nand_Gate_4.B EN 1.52428f
C2276 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_32749_13083# 0.04444f
C2277 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout a_30647_13083# 0.04995f
C2278 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_120325_49858# 0.05964f
C2279 RingCounter_0.D_FlipFlop_5.Qbar Nand_Gate_2.B 1.10693f
C2280 RingCounter_0.D_FlipFlop_14.Qbar RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.07122f
C2281 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.3-input-nand_2.Vout 0.16429f
C2282 D_FlipFlop_4.3-input-nand_1.Vout a_134897_27764# 0.01335f
C2283 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.04109f
C2284 RingCounter_0.D_FlipFlop_4.Qbar RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.11654f
C2285 D_FlipFlop_4.3-input-nand_0.Vout a_132925_30478# 0.04995f
C2286 RingCounter_0.D_FlipFlop_16.Q a_28675_13083# 0.04443f
C2287 D_FlipFlop_5.Qbar a_128237_24200# 0.06113f
C2288 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_97631_49858# 0.04543f
C2289 Nand_Gate_2.B RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.08377f
C2290 Nand_Gate_6.B Q1 0.06203f
C2291 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD 1.56255f
C2292 Nand_Gate_1.B RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0839f
C2293 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_64511_52572# 0.04995f
C2294 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout VDD 2.88547f
C2295 CDAC8_0.switch_5.Z Q2 0.06367f
C2296 CDAC8_0.switch_9.Z CLK 0.19385f
C2297 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_2.C 0.29677f
C2298 a_75898_42964# VDD 1.30491f
C2299 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_54085_49858# 0.04444f
C2300 a_107313_49858# EN 0.01149f
C2301 a_134283_26914# VDD 0.02521f
C2302 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_47119_49858# 0.04444f
C2303 a_86591_49858# a_87205_49858# 0.05935f
C2304 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.06955f
C2305 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_42431_49858# 0.04543f
C2306 D_FlipFlop_6.Qbar Q1 1.06476f
C2307 VDD Q3 3.60365f
C2308 Nand_Gate_5.B Nand_Gate_4.B 0.06408f
C2309 a_45147_49858# VDD 0.04055f
C2310 a_32749_15797# VDD 0.02793f
C2311 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout CLK 0.71127f
C2312 CDAC8_0.switch_9.Z CDAC8_0.switch_1.Z 0.14339f
C2313 EN Q4 0.2481f
C2314 Nand_Gate_7.B CDAC8_0.switch_2.Z 0.33658f
C2315 a_78881_13083# VDD 0.02865f
C2316 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_0.Vout 1.0061f
C2317 Nand_Gate_0.A a_71017_47663# 0.04705f
C2318 CDAC8_0.switch_8.Z CDAC8_0.switch_6.Z 3.59863f
C2319 RingCounter_0.D_FlipFlop_14.Qbar a_62409_13083# 0.01335f
C2320 a_121069_13083# a_121683_13083# 0.05935f
C2321 a_74193_52572# CLK 0.04619f
C2322 RingCounter_0.D_FlipFlop_2.Qbar CLK 0.09276f
C2323 a_73579_52572# VDD 0.0564f
C2324 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.06993f
C2325 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout EN 0.61318f
C2326 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout VDD 2.31704f
C2327 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B EN 0.26843f
C2328 a_51499_52572# a_52113_52572# 0.05935f
C2329 a_132311_40571# a_132925_40571# 0.05935f
C2330 Nand_Gate_6.B Nand_Gate_6.Vout 2.38777f
C2331 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD 1.48368f
C2332 CDAC8_0.switch_7.Z Q7 1.88958f
C2333 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.3-input-nand_2.C 0.26069f
C2334 D_FlipFlop_7.Inverter_1.Vout a_130209_19786# 0.04443f
C2335 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout EN 0.78747f
C2336 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_1.B 0.06986f
C2337 a_112745_49858# VDD 0.06015f
C2338 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.06955f
C2339 Nand_Gate_5.A a_117739_52572# 0.04995f
C2340 FFCLR D_FlipFlop_7.3-input-nand_1.B 0.40157f
C2341 RingCounter_0.D_FlipFlop_16.Q VDD 3.42681f
C2342 a_132311_19786# VDD 0.02521f
C2343 RingCounter_0.D_FlipFlop_7.Qbar a_113359_52572# 0.04443f
C2344 CDAC8_0.switch_9.Z Q0 0.14628f
C2345 Nand_Gate_5.B Q4 0.06203f
C2346 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.06955f
C2347 D_FlipFlop_1.3-input-nand_2.C EN 0.79121f
C2348 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.06993f
C2349 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110029_13083# 0.05964f
C2350 a_63153_49858# EN 0.01149f
C2351 FFCLR a_132925_20636# 0.045f
C2352 FFCLR D_FlipFlop_2.Inverter_1.Vout 0.57257f
C2353 a_64511_49858# a_65125_49858# 0.05935f
C2354 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_101705_49858# 0.04995f
C2355 Nand_Gate_1.B a_112615_15797# 0.04995f
C2356 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.09975f
C2357 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout CLK 0.20785f
C2358 D_FlipFlop_2.3-input-nand_1.Vout a_132311_37007# 0.04444f
C2359 D_FlipFlop_3.Qbar a_128237_40571# 0.06113f
C2360 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_2.B 0.12214f
C2361 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_110029_13083# 0.04444f
C2362 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_2.C 0.15106f
C2363 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout EN 0.78668f
C2364 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout CLK 0.23507f
C2365 a_43045_52572# VDD 0.02865f
C2366 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_58159_49858# 0.04444f
C2367 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.08641f
C2368 a_34721_13083# VDD 0.02865f
C2369 Nand_Gate_0.A VDD 8.22095f
C2370 RingCounter_0.D_FlipFlop_8.Qbar CLK 0.09276f
C2371 a_98989_13083# a_99603_13083# 0.05935f
C2372 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.04109f
C2373 FFCLR a_132925_27764# 0.045f
C2374 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Nand_Gate_1.Vout 0.04109f
C2375 a_125845_47663# VDD 0.02521f
C2376 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_117609_15797# 0.04995f
C2377 D_FlipFlop_3.3-input-nand_1.B a_134283_40571# 0.04443f
C2378 And_Gate_7.Nand_Gate_0.Vout VDD 1.43162f
C2379 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.04109f
C2380 a_92725_16975# CLK 0.04479f
C2381 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout a_41687_15797# 0.04443f
C2382 FFCLR a_128851_17072# 0.04443f
C2383 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_1.Vout 0.70307f
C2384 a_82057_16975# VDD 0.02521f
C2385 a_73449_15797# EN 0.04443f
C2386 RingCounter_0.D_FlipFlop_6.Qbar VDD 1.93578f
C2387 Nand_Gate_1.A a_104137_16975# 0.0476f
C2388 CDAC8_0.switch_6.Z Nand_Gate_6.B 4.08114f
C2389 CLK Q1 0.1175f
C2390 a_134283_44135# a_134897_44135# 0.05935f
C2391 a_68585_49858# VDD 0.06015f
C2392 D_FlipFlop_1.3-input-nand_0.Vout a_134897_36157# 0.01335f
C2393 a_75551_52572# EN 0.045f
C2394 Nand_Gate_5.B RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.07663f
C2395 a_78881_15797# CLK 0.04619f
C2396 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.07084f
C2397 D_FlipFlop_5.Nand_Gate_1.Vout Q2 0.06993f
C2398 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_2.Vout 0.88509f
C2399 D_FlipFlop_0.CLK D_FlipFlop_3.3-input-nand_0.Vout 0.04612f
C2400 D_FlipFlop_1.Nand_Gate_0.Vout a_128237_36157# 0.04444f
C2401 a_77523_15797# VDD 0.03339f
C2402 CDAC8_0.switch_9.Z Nand_Gate_4.B 1.76363f
C2403 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B EN 0.43216f
C2404 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_0.Vout 1.00694f
C2405 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout CLK 0.03574f
C2406 a_101575_13083# VDD 0.01327f
C2407 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout EN 0.62384f
C2408 a_134897_23350# VDD 0.01186f
C2409 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout EN 0.80245f
C2410 a_110029_15797# VDD 0.03178f
C2411 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout VDD 2.31704f
C2412 FFCLR D_FlipFlop_3.3-input-nand_2.Vout 0.06105f
C2413 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.3-input-nand_2.C 0.26069f
C2414 a_100347_52572# RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.05964f
C2415 a_42431_49858# a_43045_49858# 0.05935f
C2416 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0846f
C2417 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_88563_13083# 0.01335f
C2418 CDAC8_0.switch_7.Z Nand_Gate_1.B 4.80579f
C2419 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout CLK 0.03479f
C2420 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B VDD 1.79521f
C2421 FFCLR D_FlipFlop_1.Nand_Gate_0.Vout 0.65313f
C2422 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B VDD 1.73782f
C2423 And_Gate_4.Nand_Gate_0.Vout a_81685_47663# 0.05964f
C2424 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD 2.04843f
C2425 a_67227_52572# VDD 0.02521f
C2426 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.30154f
C2427 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_73449_15797# 0.04995f
C2428 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_67841_15797# 0.05964f
C2429 a_134897_30478# VDD 0.01186f
C2430 a_128237_36157# Q7 0.06113f
C2431 a_76909_13083# a_77523_13083# 0.05935f
C2432 a_123785_52572# a_124399_52572# 0.05935f
C2433 a_90665_52572# VDD 0.01186f
C2434 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_121069_13083# 0.04444f
C2435 FFCLR a_134897_33443# 0.0607f
C2436 Nand_Gate_6.Vout CLK 2.60891f
C2437 a_128851_33443# VDD 0.01186f
C2438 CDAC8_0.switch_0.Z CLK 0.16657f
C2439 a_75898_25104# VDD 1.30969f
C2440 a_76165_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.05964f
C2441 Nand_Gate_5.A RingCounter_0.D_FlipFlop_6.3-input-nand_1.B 0.29683f
C2442 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.07084f
C2443 FFCLR Q7 0.77041f
C2444 D_FlipFlop_7.3-input-nand_0.Vout VDD 1.77946f
C2445 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.07084f
C2446 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_113359_52572# 0.04444f
C2447 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C CLK 0.30901f
C2448 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout a_45147_49858# 0.04995f
C2449 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C EN 0.07664f
C2450 CDAC8_0.switch_9.Z Q4 0.29232f
C2451 Q1 Q0 0.01156f
C2452 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.16429f
C2453 D_FlipFlop_6.Qbar D_FlipFlop_6.Nand_Gate_1.Vout 0.11654f
C2454 a_39715_15797# a_40329_15797# 0.05935f
C2455 Nand_Gate_4.B a_132925_19786# 0.04741f
C2456 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_101575_13083# 0.01335f
C2457 a_57415_13083# VDD 0.01327f
C2458 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C CLK 0.30966f
C2459 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_96887_13083# 0.05964f
C2460 a_57545_52572# Nand_Gate_3.B 0.01335f
C2461 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_89921_13083# 0.05964f
C2462 a_96887_15797# VDD 0.02906f
C2463 Nand_Gate_7.B And_Gate_0.Nand_Gate_0.Vout 0.04751f
C2464 Nand_Gate_5.Vout a_125845_47663# 0.04443f
C2465 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_84489_13083# 0.04995f
C2466 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_77523_13083# 0.04543f
C2467 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_29289_15797# 0.04995f
C2468 Nand_Gate_5.Vout And_Gate_7.Nand_Gate_0.Vout 0.10129f
C2469 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_72835_13083# 0.04444f
C2470 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121683_15797# 0.01335f
C2471 a_134283_37007# VDD 0.02521f
C2472 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B a_112001_13083# 0.04443f
C2473 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_65869_13083# 0.04444f
C2474 RingCounter_0.D_FlipFlop_15.Qbar a_50755_15797# 0.04443f
C2475 a_128237_46849# VDD 0.02521f
C2476 RingCounter_0.D_FlipFlop_12.Qbar VDD 1.95446f
C2477 D_FlipFlop_5.Qbar D_FlipFlop_5.Nand_Gate_1.Vout 0.11654f
C2478 D_FlipFlop_6.3-input-nand_0.Vout a_134283_23350# 0.05964f
C2479 RingCounter_0.D_FlipFlop_9.Qbar a_105955_13083# 0.06113f
C2480 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.26069f
C2481 D_FlipFlop_0.CLK D_FlipFlop_0.Nand_Gate_1.Vout 0.04199f
C2482 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.08671f
C2483 RingCounter_0.D_FlipFlop_16.Q a_29289_15797# 0.0156f
C2484 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout EN 0.13192f
C2485 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.48398f
C2486 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout EN 0.09065f
C2487 a_54829_13083# a_55443_13083# 0.05935f
C2488 a_91279_49858# VDD 0.02906f
C2489 a_128237_24200# VDD 0.02521f
C2490 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.08671f
C2491 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.07084f
C2492 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_1.Vout 0.08671f
C2493 FFCLR a_134897_46849# 0.04454f
C2494 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.3-input-nand_2.Vout 0.16429f
C2495 Nand_Gate_6.Vout Q0 0.05048f
C2496 m3_125329_49141# VDD 0.10297f
C2497 D_FlipFlop_5.3-input-nand_0.Vout a_134283_26914# 0.05964f
C2498 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout VDD 2.8604f
C2499 CDAC8_0.switch_6.Z CLK 0.21538f
C2500 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_106699_49858# 0.01335f
C2501 a_123041_15797# VDD 0.02734f
C2502 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_41687_13083# 0.05964f
C2503 a_75898_39392# VDD 1.30474f
C2504 Nand_Gate_4.B a_50755_15797# 0.06113f
C2505 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_1.Vout 0.07775f
C2506 a_42431_49858# EN 0.04775f
C2507 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_34721_13083# 0.05964f
C2508 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_29289_13083# 0.04995f
C2509 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout CLK 0.23566f
C2510 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_63153_49858# 0.05964f
C2511 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_54829_13083# 0.05964f
C2512 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_77523_15797# 0.01335f
C2513 D_FlipFlop_4.3-input-nand_0.Vout a_134283_30478# 0.05964f
C2514 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.06935f
C2515 CDAC8_0.switch_8.Z CDAC8_0.switch_7.Z 1.87529f
C2516 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.30154f
C2517 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.26069f
C2518 D_FlipFlop_1.Nand_Gate_0.Vout Q7 0.11443f
C2519 a_86591_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.01335f
C2520 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout EN 0.10495f
C2521 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0846f
C2522 FFCLR Nand_Gate_1.B 0.91553f
C2523 D_FlipFlop_0.Qbar Q4 1.06174f
C2524 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.25963f
C2525 D_FlipFlop_3.Qbar VDD 1.89796f
C2526 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.07084f
C2527 a_117739_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.01335f
C2528 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout 0.01681f
C2529 D_FlipFlop_5.3-input-nand_1.B VDD 1.32727f
C2530 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.0846f
C2531 a_134283_36157# a_134897_36157# 0.05935f
C2532 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout VDD 2.46653f
C2533 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_1.Vout 0.08671f
C2534 a_32749_13083# a_33363_13083# 0.05935f
C2535 a_47119_49858# VDD 0.02906f
C2536 a_34721_15797# VDD 0.03119f
C2537 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout EN 1.03583f
C2538 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110029_13083# 0.04443f
C2539 a_68585_52572# a_69199_52572# 0.05935f
C2540 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout EN 0.06649f
C2541 CDAC8_0.switch_2.Z VDD 1.31298f
C2542 a_83875_13083# VDD 0.02521f
C2543 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_40329_15797# 0.04995f
C2544 D_FlipFlop_3.Qbar D_FlipFlop_3.Nand_Gate_1.Vout 0.11654f
C2545 CDAC8_0.switch_6.Z Q0 0.28955f
C2546 a_119711_52572# VDD 0.01186f
C2547 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B EN 0.43213f
C2548 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout 0.01681f
C2549 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_33363_15797# 0.01335f
C2550 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD 1.86552f
C2551 FFCLR D_FlipFlop_1.Inverter_1.Vout 0.16183f
C2552 a_52113_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.05964f
C2553 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.30154f
C2554 D_FlipFlop_0.Nand_Gate_0.Vout VDD 1.48313f
C2555 a_68585_52572# EN 0.04443f
C2556 D_FlipFlop_0.Inverter_1.Vout a_130209_44135# 0.04995f
C2557 CDAC8_0.switch_5.Z VDD 1.39285f
C2558 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout CLK 0.29759f
C2559 a_118353_49858# CLK 0.04619f
C2560 a_75898_42964# Comparator_0.Vinm 0.0371f
C2561 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_85847_15797# 0.04443f
C2562 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_1.Inverter_1.Vout 0.01422f
C2563 a_117739_49858# VDD 0.01712f
C2564 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.08671f
C2565 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_67227_49858# 0.05964f
C2566 Comparator_0.Vinm Q3 1.64937f
C2567 D_FlipFlop_5.3-input-nand_1.Vout VDD 1.78032f
C2568 Nand_Gate_5.A RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.08377f
C2569 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1541f
C2570 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.Nand_Gate_1.Vout 0.1541f
C2571 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout VDD 2.07863f
C2572 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_1.Vout 0.07758f
C2573 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_2.C 0.14342f
C2574 FFCLR a_134897_20636# 0.04023f
C2575 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout VDD 2.74107f
C2576 a_128851_20636# VDD 0.01186f
C2577 D_FlipFlop_4.Qbar a_128237_30478# 0.04443f
C2578 CDAC8_0.switch_7.Z Nand_Gate_6.B 7.53946f
C2579 D_FlipFlop_7.3-input-nand_2.Vout a_130209_19786# 0.04443f
C2580 D_FlipFlop_2.3-input-nand_1.Vout a_134283_37007# 0.05964f
C2581 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.C 1.09975f
C2582 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_112001_13083# 0.05964f
C2583 FFCLR D_FlipFlop_3.3-input-nand_2.C 0.76213f
C2584 RingCounter_0.D_FlipFlop_17.Qbar FFCLR 1.10693f
C2585 a_39715_13083# VDD 0.02521f
C2586 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout CLK 0.03574f
C2587 CDAC8_0.switch_6.Z Nand_Gate_4.B 3.52726f
C2588 FFCLR D_FlipFlop_5.Inverter_1.Vout 0.56927f
C2589 RingCounter_0.D_FlipFlop_10.Qbar a_116995_13083# 0.06113f
C2590 FFCLR a_134897_27764# 0.04023f
C2591 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout a_111387_52572# 0.04443f
C2592 a_96273_52572# CLK 0.04619f
C2593 FFCLR D_FlipFlop_2.3-input-nand_2.Vout 0.06399f
C2594 a_128851_27764# VDD 0.01186f
C2595 a_95659_52572# VDD 0.0564f
C2596 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout EN 0.62384f
C2597 RingCounter_0.D_FlipFlop_4.Qbar CLK 0.09276f
C2598 Nand_Gate_0.A Q6 1.38518f
C2599 a_114805_16975# CLK 0.06046f
C2600 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout EN 0.61318f
C2601 Nand_Gate_7.B a_67841_15797# 0.04443f
C2602 a_65869_15797# VDD 0.03178f
C2603 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.06955f
C2604 a_104137_16975# VDD 0.02521f
C2605 a_61795_15797# a_62409_15797# 0.05935f
C2606 a_128851_46849# Q4 0.01335f
C2607 RingCounter_0.D_FlipFlop_16.Q Comparator_0.Vinm 0.02272f
C2608 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C CLK 0.30862f
C2609 a_128851_43285# VDD 0.01186f
C2610 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout CLK 0.30735f
C2611 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.16415f
C2612 a_74193_49858# CLK 0.04619f
C2613 a_51369_15797# VDD 0.01571f
C2614 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Qbar 1.05791f
C2615 D_FlipFlop_1.3-input-nand_2.C a_130209_33443# 0.04443f
C2616 FFCLR CDAC8_0.switch_8.Z 2.17565f
C2617 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.08641f
C2618 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.3-input-nand_2.Vout 0.06935f
C2619 a_73579_49858# VDD 0.01712f
C2620 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 1.09975f
C2621 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.04107f
C2622 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout EN 0.78747f
C2623 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.Nand_Gate_1.Vout 0.1541f
C2624 FFCLR D_FlipFlop_0.3-input-nand_0.Vout 0.08617f
C2625 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Qbar 0.07122f
C2626 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_1.B 0.28364f
C2627 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B CLK 0.16274f
C2628 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout CLK 0.29759f
C2629 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_94915_15797# 0.04444f
C2630 a_79495_15797# VDD 0.06072f
C2631 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Inverter_1.Vout 0.25963f
C2632 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout EN 0.78734f
C2633 a_106569_13083# VDD 0.0563f
C2634 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_44403_13083# 0.04543f
C2635 a_89921_15797# a_90535_15797# 0.05935f
C2636 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_88563_15797# 0.04995f
C2637 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B a_101575_13083# 0.04995f
C2638 a_112001_15797# VDD 0.03119f
C2639 a_62539_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.01335f
C2640 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD 1.56255f
C2641 Nand_Gate_0.A Comparator_0.Vinm 4.9842f
C2642 RingCounter_0.D_FlipFlop_1.Qbar a_58159_52572# 0.04443f
C2643 CDAC8_0.switch_6.Z Q4 0.65162f
C2644 a_128237_40571# Q5 0.04443f
C2645 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.04109f
C2646 D_FlipFlop_0.CLK VDD 2.87464f
C2647 Nand_Gate_2.A VDD 7.92635f
C2648 a_124399_52572# Nand_Gate_5.B 0.06113f
C2649 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_123041_13083# 0.05964f
C2650 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_117609_13083# 0.04995f
C2651 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_96887_13083# 0.04443f
C2652 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.09975f
C2653 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.C 1.09975f
C2654 a_132311_33443# VDD 0.02521f
C2655 Nand_Gate_3.B a_63153_52572# 0.04443f
C2656 FFCLR a_128851_44135# 0.04443f
C2657 D_FlipFlop_5.Nand_Gate_1.Vout VDD 1.46545f
C2658 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_87949_13083# 0.04443f
C2659 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.06955f
C2660 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C EN 0.07664f
C2661 a_40459_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.01335f
C2662 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_1.Vout 0.0775f
C2663 a_134897_36157# EN 0.04443f
C2664 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout CLK 0.03574f
C2665 Nand_Gate_5.A a_132925_46849# 0.04685f
C2666 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout VDD 2.16852f
C2667 RingCounter_0.D_FlipFlop_13.Qbar CLK 0.09276f
C2668 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.06955f
C2669 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_65869_15797# 0.04443f
C2670 Nand_Gate_1.B a_128851_30478# 0.04732f
C2671 a_97631_52572# EN 0.045f
C2672 D_FlipFlop_7.3-input-nand_2.Vout a_132311_19786# 0.05964f
C2673 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_1.B 0.28385f
C2674 D_FlipFlop_0.3-input-nand_2.Vout a_132925_46849# 0.01335f
C2675 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout a_85847_15797# 0.04443f
C2676 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout EN 1.03583f
C2677 a_62409_13083# VDD 0.0563f
C2678 And_Gate_0.Nand_Gate_0.Vout VDD 1.38853f
C2679 CDAC8_0.switch_7.Z CLK 5.70593f
C2680 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.30154f
C2681 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_79495_13083# 0.01335f
C2682 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_74807_13083# 0.05964f
C2683 a_75898_35820# VDD 1.30478f
C2684 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_67841_13083# 0.05964f
C2685 FFCLR Nand_Gate_6.B 0.93965f
C2686 D_FlipFlop_0.Inverter_1.Vout VDD 1.73058f
C2687 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_62409_13083# 0.04995f
C2688 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_55443_13083# 0.04543f
C2689 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_50755_13083# 0.04444f
C2690 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B VDD 1.79521f
C2691 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout CLK 0.03479f
C2692 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_87205_52572# 0.04443f
C2693 a_89307_52572# VDD 0.02521f
C2694 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_123785_52572# 0.04995f
C2695 And_Gate_3.Nand_Gate_0.Vout a_114805_16975# 0.05964f
C2696 a_75898_25104# Comparator_0.Vinm 0.03584f
C2697 a_97631_49858# CLK 0.03129f
C2698 FFCLR D_FlipFlop_6.Qbar 0.03748f
C2699 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout EN 0.62384f
C2700 a_96273_49858# VDD 0.0325f
C2701 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout a_100347_52572# 0.04443f
C2702 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_105955_15797# 0.04444f
C2703 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout EN 0.78734f
C2704 a_130209_24200# VDD 0.02521f
C2705 a_112745_52572# VDD 0.01186f
C2706 Nand_Gate_4.A CLK 0.20894f
C2707 And_Gate_1.Nand_Gate_0.Vout VDD 1.39208f
C2708 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout CLK 0.23566f
C2709 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout CLK 0.71245f
C2710 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_98989_15797# 0.05964f
C2711 a_65125_52572# VDD 0.02521f
C2712 EN Q3 0.2481f
C2713 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_108671_49858# 0.04543f
C2714 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B VDD 1.73599f
C2715 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.08671f
C2716 CDAC8_0.switch_8.Z Q7 0.29972f
C2717 Nand_Gate_6.B a_95529_15797# 0.01335f
C2718 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD 2.01968f
C2719 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B a_67841_13083# 0.04443f
C2720 D_FlipFlop_2.Qbar VDD 1.89795f
C2721 a_132311_37007# a_132925_37007# 0.05935f
C2722 RingCounter_0.D_FlipFlop_8.Qbar a_39715_15797# 0.04443f
C2723 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C CLK 0.19377f
C2724 RingCounter_0.D_FlipFlop_2.Qbar RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.11654f
C2725 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_65125_49858# 0.04444f
C2726 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_58159_52572# 0.04444f
C2727 a_75898_39392# Q6 0.5017f
C2728 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout 0.01681f
C2729 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.04109f
C2730 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.16429f
C2731 D_FlipFlop_6.3-input-nand_2.Vout a_132311_20636# 0.04443f
C2732 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.04107f
C2733 Nand_Gate_6.A a_84489_15797# 0.01335f
C2734 CDAC8_0.switch_7.Z Q0 0.57741f
C2735 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout EN 0.09127f
C2736 Nand_Gate_2.Vout VDD 1.37836f
C2737 RingCounter_0.D_FlipFlop_15.Qbar RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.11654f
C2738 D_FlipFlop_0.CLK a_132925_44135# 0.0315f
C2739 D_FlipFlop_3.3-input-nand_2.Vout a_132925_43285# 0.01335f
C2740 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout EN 0.64916f
C2741 RingCounter_0.D_FlipFlop_16.Qbar a_28675_13083# 0.06113f
C2742 D_FlipFlop_2.Qbar a_128237_37007# 0.06113f
C2743 Nand_Gate_7.B Nand_Gate_7.A 0.08001f
C2744 a_42431_52572# a_43045_52572# 0.05935f
C2745 Nand_Gate_5.B Q3 0.06203f
C2746 a_53471_49858# CLK 0.03129f
C2747 a_52113_49858# VDD 0.0325f
C2748 RingCounter_0.D_FlipFlop_16.Q EN 0.26389f
C2749 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.04107f
C2750 a_75898_39392# Comparator_0.Vinm 0.03741f
C2751 D_FlipFlop_5.3-input-nand_2.Vout a_132311_24200# 0.04443f
C2752 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B VDD 1.73782f
C2753 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD 1.99837f
C2754 a_69199_52572# Nand_Gate_0.A 0.06113f
C2755 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_1.B 0.28371f
C2756 D_FlipFlop_0.3-input-nand_0.Vout a_134897_46849# 0.01335f
C2757 a_87949_13083# CLK 0.03129f
C2758 D_FlipFlop_4.Nand_Gate_0.Vout a_128851_30478# 0.04995f
C2759 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_0.Vout 0.0846f
C2760 a_85847_13083# VDD 0.02578f
C2761 RingCounter_0.D_FlipFlop_10.Qbar VDD 1.96961f
C2762 D_FlipFlop_2.3-input-nand_1.B a_134283_37007# 0.04443f
C2763 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.26069f
C2764 a_123041_13083# a_123655_13083# 0.05935f
C2765 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout VDD 2.8604f
C2766 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.06993f
C2767 a_97631_52572# a_98245_52572# 0.05935f
C2768 Nand_Gate_7.A a_57415_15797# 0.04995f
C2769 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_76165_52572# 0.04444f
C2770 a_121069_15797# a_121683_15797# 0.05935f
C2771 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.04107f
C2772 D_FlipFlop_4.3-input-nand_2.Vout a_132311_27764# 0.04443f
C2773 Nand_Gate_1.B a_134897_27764# 0.04544f
C2774 Nand_Gate_0.A EN 0.7382f
C2775 a_134283_40571# a_134897_40571# 0.05935f
C2776 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_112745_49858# 0.04995f
C2777 FFCLR D_FlipFlop_2.3-input-nand_2.C 0.76542f
C2778 RingCounter_0.D_FlipFlop_13.Qbar a_73449_13083# 0.01335f
C2779 a_128851_26914# Q2 0.01335f
C2780 a_120325_49858# CLK 0.02953f
C2781 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout VDD 2.74107f
C2782 D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_1.B 0.68045f
C2783 FFCLR CLK 0.38952f
C2784 a_119711_49858# VDD 0.06071f
C2785 CDAC8_0.switch_7.Z Nand_Gate_4.B 4.09248f
C2786 D_FlipFlop_6.Nand_Gate_0.Vout a_128237_23350# 0.04444f
C2787 a_47119_52572# VDD 0.02521f
C2788 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_69199_49858# 0.04444f
C2789 Nand_Gate_1.A Nand_Gate_1.Vout 0.0689f
C2790 Nand_Gate_3.B a_48937_47663# 0.04443f
C2791 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.30154f
C2792 FFCLR D_FlipFlop_1.3-input-nand_2.Vout 0.88667f
C2793 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.3-input-nand_2.C 0.26069f
C2794 a_134897_19786# VDD 0.01186f
C2795 CDAC8_0.switch_2.Z Comparator_0.Vinm 14.3922f
C2796 VDD Q5 3.80049f
C2797 a_128851_39721# VDD 0.01186f
C2798 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_68585_52572# 0.04995f
C2799 a_132311_20636# VDD 0.02521f
C2800 RingCounter_0.D_FlipFlop_16.Qbar VDD 1.93566f
C2801 D_FlipFlop_0.3-input-nand_0.Vout a_132311_46849# 0.04444f
C2802 a_77523_15797# EN 0.045f
C2803 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout VDD 2.46653f
C2804 Nand_Gate_4.B Nand_Gate_4.A 0.08028f
C2805 a_101575_13083# EN 0.0452f
C2806 D_FlipFlop_5.Nand_Gate_0.Vout a_128237_26914# 0.04444f
C2807 RingCounter_0.D_FlipFlop_8.Qbar RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.07122f
C2808 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.16429f
C2809 a_43789_13083# CLK 0.03129f
C2810 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout a_46505_52572# 0.04995f
C2811 Nand_Gate_1.A a_105955_15797# 0.06113f
C2812 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.06935f
C2813 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.04109f
C2814 Nand_Gate_0.A Nand_Gate_5.B 0.06463f
C2815 Nand_Gate_2.A Nand_Gate_2.B 0.08217f
C2816 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout EN 0.09127f
C2817 a_41687_13083# VDD 0.02578f
C2818 a_76909_15797# a_77523_15797# 0.05935f
C2819 a_94915_15797# VDD 0.02906f
C2820 Nand_Gate_2.A a_93097_47663# 0.04705f
C2821 D_FlipFlop_3.Nand_Gate_1.Vout Q5 0.06993f
C2822 a_100961_13083# a_101575_13083# 0.05935f
C2823 CDAC8_0.switch_5.Z Comparator_0.Vinm 52.8265f
C2824 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B EN 0.43213f
C2825 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout CLK 0.71127f
C2826 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B EN 0.26843f
C2827 a_132311_27764# VDD 0.02521f
C2828 a_134283_23350# a_134897_23350# 0.05935f
C2829 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD 1.86552f
C2830 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout EN 0.97979f
C2831 RingCounter_0.D_FlipFlop_6.Qbar Nand_Gate_5.B 1.06171f
C2832 Nand_Gate_7.B RingCounter_0.D_FlipFlop_14.3-input-nand_1.B 0.2969f
C2833 a_67841_15797# VDD 0.03119f
C2834 Nand_Gate_7.B RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0839f
C2835 a_128237_17072# VDD 0.02521f
C2836 CDAC8_0.switch_7.Z Q4 1.28022f
C2837 a_90665_52572# EN 0.04443f
C2838 Nand_Gate_2.B RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.08524f
C2839 D_FlipFlop_7.3-input-nand_1.B a_134283_17072# 0.04443f
C2840 a_76165_49858# CLK 0.03129f
C2841 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout CLK 0.03479f
C2842 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_54829_15797# 0.04444f
C2843 a_75898_42964# CDAC8_0.switch_9.Z 0.29299f
C2844 D_FlipFlop_1.3-input-nand_2.C a_132925_33443# 0.01335f
C2845 a_75551_49858# VDD 0.06071f
C2846 a_128851_33443# EN 0.05028f
C2847 FFCLR D_FlipFlop_5.3-input-nand_2.Vout 0.06105f
C2848 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.06993f
C2849 D_FlipFlop_7.Qbar a_128237_17072# 0.06113f
C2850 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.25963f
C2851 a_110643_13083# CLK 0.03129f
C2852 a_134283_26914# a_134897_26914# 0.05935f
C2853 CDAC8_0.switch_9.Z Q3 0.36261f
C2854 a_57545_52572# VDD 0.01186f
C2855 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.Vout 0.01194f
C2856 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.C 0.01194f
C2857 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_1.Vout 0.08671f
C2858 a_110029_13083# VDD 0.02578f
C2859 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_46375_13083# 0.01335f
C2860 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_90535_15797# 0.01335f
C2861 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_86591_52572# 0.04995f
C2862 FFCLR a_128851_40571# 0.04443f
C2863 D_FlipFlop_7.3-input-nand_2.C a_132311_19786# 0.04443f
C2864 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B VDD 1.73782f
C2865 a_32749_15797# a_33363_15797# 0.05935f
C2866 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout a_52727_13083# 0.04995f
C2867 a_57415_13083# EN 0.0452f
C2868 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.30154f
C2869 a_134283_30478# a_134897_30478# 0.05935f
C2870 Nand_Gate_1.B Nand_Gate_6.B 0.05373f
C2871 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.3-input-nand_2.Vout 0.16429f
C2872 a_78881_13083# a_79495_13083# 0.05935f
C2873 D_FlipFlop_3.3-input-nand_0.Vout a_132311_43285# 0.04444f
C2874 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_99603_13083# 0.01335f
C2875 a_118353_52572# CLK 0.04619f
C2876 a_134283_33443# VDD 0.02521f
C2877 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.08641f
C2878 a_75898_28676# Q3 0.50347f
C2879 RingCounter_0.D_FlipFlop_7.Qbar CLK 0.09401f
C2880 a_128237_33443# a_128851_33443# 0.05935f
C2881 a_117739_52572# VDD 0.0564f
C2882 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.04107f
C2883 And_Gate_1.Nand_Gate_0.Vout a_48565_16975# 0.05964f
C2884 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout EN 0.61318f
C2885 Nand_Gate_4.A a_37897_16975# 0.0476f
C2886 CLK Q7 0.1175f
C2887 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout a_56187_52572# 0.04443f
C2888 a_73579_52572# a_74193_52572# 0.05935f
C2889 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C VDD 3.56545f
C2890 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C VDD 3.61245f
C2891 D_FlipFlop_0.3-input-nand_1.B D_FlipFlop_0.3-input-nand_1.Vout 0.08641f
C2892 FFCLR Nand_Gate_4.B 0.89748f
C2893 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout EN 0.78747f
C2894 FFCLR a_134897_43285# 0.08436f
C2895 a_66483_13083# CLK 0.03129f
C2896 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_1.B 0.27867f
C2897 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_85847_15797# 0.05964f
C2898 a_65869_13083# VDD 0.02578f
C2899 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.30154f
C2900 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.1182f
C2901 Nand_Gate_2.B Nand_Gate_2.Vout 2.18021f
C2902 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Qbar 0.07122f
C2903 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B a_51499_49858# 0.04995f
C2904 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.04109f
C2905 D_FlipFlop_1.Qbar VDD 1.89794f
C2906 Nand_Gate_2.Vout a_93097_47663# 0.05964f
C2907 Nand_Gate_0.A CDAC8_0.switch_9.Z 0.22762f
C2908 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B CLK 0.16166f
C2909 RingCounter_0.D_FlipFlop_15.Qbar RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.07122f
C2910 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_117739_49858# 0.01335f
C2911 Nand_Gate_2.A Comparator_0.Vinm 4.04825f
C2912 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.08671f
C2913 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout CLK 0.03574f
C2914 D_FlipFlop_6.3-input-nand_2.C a_132311_20636# 0.05964f
C2915 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_57415_13083# 0.01335f
C2916 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1541f
C2917 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_52727_13083# 0.05964f
C2918 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_5.B 0.11443f
C2919 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.06993f
C2920 a_112745_49858# a_113359_49858# 0.05935f
C2921 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.04107f
C2922 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_74193_49858# 0.05964f
C2923 a_128237_23350# VDD 0.02521f
C2924 Nand_Gate_7.B D_FlipFlop_6.Inverter_1.Vout 0.12286f
C2925 a_128237_27764# Q3 0.04443f
C2926 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.25963f
C2927 a_98245_49858# VDD 0.0301f
C2928 a_56801_13083# a_57415_13083# 0.05935f
C2929 a_132925_24200# VDD 0.01186f
C2930 Nand_Gate_5.A VDD 7.74175f
C2931 D_FlipFlop_2.Qbar D_FlipFlop_2.Nand_Gate_1.Vout 0.11654f
C2932 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout VDD 2.88547f
C2933 a_134283_46849# VDD 0.02521f
C2934 Nand_Gate_5.B m3_125329_49141# 0.18891f
C2935 D_FlipFlop_0.Nand_Gate_1.Vout a_128237_44135# 0.04444f
C2936 D_FlipFlop_0.3-input-nand_2.Vout VDD 2.77266f
C2937 D_FlipFlop_5.3-input-nand_2.C a_132311_24200# 0.05964f
C2938 Nand_Gate_0.A a_74193_52572# 0.04443f
C2939 Nand_Gate_5.B a_123041_15797# 0.04443f
C2940 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout EN 0.08852f
C2941 RingCounter_0.D_FlipFlop_2.Qbar Nand_Gate_0.A 1.10693f
C2942 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_42431_49858# 0.01335f
C2943 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.Nand_Gate_1.Vout 0.1541f
C2944 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout a_67227_49858# 0.04995f
C2945 a_132311_19786# a_132925_19786# 0.05935f
C2946 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.1182f
C2947 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_0.Vout 0.07084f
C2948 a_128237_30478# VDD 0.02521f
C2949 Nand_Gate_6.B D_FlipFlop_5.Inverter_1.Vout 0.12143f
C2950 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.06935f
C2951 CDAC8_0.switch_2.Z EN 0.26953f
C2952 a_75898_35820# Comparator_0.Vinm 0.04019f
C2953 Nand_Gate_6.A VDD 4.17892f
C2954 D_FlipFlop_2.Qbar Q6 1.06174f
C2955 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_3.3-input-nand_0.Vout 0.01418f
C2956 a_119711_52572# EN 0.045f
C2957 D_FlipFlop_4.3-input-nand_2.C a_132311_27764# 0.05964f
C2958 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.07084f
C2959 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout EN 1.03583f
C2960 RingCounter_0.D_FlipFlop_2.Qbar a_68585_49858# 0.01335f
C2961 Nand_Gate_1.B CLK 0.67228f
C2962 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_65869_13083# 0.05964f
C2963 CDAC8_0.switch_5.Z EN 1.03162f
C2964 a_122427_52572# RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.05964f
C2965 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C VDD 3.56545f
C2966 Comparator_0.Vinm Vin 0.01779f
C2967 And_Gate_2.Nand_Gate_0.Vout VDD 1.38853f
C2968 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B VDD 1.79529f
C2969 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout CLK 0.03479f
C2970 a_117739_49858# EN 0.07058f
C2971 FFCLR D_FlipFlop_1.3-input-nand_2.C 0.14795f
C2972 a_43045_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.05964f
C2973 a_90665_49858# a_91279_49858# 0.05935f
C2974 Nand_Gate_7.A VDD 4.17892f
C2975 a_111387_52572# VDD 0.02521f
C2976 CDAC8_0.switch_9.Z a_75898_25104# 0.01232f
C2977 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout VDD 2.73822f
C2978 a_34721_13083# a_35335_13083# 0.05935f
C2979 a_54085_49858# VDD 0.0301f
C2980 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.06955f
C2981 D_FlipFlop_0.3-input-nand_2.C a_130209_44135# 0.04443f
C2982 a_89921_13083# CLK 0.04619f
C2983 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.06993f
C2984 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout CLK 0.23566f
C2985 a_88563_13083# VDD 0.05686f
C2986 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout EN 0.13192f
C2987 a_87205_52572# VDD 0.02521f
C2988 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_78267_49858# 0.05964f
C2989 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.08641f
C2990 RingCounter_0.D_FlipFlop_1.Qbar a_58159_49858# 0.06113f
C2991 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.04107f
C2992 a_98245_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.05964f
C2993 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.30154f
C2994 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.09975f
C2995 a_128851_36157# VDD 0.01186f
C2996 Nand_Gate_2.Vout Comparator_0.Vinm 0.04618f
C2997 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.16429f
C2998 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.3-input-nand_2.Vout 0.06935f
C2999 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.08671f
C3000 Nand_Gate_0.A a_69199_49858# 0.04741f
C3001 D_FlipFlop_5.Qbar Q2 1.06526f
C3002 Nand_Gate_5.A Nand_Gate_5.Vout 0.1063f
C3003 a_122427_49858# VDD 0.03726f
C3004 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Inverter_1.Vout 0.25963f
C3005 Nand_Gate_1.Vout VDD 1.40515f
C3006 a_79625_52572# Nand_Gate_0.B 0.01335f
C3007 Nand_Gate_1.B Q0 0.06233f
C3008 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.04109f
C3009 FFCLR D_FlipFlop_5.3-input-nand_2.C 0.76213f
C3010 a_51369_15797# EN 0.04443f
C3011 a_73579_49858# EN 0.07058f
C3012 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout VDD 2.73822f
C3013 RingCounter_0.D_FlipFlop_1.Qbar CLK 0.09276f
C3014 a_68585_49858# a_69199_49858# 0.05935f
C3015 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout Nand_Gate_0.A 0.12214f
C3016 a_134283_20636# VDD 0.02521f
C3017 D_FlipFlop_7.3-input-nand_0.Vout a_132925_19786# 0.04995f
C3018 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Inverter_1.Vout 0.25963f
C3019 RingCounter_0.D_FlipFlop_17.Qbar CLK 0.09276f
C3020 a_56801_15797# CLK 0.04619f
C3021 a_130209_43285# VDD 0.02521f
C3022 a_45761_13083# CLK 0.04619f
C3023 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout FFCLR 0.12214f
C3024 a_105955_15797# VDD 0.02906f
C3025 a_55443_15797# VDD 0.03339f
C3026 CDAC8_0.switch_6.Z Q3 0.78009f
C3027 a_128851_39721# Q6 0.01335f
C3028 a_44403_13083# VDD 0.05686f
C3029 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout VDD 2.31704f
C3030 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.C 1.09975f
C3031 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout EN 0.62384f
C3032 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK 0.29644f
C3033 a_128851_26914# VDD 0.01186f
C3034 FFCLR a_128851_37007# 0.04443f
C3035 a_63153_52572# VDD 0.02521f
C3036 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout VDD 2.73822f
C3037 a_134283_27764# VDD 0.02521f
C3038 And_Gate_6.Nand_Gate_0.Vout CLK 0.50205f
C3039 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_44403_15797# 0.04995f
C3040 Nand_Gate_4.A a_39715_15797# 0.06113f
C3041 Nand_Gate_1.B a_116995_15797# 0.06113f
C3042 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B VDD 1.73782f
C3043 a_110029_15797# a_110643_15797# 0.05935f
C3044 a_130209_17072# VDD 0.02521f
C3045 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD 2.04843f
C3046 Nand_Gate_1.B And_Gate_3.Nand_Gate_0.Vout 0.03063f
C3047 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_62409_15797# 0.04995f
C3048 FFCLR D_FlipFlop_7.3-input-nand_1.Vout 0.95741f
C3049 Nand_Gate_2.A EN 0.6104f
C3050 Nand_Gate_6.Vout a_82057_16975# 0.05964f
C3051 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout CLK 0.28425f
C3052 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_56801_15797# 0.05964f
C3053 CDAC8_0.switch_8.Z CLK 0.35798f
C3054 FFCLR a_132925_36157# 0.0468f
C3055 D_FlipFlop_1.Nand_Gate_1.Vout a_128851_33443# 0.04995f
C3056 a_41073_52572# VDD 0.02865f
C3057 Comparator_0.Vinm Q5 0.78241f
C3058 a_78267_49858# VDD 0.04111f
C3059 D_FlipFlop_7.3-input-nand_1.B D_FlipFlop_7.3-input-nand_1.Vout 0.08641f
C3060 a_75898_46095# VDD 1.30093f
C3061 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout VDD 2.07863f
C3062 Nand_Gate_3.B And_Gate_5.Nand_Gate_0.Vout 0.02391f
C3063 Nand_Gate_1.B Nand_Gate_4.B 0.05965f
C3064 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.26069f
C3065 Nand_Gate_3.B VDD 4.34021f
C3066 a_108671_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.01335f
C3067 a_112001_13083# VDD 0.02865f
C3068 Nand_Gate_0.A a_134897_37007# 0.04682f
C3069 a_67227_52572# RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.05964f
C3070 FFCLR a_51499_52572# 0.04995f
C3071 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0846f
C3072 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_64511_49858# 0.01335f
C3073 FFCLR D_FlipFlop_6.3-input-nand_0.Vout 0.1261f
C3074 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.3-input-nand_2.Vout 0.06935f
C3075 CDAC8_0.switch_9.Z CDAC8_0.switch_2.Z 0.28677f
C3076 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.25963f
C3077 a_46505_49858# a_47119_49858# 0.05935f
C3078 D_FlipFlop_0.Qbar a_128237_46849# 0.04443f
C3079 And_Gate_0.Nand_Gate_0.Vout a_70645_16975# 0.05964f
C3080 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout VDD 2.46653f
C3081 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.08671f
C3082 And_Gate_0.Nand_Gate_0.Vout EN 0.01805f
C3083 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_43789_13083# 0.05964f
C3084 FFCLR a_134897_39721# 0.08436f
C3085 a_90665_52572# a_91279_52572# 0.05935f
C3086 a_75898_21528# CDAC8_0.switch_2.Z 0.29774f
C3087 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C CLK 0.30966f
C3088 RingCounter_0.D_FlipFlop_11.Qbar a_94915_15797# 0.04443f
C3089 Nand_Gate_2.A Nand_Gate_5.B 0.06495f
C3090 a_74807_15797# VDD 0.02906f
C3091 FFCLR D_FlipFlop_4.3-input-nand_0.Vout 0.12261f
C3092 CDAC8_0.switch_9.Z CDAC8_0.switch_5.Z 1.1471f
C3093 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.3-input-nand_2.Vout 0.06935f
C3094 D_FlipFlop_3.3-input-nand_0.Vout a_134283_43285# 0.05964f
C3095 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B a_63153_49858# 0.04443f
C3096 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.08641f
C3097 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B EN 0.43213f
C3098 D_FlipFlop_4.Qbar VDD 1.89806f
C3099 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.04107f
C3100 D_FlipFlop_4.Nand_Gate_1.Vout Q3 0.06993f
C3101 RingCounter_0.D_FlipFlop_14.Qbar VDD 1.95446f
C3102 Nand_Gate_0.A CDAC8_0.switch_6.Z 9.49208f
C3103 D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_7.B 0.67985f
C3104 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD 1.86552f
C3105 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_54085_49858# 0.05964f
C3106 a_128237_44135# VDD 0.02521f
C3107 Nand_Gate_6.B a_94915_13083# 0.04443f
C3108 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.26069f
C3109 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout a_78267_49858# 0.04995f
C3110 a_96273_49858# EN 0.01149f
C3111 a_74193_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.05964f
C3112 a_112745_52572# EN 0.04443f
C3113 a_75898_25104# CDAC8_0.switch_0.Z 0.29672f
C3114 D_FlipFlop_0.3-input-nand_2.C VDD 2.74431f
C3115 And_Gate_1.Nand_Gate_0.Vout EN 0.01805f
C3116 RingCounter_0.D_FlipFlop_14.Qbar RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.11654f
C3117 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout CLK 0.03479f
C3118 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.06955f
C3119 a_56187_52572# VDD 0.02521f
C3120 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.3-input-nand_2.Vout 0.06935f
C3121 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.07084f
C3122 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout a_65125_49858# 0.04443f
C3123 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B EN 0.26841f
C3124 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_98989_13083# 0.04443f
C3125 a_132311_43285# VDD 0.02521f
C3126 Nand_Gate_7.B a_72835_13083# 0.04443f
C3127 a_67841_13083# VDD 0.02865f
C3128 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout EN 0.97916f
C3129 D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_6.B 0.68025f
C3130 a_79625_52572# VDD 0.01186f
C3131 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD 1.56255f
C3132 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.04109f
C3133 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_7.3-input-nand_0.Vout 0.01418f
C3134 D_FlipFlop_2.3-input-nand_2.Vout a_132925_39721# 0.01335f
C3135 RingCounter_0.D_FlipFlop_3.Qbar a_79625_49858# 0.01335f
C3136 D_FlipFlop_7.Inverter_1.Vout a_130209_17072# 0.04995f
C3137 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout CLK 0.23566f
C3138 a_75898_28676# CDAC8_0.switch_5.Z 0.29667f
C3139 Nand_Gate_6.B CLK 0.52757f
C3140 Vin GND 0.55041f
C3141 Q0 GND 16.44317f
C3142 Q1 GND 20.25822f
C3143 Q2 GND 20.04616f
C3144 Q3 GND 19.81573f
C3145 Q7 GND 22.19323f
C3146 Q6 GND 22.18259f
C3147 Q5 GND 22.18194f
C3148 Q4 GND 22.16874f
C3149 CLK GND 0.15559p
C3150 EN GND 0.20021p
C3151 Vbias GND 30.04625f
C3152 VDD GND 2.38329p
C3153 m3_125329_49141# GND 0.68263f $ **FLOATING
C3154 a_123655_13083# GND 0.31947f
C3155 a_123041_13083# GND 0.25914f
C3156 a_121683_13083# GND 0.3185f
C3157 a_121069_13083# GND 0.25914f
C3158 a_118967_13083# GND 0.3185f
C3159 a_117609_13083# GND 0.3185f
C3160 a_116995_13083# GND 0.25913f
C3161 a_112615_13083# GND 0.31947f
C3162 a_112001_13083# GND 0.25914f
C3163 a_110643_13083# GND 0.3185f
C3164 a_110029_13083# GND 0.25914f
C3165 a_107927_13083# GND 0.3185f
C3166 a_106569_13083# GND 0.3185f
C3167 a_105955_13083# GND 0.25913f
C3168 a_101575_13083# GND 0.31947f
C3169 a_100961_13083# GND 0.25914f
C3170 a_99603_13083# GND 0.3185f
C3171 a_98989_13083# GND 0.25914f
C3172 a_96887_13083# GND 0.3185f
C3173 a_95529_13083# GND 0.3185f
C3174 a_94915_13083# GND 0.25913f
C3175 a_90535_13083# GND 0.31947f
C3176 a_89921_13083# GND 0.25914f
C3177 a_88563_13083# GND 0.3185f
C3178 a_87949_13083# GND 0.25914f
C3179 a_85847_13083# GND 0.3185f
C3180 a_84489_13083# GND 0.3185f
C3181 a_83875_13083# GND 0.25913f
C3182 a_79495_13083# GND 0.31947f
C3183 a_78881_13083# GND 0.25914f
C3184 a_77523_13083# GND 0.3185f
C3185 a_76909_13083# GND 0.25914f
C3186 a_74807_13083# GND 0.3185f
C3187 a_73449_13083# GND 0.3185f
C3188 a_72835_13083# GND 0.25913f
C3189 a_68455_13083# GND 0.31947f
C3190 a_67841_13083# GND 0.25914f
C3191 a_66483_13083# GND 0.3185f
C3192 a_65869_13083# GND 0.25914f
C3193 a_63767_13083# GND 0.3185f
C3194 a_62409_13083# GND 0.3185f
C3195 a_61795_13083# GND 0.25913f
C3196 a_57415_13083# GND 0.31947f
C3197 a_56801_13083# GND 0.25914f
C3198 a_55443_13083# GND 0.3185f
C3199 a_54829_13083# GND 0.25914f
C3200 a_52727_13083# GND 0.3185f
C3201 a_51369_13083# GND 0.3185f
C3202 a_50755_13083# GND 0.25913f
C3203 a_46375_13083# GND 0.31947f
C3204 a_45761_13083# GND 0.25914f
C3205 a_44403_13083# GND 0.3185f
C3206 a_43789_13083# GND 0.25914f
C3207 a_41687_13083# GND 0.3185f
C3208 a_40329_13083# GND 0.3185f
C3209 a_39715_13083# GND 0.25913f
C3210 a_35335_13083# GND 0.31947f
C3211 a_34721_13083# GND 0.25914f
C3212 a_33363_13083# GND 0.3185f
C3213 a_32749_13083# GND 0.25914f
C3214 a_30647_13083# GND 0.3185f
C3215 a_29289_13083# GND 0.3185f
C3216 a_28675_13083# GND 0.25913f
C3217 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout GND 1.02192f
C3218 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout GND 1.20008f
C3219 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout GND 1.02192f
C3220 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout GND 1.20008f
C3221 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout GND 1.02192f
C3222 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout GND 1.20008f
C3223 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout GND 1.02192f
C3224 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout GND 1.20008f
C3225 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout GND 1.02192f
C3226 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout GND 1.20008f
C3227 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout GND 1.02192f
C3228 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout GND 1.20008f
C3229 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout GND 1.02192f
C3230 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout GND 1.20008f
C3231 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout GND 1.02192f
C3232 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout GND 1.20008f
C3233 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout GND 1.02192f
C3234 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout GND 1.20008f
C3235 RingCounter_0.D_FlipFlop_10.3-input-nand_1.B GND 1.86871f
C3236 a_123655_15797# GND 0.31947f
C3237 a_123041_15797# GND 0.25914f
C3238 a_121683_15797# GND 0.3185f
C3239 a_121069_15797# GND 0.25913f
C3240 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout GND 1.11634f
C3241 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C GND 1.93731f
C3242 a_118967_15797# GND 0.3185f
C3243 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout GND 2.14781f
C3244 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout GND 2.1681f
C3245 a_117609_15797# GND 0.3185f
C3246 a_116995_15797# GND 0.25913f
C3247 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout GND 1.53057f
C3248 RingCounter_0.D_FlipFlop_10.Qbar GND 1.69483f
C3249 RingCounter_0.D_FlipFlop_9.3-input-nand_1.B GND 1.86853f
C3250 a_112615_15797# GND 0.31947f
C3251 a_112001_15797# GND 0.25914f
C3252 a_110643_15797# GND 0.3185f
C3253 a_110029_15797# GND 0.25913f
C3254 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout GND 1.08165f
C3255 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C GND 1.9378f
C3256 a_107927_15797# GND 0.3185f
C3257 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout GND 2.1482f
C3258 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout GND 2.16859f
C3259 a_106569_15797# GND 0.3185f
C3260 a_105955_15797# GND 0.25913f
C3261 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout GND 1.53106f
C3262 RingCounter_0.D_FlipFlop_9.Qbar GND 1.69532f
C3263 RingCounter_0.D_FlipFlop_11.3-input-nand_1.B GND 1.86853f
C3264 a_101575_15797# GND 0.31947f
C3265 a_100961_15797# GND 0.25914f
C3266 a_99603_15797# GND 0.3185f
C3267 a_98989_15797# GND 0.25913f
C3268 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout GND 1.08165f
C3269 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C GND 1.9378f
C3270 a_96887_15797# GND 0.3185f
C3271 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout GND 2.1482f
C3272 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout GND 2.16859f
C3273 a_95529_15797# GND 0.3185f
C3274 a_94915_15797# GND 0.25913f
C3275 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout GND 1.53106f
C3276 RingCounter_0.D_FlipFlop_11.Qbar GND 1.69532f
C3277 RingCounter_0.D_FlipFlop_12.3-input-nand_1.B GND 1.86853f
C3278 a_90535_15797# GND 0.31947f
C3279 a_89921_15797# GND 0.25914f
C3280 a_88563_15797# GND 0.3185f
C3281 a_87949_15797# GND 0.25913f
C3282 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout GND 1.08165f
C3283 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C GND 1.9378f
C3284 a_85847_15797# GND 0.3185f
C3285 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout GND 2.1482f
C3286 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout GND 2.16859f
C3287 a_84489_15797# GND 0.3185f
C3288 a_83875_15797# GND 0.25913f
C3289 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout GND 1.53106f
C3290 RingCounter_0.D_FlipFlop_12.Qbar GND 1.69532f
C3291 RingCounter_0.D_FlipFlop_13.3-input-nand_1.B GND 1.86853f
C3292 a_79495_15797# GND 0.31947f
C3293 a_78881_15797# GND 0.25914f
C3294 a_77523_15797# GND 0.31884f
C3295 a_76909_15797# GND 0.25913f
C3296 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout GND 1.08171f
C3297 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C GND 1.9378f
C3298 a_74807_15797# GND 0.3185f
C3299 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout GND 2.1482f
C3300 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout GND 2.16859f
C3301 a_73449_15797# GND 0.3185f
C3302 a_72835_15797# GND 0.25913f
C3303 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout GND 1.53106f
C3304 RingCounter_0.D_FlipFlop_13.Qbar GND 1.69532f
C3305 RingCounter_0.D_FlipFlop_14.3-input-nand_1.B GND 1.86853f
C3306 a_68455_15797# GND 0.31947f
C3307 a_67841_15797# GND 0.25914f
C3308 a_66483_15797# GND 0.3185f
C3309 a_65869_15797# GND 0.25913f
C3310 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout GND 1.08165f
C3311 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C GND 1.9378f
C3312 a_63767_15797# GND 0.3185f
C3313 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout GND 2.1482f
C3314 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout GND 2.16859f
C3315 a_62409_15797# GND 0.3185f
C3316 a_61795_15797# GND 0.25913f
C3317 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout GND 1.53106f
C3318 RingCounter_0.D_FlipFlop_14.Qbar GND 1.69532f
C3319 RingCounter_0.D_FlipFlop_15.3-input-nand_1.B GND 1.86853f
C3320 a_57415_15797# GND 0.31947f
C3321 a_56801_15797# GND 0.25914f
C3322 a_55443_15797# GND 0.3185f
C3323 a_54829_15797# GND 0.25913f
C3324 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout GND 1.08165f
C3325 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C GND 1.9378f
C3326 a_52727_15797# GND 0.3185f
C3327 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout GND 2.1482f
C3328 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout GND 2.16859f
C3329 a_51369_15797# GND 0.3185f
C3330 a_50755_15797# GND 0.25913f
C3331 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout GND 1.53106f
C3332 RingCounter_0.D_FlipFlop_15.Qbar GND 1.69532f
C3333 RingCounter_0.D_FlipFlop_8.3-input-nand_1.B GND 1.86853f
C3334 a_46375_15797# GND 0.31947f
C3335 a_45761_15797# GND 0.25914f
C3336 a_44403_15797# GND 0.3185f
C3337 a_43789_15797# GND 0.25913f
C3338 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout GND 1.08165f
C3339 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C GND 1.9378f
C3340 a_41687_15797# GND 0.3185f
C3341 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout GND 2.1482f
C3342 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout GND 2.16859f
C3343 a_40329_15797# GND 0.3185f
C3344 a_39715_15797# GND 0.25913f
C3345 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout GND 1.53106f
C3346 RingCounter_0.D_FlipFlop_8.Qbar GND 1.69532f
C3347 RingCounter_0.D_FlipFlop_16.3-input-nand_1.B GND 1.86853f
C3348 a_35335_15797# GND 0.31947f
C3349 a_34721_15797# GND 0.25914f
C3350 a_33363_15797# GND 0.3185f
C3351 a_32749_15797# GND 0.25913f
C3352 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout GND 1.55623f
C3353 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C GND 1.95415f
C3354 a_30647_15797# GND 0.3185f
C3355 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout GND 2.14783f
C3356 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout GND 2.16819f
C3357 a_29289_15797# GND 0.3185f
C3358 a_28675_15797# GND 0.25913f
C3359 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout GND 1.57941f
C3360 RingCounter_0.D_FlipFlop_16.Qbar GND 1.69505f
C3361 Comparator_0.Vinm GND 0.48681p
C3362 a_134897_17072# GND 0.31947f
C3363 a_134283_17072# GND 0.25914f
C3364 a_132925_17072# GND 0.3185f
C3365 a_132311_17072# GND 0.25914f
C3366 a_130209_17072# GND 0.3185f
C3367 a_128851_17072# GND 0.3185f
C3368 a_128237_17072# GND 0.25913f
C3369 a_114805_16975# GND 0.35808f
C3370 a_104137_16975# GND 0.3185f
C3371 a_92725_16975# GND 0.3185f
C3372 a_82057_16975# GND 0.3185f
C3373 a_70645_16975# GND 0.3185f
C3374 a_59977_16975# GND 0.3185f
C3375 a_48565_16975# GND 0.3185f
C3376 a_37897_16975# GND 0.3185f
C3377 D_FlipFlop_7.3-input-nand_1.Vout GND 1.49356f
C3378 D_FlipFlop_7.Nand_Gate_1.Vout GND 1.60757f
C3379 And_Gate_3.Nand_Gate_0.Vout GND 1.68726f
C3380 Nand_Gate_1.Vout GND 2.2865f
C3381 Nand_Gate_1.A GND 6.41534f
C3382 And_Gate_2.Nand_Gate_0.Vout GND 1.632f
C3383 Nand_Gate_6.Vout GND 2.23235f
C3384 Nand_Gate_6.A GND 6.41534f
C3385 And_Gate_0.Nand_Gate_0.Vout GND 1.69185f
C3386 Nand_Gate_7.A GND 6.45096f
C3387 And_Gate_1.Nand_Gate_0.Vout GND 1.69181f
C3388 Nand_Gate_4.A GND 6.44589f
C3389 D_FlipFlop_7.3-input-nand_1.B GND 1.85534f
C3390 a_134897_19786# GND 0.3185f
C3391 a_134283_19786# GND 0.25914f
C3392 a_132925_19786# GND 0.3185f
C3393 a_132311_19786# GND 0.25913f
C3394 D_FlipFlop_7.3-input-nand_0.Vout GND 1.55899f
C3395 D_FlipFlop_7.3-input-nand_2.C GND 2.11385f
C3396 a_130209_19786# GND 0.3185f
C3397 D_FlipFlop_7.3-input-nand_2.Vout GND 2.16307f
C3398 D_FlipFlop_7.Inverter_1.Vout GND 2.73247f
C3399 a_128851_19786# GND 0.3185f
C3400 a_128237_19786# GND 0.25913f
C3401 Nand_Gate_4.B GND 17.04609f
C3402 D_FlipFlop_7.Nand_Gate_0.Vout GND 1.59582f
C3403 D_FlipFlop_7.Qbar GND 1.67874f
C3404 CDAC8_0.switch_1.Z GND 2.54829f
C3405 a_75898_18814# GND 2.04129f
C3406 a_134897_20636# GND 0.3185f
C3407 a_134283_20636# GND 0.25914f
C3408 a_132925_20636# GND 0.3185f
C3409 a_132311_20636# GND 0.25914f
C3410 a_130209_20636# GND 0.3185f
C3411 a_128851_20636# GND 0.3185f
C3412 a_128237_20636# GND 0.25913f
C3413 D_FlipFlop_6.3-input-nand_1.Vout GND 1.48407f
C3414 D_FlipFlop_6.Nand_Gate_1.Vout GND 1.58498f
C3415 CDAC8_0.switch_2.Z GND 4.74084f
C3416 a_75898_21528# GND 2.05447f
C3417 D_FlipFlop_6.3-input-nand_1.B GND 1.67554f
C3418 a_134897_23350# GND 0.3185f
C3419 a_134283_23350# GND 0.25914f
C3420 a_132925_23350# GND 0.3185f
C3421 a_132311_23350# GND 0.25913f
C3422 D_FlipFlop_6.3-input-nand_0.Vout GND 1.55854f
C3423 D_FlipFlop_6.3-input-nand_2.C GND 2.1043f
C3424 a_130209_23350# GND 0.3185f
C3425 D_FlipFlop_6.3-input-nand_2.Vout GND 2.15354f
C3426 D_FlipFlop_6.Inverter_1.Vout GND 2.71067f
C3427 a_128851_23350# GND 0.3185f
C3428 a_128237_23350# GND 0.25913f
C3429 Nand_Gate_7.B GND 15.4413f
C3430 D_FlipFlop_6.Nand_Gate_0.Vout GND 1.59582f
C3431 D_FlipFlop_6.Qbar GND 1.68185f
C3432 a_134897_24200# GND 0.3185f
C3433 a_134283_24200# GND 0.25914f
C3434 a_132925_24200# GND 0.3185f
C3435 a_132311_24200# GND 0.25914f
C3436 a_130209_24200# GND 0.3185f
C3437 a_128851_24200# GND 0.3185f
C3438 a_128237_24200# GND 0.25913f
C3439 D_FlipFlop_5.3-input-nand_1.Vout GND 1.48407f
C3440 D_FlipFlop_5.Nand_Gate_1.Vout GND 1.58498f
C3441 CDAC8_0.switch_0.Z GND 8.76943f
C3442 a_75898_25104# GND 2.08821f
C3443 D_FlipFlop_5.3-input-nand_1.B GND 1.67554f
C3444 a_134897_26914# GND 0.3185f
C3445 a_134283_26914# GND 0.25914f
C3446 a_132925_26914# GND 0.3185f
C3447 a_132311_26914# GND 0.25913f
C3448 D_FlipFlop_5.3-input-nand_0.Vout GND 1.55854f
C3449 D_FlipFlop_5.3-input-nand_2.C GND 2.1043f
C3450 a_130209_26914# GND 0.3185f
C3451 D_FlipFlop_5.3-input-nand_2.Vout GND 2.15354f
C3452 D_FlipFlop_5.Inverter_1.Vout GND 2.71067f
C3453 a_128851_26914# GND 0.3185f
C3454 a_128237_26914# GND 0.25913f
C3455 Nand_Gate_6.B GND 15.91091f
C3456 D_FlipFlop_5.Nand_Gate_0.Vout GND 1.59582f
C3457 D_FlipFlop_5.Qbar GND 1.68185f
C3458 a_134897_27764# GND 0.3185f
C3459 a_134283_27764# GND 0.25914f
C3460 a_132925_27764# GND 0.3185f
C3461 a_132311_27764# GND 0.25914f
C3462 a_130209_27764# GND 0.3185f
C3463 a_128851_27764# GND 0.3185f
C3464 a_128237_27764# GND 0.25913f
C3465 D_FlipFlop_4.3-input-nand_1.Vout GND 1.48407f
C3466 D_FlipFlop_4.Nand_Gate_1.Vout GND 1.58498f
C3467 CDAC8_0.switch_5.Z GND 16.28138f
C3468 a_75898_28676# GND 2.08822f
C3469 D_FlipFlop_4.3-input-nand_1.B GND 1.67554f
C3470 a_134897_30478# GND 0.3185f
C3471 a_134283_30478# GND 0.25914f
C3472 a_132925_30478# GND 0.3185f
C3473 a_132311_30478# GND 0.25913f
C3474 D_FlipFlop_4.3-input-nand_0.Vout GND 1.63441f
C3475 D_FlipFlop_4.3-input-nand_2.C GND 2.11383f
C3476 a_130209_30478# GND 0.3185f
C3477 D_FlipFlop_4.3-input-nand_2.Vout GND 2.16272f
C3478 D_FlipFlop_4.Inverter_1.Vout GND 2.72021f
C3479 a_128851_30478# GND 0.3185f
C3480 a_128237_30478# GND 0.25913f
C3481 Nand_Gate_1.B GND 17.9523f
C3482 D_FlipFlop_4.Nand_Gate_0.Vout GND 1.61842f
C3483 D_FlipFlop_4.Qbar GND 1.69138f
C3484 a_134897_33443# GND 0.3185f
C3485 a_134283_33443# GND 0.25914f
C3486 a_132925_33443# GND 0.3185f
C3487 a_132311_33443# GND 0.25914f
C3488 a_130209_33443# GND 0.3185f
C3489 a_128851_33443# GND 0.3185f
C3490 a_128237_33443# GND 0.25913f
C3491 D_FlipFlop_1.3-input-nand_1.Vout GND 1.49356f
C3492 D_FlipFlop_1.Nand_Gate_1.Vout GND 1.60757f
C3493 D_FlipFlop_1.3-input-nand_1.B GND 1.68455f
C3494 a_134897_36157# GND 0.3185f
C3495 a_134283_36157# GND 0.25914f
C3496 a_132925_36157# GND 0.3185f
C3497 a_132311_36157# GND 0.25913f
C3498 D_FlipFlop_1.3-input-nand_0.Vout GND 1.56104f
C3499 D_FlipFlop_1.3-input-nand_2.C GND 2.11385f
C3500 a_130209_36157# GND 0.3185f
C3501 D_FlipFlop_1.3-input-nand_2.Vout GND 2.16307f
C3502 D_FlipFlop_1.Inverter_1.Vout GND 2.73247f
C3503 a_128851_36157# GND 0.3185f
C3504 a_128237_36157# GND 0.25913f
C3505 D_FlipFlop_1.Nand_Gate_0.Vout GND 1.59582f
C3506 D_FlipFlop_1.Qbar GND 1.6856f
C3507 CDAC8_0.switch_7.Z GND 0.26711p
C3508 a_75898_35820# GND 2.09412f
C3509 a_134897_37007# GND 0.3185f
C3510 a_134283_37007# GND 0.25914f
C3511 a_132925_37007# GND 0.3185f
C3512 a_132311_37007# GND 0.25914f
C3513 a_130209_37007# GND 0.3185f
C3514 a_128851_37007# GND 0.3185f
C3515 a_128237_37007# GND 0.25913f
C3516 D_FlipFlop_2.3-input-nand_1.Vout GND 1.48407f
C3517 D_FlipFlop_2.Nand_Gate_1.Vout GND 1.58498f
C3518 D_FlipFlop_2.3-input-nand_1.B GND 1.67684f
C3519 a_134897_39721# GND 0.3185f
C3520 a_134283_39721# GND 0.25914f
C3521 a_132925_39721# GND 0.3185f
C3522 a_132311_39721# GND 0.25913f
C3523 D_FlipFlop_2.3-input-nand_0.Vout GND 1.55854f
C3524 D_FlipFlop_2.3-input-nand_2.C GND 2.1043f
C3525 a_130209_39721# GND 0.3185f
C3526 D_FlipFlop_2.3-input-nand_2.Vout GND 2.15354f
C3527 D_FlipFlop_2.Inverter_1.Vout GND 2.71067f
C3528 a_128851_39721# GND 0.3185f
C3529 a_128237_39721# GND 0.25913f
C3530 D_FlipFlop_2.Nand_Gate_0.Vout GND 1.59582f
C3531 D_FlipFlop_2.Qbar GND 1.68185f
C3532 CDAC8_0.switch_6.Z GND 0.12215p
C3533 a_75898_39392# GND 2.09412f
C3534 a_134897_40571# GND 0.3185f
C3535 a_134283_40571# GND 0.25914f
C3536 a_132925_40571# GND 0.3185f
C3537 a_132311_40571# GND 0.25914f
C3538 a_130209_40571# GND 0.3185f
C3539 a_128851_40571# GND 0.3185f
C3540 a_128237_40571# GND 0.25913f
C3541 D_FlipFlop_3.3-input-nand_1.Vout GND 1.48407f
C3542 D_FlipFlop_3.Nand_Gate_1.Vout GND 1.58498f
C3543 D_FlipFlop_3.3-input-nand_1.B GND 1.67684f
C3544 a_134897_43285# GND 0.3185f
C3545 a_134283_43285# GND 0.25914f
C3546 a_132925_43285# GND 0.3185f
C3547 a_132311_43285# GND 0.25913f
C3548 D_FlipFlop_3.3-input-nand_0.Vout GND 1.55854f
C3549 D_FlipFlop_3.3-input-nand_2.C GND 2.1043f
C3550 a_130209_43285# GND 0.3185f
C3551 D_FlipFlop_3.3-input-nand_2.Vout GND 2.15354f
C3552 D_FlipFlop_3.Inverter_1.Vout GND 2.71067f
C3553 a_128851_43285# GND 0.3185f
C3554 a_128237_43285# GND 0.25913f
C3555 D_FlipFlop_3.Nand_Gate_0.Vout GND 1.59582f
C3556 D_FlipFlop_3.Qbar GND 1.68185f
C3557 CDAC8_0.switch_9.Z GND 56.85815f
C3558 a_75898_42964# GND 2.09405f
C3559 a_134897_44135# GND 0.3185f
C3560 a_134283_44135# GND 0.25914f
C3561 a_132925_44135# GND 0.3185f
C3562 a_132311_44135# GND 0.25914f
C3563 a_130209_44135# GND 0.3185f
C3564 a_128851_44135# GND 0.3185f
C3565 a_128237_44135# GND 0.25913f
C3566 D_FlipFlop_0.3-input-nand_1.Vout GND 1.48407f
C3567 D_FlipFlop_0.Nand_Gate_1.Vout GND 1.58498f
C3568 CDAC8_0.switch_8.Z GND 30.02871f
C3569 a_75898_46095# GND 2.08841f
C3570 D_FlipFlop_0.3-input-nand_1.B GND 1.68026f
C3571 a_134897_46849# GND 0.31947f
C3572 a_134283_46849# GND 0.25914f
C3573 a_132925_46849# GND 0.3185f
C3574 a_132311_46849# GND 0.25913f
C3575 D_FlipFlop_0.3-input-nand_0.Vout GND 1.63441f
C3576 D_FlipFlop_0.3-input-nand_2.C GND 2.11383f
C3577 a_130209_46849# GND 0.3185f
C3578 D_FlipFlop_0.3-input-nand_2.Vout GND 2.16272f
C3579 D_FlipFlop_0.Inverter_1.Vout GND 2.72021f
C3580 a_128851_46849# GND 0.3185f
C3581 a_128237_46849# GND 0.25913f
C3582 D_FlipFlop_0.Nand_Gate_0.Vout GND 1.61842f
C3583 D_FlipFlop_0.Qbar GND 1.69138f
C3584 a_125845_47663# GND 0.3185f
C3585 a_115177_47663# GND 0.32117f
C3586 a_103765_47663# GND 0.3185f
C3587 a_93097_47663# GND 0.3185f
C3588 a_81685_47663# GND 0.3185f
C3589 a_71017_47663# GND 0.3185f
C3590 a_59605_47663# GND 0.3185f
C3591 a_48937_47663# GND 0.3185f
C3592 D_FlipFlop_0.CLK GND 5.13796f
C3593 And_Gate_7.Nand_Gate_0.Vout GND 1.71608f
C3594 Nand_Gate_5.Vout GND 2.5275f
C3595 And_Gate_6.Nand_Gate_0.Vout GND 1.6478f
C3596 Nand_Gate_2.Vout GND 2.35535f
C3597 And_Gate_4.Nand_Gate_0.Vout GND 1.6478f
C3598 And_Gate_5.Nand_Gate_0.Vout GND 1.68293f
C3599 a_124399_49858# GND 0.25913f
C3600 a_123785_49858# GND 0.3185f
C3601 a_122427_49858# GND 0.3185f
C3602 a_120325_49858# GND 0.25914f
C3603 a_119711_49858# GND 0.3185f
C3604 a_118353_49858# GND 0.25914f
C3605 a_117739_49858# GND 0.31947f
C3606 a_113359_49858# GND 0.25913f
C3607 a_112745_49858# GND 0.3185f
C3608 a_111387_49858# GND 0.3185f
C3609 a_109285_49858# GND 0.25914f
C3610 a_108671_49858# GND 0.3185f
C3611 a_107313_49858# GND 0.25914f
C3612 a_106699_49858# GND 0.31947f
C3613 a_102319_49858# GND 0.25913f
C3614 a_101705_49858# GND 0.3185f
C3615 a_100347_49858# GND 0.3185f
C3616 a_98245_49858# GND 0.25914f
C3617 a_97631_49858# GND 0.3185f
C3618 a_96273_49858# GND 0.25914f
C3619 a_95659_49858# GND 0.31947f
C3620 a_91279_49858# GND 0.25913f
C3621 a_90665_49858# GND 0.3185f
C3622 a_89307_49858# GND 0.3185f
C3623 a_87205_49858# GND 0.25914f
C3624 a_86591_49858# GND 0.3185f
C3625 a_85233_49858# GND 0.25914f
C3626 a_84619_49858# GND 0.31947f
C3627 a_80239_49858# GND 0.25913f
C3628 a_79625_49858# GND 0.3185f
C3629 a_78267_49858# GND 0.3185f
C3630 a_76165_49858# GND 0.25914f
C3631 a_75551_49858# GND 0.3185f
C3632 a_74193_49858# GND 0.25914f
C3633 a_73579_49858# GND 0.31947f
C3634 a_69199_49858# GND 0.25913f
C3635 a_68585_49858# GND 0.3185f
C3636 a_67227_49858# GND 0.3185f
C3637 a_65125_49858# GND 0.25914f
C3638 a_64511_49858# GND 0.3185f
C3639 a_63153_49858# GND 0.25914f
C3640 a_62539_49858# GND 0.31947f
C3641 a_58159_49858# GND 0.25913f
C3642 a_57545_49858# GND 0.3185f
C3643 a_56187_49858# GND 0.3185f
C3644 a_54085_49858# GND 0.25914f
C3645 a_53471_49858# GND 0.3185f
C3646 a_52113_49858# GND 0.25914f
C3647 a_51499_49858# GND 0.31947f
C3648 a_47119_49858# GND 0.25913f
C3649 a_46505_49858# GND 0.3185f
C3650 a_45147_49858# GND 0.3185f
C3651 a_43045_49858# GND 0.25914f
C3652 a_42431_49858# GND 0.3185f
C3653 a_41073_49858# GND 0.25914f
C3654 a_40459_49858# GND 0.31947f
C3655 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout GND 1.30196f
C3656 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout GND 1.14219f
C3657 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout GND 1.2078f
C3658 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout GND 1.14219f
C3659 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout GND 1.2078f
C3660 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout GND 1.14219f
C3661 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout GND 1.2078f
C3662 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout GND 1.14219f
C3663 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout GND 1.2078f
C3664 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout GND 1.14219f
C3665 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout GND 1.2078f
C3666 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout GND 1.14219f
C3667 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout GND 1.2078f
C3668 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout GND 1.14219f
C3669 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout GND 1.52583f
C3670 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout GND 1.49356f
C3671 Nand_Gate_5.B GND 21.15988f
C3672 a_124399_52572# GND 0.25913f
C3673 a_123785_52572# GND 0.3185f
C3674 RingCounter_0.D_FlipFlop_6.Qbar GND 1.67467f
C3675 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout GND 1.61842f
C3676 a_122427_52572# GND 0.3185f
C3677 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout GND 2.19271f
C3678 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout GND 2.16268f
C3679 a_120325_52572# GND 0.25913f
C3680 a_119711_52572# GND 0.3185f
C3681 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C GND 2.0746f
C3682 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout GND 1.63487f
C3683 a_118353_52572# GND 0.25914f
C3684 a_117739_52572# GND 0.31947f
C3685 RingCounter_0.D_FlipFlop_6.3-input-nand_1.B GND 1.77816f
C3686 Nand_Gate_5.A GND 14.16197f
C3687 a_113359_52572# GND 0.25913f
C3688 a_112745_52572# GND 0.3185f
C3689 RingCounter_0.D_FlipFlop_7.Qbar GND 1.64558f
C3690 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout GND 1.61379f
C3691 a_111387_52572# GND 0.3185f
C3692 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout GND 2.12198f
C3693 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout GND 2.16268f
C3694 a_109285_52572# GND 0.25913f
C3695 a_108671_52572# GND 0.3185f
C3696 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C GND 2.07451f
C3697 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout GND 1.63487f
C3698 a_107313_52572# GND 0.25914f
C3699 a_106699_52572# GND 0.31947f
C3700 RingCounter_0.D_FlipFlop_7.3-input-nand_1.B GND 1.77816f
C3701 Nand_Gate_2.B GND 8.26839f
C3702 a_102319_52572# GND 0.25913f
C3703 a_101705_52572# GND 0.3185f
C3704 RingCounter_0.D_FlipFlop_5.Qbar GND 1.64558f
C3705 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout GND 1.61379f
C3706 a_100347_52572# GND 0.3185f
C3707 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout GND 2.12198f
C3708 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout GND 2.16268f
C3709 a_98245_52572# GND 0.25913f
C3710 a_97631_52572# GND 0.3185f
C3711 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C GND 2.07451f
C3712 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout GND 1.63487f
C3713 a_96273_52572# GND 0.25914f
C3714 a_95659_52572# GND 0.31947f
C3715 RingCounter_0.D_FlipFlop_5.3-input-nand_1.B GND 1.77816f
C3716 Nand_Gate_2.A GND 14.52792f
C3717 a_91279_52572# GND 0.25913f
C3718 a_90665_52572# GND 0.3185f
C3719 RingCounter_0.D_FlipFlop_4.Qbar GND 1.64558f
C3720 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout GND 1.61379f
C3721 a_89307_52572# GND 0.3185f
C3722 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout GND 2.12198f
C3723 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout GND 2.16268f
C3724 a_87205_52572# GND 0.25913f
C3725 a_86591_52572# GND 0.3185f
C3726 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C GND 2.07451f
C3727 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout GND 1.63487f
C3728 a_85233_52572# GND 0.25914f
C3729 a_84619_52572# GND 0.31947f
C3730 RingCounter_0.D_FlipFlop_4.3-input-nand_1.B GND 1.77816f
C3731 Nand_Gate_0.B GND 8.26839f
C3732 a_80239_52572# GND 0.25913f
C3733 a_79625_52572# GND 0.3185f
C3734 RingCounter_0.D_FlipFlop_3.Qbar GND 1.64558f
C3735 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout GND 1.61379f
C3736 a_78267_52572# GND 0.3185f
C3737 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout GND 2.12198f
C3738 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout GND 2.16268f
C3739 a_76165_52572# GND 0.25913f
C3740 a_75551_52572# GND 0.3185f
C3741 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C GND 2.07451f
C3742 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout GND 1.63487f
C3743 a_74193_52572# GND 0.25914f
C3744 a_73579_52572# GND 0.31947f
C3745 RingCounter_0.D_FlipFlop_3.3-input-nand_1.B GND 1.77816f
C3746 Nand_Gate_0.A GND 16.27577f
C3747 a_69199_52572# GND 0.25913f
C3748 a_68585_52572# GND 0.3185f
C3749 RingCounter_0.D_FlipFlop_2.Qbar GND 1.64558f
C3750 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout GND 1.61379f
C3751 a_67227_52572# GND 0.3185f
C3752 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout GND 2.12198f
C3753 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout GND 2.16268f
C3754 a_65125_52572# GND 0.25913f
C3755 a_64511_52572# GND 0.3185f
C3756 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C GND 2.07451f
C3757 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout GND 1.63487f
C3758 a_63153_52572# GND 0.25914f
C3759 a_62539_52572# GND 0.31947f
C3760 RingCounter_0.D_FlipFlop_2.3-input-nand_1.B GND 1.77816f
C3761 Nand_Gate_3.B GND 8.28148f
C3762 a_58159_52572# GND 0.25913f
C3763 a_57545_52572# GND 0.3185f
C3764 RingCounter_0.D_FlipFlop_1.Qbar GND 1.64558f
C3765 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout GND 1.61379f
C3766 a_56187_52572# GND 0.3185f
C3767 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout GND 2.12198f
C3768 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout GND 2.16268f
C3769 a_54085_52572# GND 0.25913f
C3770 a_53471_52572# GND 0.3185f
C3771 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C GND 2.07451f
C3772 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout GND 1.63487f
C3773 a_52113_52572# GND 0.25914f
C3774 a_51499_52572# GND 0.31947f
C3775 RingCounter_0.D_FlipFlop_1.3-input-nand_1.B GND 1.77816f
C3776 FFCLR GND 33.20392f
C3777 a_47119_52572# GND 0.25913f
C3778 a_46505_52572# GND 0.3185f
C3779 RingCounter_0.D_FlipFlop_17.Qbar GND 1.64558f
C3780 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout GND 1.07087f
C3781 a_45147_52572# GND 0.3185f
C3782 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout GND 2.19633f
C3783 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout GND 2.00038f
C3784 a_43045_52572# GND 0.25913f
C3785 a_42431_52572# GND 0.3185f
C3786 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C GND 2.15216f
C3787 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout GND 0.9832f
C3788 a_41073_52572# GND 0.25914f
C3789 a_40459_52572# GND 0.31947f
C3790 RingCounter_0.D_FlipFlop_17.3-input-nand_1.B GND 1.84792f
C3791 RingCounter_0.D_FlipFlop_16.Q GND 24.41932f
C3792 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 GND 0.45666f
C3793 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 GND 0.47347f
C3794 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 GND 0.05122f
C3795 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 GND 0.05958f
C3796 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 GND 0.0577f
C3797 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 GND 0.12257f
C3798 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 GND 0.23742f
C3799 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 GND 0.45664f
C3800 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 GND 0.1334f
C3801 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 GND 0.05705f
C3802 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 GND 0.10533f
C3803 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 GND 0.18236f
C3804 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 GND 0.13574f
C3805 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 GND 0.06431f
C3806 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 GND 0.16533f
C3807 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 GND 0.06323f
C3808 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 GND 0.06194f
C3809 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 GND 0.35224f
C3810 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 GND 0.11629f
C3811 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 GND 0.06194f
C3812 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 GND 0.39067f
C3813 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 GND 0.22727f
C3814 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 GND 0.06839f
C3815 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 GND 0.06358f
C3816 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 GND 0.03611f
C3817 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 GND 0.06992f
C3818 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 GND 0.25335f
C3819 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 GND 0.24817f
C3820 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 GND 0.05234f
C3821 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 GND 0.48726f
C3822 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 GND 0.14234f
C3823 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 GND 0.03542f
C3824 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 GND 0.05152f
C3825 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 GND 0.13202f
C3826 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 GND 0.13202f
C3827 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 GND 0.06862f
C3828 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 GND 0.06624f
C3829 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 GND 0.07883f
C3830 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 GND 0.39844f
C3831 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 GND 0.20187f
C3832 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 GND 0.45666f
C3833 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 GND 0.47347f
C3834 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 GND 0.05122f
C3835 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 GND 0.05958f
C3836 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 GND 0.0577f
C3837 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 GND 0.12257f
C3838 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 GND 0.23742f
C3839 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 GND 0.45664f
C3840 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 GND 0.1334f
C3841 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 GND 0.05705f
C3842 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 GND 0.10533f
C3843 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 GND 0.18236f
C3844 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 GND 0.13574f
C3845 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 GND 0.06431f
C3846 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 GND 0.16533f
C3847 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 GND 0.06323f
C3848 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 GND 0.06194f
C3849 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 GND 0.35224f
C3850 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 GND 0.11629f
C3851 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 GND 0.06194f
C3852 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 GND 0.39067f
C3853 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 GND 0.22727f
C3854 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 GND 0.06839f
C3855 a_139663_37417.t2 GND 0.74021f
C3856 a_139663_37417.t3 GND 2.25506f
C3857 a_139663_37417.t0 GND 2.25426f
C3858 a_139663_37417.n0 GND 1.45916f
C3859 a_139663_37417.n1 GND 0.92425f
C3860 a_139663_37417.t1 GND 1.56705f
C3861 And_Gate_0.B.t2 GND 0.07874f
C3862 Nand_Gate_7.Vout GND -0.158f
C3863 And_Gate_0.B.n0 GND 0.04472f
C3864 And_Gate_0.B.n1 GND 0.0866f
C3865 And_Gate_0.B.t3 GND 0.31378f
C3866 And_Gate_0.Nand_Gate_0.B GND -0.2359f
C3867 And_Gate_0.B.n2 GND 0.30737f
C3868 And_Gate_0.B.n3 GND 0.06483f
C3869 And_Gate_0.B.t4 GND 0.60348f
C3870 And_Gate_0.B.n4 GND 0.17629f
C3871 And_Gate_0.B.n5 GND 0.04387f
C3872 And_Gate_0.B.n6 GND 0.06381f
C3873 And_Gate_0.B.n7 GND 1.30112f
C3874 And_Gate_0.B.n8 GND 1.30112f
C3875 And_Gate_0.B.n9 GND 0.08499f
C3876 And_Gate_0.B.t1 GND 0.08204f
C3877 And_Gate_0.B.t0 GND 0.09763f
C3878 And_Gate_0.B.n10 GND 0.49348f
C3879 And_Gate_0.B.n11 GND 0.25003f
C3880 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 GND 0.05201f
C3881 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 GND 0.22649f
C3882 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 GND 0.05616f
C3883 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 GND 0.39877f
C3884 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 GND 0.39189f
C3885 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 GND 0.04283f
C3886 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 GND 0.20732f
C3887 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 GND 0.05972f
C3888 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 GND 0.02559f
C3889 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 GND 0.04796f
C3890 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 GND 0.10804f
C3891 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 GND 0.10804f
C3892 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 GND 0.06475f
C3893 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 GND 0.05421f
C3894 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 GND 0.05522f
C3895 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 GND 0.05409f
C3896 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 GND 0.30759f
C3897 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 GND 0.17406f
C3898 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 GND 0.03715f
C3899 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 GND 0.07037f
C3900 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 GND 0.16004f
C3901 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 GND 0.07725f
C3902 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 GND 0.2799f
C3903 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 GND 0.27418f
C3904 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 GND 0.05783f
C3905 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 GND 0.53832f
C3906 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 GND 0.15726f
C3907 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 GND 0.03913f
C3908 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 GND 0.05692f
C3909 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 GND 0.14585f
C3910 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 GND 0.14585f
C3911 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 GND 0.07581f
C3912 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 GND 0.07318f
C3913 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 GND 0.07454f
C3914 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 GND 0.07302f
C3915 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 GND 0.41525f
C3916 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 GND 0.23391f
C3917 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 GND 0.22303f
C3918 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 GND 0.05201f
C3919 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 GND 0.22649f
C3920 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 GND 0.05616f
C3921 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 GND 0.39877f
C3922 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 GND 0.39189f
C3923 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 GND 0.04283f
C3924 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 GND 0.20732f
C3925 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 GND 0.05972f
C3926 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 GND 0.02559f
C3927 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 GND 0.04796f
C3928 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 GND 0.10804f
C3929 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 GND 0.10804f
C3930 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 GND 0.06475f
C3931 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 GND 0.05421f
C3932 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 GND 0.05522f
C3933 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 GND 0.05409f
C3934 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 GND 0.30759f
C3935 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 GND 0.17406f
C3936 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 GND 0.03715f
C3937 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 GND 0.07037f
C3938 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 GND 0.16004f
C3939 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 GND 0.07725f
C3940 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 GND 0.2799f
C3941 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 GND 0.27418f
C3942 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 GND 0.05783f
C3943 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 GND 0.53832f
C3944 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 GND 0.15726f
C3945 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 GND 0.03913f
C3946 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 GND 0.05692f
C3947 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 GND 0.14585f
C3948 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 GND 0.14585f
C3949 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 GND 0.07581f
C3950 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 GND 0.07318f
C3951 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 GND 0.07454f
C3952 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 GND 0.07302f
C3953 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 GND 0.41525f
C3954 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 GND 0.23391f
C3955 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 GND 0.22303f
C3956 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 GND 0.07024f
C3957 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 GND 0.03989f
C3958 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 GND 0.07725f
C3959 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 GND 0.2799f
C3960 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 GND 0.27418f
C3961 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 GND 0.05783f
C3962 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 GND 0.53832f
C3963 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 GND 0.15726f
C3964 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 GND 0.03913f
C3965 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 GND 0.05692f
C3966 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 GND 0.14585f
C3967 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 GND 0.14585f
C3968 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 GND 0.07581f
C3969 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 GND 0.07318f
C3970 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 GND 0.07454f
C3971 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 GND 0.07302f
C3972 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 GND 0.41525f
C3973 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 GND 0.23391f
C3974 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 GND 0.22303f
C3975 Nand_Gate_0.B.t11 GND 0.33127f
C3976 Nand_Gate_0.B.n0 GND 0.09677f
C3977 Nand_Gate_0.B.n1 GND 0.04199f
C3978 Nand_Gate_0.B.n2 GND 0.18462f
C3979 Nand_Gate_0.B.t5 GND 0.15408f
C3980 Nand_Gate_0.B.n3 GND 0.04834f
C3981 Nand_Gate_0.B.n4 GND 0.12256f
C3982 Nand_Gate_0.B.t1 GND 0.04493f
C3983 Nand_Gate_0.B.n5 GND 0.06922f
C3984 Nand_Gate_0.B.t3 GND 0.04587f
C3985 Nand_Gate_0.B.t2 GND 0.04493f
C3986 Nand_Gate_0.B.n6 GND 0.25554f
C3987 Nand_Gate_0.B.n7 GND 0.08338f
C3988 Nand_Gate_0.B.n8 GND 0.02717f
C3989 Nand_Gate_0.B.n9 GND 0.05379f
C3990 Nand_Gate_0.B.t9 GND 0.33129f
C3991 Nand_Gate_0.B.n10 GND 0.32557f
C3992 Nand_Gate_0.B.n11 GND 0.03558f
C3993 Nand_Gate_0.B.t10 GND 0.17224f
C3994 Nand_Gate_0.B.n12 GND 0.04961f
C3995 Nand_Gate_0.B.n13 GND 0.02126f
C3996 Nand_Gate_0.B.n14 GND 0.03984f
C3997 Nand_Gate_0.B.n15 GND 0.05014f
C3998 Nand_Gate_0.B.t6 GND 0.33129f
C3999 Nand_Gate_0.B.n16 GND 0.32557f
C4000 Nand_Gate_0.B.n17 GND 0.03558f
C4001 Nand_Gate_0.B.t7 GND 0.17224f
C4002 Nand_Gate_0.B.n18 GND 0.04961f
C4003 Nand_Gate_0.B.n19 GND 0.02126f
C4004 Nand_Gate_0.B.n20 GND 0.03984f
C4005 Nand_Gate_0.B.n22 GND 0.15033f
C4006 Nand_Gate_0.B.n23 GND 0.41862f
C4007 Nand_Gate_0.B.n24 GND 0.18785f
C4008 Nand_Gate_0.B.t4 GND 0.17224f
C4009 Nand_Gate_0.B.t8 GND 0.33127f
C4010 Nand_Gate_0.B.n25 GND 0.09677f
C4011 Nand_Gate_0.B.n26 GND 0.04139f
C4012 Nand_Gate_0.B.n27 GND 0.07641f
C4013 Nand_Gate_0.B.n28 GND 0.87221f
C4014 Nand_Gate_0.B.n29 GND 1.18609f
C4015 Nand_Gate_0.B.n30 GND 0.05328f
C4016 Nand_Gate_0.B.n31 GND 0.01961f
C4017 Nand_Gate_0.B.n33 GND 0.04665f
C4018 Nand_Gate_0.B.t0 GND 0.04321f
C4019 Nand_Gate_0.B.n34 GND 0.18816f
C4020 a_139804_27676.t2 GND 1.19983f
C4021 a_139804_27676.t1 GND 1.19983f
C4022 a_139804_27676.n0 GND 2.49728f
C4023 a_139804_27676.t0 GND 2.30305f
C4024 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 GND 0.0608f
C4025 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 GND 0.13827f
C4026 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 GND 0.06674f
C4027 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 GND 0.24183f
C4028 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 GND 0.23689f
C4029 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 GND 0.04996f
C4030 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 GND 0.46511f
C4031 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 GND 0.13587f
C4032 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 GND 0.03381f
C4033 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 GND 0.04918f
C4034 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 GND 0.12602f
C4035 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 GND 0.12602f
C4036 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 GND 0.0655f
C4037 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 GND 0.06323f
C4038 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 GND 0.07525f
C4039 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 GND 0.38033f
C4040 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 GND 0.1927f
C4041 Q0.t6 GND 0.14104f
C4042 Q0.n0 GND 0.0412f
C4043 Q0.n1 GND 0.01788f
C4044 Q0.n2 GND 0.0786f
C4045 Q0.t9 GND 0.0656f
C4046 Q0.n3 GND 0.0176f
C4047 Q0.n4 GND 0.04807f
C4048 Q0.t2 GND 0.0184f
C4049 Q0.n5 GND 0.09022f
C4050 Q0.n6 GND 0.02214f
C4051 Q0.t1 GND 0.01953f
C4052 Q0.t0 GND 0.01913f
C4053 Q0.n7 GND 0.10879f
C4054 Q0.n8 GND 0.0362f
C4055 Q0.t3 GND 0.01913f
C4056 Q0.n9 GND 0.02645f
C4057 Q0.n10 GND 0.01124f
C4058 Q0.n11 GND 6.2933f
C4059 Q0.t7 GND 0.07345f
C4060 Q0.t8 GND 0.07345f
C4061 Q0.t5 GND 0.14141f
C4062 Q0.n12 GND 0.11441f
C4063 Q0.n13 GND 0.11507f
C4064 Q0.t4 GND 0.12571f
C4065 Q0.n14 GND 1.44692f
C4066 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 GND 0.04607f
C4067 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 GND 0.10477f
C4068 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 GND 0.05057f
C4069 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 GND 0.35243f
C4070 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 GND 0.3654f
C4071 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 GND 0.03953f
C4072 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 GND 0.05278f
C4073 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 GND 0.27708f
C4074 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 GND 0.27709f
C4075 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 GND 0.17949f
C4076 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 GND 0.03786f
C4077 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 GND 0.35241f
C4078 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 GND 0.10295f
C4079 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 GND 0.02562f
C4080 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 GND 0.03726f
C4081 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 GND 0.09548f
C4082 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 GND 0.09548f
C4083 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 GND 0.04963f
C4084 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 GND 0.04792f
C4085 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 GND 0.28399f
C4086 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 GND 0.04998f
C4087 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 GND 0.02839f
C4088 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 GND 0.05497f
C4089 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 GND 0.38308f
C4090 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 GND 0.39717f
C4091 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 GND 0.04297f
C4092 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 GND 0.05737f
C4093 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 GND 0.30118f
C4094 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 GND 0.30119f
C4095 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 GND 0.1951f
C4096 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 GND 0.04115f
C4097 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 GND 0.38306f
C4098 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 GND 0.1119f
C4099 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 GND 0.02784f
C4100 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 GND 0.0405f
C4101 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 GND 0.10379f
C4102 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 GND 0.10379f
C4103 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 GND 0.05395f
C4104 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 GND 0.05208f
C4105 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 GND 0.30868f
C4106 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 GND 0.36784f
C4107 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 GND 0.10746f
C4108 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 GND 0.04662f
C4109 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 GND 0.04798f
C4110 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 GND 0.22815f
C4111 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 GND 0.0518f
C4112 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 GND 0.36785f
C4113 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 GND 0.38072f
C4114 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 GND 0.19125f
C4115 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 GND 0.18752f
C4116 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 GND 0.10934f
C4117 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 GND 0.01378f
C4118 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 GND 0.01095f
C4119 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 GND 0.05094f
C4120 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 GND 0.04989f
C4121 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 GND 0.28374f
C4122 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 GND 0.09258f
C4123 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 GND 0.04989f
C4124 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 GND 0.31407f
C4125 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 GND 0.1838f
C4126 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 GND 0.205f
C4127 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 GND 0.36784f
C4128 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 GND 0.10746f
C4129 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 GND 0.04662f
C4130 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 GND 0.04798f
C4131 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 GND 0.22815f
C4132 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 GND 0.0518f
C4133 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 GND 0.36785f
C4134 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 GND 0.38072f
C4135 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 GND 0.19125f
C4136 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 GND 0.18752f
C4137 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 GND 0.10934f
C4138 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 GND 0.01378f
C4139 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 GND 0.01506f
C4140 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 GND 0.05094f
C4141 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 GND 0.04989f
C4142 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 GND 0.28374f
C4143 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 GND 0.09441f
C4144 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 GND 0.04989f
C4145 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 GND 0.31407f
C4146 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 GND 0.1838f
C4147 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 GND 0.205f
C4148 Nand_Gate_6.Vout.t1 GND 0.07874f
C4149 Nand_Gate_6.Vout.n0 GND 0.04472f
C4150 Nand_Gate_6.Vout.n1 GND 0.0866f
C4151 Nand_Gate_6.Vout.t3 GND 0.31378f
C4152 Nand_Gate_6.Vout.n2 GND 0.30737f
C4153 Nand_Gate_6.Vout.n3 GND 0.06483f
C4154 Nand_Gate_6.Vout.t4 GND 0.60348f
C4155 Nand_Gate_6.Vout.n4 GND 0.17629f
C4156 Nand_Gate_6.Vout.n5 GND 0.04387f
C4157 Nand_Gate_6.Vout.n6 GND 0.06381f
C4158 Nand_Gate_6.Vout.n7 GND 1.30112f
C4159 Nand_Gate_6.Vout.n8 GND 1.30112f
C4160 Nand_Gate_6.Vout.n9 GND 0.08499f
C4161 Nand_Gate_6.Vout.t2 GND 0.08204f
C4162 Nand_Gate_6.Vout.t0 GND 0.09763f
C4163 Nand_Gate_6.Vout.n10 GND 0.49348f
C4164 Nand_Gate_6.Vout.n11 GND 0.25003f
C4165 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 GND 0.36784f
C4166 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 GND 0.10746f
C4167 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 GND 0.04662f
C4168 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 GND 0.04798f
C4169 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 GND 0.22815f
C4170 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 GND 0.0518f
C4171 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 GND 0.36785f
C4172 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 GND 0.38072f
C4173 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 GND 0.19125f
C4174 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 GND 0.18752f
C4175 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 GND 0.10934f
C4176 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 GND 0.01378f
C4177 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 GND 0.01506f
C4178 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 GND 0.05094f
C4179 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 GND 0.04989f
C4180 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 GND 0.28374f
C4181 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 GND 0.09441f
C4182 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 GND 0.04989f
C4183 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 GND 0.31407f
C4184 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 GND 0.1838f
C4185 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 GND 0.205f
C4186 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 GND 0.36784f
C4187 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 GND 0.10746f
C4188 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 GND 0.04662f
C4189 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 GND 0.04798f
C4190 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 GND 0.22815f
C4191 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 GND 0.0518f
C4192 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 GND 0.36785f
C4193 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 GND 0.38072f
C4194 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 GND 0.19125f
C4195 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 GND 0.18752f
C4196 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 GND 0.10934f
C4197 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 GND 0.01378f
C4198 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 GND 0.01506f
C4199 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 GND 0.05094f
C4200 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 GND 0.04989f
C4201 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 GND 0.28374f
C4202 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 GND 0.09441f
C4203 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 GND 0.04989f
C4204 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 GND 0.31407f
C4205 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 GND 0.1838f
C4206 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 GND 0.205f
C4207 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 GND 0.04607f
C4208 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 GND 0.10477f
C4209 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 GND 0.05057f
C4210 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 GND 0.35243f
C4211 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 GND 0.3654f
C4212 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 GND 0.03953f
C4213 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 GND 0.05278f
C4214 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 GND 0.27708f
C4215 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 GND 0.27709f
C4216 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 GND 0.17949f
C4217 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 GND 0.03786f
C4218 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 GND 0.35241f
C4219 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 GND 0.10295f
C4220 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 GND 0.02562f
C4221 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 GND 0.03726f
C4222 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 GND 0.09548f
C4223 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 GND 0.09548f
C4224 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 GND 0.04963f
C4225 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 GND 0.04792f
C4226 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 GND 0.28399f
C4227 D_FlipFlop_6.3-input-nand_2.Vout.t5 GND 0.35515f
C4228 D_FlipFlop_6.3-input-nand_2.Vout.n0 GND 0.10375f
C4229 D_FlipFlop_6.3-input-nand_2.Vout.n1 GND 0.04502f
C4230 D_FlipFlop_6.3-input-nand_2.Vout.n2 GND 0.19793f
C4231 D_FlipFlop_6.3-input-nand_2.Vout.t7 GND 0.17747f
C4232 D_FlipFlop_6.3-input-nand_2.Vout.t1 GND 0.04817f
C4233 D_FlipFlop_6.3-input-nand_2.Vout.n3 GND 0.30324f
C4234 D_FlipFlop_6.3-input-nand_2.Vout.t3 GND 0.04918f
C4235 D_FlipFlop_6.3-input-nand_2.Vout.t2 GND 0.04817f
C4236 D_FlipFlop_6.3-input-nand_2.Vout.n4 GND 0.27396f
C4237 D_FlipFlop_6.3-input-nand_2.Vout.n5 GND 0.09115f
C4238 D_FlipFlop_6.3-input-nand_2.Vout.n6 GND 0.01454f
C4239 D_FlipFlop_6.3-input-nand_2.Vout.n7 GND 0.01331f
C4240 D_FlipFlop_6.3-input-nand_2.Vout.t4 GND 0.35517f
C4241 D_FlipFlop_6.3-input-nand_2.Vout.n8 GND 0.36759f
C4242 D_FlipFlop_6.3-input-nand_2.Vout.t6 GND 0.18465f
C4243 D_FlipFlop_6.3-input-nand_2.Vout.n9 GND 0.18106f
C4244 D_FlipFlop_6.3-input-nand_2.Vout.n10 GND 0.10557f
C4245 D_FlipFlop_6.3-input-nand_2.Vout.n11 GND 0.05002f
C4246 D_FlipFlop_6.3-input-nand_2.Vout.t0 GND 0.04632f
C4247 D_FlipFlop_6.3-input-nand_2.Vout.n12 GND 0.22028f
C4248 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 GND 0.06069f
C4249 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 GND 0.03447f
C4250 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 GND 0.06674f
C4251 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 GND 0.24183f
C4252 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 GND 0.23689f
C4253 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 GND 0.04996f
C4254 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 GND 0.46511f
C4255 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 GND 0.13587f
C4256 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 GND 0.03381f
C4257 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 GND 0.04918f
C4258 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 GND 0.12602f
C4259 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 GND 0.12602f
C4260 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 GND 0.0655f
C4261 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 GND 0.06323f
C4262 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 GND 0.07525f
C4263 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 GND 0.38033f
C4264 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 GND 0.1927f
C4265 D_FlipFlop_2.3-input-nand_2.Vout.t5 GND 0.35515f
C4266 D_FlipFlop_2.3-input-nand_2.Vout.n0 GND 0.10375f
C4267 D_FlipFlop_2.3-input-nand_2.Vout.n1 GND 0.04502f
C4268 D_FlipFlop_2.3-input-nand_2.Vout.n2 GND 0.19793f
C4269 D_FlipFlop_2.3-input-nand_2.Vout.t7 GND 0.17747f
C4270 D_FlipFlop_2.3-input-nand_2.Vout.t1 GND 0.04817f
C4271 D_FlipFlop_2.3-input-nand_2.Vout.n3 GND 0.30324f
C4272 D_FlipFlop_2.3-input-nand_2.Vout.t2 GND 0.04918f
C4273 D_FlipFlop_2.3-input-nand_2.Vout.t3 GND 0.04817f
C4274 D_FlipFlop_2.3-input-nand_2.Vout.n4 GND 0.27396f
C4275 D_FlipFlop_2.3-input-nand_2.Vout.n5 GND 0.09115f
C4276 D_FlipFlop_2.3-input-nand_2.Vout.n6 GND 0.01454f
C4277 D_FlipFlop_2.3-input-nand_2.Vout.n7 GND 0.01331f
C4278 D_FlipFlop_2.3-input-nand_2.Vout.t4 GND 0.35517f
C4279 D_FlipFlop_2.3-input-nand_2.Vout.n8 GND 0.36759f
C4280 D_FlipFlop_2.3-input-nand_2.Vout.t6 GND 0.18465f
C4281 D_FlipFlop_2.3-input-nand_2.Vout.n9 GND 0.18106f
C4282 D_FlipFlop_2.3-input-nand_2.Vout.n10 GND 0.10557f
C4283 D_FlipFlop_2.3-input-nand_2.Vout.n11 GND 0.05002f
C4284 D_FlipFlop_2.3-input-nand_2.Vout.t0 GND 0.04632f
C4285 D_FlipFlop_2.3-input-nand_2.Vout.n12 GND 0.22028f
C4286 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 GND 0.06358f
C4287 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 GND 0.03611f
C4288 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 GND 0.06992f
C4289 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 GND 0.25335f
C4290 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 GND 0.24817f
C4291 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 GND 0.05234f
C4292 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 GND 0.48726f
C4293 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 GND 0.14234f
C4294 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 GND 0.03542f
C4295 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 GND 0.05152f
C4296 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 GND 0.13202f
C4297 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 GND 0.13202f
C4298 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 GND 0.06862f
C4299 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 GND 0.06624f
C4300 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 GND 0.07883f
C4301 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 GND 0.39844f
C4302 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 GND 0.20187f
C4303 And_Gate_1.B.t1 GND 0.03938f
C4304 And_Gate_1.B.t2 GND 0.04686f
C4305 And_Gate_1.B.n0 GND 0.23687f
C4306 Nand_Gate_4.Vout GND -0.07584f
C4307 And_Gate_1.B.n1 GND 0.12001f
C4308 And_Gate_1.B.n2 GND 0.04079f
C4309 And_Gate_1.B.t3 GND 0.15061f
C4310 And_Gate_1.Nand_Gate_0.B GND -0.11323f
C4311 And_Gate_1.B.n3 GND 0.14754f
C4312 And_Gate_1.B.n4 GND 0.03112f
C4313 And_Gate_1.B.t4 GND 0.28967f
C4314 And_Gate_1.B.n5 GND 0.08462f
C4315 And_Gate_1.B.n6 GND 0.02106f
C4316 And_Gate_1.B.n7 GND 0.03063f
C4317 And_Gate_1.B.n8 GND 0.62454f
C4318 And_Gate_1.B.n9 GND 0.62454f
C4319 And_Gate_1.B.n10 GND 0.04157f
C4320 And_Gate_1.B.n11 GND 0.02147f
C4321 And_Gate_1.B.t0 GND 0.0378f
C4322 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 GND 0.05803f
C4323 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 GND 0.15518f
C4324 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 GND 0.11917f
C4325 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 GND 0.23082f
C4326 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 GND 0.44396f
C4327 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 GND 0.12969f
C4328 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 GND 0.05546f
C4329 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 GND 0.1024f
C4330 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 GND 0.1773f
C4331 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 GND 0.13197f
C4332 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 GND 0.06252f
C4333 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 GND 0.44398f
C4334 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 GND 0.46032f
C4335 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 GND 0.0498f
C4336 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 GND 0.06649f
C4337 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 GND 0.22095f
C4338 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 GND 0.06022f
C4339 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 GND 0.37982f
C4340 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 GND 0.06148f
C4341 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 GND 0.06022f
C4342 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 GND 0.34246f
C4343 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 GND 0.11306f
C4344 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 GND 0.16074f
C4345 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 GND 0.36784f
C4346 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 GND 0.10746f
C4347 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 GND 0.04662f
C4348 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 GND 0.04798f
C4349 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 GND 0.22815f
C4350 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 GND 0.0518f
C4351 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 GND 0.36785f
C4352 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 GND 0.38072f
C4353 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 GND 0.19125f
C4354 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 GND 0.18752f
C4355 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 GND 0.10934f
C4356 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 GND 0.01378f
C4357 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 GND 0.01095f
C4358 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 GND 0.05094f
C4359 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 GND 0.04989f
C4360 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 GND 0.28374f
C4361 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 GND 0.09258f
C4362 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 GND 0.04989f
C4363 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 GND 0.31407f
C4364 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 GND 0.1838f
C4365 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 GND 0.205f
C4366 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 GND 0.04607f
C4367 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 GND 0.10477f
C4368 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 GND 0.05057f
C4369 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 GND 0.35243f
C4370 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 GND 0.3654f
C4371 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 GND 0.03953f
C4372 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 GND 0.05278f
C4373 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 GND 0.27708f
C4374 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 GND 0.27709f
C4375 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 GND 0.17949f
C4376 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 GND 0.03786f
C4377 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 GND 0.35241f
C4378 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 GND 0.10295f
C4379 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 GND 0.02562f
C4380 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 GND 0.03726f
C4381 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 GND 0.09548f
C4382 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 GND 0.09548f
C4383 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 GND 0.04963f
C4384 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 GND 0.04792f
C4385 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 GND 0.28399f
C4386 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 GND 0.06323f
C4387 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 GND 0.07525f
C4388 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 GND 0.38033f
C4389 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 GND 0.1927f
C4390 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 GND 0.0655f
C4391 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 GND 0.24183f
C4392 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 GND 0.23689f
C4393 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 GND 0.04996f
C4394 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 GND 0.46511f
C4395 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 GND 0.13587f
C4396 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 GND 0.03381f
C4397 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 GND 0.04918f
C4398 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 GND 0.12602f
C4399 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 GND 0.12602f
C4400 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 GND 0.06674f
C4401 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 GND 0.0608f
C4402 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 GND 0.13827f
C4403 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 GND 0.05969f
C4404 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 GND 0.15961f
C4405 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 GND 0.12257f
C4406 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 GND 0.23742f
C4407 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 GND 0.45664f
C4408 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 GND 0.1334f
C4409 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 GND 0.05705f
C4410 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 GND 0.10533f
C4411 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 GND 0.18236f
C4412 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 GND 0.13574f
C4413 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 GND 0.06431f
C4414 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 GND 0.45666f
C4415 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 GND 0.47347f
C4416 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 GND 0.05122f
C4417 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 GND 0.06839f
C4418 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 GND 0.22727f
C4419 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 GND 0.06194f
C4420 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 GND 0.39067f
C4421 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 GND 0.06323f
C4422 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 GND 0.06194f
C4423 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 GND 0.35224f
C4424 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 GND 0.11629f
C4425 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 GND 0.16533f
C4426 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 GND 0.07037f
C4427 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 GND 0.16004f
C4428 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 GND 0.07725f
C4429 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 GND 0.2799f
C4430 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 GND 0.27418f
C4431 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 GND 0.05783f
C4432 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 GND 0.53832f
C4433 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 GND 0.15726f
C4434 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 GND 0.03913f
C4435 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 GND 0.05692f
C4436 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 GND 0.14585f
C4437 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 GND 0.14585f
C4438 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 GND 0.07581f
C4439 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 GND 0.07318f
C4440 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 GND 0.07454f
C4441 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 GND 0.07302f
C4442 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 GND 0.41525f
C4443 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 GND 0.23391f
C4444 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 GND 0.22303f
C4445 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 GND 0.07024f
C4446 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 GND 0.03989f
C4447 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 GND 0.07725f
C4448 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 GND 0.2799f
C4449 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 GND 0.27418f
C4450 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 GND 0.05783f
C4451 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 GND 0.53832f
C4452 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 GND 0.15726f
C4453 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 GND 0.03913f
C4454 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 GND 0.05692f
C4455 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 GND 0.14585f
C4456 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 GND 0.14585f
C4457 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 GND 0.07581f
C4458 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 GND 0.07318f
C4459 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 GND 0.07454f
C4460 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 GND 0.07302f
C4461 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 GND 0.41525f
C4462 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 GND 0.23391f
C4463 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 GND 0.22303f
C4464 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 GND 0.45666f
C4465 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 GND 0.47347f
C4466 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 GND 0.05122f
C4467 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 GND 0.05969f
C4468 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 GND 0.15961f
C4469 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 GND 0.12257f
C4470 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 GND 0.23742f
C4471 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 GND 0.45664f
C4472 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 GND 0.1334f
C4473 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 GND 0.05705f
C4474 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 GND 0.10533f
C4475 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 GND 0.18236f
C4476 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 GND 0.13574f
C4477 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 GND 0.06431f
C4478 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 GND 0.16533f
C4479 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 GND 0.06323f
C4480 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 GND 0.06194f
C4481 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 GND 0.35224f
C4482 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 GND 0.11629f
C4483 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 GND 0.06194f
C4484 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 GND 0.39067f
C4485 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 GND 0.22727f
C4486 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 GND 0.06839f
C4487 Vbias.t6 GND 1.28887f
C4488 Vbias.n0 GND 0.48561f
C4489 Vbias.t0 GND 4.62462f
C4490 Vbias.t4 GND 1.27672f
C4491 Vbias.n1 GND 0.43915f
C4492 Vbias.t8 GND 0.5558f
C4493 Vbias.n2 GND 0.39434f
C4494 Vbias.n3 GND 1.06417f
C4495 Vbias.n4 GND 0.17495f
C4496 Vbias.n5 GND 0.20178f
C4497 Vbias.n6 GND 0.23277f
C4498 Vbias.n7 GND 0.2392f
C4499 Vbias.n8 GND 0.4184f
C4500 Vbias.n9 GND 0.4184f
C4501 Vbias.n10 GND 6.1943f
C4502 Vbias.n11 GND 0.33996f
C4503 Vbias.n12 GND 0.33996f
C4504 Vbias.n13 GND 0.19841f
C4505 Vbias.t5 GND 6.31206f
C4506 Vbias.t9 GND 2.77919f
C4507 Vbias.n14 GND 0.42621f
C4508 Vbias.n15 GND 0.42621f
C4509 Vbias.n16 GND 0.29344f
C4510 Vbias.n17 GND 53.2923f
C4511 Vbias.n18 GND 38.8878f
C4512 Vbias.n19 GND 1.636f
C4513 Vbias.n20 GND 1.636f
C4514 Vbias.t2 GND 16.0547f
C4515 Vbias.n22 GND 22.7341f
C4516 Vbias.n23 GND 1.6091f
C4517 Vbias.n24 GND 2.43126f
C4518 Vbias.n25 GND 1.6091f
C4519 Vbias.n26 GND 1.63286f
C4520 Vbias.n27 GND 41.1226f
C4521 Vbias.n28 GND 31.4425f
C4522 Vbias.n29 GND 0.4184f
C4523 Vbias.n30 GND 0.2392f
C4524 Vbias.n31 GND 0.2489f
C4525 Vbias.n32 GND 0.23277f
C4526 Vbias.n33 GND 0.4184f
C4527 Vbias.n34 GND 6.1943f
C4528 Vbias.n35 GND 6.1943f
C4529 Vbias.n36 GND 0.3327f
C4530 Vbias.n37 GND 0.19591f
C4531 Vbias.n38 GND 0.19841f
C4532 Vbias.n39 GND 0.19591f
C4533 Vbias.n40 GND 0.3327f
C4534 Vbias.n41 GND 6.1943f
C4535 Vbias.n42 GND 6.1943f
C4536 Vbias.n43 GND 0.33996f
C4537 Vbias.n44 GND 0.33996f
C4538 Vbias.n45 GND 0.19841f
C4539 Vbias.t1 GND 6.31206f
C4540 Vbias.t7 GND 19.89f
C4541 Vbias.n46 GND 0.2535f
C4542 Vbias.n47 GND 0.2535f
C4543 Vbias.n48 GND 0.14785f
C4544 Vbias.n50 GND 31.0657f
C4545 Vbias.n51 GND 0.13915f
C4546 Vbias.n52 GND 0.37755f
C4547 Vbias.n53 GND 0.13915f
C4548 Vbias.n54 GND 0.24721f
C4549 Vbias.n55 GND 20.1609f
C4550 Vbias.n56 GND 20.1609f
C4551 Vbias.n57 GND 0.3327f
C4552 Vbias.n58 GND 0.19591f
C4553 Vbias.n59 GND 0.19841f
C4554 Vbias.n60 GND 0.19591f
C4555 Vbias.n61 GND 0.3327f
C4556 Vbias.n62 GND 6.1943f
C4557 Vbias.n63 GND 0.2489f
C4558 Vbias.n64 GND 0.42621f
C4559 Vbias.t3 GND 2.77919f
C4560 Vbias.n65 GND 0.42621f
C4561 Vbias.n66 GND 0.29344f
C4562 Vbias.n67 GND 0.20178f
C4563 Vbias.n68 GND 0.03376f
C4564 Vbias.n69 GND 0.1106f
C4565 a_138485_16882.t2 GND 0.70901f
C4566 a_138485_16882.t3 GND 0.66541f
C4567 a_138485_16882.t4 GND 1.2388f
C4568 a_138485_16882.n0 GND 0.6901f
C4569 a_138485_16882.t1 GND 1.2388f
C4570 a_138485_16882.n1 GND 0.3967f
C4571 a_138485_16882.n2 GND 0.44526f
C4572 a_138485_16882.t0 GND 2.81593f
C4573 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 GND 0.04998f
C4574 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 GND 0.02839f
C4575 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 GND 0.05497f
C4576 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 GND 0.38308f
C4577 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 GND 0.39717f
C4578 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 GND 0.04297f
C4579 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 GND 0.05737f
C4580 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 GND 0.30118f
C4581 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 GND 0.30119f
C4582 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 GND 0.1951f
C4583 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 GND 0.04115f
C4584 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 GND 0.38306f
C4585 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 GND 0.1119f
C4586 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 GND 0.02784f
C4587 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 GND 0.0405f
C4588 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 GND 0.10379f
C4589 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 GND 0.10379f
C4590 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 GND 0.05395f
C4591 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 GND 0.05208f
C4592 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 GND 0.30868f
C4593 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 GND 0.06067f
C4594 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 GND 0.26418f
C4595 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 GND 0.0655f
C4596 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 GND 0.46513f
C4597 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 GND 0.4571f
C4598 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 GND 0.04996f
C4599 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 GND 0.24182f
C4600 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 GND 0.06966f
C4601 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 GND 0.02985f
C4602 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 GND 0.05594f
C4603 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 GND 0.12602f
C4604 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 GND 0.12602f
C4605 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 GND 0.07553f
C4606 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 GND 0.03814f
C4607 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 GND 0.06323f
C4608 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 GND 0.07525f
C4609 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 GND 0.37895f
C4610 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 GND 0.03999f
C4611 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 GND 0.02271f
C4612 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 GND 0.04398f
C4613 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 GND 0.30646f
C4614 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 GND 0.31774f
C4615 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 GND 0.03438f
C4616 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 GND 0.0459f
C4617 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 GND 0.24094f
C4618 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 GND 0.24095f
C4619 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 GND 0.15608f
C4620 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 GND 0.03292f
C4621 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 GND 0.30645f
C4622 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 GND 0.08952f
C4623 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 GND 0.02228f
C4624 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 GND 0.0324f
C4625 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 GND 0.08303f
C4626 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 GND 0.08303f
C4627 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 GND 0.04316f
C4628 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 GND 0.04167f
C4629 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 GND 0.24695f
C4630 RingCounter_0.D_FlipFlop_16.Q.t4 GND 0.09863f
C4631 RingCounter_0.D_FlipFlop_16.Q.n0 GND 0.09693f
C4632 RingCounter_0.D_FlipFlop_16.Q.n1 GND 0.01059f
C4633 RingCounter_0.D_FlipFlop_16.Q.t6 GND 0.05128f
C4634 RingCounter_0.D_FlipFlop_16.Q.n2 GND 0.01477f
C4635 RingCounter_0.D_FlipFlop_16.Q.n4 GND 0.01186f
C4636 RingCounter_0.D_FlipFlop_16.Q.n5 GND 0.01493f
C4637 RingCounter_0.D_FlipFlop_16.Q.t9 GND 0.09863f
C4638 RingCounter_0.D_FlipFlop_16.Q.n6 GND 0.09693f
C4639 RingCounter_0.D_FlipFlop_16.Q.n7 GND 0.01059f
C4640 RingCounter_0.D_FlipFlop_16.Q.t7 GND 0.05128f
C4641 RingCounter_0.D_FlipFlop_16.Q.n8 GND 0.01477f
C4642 RingCounter_0.D_FlipFlop_16.Q.n10 GND 0.01186f
C4643 RingCounter_0.D_FlipFlop_16.Q.n12 GND 0.83774f
C4644 RingCounter_0.D_FlipFlop_16.Q.t5 GND 0.09863f
C4645 RingCounter_0.D_FlipFlop_16.Q.n13 GND 0.02881f
C4646 RingCounter_0.D_FlipFlop_16.Q.n14 GND 0.0125f
C4647 RingCounter_0.D_FlipFlop_16.Q.n15 GND 0.05497f
C4648 RingCounter_0.D_FlipFlop_16.Q.t8 GND 0.04587f
C4649 RingCounter_0.D_FlipFlop_16.Q.n16 GND 0.01439f
C4650 RingCounter_0.D_FlipFlop_16.Q.n17 GND 0.03074f
C4651 RingCounter_0.D_FlipFlop_16.Q.n18 GND 1.6069f
C4652 RingCounter_0.D_FlipFlop_16.Q.t1 GND 0.01338f
C4653 RingCounter_0.D_FlipFlop_16.Q.n19 GND 0.02059f
C4654 RingCounter_0.D_FlipFlop_16.Q.t3 GND 0.01366f
C4655 RingCounter_0.D_FlipFlop_16.Q.t2 GND 0.01338f
C4656 RingCounter_0.D_FlipFlop_16.Q.n20 GND 0.07608f
C4657 RingCounter_0.D_FlipFlop_16.Q.n21 GND 0.02531f
C4658 RingCounter_0.D_FlipFlop_16.Q.n22 GND 0.01548f
C4659 RingCounter_0.D_FlipFlop_16.Q.t0 GND 0.01286f
C4660 RingCounter_0.D_FlipFlop_16.Q.n23 GND 0.06309f
C4661 CDAC8_0.switch_0.Z.t2 GND 0.03316f
C4662 CDAC8_0.switch_0.Z.t1 GND 0.03316f
C4663 CDAC8_0.switch_0.Z.n0 GND 0.11982f
C4664 CDAC8_0.switch_0.Z.n1 GND 0.27578f
C4665 CDAC8_0.switch_0.Z.t3 GND 0.03482f
C4666 CDAC8_0.switch_0.Z.t5 GND 5.94383f
C4667 CDAC8_0.switch_0.Z.n2 GND 2.04684f
C4668 CDAC8_0.switch_0.Z.t7 GND 5.94383f
C4669 CDAC8_0.switch_0.Z.t6 GND 5.85885f
C4670 CDAC8_0.switch_0.Z.n3 GND 2.17361f
C4671 CDAC8_0.switch_0.Z.t4 GND 5.85885f
C4672 CDAC8_0.switch_0.Z.n4 GND 2.17361f
C4673 CDAC8_0.switch_0.Z.n5 GND 2.00334f
C4674 CDAC8_0.switch_0.Z.n6 GND 0.50573f
C4675 CDAC8_0.switch_0.Z.n7 GND 0.11883f
C4676 CDAC8_0.switch_0.Z.t0 GND 0.0348f
C4677 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 GND 0.06323f
C4678 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 GND 0.07525f
C4679 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 GND 0.38033f
C4680 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 GND 0.1927f
C4681 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 GND 0.0655f
C4682 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 GND 0.24183f
C4683 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 GND 0.23689f
C4684 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 GND 0.04996f
C4685 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 GND 0.46511f
C4686 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 GND 0.13587f
C4687 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 GND 0.03381f
C4688 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 GND 0.04918f
C4689 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 GND 0.12602f
C4690 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 GND 0.12602f
C4691 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 GND 0.06674f
C4692 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 GND 0.0608f
C4693 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 GND 0.13827f
C4694 D_FlipFlop_4.3-input-nand_2.C.t5 GND 0.3425f
C4695 D_FlipFlop_4.3-input-nand_2.C.n0 GND 0.3551f
C4696 D_FlipFlop_4.3-input-nand_2.C.n1 GND 0.03842f
C4697 D_FlipFlop_4.3-input-nand_2.C.t2 GND 0.04477f
C4698 D_FlipFlop_4.3-input-nand_2.C.n2 GND 0.11971f
C4699 D_FlipFlop_4.3-input-nand_2.C.n3 GND 0.09193f
C4700 D_FlipFlop_4.3-input-nand_2.C.t6 GND 0.17806f
C4701 D_FlipFlop_4.3-input-nand_2.C.t7 GND 0.34248f
C4702 D_FlipFlop_4.3-input-nand_2.C.n4 GND 0.10005f
C4703 D_FlipFlop_4.3-input-nand_2.C.n5 GND 0.04279f
C4704 D_FlipFlop_4.3-input-nand_2.C.n6 GND 0.079f
C4705 D_FlipFlop_4.3-input-nand_2.C.n7 GND 0.13677f
C4706 D_FlipFlop_4.3-input-nand_2.C.n8 GND 0.10181f
C4707 D_FlipFlop_4.3-input-nand_2.C.n9 GND 0.04823f
C4708 D_FlipFlop_4.3-input-nand_2.C.n10 GND 0.124f
C4709 D_FlipFlop_4.3-input-nand_2.C.t1 GND 0.04742f
C4710 D_FlipFlop_4.3-input-nand_2.C.t0 GND 0.04645f
C4711 D_FlipFlop_4.3-input-nand_2.C.n11 GND 0.26418f
C4712 D_FlipFlop_4.3-input-nand_2.C.n12 GND 0.08722f
C4713 D_FlipFlop_4.3-input-nand_2.C.t3 GND 0.04645f
C4714 D_FlipFlop_4.3-input-nand_2.C.n13 GND 0.293f
C4715 D_FlipFlop_4.3-input-nand_2.C.t4 GND 0.17045f
C4716 D_FlipFlop_4.3-input-nand_2.C.n14 GND 0.05129f
C4717 D_FlipFlop_4.3-input-nand_2.Vout.t4 GND 0.35515f
C4718 D_FlipFlop_4.3-input-nand_2.Vout.n0 GND 0.10375f
C4719 D_FlipFlop_4.3-input-nand_2.Vout.n1 GND 0.04502f
C4720 D_FlipFlop_4.3-input-nand_2.Vout.t3 GND 0.04632f
C4721 D_FlipFlop_4.3-input-nand_2.Vout.n2 GND 0.22028f
C4722 D_FlipFlop_4.3-input-nand_2.Vout.n3 GND 0.05002f
C4723 D_FlipFlop_4.3-input-nand_2.Vout.t6 GND 0.35517f
C4724 D_FlipFlop_4.3-input-nand_2.Vout.n4 GND 0.36759f
C4725 D_FlipFlop_4.3-input-nand_2.Vout.t5 GND 0.18465f
C4726 D_FlipFlop_4.3-input-nand_2.Vout.n5 GND 0.18106f
C4727 D_FlipFlop_4.3-input-nand_2.Vout.n6 GND 0.10557f
C4728 D_FlipFlop_4.3-input-nand_2.Vout.n7 GND 0.01331f
C4729 D_FlipFlop_4.3-input-nand_2.Vout.n8 GND 0.01454f
C4730 D_FlipFlop_4.3-input-nand_2.Vout.t1 GND 0.04918f
C4731 D_FlipFlop_4.3-input-nand_2.Vout.t0 GND 0.04817f
C4732 D_FlipFlop_4.3-input-nand_2.Vout.n9 GND 0.27396f
C4733 D_FlipFlop_4.3-input-nand_2.Vout.n10 GND 0.09115f
C4734 D_FlipFlop_4.3-input-nand_2.Vout.t2 GND 0.04817f
C4735 D_FlipFlop_4.3-input-nand_2.Vout.n11 GND 0.30324f
C4736 D_FlipFlop_4.3-input-nand_2.Vout.t7 GND 0.17747f
C4737 D_FlipFlop_4.3-input-nand_2.Vout.n12 GND 0.19793f
C4738 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 GND 0.07024f
C4739 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 GND 0.03989f
C4740 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 GND 0.07725f
C4741 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 GND 0.2799f
C4742 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 GND 0.27418f
C4743 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 GND 0.05783f
C4744 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 GND 0.53832f
C4745 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 GND 0.15726f
C4746 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 GND 0.03913f
C4747 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 GND 0.05692f
C4748 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 GND 0.14585f
C4749 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 GND 0.14585f
C4750 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 GND 0.07581f
C4751 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 GND 0.07318f
C4752 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 GND 0.07454f
C4753 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 GND 0.07302f
C4754 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 GND 0.41525f
C4755 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 GND 0.23391f
C4756 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 GND 0.22303f
C4757 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 GND 0.05201f
C4758 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 GND 0.22649f
C4759 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 GND 0.05616f
C4760 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 GND 0.39877f
C4761 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 GND 0.39189f
C4762 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 GND 0.04283f
C4763 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 GND 0.20732f
C4764 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 GND 0.05972f
C4765 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 GND 0.02559f
C4766 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 GND 0.04796f
C4767 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 GND 0.10804f
C4768 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 GND 0.10804f
C4769 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 GND 0.06475f
C4770 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 GND 0.05421f
C4771 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 GND 0.05522f
C4772 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 GND 0.05409f
C4773 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 GND 0.30759f
C4774 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 GND 0.17406f
C4775 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 GND 0.03715f
C4776 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 GND 0.05201f
C4777 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 GND 0.22649f
C4778 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 GND 0.05616f
C4779 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 GND 0.39877f
C4780 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 GND 0.39189f
C4781 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 GND 0.04283f
C4782 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 GND 0.20732f
C4783 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 GND 0.05972f
C4784 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 GND 0.02559f
C4785 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 GND 0.04796f
C4786 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 GND 0.10804f
C4787 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 GND 0.10804f
C4788 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 GND 0.06475f
C4789 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 GND 0.05421f
C4790 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 GND 0.05522f
C4791 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 GND 0.05409f
C4792 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 GND 0.30759f
C4793 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 GND 0.17406f
C4794 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 GND 0.03715f
C4795 And_Gate_5.A.t1 GND 0.03572f
C4796 Nand_Gate_3.Vout GND -0.07167f
C4797 And_Gate_5.A.n0 GND 0.02029f
C4798 And_Gate_5.A.n1 GND 0.03928f
C4799 And_Gate_5.A.t4 GND 0.14233f
C4800 And_Gate_5.Nand_Gate_0.A GND -0.10701f
C4801 And_Gate_5.A.n2 GND 0.13943f
C4802 And_Gate_5.A.n3 GND 0.02941f
C4803 And_Gate_5.A.t3 GND 0.27375f
C4804 And_Gate_5.A.n4 GND 0.07997f
C4805 And_Gate_5.A.n5 GND 0.0199f
C4806 And_Gate_5.A.n6 GND 0.02895f
C4807 And_Gate_5.A.n7 GND 0.55617f
C4808 And_Gate_5.A.n8 GND 0.55617f
C4809 And_Gate_5.A.n9 GND 0.03855f
C4810 And_Gate_5.A.t2 GND 0.03721f
C4811 And_Gate_5.A.t0 GND 0.04429f
C4812 And_Gate_5.A.n10 GND 0.22385f
C4813 And_Gate_5.A.n11 GND 0.11341f
C4814 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 GND 0.05969f
C4815 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 GND 0.15961f
C4816 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 GND 0.12257f
C4817 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 GND 0.23742f
C4818 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 GND 0.45664f
C4819 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 GND 0.1334f
C4820 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 GND 0.05705f
C4821 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 GND 0.10533f
C4822 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 GND 0.18236f
C4823 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 GND 0.13574f
C4824 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 GND 0.06431f
C4825 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 GND 0.45666f
C4826 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 GND 0.47347f
C4827 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 GND 0.05122f
C4828 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 GND 0.06839f
C4829 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 GND 0.22727f
C4830 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 GND 0.06194f
C4831 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 GND 0.39067f
C4832 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 GND 0.06323f
C4833 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 GND 0.06194f
C4834 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 GND 0.35224f
C4835 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 GND 0.11629f
C4836 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 GND 0.16533f
C4837 And_Gate_0.Vout.t1 GND 0.12492f
C4838 And_Gate_0.Inverter_0.Vout GND 0.03629f
C4839 And_Gate_0.Vout.n0 GND 0.13783f
C4840 And_Gate_0.Vout.t4 GND 0.95742f
C4841 D_FlipFlop_6.3-input-nand_0.C GND -0.56919f
C4842 And_Gate_0.Vout.n1 GND 0.99266f
C4843 And_Gate_0.Vout.n2 GND 0.10739f
C4844 And_Gate_0.Vout.n3 GND 0.14338f
C4845 And_Gate_0.Vout.t5 GND 0.44073f
C4846 D_FlipFlop_6.CLK GND -0.01479f
C4847 And_Gate_0.Vout.n4 GND 0.35269f
C4848 And_Gate_0.Vout.t3 GND 0.95737f
C4849 D_FlipFlop_6.3-input-nand_1.C GND -0.32001f
C4850 And_Gate_0.Vout.t6 GND 0.49778f
C4851 D_FlipFlop_6.Inverter_1.Vin GND -0.3108f
C4852 And_Gate_0.Vout.n5 GND 0.52493f
C4853 And_Gate_0.Vout.t2 GND 0.95737f
C4854 And_Gate_0.Vout.n6 GND 0.84748f
C4855 And_Gate_0.Vout.n7 GND 0.84981f
C4856 And_Gate_0.Vout.n8 GND 0.53181f
C4857 And_Gate_0.Vout.t7 GND 0.44069f
C4858 And_Gate_0.Vout.n9 GND 0.0818f
C4859 And_Gate_0.Vout.n10 GND 0.19316f
C4860 And_Gate_0.Vout.n11 GND 18.7304f
C4861 And_Gate_0.Vout.t0 GND 0.13044f
C4862 And_Gate_0.Vout.n12 GND 15.2812f
C4863 And_Gate_0.Vout.n13 GND 0.29731f
C4864 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 GND 0.05201f
C4865 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 GND 0.22649f
C4866 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 GND 0.05616f
C4867 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 GND 0.39877f
C4868 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 GND 0.39189f
C4869 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 GND 0.04283f
C4870 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 GND 0.20732f
C4871 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 GND 0.05972f
C4872 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 GND 0.02559f
C4873 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 GND 0.04796f
C4874 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 GND 0.10804f
C4875 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 GND 0.10804f
C4876 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 GND 0.06475f
C4877 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 GND 0.05421f
C4878 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 GND 0.05522f
C4879 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 GND 0.05409f
C4880 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 GND 0.30759f
C4881 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 GND 0.17406f
C4882 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 GND 0.03715f
C4883 And_Gate_6.Vout.t1 GND 0.09234f
C4884 And_Gate_6.Inverter_0.Vout GND -0.29682f
C4885 And_Gate_6.Vout.n0 GND 0.05245f
C4886 And_Gate_6.Vout.n1 GND 0.10156f
C4887 And_Gate_6.Vout.t5 GND 0.70775f
C4888 D_FlipFlop_3.3-input-nand_0.C GND -0.42076f
C4889 And_Gate_6.Vout.n2 GND 0.7338f
C4890 And_Gate_6.Vout.n3 GND 0.07939f
C4891 And_Gate_6.Vout.n4 GND 0.10599f
C4892 And_Gate_6.Vout.t2 GND 0.32576f
C4893 D_FlipFlop_3.CLK GND 0.04733f
C4894 And_Gate_6.Vout.n5 GND 0.31014f
C4895 And_Gate_6.Vout.n6 GND 0.09329f
C4896 And_Gate_6.Vout.t7 GND 0.70772f
C4897 D_FlipFlop_3.3-input-nand_1.C GND -0.23656f
C4898 And_Gate_6.Vout.t3 GND 0.36798f
C4899 D_FlipFlop_3.Inverter_1.Vin GND -0.22976f
C4900 And_Gate_6.Vout.n7 GND 0.38805f
C4901 And_Gate_6.Vout.t6 GND 0.70772f
C4902 And_Gate_6.Vout.n8 GND 0.62648f
C4903 And_Gate_6.Vout.n9 GND 0.6282f
C4904 And_Gate_6.Vout.n10 GND 0.39313f
C4905 And_Gate_6.Vout.t4 GND 0.32577f
C4906 And_Gate_6.Vout.n11 GND 7.68586f
C4907 And_Gate_6.Vout.n12 GND 5.63698f
C4908 And_Gate_6.Vout.n13 GND 0.09967f
C4909 And_Gate_6.Vout.t0 GND 0.09623f
C4910 And_Gate_6.Vout.n14 GND 0.57031f
C4911 Q4.t0 GND 0.01589f
C4912 Q4.n0 GND 0.07793f
C4913 Q4.n1 GND 0.01912f
C4914 Q4.t3 GND 0.01687f
C4915 Q4.t2 GND 0.01653f
C4916 Q4.n2 GND 0.09398f
C4917 Q4.n3 GND 0.03127f
C4918 Q4.t1 GND 0.01653f
C4919 Q4.n4 GND 0.02546f
C4920 Q4.n5 GND 0.03664f
C4921 Q4.n6 GND 0.01877f
C4922 Q4.t5 GND 0.12183f
C4923 Q4.n7 GND 0.03559f
C4924 Q4.n8 GND 0.01544f
C4925 Q4.n9 GND 0.0679f
C4926 Q4.t9 GND 0.05667f
C4927 Q4.n11 GND 0.01459f
C4928 Q4.n13 GND 3.26567f
C4929 Q4.n14 GND 1.24988f
C4930 Q4.t4 GND 0.12215f
C4931 Q4.t6 GND 0.12215f
C4932 Q4.t8 GND 0.06345f
C4933 Q4.n15 GND 0.09883f
C4934 Q4.n16 GND 0.07245f
C4935 Q4.t7 GND 0.06334f
C4936 Q4.n17 GND 0.02077f
C4937 Nand_Gate_1.A.t10 GND 0.27993f
C4938 Nand_Gate_1.A.n0 GND 0.08177f
C4939 Nand_Gate_1.A.n1 GND 0.03548f
C4940 Nand_Gate_1.A.n2 GND 0.15601f
C4941 Nand_Gate_1.A.t6 GND 0.1302f
C4942 Nand_Gate_1.A.n3 GND 0.04085f
C4943 Nand_Gate_1.A.t1 GND 0.03651f
C4944 Nand_Gate_1.A.n4 GND 0.159f
C4945 Nand_Gate_1.A.n5 GND 0.03942f
C4946 Nand_Gate_1.A.t7 GND 0.27994f
C4947 Nand_Gate_1.A.n6 GND 0.27511f
C4948 Nand_Gate_1.A.n7 GND 0.03007f
C4949 Nand_Gate_1.A.t11 GND 0.14554f
C4950 Nand_Gate_1.A.n8 GND 0.04192f
C4951 Nand_Gate_1.A.n9 GND 0.01797f
C4952 Nand_Gate_1.A.n10 GND 0.03367f
C4953 Nand_Gate_1.A.n11 GND 0.04236f
C4954 Nand_Gate_1.A.t9 GND 0.27994f
C4955 Nand_Gate_1.A.n12 GND 0.27511f
C4956 Nand_Gate_1.A.n13 GND 0.03007f
C4957 Nand_Gate_1.A.t4 GND 0.14554f
C4958 Nand_Gate_1.A.n14 GND 0.04192f
C4959 Nand_Gate_1.A.n15 GND 0.01797f
C4960 Nand_Gate_1.A.n16 GND 0.03367f
C4961 Nand_Gate_1.A.n18 GND 0.12656f
C4962 Nand_Gate_1.A.n19 GND 0.03459f
C4963 Nand_Gate_1.A.n20 GND 0.09204f
C4964 Nand_Gate_1.A.t5 GND 0.14555f
C4965 Nand_Gate_1.A.n21 GND 0.14257f
C4966 Nand_Gate_1.A.n22 GND 0.03007f
C4967 Nand_Gate_1.A.t8 GND 0.27993f
C4968 Nand_Gate_1.A.n23 GND 0.08177f
C4969 Nand_Gate_1.A.n24 GND 0.02035f
C4970 Nand_Gate_1.A.n25 GND 0.0296f
C4971 Nand_Gate_1.A.n26 GND 0.14551f
C4972 Nand_Gate_1.A.n27 GND 0.25531f
C4973 Nand_Gate_1.A.n28 GND 0.15873f
C4974 Nand_Gate_1.A.n29 GND 0.34318f
C4975 Nand_Gate_1.A.n31 GND 0.04546f
C4976 Nand_Gate_1.A.n32 GND 0.02608f
C4977 Nand_Gate_1.A.t0 GND 0.03876f
C4978 Nand_Gate_1.A.t3 GND 0.03797f
C4979 Nand_Gate_1.A.n33 GND 0.21593f
C4980 Nand_Gate_1.A.n34 GND 0.07184f
C4981 Nand_Gate_1.A.t2 GND 0.03797f
C4982 Nand_Gate_1.A.n35 GND 0.05849f
C4983 Nand_Gate_1.A.n36 GND 0.10356f
C4984 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 GND 0.0608f
C4985 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 GND 0.13827f
C4986 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 GND 0.06674f
C4987 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 GND 0.24183f
C4988 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 GND 0.23689f
C4989 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 GND 0.04996f
C4990 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 GND 0.46511f
C4991 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 GND 0.13587f
C4992 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 GND 0.03381f
C4993 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 GND 0.04918f
C4994 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 GND 0.12602f
C4995 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 GND 0.12602f
C4996 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 GND 0.0655f
C4997 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 GND 0.06323f
C4998 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 GND 0.07525f
C4999 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 GND 0.38033f
C5000 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 GND 0.1927f
C5001 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 GND 0.0608f
C5002 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 GND 0.13827f
C5003 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 GND 0.06674f
C5004 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 GND 0.24183f
C5005 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 GND 0.23689f
C5006 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 GND 0.04996f
C5007 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 GND 0.46511f
C5008 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 GND 0.13587f
C5009 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 GND 0.03381f
C5010 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 GND 0.04918f
C5011 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 GND 0.12602f
C5012 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 GND 0.12602f
C5013 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 GND 0.0655f
C5014 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 GND 0.06323f
C5015 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 GND 0.07525f
C5016 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 GND 0.38033f
C5017 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 GND 0.1927f
C5018 Q2.t9 GND 0.11806f
C5019 Q2.n0 GND 0.03449f
C5020 Q2.n1 GND 0.01496f
C5021 Q2.n2 GND 0.06579f
C5022 Q2.t8 GND 0.05415f
C5023 Q2.t1 GND 0.0154f
C5024 Q2.n3 GND 0.07552f
C5025 Q2.n4 GND 0.01853f
C5026 Q2.t3 GND 0.01635f
C5027 Q2.t2 GND 0.01601f
C5028 Q2.n5 GND 0.09106f
C5029 Q2.n6 GND 0.0303f
C5030 Q2.t0 GND 0.01601f
C5031 Q2.n7 GND 0.02467f
C5032 Q2.n8 GND 0.0409f
C5033 Q2.n9 GND 0.01975f
C5034 Q2.n11 GND 0.03836f
C5035 Q2.n12 GND 5.50481f
C5036 Q2.t4 GND 0.06148f
C5037 Q2.t7 GND 0.11836f
C5038 Q2.t5 GND 0.06148f
C5039 Q2.n13 GND 0.09576f
C5040 Q2.n14 GND 0.09631f
C5041 Q2.t6 GND 0.10522f
C5042 Q2.n15 GND 1.21113f
C5043 And_Gate_4.A.t1 GND 0.07612f
C5044 And_Gate_4.A.t2 GND 0.09059f
C5045 And_Gate_4.A.n0 GND 0.45787f
C5046 Nand_Gate_0.Vout GND -0.1466f
C5047 And_Gate_4.A.n1 GND 0.23199f
C5048 And_Gate_4.A.n2 GND 0.07886f
C5049 And_Gate_4.A.t3 GND 0.29114f
C5050 And_Gate_4.Nand_Gate_0.A GND -0.21888f
C5051 And_Gate_4.A.n3 GND 0.28519f
C5052 And_Gate_4.A.n4 GND 0.06015f
C5053 And_Gate_4.A.t4 GND 0.55994f
C5054 And_Gate_4.A.n5 GND 0.16357f
C5055 And_Gate_4.A.n6 GND 0.0407f
C5056 And_Gate_4.A.n7 GND 0.05921f
C5057 And_Gate_4.A.n8 GND 1.13762f
C5058 And_Gate_4.A.n9 GND 1.13762f
C5059 And_Gate_4.A.n10 GND 0.08035f
C5060 And_Gate_4.A.n11 GND 0.0415f
C5061 And_Gate_4.A.t0 GND 0.07306f
C5062 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 GND 0.06358f
C5063 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 GND 0.03611f
C5064 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 GND 0.06992f
C5065 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 GND 0.25335f
C5066 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 GND 0.24817f
C5067 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 GND 0.05234f
C5068 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 GND 0.48726f
C5069 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 GND 0.14234f
C5070 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 GND 0.03542f
C5071 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 GND 0.05152f
C5072 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 GND 0.13202f
C5073 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 GND 0.13202f
C5074 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 GND 0.06862f
C5075 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 GND 0.06624f
C5076 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 GND 0.07883f
C5077 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 GND 0.39844f
C5078 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 GND 0.20187f
C5079 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 GND 0.05958f
C5080 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 GND 0.0577f
C5081 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 GND 0.12257f
C5082 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 GND 0.23742f
C5083 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 GND 0.45664f
C5084 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 GND 0.1334f
C5085 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 GND 0.05705f
C5086 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 GND 0.10533f
C5087 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 GND 0.18236f
C5088 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 GND 0.13574f
C5089 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 GND 0.06431f
C5090 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 GND 0.45666f
C5091 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 GND 0.47347f
C5092 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 GND 0.05122f
C5093 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 GND 0.06839f
C5094 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 GND 0.22727f
C5095 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 GND 0.06194f
C5096 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 GND 0.39067f
C5097 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 GND 0.06323f
C5098 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 GND 0.06194f
C5099 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 GND 0.35224f
C5100 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 GND 0.11629f
C5101 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 GND 0.16533f
C5102 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 GND 0.07037f
C5103 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 GND 0.16004f
C5104 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 GND 0.07725f
C5105 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 GND 0.2799f
C5106 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 GND 0.27418f
C5107 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 GND 0.05783f
C5108 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 GND 0.53832f
C5109 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 GND 0.15726f
C5110 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 GND 0.03913f
C5111 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 GND 0.05692f
C5112 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 GND 0.14585f
C5113 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 GND 0.14585f
C5114 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 GND 0.07581f
C5115 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 GND 0.07318f
C5116 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 GND 0.07454f
C5117 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 GND 0.07302f
C5118 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 GND 0.41525f
C5119 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 GND 0.23391f
C5120 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 GND 0.22303f
C5121 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 GND 0.07024f
C5122 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 GND 0.03989f
C5123 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 GND 0.07725f
C5124 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 GND 0.2799f
C5125 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 GND 0.27418f
C5126 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 GND 0.05783f
C5127 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 GND 0.53832f
C5128 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 GND 0.15726f
C5129 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 GND 0.03913f
C5130 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 GND 0.05692f
C5131 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 GND 0.14585f
C5132 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 GND 0.14585f
C5133 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 GND 0.07581f
C5134 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 GND 0.07318f
C5135 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 GND 0.07454f
C5136 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 GND 0.07302f
C5137 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 GND 0.41525f
C5138 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 GND 0.23391f
C5139 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 GND 0.22303f
C5140 And_Gate_2.Vout.t1 GND 0.10621f
C5141 And_Gate_2.Inverter_0.Vout GND 0.03085f
C5142 And_Gate_2.Vout.n0 GND 0.11719f
C5143 And_Gate_2.Vout.t7 GND 0.81407f
C5144 D_FlipFlop_5.3-input-nand_0.C GND -0.48397f
C5145 And_Gate_2.Vout.n1 GND 0.84403f
C5146 And_Gate_2.Vout.n2 GND 0.09131f
C5147 And_Gate_2.Vout.n3 GND 0.12192f
C5148 And_Gate_2.Vout.t4 GND 0.37472f
C5149 D_FlipFlop_5.CLK GND -0.0253f
C5150 And_Gate_2.Vout.n4 GND 0.294f
C5151 And_Gate_2.Vout.t3 GND 0.81403f
C5152 D_FlipFlop_5.3-input-nand_1.C GND -0.2721f
C5153 And_Gate_2.Vout.t5 GND 0.42325f
C5154 D_FlipFlop_5.Inverter_1.Vin GND -0.26427f
C5155 And_Gate_2.Vout.n5 GND 0.44634f
C5156 And_Gate_2.Vout.t2 GND 0.81403f
C5157 And_Gate_2.Vout.n6 GND 0.72059f
C5158 And_Gate_2.Vout.n7 GND 0.72257f
C5159 And_Gate_2.Vout.n8 GND 0.45218f
C5160 And_Gate_2.Vout.t6 GND 0.37471f
C5161 And_Gate_2.Vout.n9 GND 0.07492f
C5162 And_Gate_2.Vout.n10 GND 0.17642f
C5163 And_Gate_2.Vout.n11 GND 11.6967f
C5164 And_Gate_2.Vout.t0 GND 0.11091f
C5165 And_Gate_2.Vout.n12 GND 9.27182f
C5166 And_Gate_2.Vout.n13 GND 0.2528f
C5167 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 GND 0.36784f
C5168 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 GND 0.10746f
C5169 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 GND 0.04662f
C5170 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 GND 0.04798f
C5171 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 GND 0.22815f
C5172 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 GND 0.0518f
C5173 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 GND 0.36785f
C5174 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 GND 0.38072f
C5175 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 GND 0.19125f
C5176 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 GND 0.18752f
C5177 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 GND 0.10934f
C5178 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 GND 0.01378f
C5179 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 GND 0.01506f
C5180 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 GND 0.05094f
C5181 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 GND 0.04989f
C5182 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 GND 0.28374f
C5183 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 GND 0.09441f
C5184 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 GND 0.04989f
C5185 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 GND 0.31407f
C5186 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 GND 0.1838f
C5187 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 GND 0.205f
C5188 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 GND 0.07037f
C5189 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 GND 0.16004f
C5190 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 GND 0.07725f
C5191 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 GND 0.2799f
C5192 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 GND 0.27418f
C5193 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 GND 0.05783f
C5194 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 GND 0.53832f
C5195 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 GND 0.15726f
C5196 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 GND 0.03913f
C5197 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 GND 0.05692f
C5198 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 GND 0.14585f
C5199 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 GND 0.14585f
C5200 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 GND 0.07581f
C5201 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 GND 0.07318f
C5202 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 GND 0.07454f
C5203 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 GND 0.07302f
C5204 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 GND 0.41525f
C5205 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 GND 0.23391f
C5206 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 GND 0.22303f
C5207 D_FlipFlop_5.3-input-nand_2.Vout.t4 GND 0.35515f
C5208 D_FlipFlop_5.3-input-nand_2.Vout.n0 GND 0.10375f
C5209 D_FlipFlop_5.3-input-nand_2.Vout.n1 GND 0.04502f
C5210 D_FlipFlop_5.3-input-nand_2.Vout.n2 GND 0.19793f
C5211 D_FlipFlop_5.3-input-nand_2.Vout.t6 GND 0.17747f
C5212 D_FlipFlop_5.3-input-nand_2.Vout.t1 GND 0.04817f
C5213 D_FlipFlop_5.3-input-nand_2.Vout.n3 GND 0.30324f
C5214 D_FlipFlop_5.3-input-nand_2.Vout.t3 GND 0.04918f
C5215 D_FlipFlop_5.3-input-nand_2.Vout.t2 GND 0.04817f
C5216 D_FlipFlop_5.3-input-nand_2.Vout.n4 GND 0.27396f
C5217 D_FlipFlop_5.3-input-nand_2.Vout.n5 GND 0.09115f
C5218 D_FlipFlop_5.3-input-nand_2.Vout.n6 GND 0.01454f
C5219 D_FlipFlop_5.3-input-nand_2.Vout.n7 GND 0.01331f
C5220 D_FlipFlop_5.3-input-nand_2.Vout.t7 GND 0.35517f
C5221 D_FlipFlop_5.3-input-nand_2.Vout.n8 GND 0.36759f
C5222 D_FlipFlop_5.3-input-nand_2.Vout.t5 GND 0.18465f
C5223 D_FlipFlop_5.3-input-nand_2.Vout.n9 GND 0.18106f
C5224 D_FlipFlop_5.3-input-nand_2.Vout.n10 GND 0.10557f
C5225 D_FlipFlop_5.3-input-nand_2.Vout.n11 GND 0.05002f
C5226 D_FlipFlop_5.3-input-nand_2.Vout.t0 GND 0.04632f
C5227 D_FlipFlop_5.3-input-nand_2.Vout.n12 GND 0.22028f
C5228 Nand_Gate_7.A.t10 GND 0.27993f
C5229 Nand_Gate_7.A.n0 GND 0.08177f
C5230 Nand_Gate_7.A.n1 GND 0.03548f
C5231 Nand_Gate_7.A.n2 GND 0.15601f
C5232 Nand_Gate_7.A.t6 GND 0.1302f
C5233 Nand_Gate_7.A.n3 GND 0.04085f
C5234 Nand_Gate_7.A.t1 GND 0.03651f
C5235 Nand_Gate_7.A.n4 GND 0.159f
C5236 Nand_Gate_7.A.n5 GND 0.03942f
C5237 Nand_Gate_7.A.t7 GND 0.27994f
C5238 Nand_Gate_7.A.n6 GND 0.27511f
C5239 Nand_Gate_7.A.n7 GND 0.03007f
C5240 Nand_Gate_7.A.t5 GND 0.14554f
C5241 Nand_Gate_7.A.n8 GND 0.04192f
C5242 Nand_Gate_7.A.n9 GND 0.01797f
C5243 Nand_Gate_7.A.n10 GND 0.03367f
C5244 Nand_Gate_7.A.n11 GND 0.04236f
C5245 Nand_Gate_7.A.t4 GND 0.27994f
C5246 Nand_Gate_7.A.n12 GND 0.27511f
C5247 Nand_Gate_7.A.n13 GND 0.03007f
C5248 Nand_Gate_7.A.t8 GND 0.14554f
C5249 Nand_Gate_7.A.n14 GND 0.04192f
C5250 Nand_Gate_7.A.n15 GND 0.01797f
C5251 Nand_Gate_7.A.n16 GND 0.03367f
C5252 Nand_Gate_7.A.n18 GND 0.12703f
C5253 Nand_Gate_7.A.n19 GND 0.0915f
C5254 Nand_Gate_7.A.t9 GND 0.14555f
C5255 Nand_Gate_7.A.n20 GND 0.14257f
C5256 Nand_Gate_7.A.n21 GND 0.03007f
C5257 Nand_Gate_7.A.t11 GND 0.27993f
C5258 Nand_Gate_7.A.n22 GND 0.08177f
C5259 Nand_Gate_7.A.n23 GND 0.02035f
C5260 Nand_Gate_7.A.n24 GND 0.0296f
C5261 Nand_Gate_7.A.n25 GND 0.14551f
C5262 Nand_Gate_7.A.n26 GND 0.25531f
C5263 Nand_Gate_7.A.n27 GND 0.15839f
C5264 Nand_Gate_7.A.n28 GND 0.34271f
C5265 Nand_Gate_7.A.n30 GND 0.04546f
C5266 Nand_Gate_7.A.n31 GND 0.02608f
C5267 Nand_Gate_7.A.t0 GND 0.03876f
C5268 Nand_Gate_7.A.t3 GND 0.03797f
C5269 Nand_Gate_7.A.n32 GND 0.21593f
C5270 Nand_Gate_7.A.n33 GND 0.07184f
C5271 Nand_Gate_7.A.t2 GND 0.03797f
C5272 Nand_Gate_7.A.n34 GND 0.05849f
C5273 Nand_Gate_7.A.n35 GND 0.10356f
C5274 Nand_Gate_1.Vout.t1 GND 0.08189f
C5275 Nand_Gate_1.Vout.n0 GND 0.04651f
C5276 Nand_Gate_1.Vout.n1 GND 0.09007f
C5277 Nand_Gate_1.Vout.t4 GND 0.32633f
C5278 Nand_Gate_1.Vout.n2 GND 0.31966f
C5279 Nand_Gate_1.Vout.n3 GND 0.06742f
C5280 Nand_Gate_1.Vout.t3 GND 0.62762f
C5281 Nand_Gate_1.Vout.n4 GND 0.18335f
C5282 Nand_Gate_1.Vout.n5 GND 0.04562f
C5283 Nand_Gate_1.Vout.n6 GND 0.06636f
C5284 Nand_Gate_1.Vout.n7 GND 1.35316f
C5285 Nand_Gate_1.Vout.n8 GND 1.35316f
C5286 Nand_Gate_1.Vout.n9 GND 0.08839f
C5287 Nand_Gate_1.Vout.t0 GND 0.08532f
C5288 Nand_Gate_1.Vout.t2 GND 0.10154f
C5289 Nand_Gate_1.Vout.n10 GND 0.51322f
C5290 Nand_Gate_1.Vout.n11 GND 0.26003f
C5291 D_FlipFlop_7.3-input-nand_2.Vout.t4 GND 0.35515f
C5292 D_FlipFlop_7.3-input-nand_2.Vout.n0 GND 0.10375f
C5293 D_FlipFlop_7.3-input-nand_2.Vout.n1 GND 0.04502f
C5294 D_FlipFlop_7.3-input-nand_2.Vout.t1 GND 0.04632f
C5295 D_FlipFlop_7.3-input-nand_2.Vout.n2 GND 0.22028f
C5296 D_FlipFlop_7.3-input-nand_2.Vout.n3 GND 0.05002f
C5297 D_FlipFlop_7.3-input-nand_2.Vout.t7 GND 0.35517f
C5298 D_FlipFlop_7.3-input-nand_2.Vout.n4 GND 0.36759f
C5299 D_FlipFlop_7.3-input-nand_2.Vout.t5 GND 0.18465f
C5300 D_FlipFlop_7.3-input-nand_2.Vout.n5 GND 0.18106f
C5301 D_FlipFlop_7.3-input-nand_2.Vout.n6 GND 0.10557f
C5302 D_FlipFlop_7.3-input-nand_2.Vout.n7 GND 0.01331f
C5303 D_FlipFlop_7.3-input-nand_2.Vout.n8 GND 0.01454f
C5304 D_FlipFlop_7.3-input-nand_2.Vout.t3 GND 0.04918f
C5305 D_FlipFlop_7.3-input-nand_2.Vout.t0 GND 0.04817f
C5306 D_FlipFlop_7.3-input-nand_2.Vout.n9 GND 0.27396f
C5307 D_FlipFlop_7.3-input-nand_2.Vout.n10 GND 0.09115f
C5308 D_FlipFlop_7.3-input-nand_2.Vout.t2 GND 0.04817f
C5309 D_FlipFlop_7.3-input-nand_2.Vout.n11 GND 0.30324f
C5310 D_FlipFlop_7.3-input-nand_2.Vout.t6 GND 0.17747f
C5311 D_FlipFlop_7.3-input-nand_2.Vout.n12 GND 0.19793f
C5312 D_FlipFlop_7.3-input-nand_2.C.t7 GND 0.3425f
C5313 D_FlipFlop_7.3-input-nand_2.C.n0 GND 0.3551f
C5314 D_FlipFlop_7.3-input-nand_2.C.n1 GND 0.03842f
C5315 D_FlipFlop_7.3-input-nand_2.C.t2 GND 0.04477f
C5316 D_FlipFlop_7.3-input-nand_2.C.n2 GND 0.11971f
C5317 D_FlipFlop_7.3-input-nand_2.C.n3 GND 0.09193f
C5318 D_FlipFlop_7.3-input-nand_2.C.t5 GND 0.17806f
C5319 D_FlipFlop_7.3-input-nand_2.C.t6 GND 0.34248f
C5320 D_FlipFlop_7.3-input-nand_2.C.n4 GND 0.10005f
C5321 D_FlipFlop_7.3-input-nand_2.C.n5 GND 0.04279f
C5322 D_FlipFlop_7.3-input-nand_2.C.n6 GND 0.079f
C5323 D_FlipFlop_7.3-input-nand_2.C.n7 GND 0.13677f
C5324 D_FlipFlop_7.3-input-nand_2.C.n8 GND 0.10181f
C5325 D_FlipFlop_7.3-input-nand_2.C.n9 GND 0.04823f
C5326 D_FlipFlop_7.3-input-nand_2.C.n10 GND 0.124f
C5327 D_FlipFlop_7.3-input-nand_2.C.t1 GND 0.04742f
C5328 D_FlipFlop_7.3-input-nand_2.C.t0 GND 0.04645f
C5329 D_FlipFlop_7.3-input-nand_2.C.n11 GND 0.26418f
C5330 D_FlipFlop_7.3-input-nand_2.C.n12 GND 0.08722f
C5331 D_FlipFlop_7.3-input-nand_2.C.t3 GND 0.04645f
C5332 D_FlipFlop_7.3-input-nand_2.C.n13 GND 0.293f
C5333 D_FlipFlop_7.3-input-nand_2.C.t4 GND 0.17045f
C5334 D_FlipFlop_7.3-input-nand_2.C.n14 GND 0.05129f
C5335 Q5.t2 GND 0.01626f
C5336 Q5.n0 GND 0.07974f
C5337 Q5.n1 GND 0.01957f
C5338 Q5.t1 GND 0.01726f
C5339 Q5.t0 GND 0.01691f
C5340 Q5.n2 GND 0.09616f
C5341 Q5.n3 GND 0.03199f
C5342 Q5.t3 GND 0.01691f
C5343 Q5.n4 GND 0.02605f
C5344 Q5.n5 GND 0.03693f
C5345 Q5.n6 GND 0.0192f
C5346 Q5.t8 GND 0.12466f
C5347 Q5.n7 GND 0.03642f
C5348 Q5.n8 GND 0.0158f
C5349 Q5.n9 GND 0.06947f
C5350 Q5.t9 GND 0.05798f
C5351 Q5.n11 GND 0.0161f
C5352 Q5.n13 GND 3.34141f
C5353 Q5.t6 GND 0.12498f
C5354 Q5.t7 GND 0.12498f
C5355 Q5.t5 GND 0.06492f
C5356 Q5.n14 GND 0.10112f
C5357 Q5.n15 GND 0.1017f
C5358 Q5.t4 GND 0.05702f
C5359 Q5.n16 GND 1.27887f
C5360 And_Gate_5.Vout.t1 GND 0.12971f
C5361 And_Gate_5.Inverter_0.Vout GND -0.41694f
C5362 And_Gate_5.Vout.n0 GND 0.07367f
C5363 And_Gate_5.Vout.n1 GND 0.14266f
C5364 And_Gate_5.Vout.t3 GND 0.99417f
C5365 D_FlipFlop_1.3-input-nand_0.C GND -0.59104f
C5366 And_Gate_5.Vout.n2 GND 1.03076f
C5367 And_Gate_5.Vout.n3 GND 0.11151f
C5368 And_Gate_5.Vout.n4 GND 0.14889f
C5369 And_Gate_5.Vout.t6 GND 0.45759f
C5370 D_FlipFlop_1.CLK GND 0.04956f
C5371 And_Gate_5.Vout.n5 GND 0.43197f
C5372 And_Gate_5.Vout.n6 GND 0.13105f
C5373 And_Gate_5.Vout.t5 GND 0.99413f
C5374 D_FlipFlop_1.3-input-nand_1.C GND -0.33229f
C5375 And_Gate_5.Vout.t7 GND 0.51689f
C5376 D_FlipFlop_1.Inverter_1.Vin GND -0.32274f
C5377 And_Gate_5.Vout.n7 GND 0.54508f
C5378 And_Gate_5.Vout.t4 GND 0.99413f
C5379 And_Gate_5.Vout.n8 GND 0.88002f
C5380 And_Gate_5.Vout.n9 GND 0.88243f
C5381 And_Gate_5.Vout.n10 GND 0.55222f
C5382 And_Gate_5.Vout.t2 GND 0.45761f
C5383 And_Gate_5.Vout.n11 GND 0.02134f
C5384 And_Gate_5.Vout.n12 GND 24.0592f
C5385 And_Gate_5.Vout.n13 GND 21.6821f
C5386 And_Gate_5.Vout.n14 GND 0.14f
C5387 And_Gate_5.Vout.t0 GND 0.13517f
C5388 And_Gate_5.Vout.n15 GND 0.8011f
C5389 Q7.t1 GND 0.01626f
C5390 Q7.n0 GND 0.07974f
C5391 Q7.n1 GND 0.01957f
C5392 Q7.t2 GND 0.01726f
C5393 Q7.t3 GND 0.01691f
C5394 Q7.n2 GND 0.09616f
C5395 Q7.n3 GND 0.03199f
C5396 Q7.t0 GND 0.01691f
C5397 Q7.n4 GND 0.02605f
C5398 Q7.n5 GND 0.03769f
C5399 Q7.n6 GND 0.0192f
C5400 Q7.t5 GND 0.12466f
C5401 Q7.n7 GND 0.03642f
C5402 Q7.n8 GND 0.0158f
C5403 Q7.n9 GND 0.06947f
C5404 Q7.t6 GND 0.05798f
C5405 Q7.n11 GND 0.01451f
C5406 Q7.n13 GND 3.34141f
C5407 Q7.t7 GND 0.12498f
C5408 Q7.t8 GND 0.12498f
C5409 Q7.t4 GND 0.06492f
C5410 Q7.n14 GND 0.10112f
C5411 Q7.n15 GND 0.1017f
C5412 Q7.t9 GND 0.05702f
C5413 Q7.n16 GND 1.27887f
C5414 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 GND 0.07024f
C5415 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 GND 0.03989f
C5416 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 GND 0.07725f
C5417 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 GND 0.2799f
C5418 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 GND 0.27418f
C5419 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 GND 0.05783f
C5420 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 GND 0.53832f
C5421 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 GND 0.15726f
C5422 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 GND 0.03913f
C5423 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 GND 0.05692f
C5424 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 GND 0.14585f
C5425 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 GND 0.14585f
C5426 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 GND 0.07581f
C5427 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 GND 0.07318f
C5428 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 GND 0.07454f
C5429 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 GND 0.07302f
C5430 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 GND 0.41525f
C5431 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 GND 0.23391f
C5432 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 GND 0.22303f
C5433 Nand_Gate_1.B.t13 GND 0.47211f
C5434 Nand_Gate_1.B.n0 GND 0.13792f
C5435 Nand_Gate_1.B.n1 GND 0.05984f
C5436 Nand_Gate_1.B.n2 GND 0.26311f
C5437 Nand_Gate_1.B.t16 GND 0.21959f
C5438 Nand_Gate_1.B.n3 GND 0.06889f
C5439 Nand_Gate_1.B.t2 GND 0.06158f
C5440 Nand_Gate_1.B.n4 GND 0.26816f
C5441 Nand_Gate_1.B.n5 GND 0.06649f
C5442 Nand_Gate_1.B.t10 GND 0.47213f
C5443 Nand_Gate_1.B.n6 GND 0.46399f
C5444 Nand_Gate_1.B.n7 GND 0.05071f
C5445 Nand_Gate_1.B.t6 GND 0.24546f
C5446 Nand_Gate_1.B.n8 GND 0.07071f
C5447 Nand_Gate_1.B.n9 GND 0.0303f
C5448 Nand_Gate_1.B.n10 GND 0.05678f
C5449 Nand_Gate_1.B.n11 GND 0.07145f
C5450 Nand_Gate_1.B.t5 GND 0.47213f
C5451 Nand_Gate_1.B.n12 GND 0.46399f
C5452 Nand_Gate_1.B.n13 GND 0.05071f
C5453 Nand_Gate_1.B.t11 GND 0.24546f
C5454 Nand_Gate_1.B.n14 GND 0.07071f
C5455 Nand_Gate_1.B.n15 GND 0.0303f
C5456 Nand_Gate_1.B.n16 GND 0.05678f
C5457 Nand_Gate_1.B.n18 GND 0.21345f
C5458 Nand_Gate_1.B.n19 GND 0.05834f
C5459 Nand_Gate_1.B.n20 GND 0.15524f
C5460 Nand_Gate_1.B.t15 GND 0.47213f
C5461 Nand_Gate_1.B.n21 GND 0.47546f
C5462 Nand_Gate_1.B.n22 GND 0.05071f
C5463 Nand_Gate_1.B.t14 GND 0.24546f
C5464 Nand_Gate_1.B.n23 GND 0.07071f
C5465 Nand_Gate_1.B.n24 GND 0.01883f
C5466 Nand_Gate_1.B.n25 GND 0.02935f
C5467 Nand_Gate_1.B.n26 GND 0.29279f
C5468 Nand_Gate_1.B.t8 GND 0.47213f
C5469 Nand_Gate_1.B.n27 GND 0.47546f
C5470 Nand_Gate_1.B.n28 GND 0.05071f
C5471 Nand_Gate_1.B.t7 GND 0.24546f
C5472 Nand_Gate_1.B.n29 GND 0.07071f
C5473 Nand_Gate_1.B.n30 GND 0.01883f
C5474 Nand_Gate_1.B.n31 GND 0.02935f
C5475 Nand_Gate_1.B.n33 GND 0.76027f
C5476 Nand_Gate_1.B.n34 GND 0.31374f
C5477 Nand_Gate_1.B.n35 GND 0.13131f
C5478 Nand_Gate_1.B.t17 GND 0.47211f
C5479 Nand_Gate_1.B.n36 GND 0.13792f
C5480 Nand_Gate_1.B.n37 GND 0.05984f
C5481 Nand_Gate_1.B.n38 GND 0.26311f
C5482 Nand_Gate_1.B.t9 GND 0.21957f
C5483 Nand_Gate_1.B.n39 GND 0.06876f
C5484 Nand_Gate_1.B.n40 GND 0.15969f
C5485 Nand_Gate_1.B.n41 GND 3.82373f
C5486 Nand_Gate_1.B.t4 GND 0.24547f
C5487 Nand_Gate_1.B.n42 GND 0.26225f
C5488 Nand_Gate_1.B.t12 GND 0.47211f
C5489 Nand_Gate_1.B.n43 GND 1.07465f
C5490 Nand_Gate_1.B.n44 GND 5.83655f
C5491 Nand_Gate_1.B.n45 GND 0.08001f
C5492 Nand_Gate_1.B.n46 GND 0.26771f
C5493 Nand_Gate_1.B.n47 GND 0.5788f
C5494 Nand_Gate_1.B.n49 GND 0.07667f
C5495 Nand_Gate_1.B.n50 GND 0.04399f
C5496 Nand_Gate_1.B.t1 GND 0.06538f
C5497 Nand_Gate_1.B.t0 GND 0.06404f
C5498 Nand_Gate_1.B.n51 GND 0.36418f
C5499 Nand_Gate_1.B.n52 GND 0.12117f
C5500 Nand_Gate_1.B.t3 GND 0.06404f
C5501 Nand_Gate_1.B.n53 GND 0.09864f
C5502 Nand_Gate_1.B.n54 GND 0.17466f
C5503 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 GND 0.04998f
C5504 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 GND 0.02839f
C5505 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 GND 0.05497f
C5506 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 GND 0.38308f
C5507 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 GND 0.39717f
C5508 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 GND 0.04297f
C5509 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 GND 0.05737f
C5510 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 GND 0.30118f
C5511 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 GND 0.30119f
C5512 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 GND 0.1951f
C5513 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 GND 0.04115f
C5514 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 GND 0.38306f
C5515 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 GND 0.1119f
C5516 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 GND 0.02784f
C5517 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 GND 0.0405f
C5518 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 GND 0.10379f
C5519 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 GND 0.10379f
C5520 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 GND 0.05395f
C5521 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 GND 0.05208f
C5522 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 GND 0.30868f
C5523 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 GND 0.36784f
C5524 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 GND 0.10746f
C5525 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 GND 0.04662f
C5526 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 GND 0.04798f
C5527 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 GND 0.22815f
C5528 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 GND 0.0518f
C5529 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 GND 0.36785f
C5530 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 GND 0.38072f
C5531 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 GND 0.19125f
C5532 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 GND 0.18752f
C5533 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 GND 0.10934f
C5534 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 GND 0.01378f
C5535 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 GND 0.01095f
C5536 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 GND 0.05094f
C5537 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 GND 0.04989f
C5538 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 GND 0.28374f
C5539 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 GND 0.09258f
C5540 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 GND 0.04989f
C5541 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 GND 0.31407f
C5542 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 GND 0.1838f
C5543 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 GND 0.205f
C5544 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 GND 0.04607f
C5545 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 GND 0.10477f
C5546 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 GND 0.05057f
C5547 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 GND 0.35243f
C5548 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 GND 0.3654f
C5549 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 GND 0.03953f
C5550 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 GND 0.05278f
C5551 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 GND 0.27708f
C5552 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 GND 0.27709f
C5553 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 GND 0.17949f
C5554 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 GND 0.03786f
C5555 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 GND 0.35241f
C5556 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 GND 0.10295f
C5557 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 GND 0.02562f
C5558 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 GND 0.03726f
C5559 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 GND 0.09548f
C5560 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 GND 0.09548f
C5561 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 GND 0.04963f
C5562 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 GND 0.04792f
C5563 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 GND 0.28399f
C5564 Nand_Gate_3.B.t9 GND 0.33127f
C5565 Nand_Gate_3.B.n0 GND 0.09677f
C5566 Nand_Gate_3.B.n1 GND 0.04199f
C5567 Nand_Gate_3.B.n2 GND 0.18462f
C5568 Nand_Gate_3.B.t7 GND 0.15408f
C5569 Nand_Gate_3.B.n3 GND 0.04834f
C5570 Nand_Gate_3.B.n4 GND 0.12256f
C5571 Nand_Gate_3.B.t1 GND 0.04493f
C5572 Nand_Gate_3.B.n5 GND 0.06922f
C5573 Nand_Gate_3.B.t3 GND 0.04587f
C5574 Nand_Gate_3.B.t2 GND 0.04493f
C5575 Nand_Gate_3.B.n6 GND 0.25554f
C5576 Nand_Gate_3.B.n7 GND 0.08338f
C5577 Nand_Gate_3.B.n8 GND 0.02717f
C5578 Nand_Gate_3.B.n9 GND 0.05379f
C5579 Nand_Gate_3.B.t11 GND 0.33129f
C5580 Nand_Gate_3.B.n10 GND 0.32557f
C5581 Nand_Gate_3.B.n11 GND 0.03558f
C5582 Nand_Gate_3.B.t5 GND 0.17224f
C5583 Nand_Gate_3.B.n12 GND 0.04961f
C5584 Nand_Gate_3.B.n13 GND 0.02126f
C5585 Nand_Gate_3.B.n14 GND 0.03984f
C5586 Nand_Gate_3.B.n15 GND 0.05014f
C5587 Nand_Gate_3.B.t4 GND 0.33129f
C5588 Nand_Gate_3.B.n16 GND 0.32557f
C5589 Nand_Gate_3.B.n17 GND 0.03558f
C5590 Nand_Gate_3.B.t10 GND 0.17224f
C5591 Nand_Gate_3.B.n18 GND 0.04961f
C5592 Nand_Gate_3.B.n19 GND 0.02126f
C5593 Nand_Gate_3.B.n20 GND 0.03984f
C5594 Nand_Gate_3.B.n22 GND 0.15033f
C5595 Nand_Gate_3.B.n23 GND 0.41862f
C5596 Nand_Gate_3.B.n24 GND 0.18785f
C5597 Nand_Gate_3.B.t6 GND 0.17224f
C5598 Nand_Gate_3.B.t8 GND 0.33127f
C5599 Nand_Gate_3.B.n25 GND 0.09677f
C5600 Nand_Gate_3.B.n26 GND 0.04139f
C5601 Nand_Gate_3.B.n27 GND 0.07641f
C5602 Nand_Gate_3.B.n28 GND 0.87221f
C5603 Nand_Gate_3.B.n29 GND 1.18609f
C5604 Nand_Gate_3.B.n30 GND 0.05328f
C5605 Nand_Gate_3.B.n31 GND 0.01961f
C5606 Nand_Gate_3.B.n33 GND 0.04665f
C5607 Nand_Gate_3.B.t0 GND 0.04321f
C5608 Nand_Gate_3.B.n34 GND 0.18816f
C5609 Nand_Gate_2.Vout.t1 GND 0.07306f
C5610 Nand_Gate_2.Vout.n0 GND 0.0415f
C5611 Nand_Gate_2.Vout.n1 GND 0.08035f
C5612 Nand_Gate_2.Vout.t4 GND 0.29114f
C5613 Nand_Gate_2.Vout.n2 GND 0.28519f
C5614 Nand_Gate_2.Vout.n3 GND 0.06015f
C5615 Nand_Gate_2.Vout.t3 GND 0.55994f
C5616 Nand_Gate_2.Vout.n4 GND 0.16357f
C5617 Nand_Gate_2.Vout.n5 GND 0.0407f
C5618 Nand_Gate_2.Vout.n6 GND 0.05921f
C5619 Nand_Gate_2.Vout.n7 GND 1.13762f
C5620 Nand_Gate_2.Vout.n8 GND 1.13762f
C5621 Nand_Gate_2.Vout.n9 GND 0.07886f
C5622 Nand_Gate_2.Vout.t2 GND 0.07612f
C5623 Nand_Gate_2.Vout.t0 GND 0.09059f
C5624 Nand_Gate_2.Vout.n10 GND 0.45787f
C5625 Nand_Gate_2.Vout.n11 GND 0.23199f
C5626 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 GND 0.36784f
C5627 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 GND 0.10746f
C5628 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 GND 0.04662f
C5629 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 GND 0.205f
C5630 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 GND 0.1838f
C5631 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 GND 0.04989f
C5632 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 GND 0.31407f
C5633 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 GND 0.05094f
C5634 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 GND 0.04989f
C5635 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 GND 0.28374f
C5636 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 GND 0.09258f
C5637 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 GND 0.01095f
C5638 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 GND 0.01378f
C5639 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 GND 0.36785f
C5640 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 GND 0.38072f
C5641 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 GND 0.19125f
C5642 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 GND 0.18752f
C5643 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 GND 0.10934f
C5644 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 GND 0.0518f
C5645 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 GND 0.04798f
C5646 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 GND 0.22815f
C5647 CDAC8_0.switch_1.Z.t3 GND 0.0253f
C5648 CDAC8_0.switch_1.Z.t1 GND 0.02525f
C5649 CDAC8_0.switch_1.Z.n0 GND 0.05629f
C5650 CDAC8_0.switch_1.Z.n1 GND 0.01036f
C5651 CDAC8_0.switch_1.Z.t4 GND 5.82511f
C5652 CDAC8_0.switch_1.Z.n2 GND 0.11275f
C5653 CDAC8_0.switch_1.Z.n3 GND 0.02706f
C5654 CDAC8_0.switch_1.Z.t2 GND 0.02612f
C5655 CDAC8_0.switch_1.Z.t0 GND 0.02612f
C5656 CDAC8_0.switch_1.Z.n4 GND 0.09382f
C5657 CDAC8_0.switch_1.Z.n5 GND 0.28853f
C5658 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 GND 0.46931f
C5659 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 GND 0.1371f
C5660 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 GND 0.05949f
C5661 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 GND 0.06121f
C5662 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 GND 0.29108f
C5663 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 GND 0.06609f
C5664 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 GND 0.46933f
C5665 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 GND 0.48575f
C5666 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 GND 0.244f
C5667 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 GND 0.23925f
C5668 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 GND 0.13951f
C5669 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 GND 0.01758f
C5670 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 GND 0.01397f
C5671 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 GND 0.06499f
C5672 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 GND 0.06366f
C5673 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 GND 0.36201f
C5674 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 GND 0.11813f
C5675 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 GND 0.06366f
C5676 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 GND 0.40071f
C5677 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 GND 0.23451f
C5678 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 GND 0.26155f
C5679 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 GND 0.45666f
C5680 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 GND 0.47347f
C5681 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 GND 0.05122f
C5682 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 GND 0.05969f
C5683 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 GND 0.15961f
C5684 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 GND 0.12257f
C5685 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 GND 0.23742f
C5686 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 GND 0.45664f
C5687 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 GND 0.1334f
C5688 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 GND 0.05705f
C5689 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 GND 0.10533f
C5690 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 GND 0.18236f
C5691 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 GND 0.13574f
C5692 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 GND 0.06431f
C5693 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 GND 0.16533f
C5694 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 GND 0.06323f
C5695 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 GND 0.06194f
C5696 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 GND 0.35224f
C5697 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 GND 0.11629f
C5698 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 GND 0.06194f
C5699 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 GND 0.39067f
C5700 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 GND 0.22727f
C5701 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 GND 0.06839f
C5702 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 GND 0.36784f
C5703 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 GND 0.10746f
C5704 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 GND 0.04662f
C5705 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 GND 0.205f
C5706 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 GND 0.1838f
C5707 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 GND 0.04989f
C5708 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 GND 0.31407f
C5709 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 GND 0.05094f
C5710 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 GND 0.04989f
C5711 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 GND 0.28374f
C5712 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 GND 0.09441f
C5713 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 GND 0.01506f
C5714 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 GND 0.01378f
C5715 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 GND 0.36785f
C5716 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 GND 0.38072f
C5717 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 GND 0.19125f
C5718 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 GND 0.18752f
C5719 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 GND 0.10934f
C5720 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 GND 0.0518f
C5721 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 GND 0.04798f
C5722 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 GND 0.22815f
C5723 Q1.t8 GND 0.11808f
C5724 Q1.n0 GND 0.03449f
C5725 Q1.n1 GND 0.01497f
C5726 Q1.n2 GND 0.06581f
C5727 Q1.t4 GND 0.05417f
C5728 Q1.t3 GND 0.0154f
C5729 Q1.n3 GND 0.07553f
C5730 Q1.n4 GND 0.01853f
C5731 Q1.t1 GND 0.01635f
C5732 Q1.t0 GND 0.01602f
C5733 Q1.n5 GND 0.09108f
C5734 Q1.n6 GND 0.03031f
C5735 Q1.t2 GND 0.01602f
C5736 Q1.n7 GND 0.02467f
C5737 Q1.n8 GND 0.04119f
C5738 Q1.n9 GND 0.01949f
C5739 Q1.n11 GND 0.03785f
C5740 Q1.n12 GND 5.26881f
C5741 Q1.t7 GND 0.06149f
C5742 Q1.t6 GND 0.11839f
C5743 Q1.t9 GND 0.06149f
C5744 Q1.n13 GND 0.09578f
C5745 Q1.n14 GND 0.09633f
C5746 Q1.t5 GND 0.10524f
C5747 Q1.n15 GND 1.21138f
C5748 Nand_Gate_7.B.t5 GND 0.74634f
C5749 Nand_Gate_7.B.n0 GND 0.21803f
C5750 Nand_Gate_7.B.n1 GND 0.0946f
C5751 Nand_Gate_7.B.n2 GND 0.41594f
C5752 Nand_Gate_7.B.t15 GND 0.34714f
C5753 Nand_Gate_7.B.n3 GND 0.1089f
C5754 Nand_Gate_7.B.n4 GND 0.27612f
C5755 Nand_Gate_7.B.t1 GND 0.10123f
C5756 Nand_Gate_7.B.n5 GND 0.15594f
C5757 Nand_Gate_7.B.t2 GND 0.10335f
C5758 Nand_Gate_7.B.t3 GND 0.10123f
C5759 Nand_Gate_7.B.n6 GND 0.57571f
C5760 Nand_Gate_7.B.n7 GND 0.19155f
C5761 Nand_Gate_7.B.n8 GND 0.06954f
C5762 Nand_Gate_7.B.n9 GND 0.1212f
C5763 Nand_Gate_7.B.t10 GND 0.74637f
C5764 Nand_Gate_7.B.n10 GND 0.73349f
C5765 Nand_Gate_7.B.n11 GND 0.08017f
C5766 Nand_Gate_7.B.t14 GND 0.38804f
C5767 Nand_Gate_7.B.n12 GND 0.11178f
C5768 Nand_Gate_7.B.n13 GND 0.0479f
C5769 Nand_Gate_7.B.n14 GND 0.08976f
C5770 Nand_Gate_7.B.n15 GND 0.11295f
C5771 Nand_Gate_7.B.t13 GND 0.74637f
C5772 Nand_Gate_7.B.n16 GND 0.73349f
C5773 Nand_Gate_7.B.n17 GND 0.08017f
C5774 Nand_Gate_7.B.t11 GND 0.38804f
C5775 Nand_Gate_7.B.n18 GND 0.11178f
C5776 Nand_Gate_7.B.n19 GND 0.0479f
C5777 Nand_Gate_7.B.n20 GND 0.08976f
C5778 Nand_Gate_7.B.n21 GND 0.01346f
C5779 Nand_Gate_7.B.n22 GND 0.33743f
C5780 Nand_Gate_7.B.n23 GND 0.09223f
C5781 Nand_Gate_7.B.n24 GND 0.24541f
C5782 Nand_Gate_7.B.t12 GND 0.74637f
C5783 Nand_Gate_7.B.n25 GND 0.75163f
C5784 Nand_Gate_7.B.n26 GND 0.08017f
C5785 Nand_Gate_7.B.t17 GND 0.38804f
C5786 Nand_Gate_7.B.n27 GND 0.11178f
C5787 Nand_Gate_7.B.n28 GND 0.02977f
C5788 Nand_Gate_7.B.n29 GND 0.04639f
C5789 Nand_Gate_7.B.n30 GND 0.46286f
C5790 Nand_Gate_7.B.t6 GND 0.74637f
C5791 Nand_Gate_7.B.n31 GND 0.75163f
C5792 Nand_Gate_7.B.n32 GND 0.08017f
C5793 Nand_Gate_7.B.t7 GND 0.38804f
C5794 Nand_Gate_7.B.n33 GND 0.11178f
C5795 Nand_Gate_7.B.n34 GND 0.02977f
C5796 Nand_Gate_7.B.n35 GND 0.04639f
C5797 Nand_Gate_7.B.n36 GND 0.01346f
C5798 Nand_Gate_7.B.n37 GND 1.20187f
C5799 Nand_Gate_7.B.n38 GND 0.49755f
C5800 Nand_Gate_7.B.n39 GND 0.20758f
C5801 Nand_Gate_7.B.t4 GND 0.74634f
C5802 Nand_Gate_7.B.n40 GND 0.21803f
C5803 Nand_Gate_7.B.n41 GND 0.0946f
C5804 Nand_Gate_7.B.n42 GND 0.41594f
C5805 Nand_Gate_7.B.t8 GND 0.3471f
C5806 Nand_Gate_7.B.n43 GND 0.10713f
C5807 Nand_Gate_7.B.n44 GND 0.24887f
C5808 Nand_Gate_7.B.n45 GND 13.7262f
C5809 Nand_Gate_7.B.t16 GND 0.38806f
C5810 Nand_Gate_7.B.n46 GND 0.41458f
C5811 Nand_Gate_7.B.t9 GND 0.74634f
C5812 Nand_Gate_7.B.n47 GND 1.69885f
C5813 Nand_Gate_7.B.n48 GND 16.1408f
C5814 Nand_Gate_7.B.n49 GND 0.12649f
C5815 Nand_Gate_7.B.n50 GND 0.42321f
C5816 Nand_Gate_7.B.n51 GND 0.91499f
C5817 Nand_Gate_7.B.n52 GND 0.01373f
C5818 Nand_Gate_7.B.n53 GND 0.10511f
C5819 Nand_Gate_7.B.t0 GND 0.09735f
C5820 Nand_Gate_7.B.n54 GND 0.42392f
C5821 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 GND 0.36784f
C5822 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 GND 0.10746f
C5823 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 GND 0.04662f
C5824 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 GND 0.04798f
C5825 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 GND 0.22815f
C5826 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 GND 0.0518f
C5827 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 GND 0.36785f
C5828 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 GND 0.38072f
C5829 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 GND 0.19125f
C5830 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 GND 0.18752f
C5831 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 GND 0.10934f
C5832 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 GND 0.01378f
C5833 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 GND 0.01506f
C5834 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 GND 0.05094f
C5835 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 GND 0.04989f
C5836 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 GND 0.28374f
C5837 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 GND 0.09441f
C5838 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 GND 0.04989f
C5839 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 GND 0.31407f
C5840 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 GND 0.1838f
C5841 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 GND 0.205f
C5842 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 GND 0.45666f
C5843 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 GND 0.47347f
C5844 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 GND 0.05122f
C5845 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 GND 0.05969f
C5846 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 GND 0.15961f
C5847 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 GND 0.12257f
C5848 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 GND 0.23742f
C5849 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 GND 0.45664f
C5850 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 GND 0.1334f
C5851 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 GND 0.05705f
C5852 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 GND 0.10533f
C5853 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 GND 0.18236f
C5854 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 GND 0.13574f
C5855 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 GND 0.06431f
C5856 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 GND 0.16533f
C5857 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 GND 0.06323f
C5858 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 GND 0.06194f
C5859 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 GND 0.35224f
C5860 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 GND 0.11629f
C5861 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 GND 0.06194f
C5862 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 GND 0.39067f
C5863 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 GND 0.22727f
C5864 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 GND 0.06839f
C5865 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 GND 0.07282f
C5866 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 GND 0.31709f
C5867 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 GND 0.07862f
C5868 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 GND 0.55828f
C5869 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 GND 0.54865f
C5870 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 GND 0.05997f
C5871 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 GND 0.29025f
C5872 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 GND 0.08361f
C5873 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 GND 0.03583f
C5874 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 GND 0.06714f
C5875 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 GND 0.15126f
C5876 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 GND 0.15126f
C5877 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 GND 0.09065f
C5878 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 GND 0.04578f
C5879 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 GND 0.07589f
C5880 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 GND 0.0773f
C5881 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 GND 0.07572f
C5882 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 GND 0.43063f
C5883 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 GND 0.24092f
C5884 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 GND 0.07037f
C5885 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 GND 0.16004f
C5886 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 GND 0.07725f
C5887 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 GND 0.2799f
C5888 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 GND 0.27418f
C5889 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 GND 0.05783f
C5890 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 GND 0.53832f
C5891 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 GND 0.15726f
C5892 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 GND 0.03913f
C5893 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 GND 0.05692f
C5894 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 GND 0.14585f
C5895 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 GND 0.14585f
C5896 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 GND 0.07581f
C5897 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 GND 0.07318f
C5898 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 GND 0.07454f
C5899 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 GND 0.07302f
C5900 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 GND 0.41525f
C5901 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 GND 0.23391f
C5902 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 GND 0.22303f
C5903 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 GND 0.07024f
C5904 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 GND 0.03989f
C5905 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 GND 0.07725f
C5906 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 GND 0.2799f
C5907 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 GND 0.27418f
C5908 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 GND 0.05783f
C5909 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 GND 0.53832f
C5910 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 GND 0.15726f
C5911 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 GND 0.03913f
C5912 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 GND 0.05692f
C5913 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 GND 0.14585f
C5914 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 GND 0.14585f
C5915 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 GND 0.07581f
C5916 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 GND 0.07318f
C5917 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 GND 0.07454f
C5918 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 GND 0.07302f
C5919 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 GND 0.41525f
C5920 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 GND 0.23391f
C5921 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 GND 0.22303f
C5922 D_FlipFlop_0.3-input-nand_2.C.t6 GND 0.3425f
C5923 D_FlipFlop_0.3-input-nand_2.C.n0 GND 0.3551f
C5924 D_FlipFlop_0.3-input-nand_2.C.n1 GND 0.03842f
C5925 D_FlipFlop_0.3-input-nand_2.C.t1 GND 0.04477f
C5926 D_FlipFlop_0.3-input-nand_2.C.n2 GND 0.11971f
C5927 D_FlipFlop_0.3-input-nand_2.C.n3 GND 0.09193f
C5928 D_FlipFlop_0.3-input-nand_2.C.t4 GND 0.17806f
C5929 D_FlipFlop_0.3-input-nand_2.C.t5 GND 0.34248f
C5930 D_FlipFlop_0.3-input-nand_2.C.n4 GND 0.10005f
C5931 D_FlipFlop_0.3-input-nand_2.C.n5 GND 0.04279f
C5932 D_FlipFlop_0.3-input-nand_2.C.n6 GND 0.079f
C5933 D_FlipFlop_0.3-input-nand_2.C.n7 GND 0.13677f
C5934 D_FlipFlop_0.3-input-nand_2.C.n8 GND 0.10181f
C5935 D_FlipFlop_0.3-input-nand_2.C.n9 GND 0.04823f
C5936 D_FlipFlop_0.3-input-nand_2.C.n10 GND 0.124f
C5937 D_FlipFlop_0.3-input-nand_2.C.t3 GND 0.04742f
C5938 D_FlipFlop_0.3-input-nand_2.C.t0 GND 0.04645f
C5939 D_FlipFlop_0.3-input-nand_2.C.n11 GND 0.26418f
C5940 D_FlipFlop_0.3-input-nand_2.C.n12 GND 0.08722f
C5941 D_FlipFlop_0.3-input-nand_2.C.t2 GND 0.04645f
C5942 D_FlipFlop_0.3-input-nand_2.C.n13 GND 0.293f
C5943 D_FlipFlop_0.3-input-nand_2.C.t7 GND 0.17045f
C5944 D_FlipFlop_0.3-input-nand_2.C.n14 GND 0.05129f
C5945 D_FlipFlop_3.3-input-nand_2.C.t7 GND 0.3425f
C5946 D_FlipFlop_3.3-input-nand_2.C.n0 GND 0.3551f
C5947 D_FlipFlop_3.3-input-nand_2.C.n1 GND 0.03842f
C5948 D_FlipFlop_3.3-input-nand_2.C.t2 GND 0.04477f
C5949 D_FlipFlop_3.3-input-nand_2.C.n2 GND 0.11971f
C5950 D_FlipFlop_3.3-input-nand_2.C.n3 GND 0.09193f
C5951 D_FlipFlop_3.3-input-nand_2.C.t5 GND 0.17806f
C5952 D_FlipFlop_3.3-input-nand_2.C.t6 GND 0.34248f
C5953 D_FlipFlop_3.3-input-nand_2.C.n4 GND 0.10005f
C5954 D_FlipFlop_3.3-input-nand_2.C.n5 GND 0.04279f
C5955 D_FlipFlop_3.3-input-nand_2.C.n6 GND 0.079f
C5956 D_FlipFlop_3.3-input-nand_2.C.n7 GND 0.13677f
C5957 D_FlipFlop_3.3-input-nand_2.C.n8 GND 0.10181f
C5958 D_FlipFlop_3.3-input-nand_2.C.n9 GND 0.04823f
C5959 D_FlipFlop_3.3-input-nand_2.C.n10 GND 0.124f
C5960 D_FlipFlop_3.3-input-nand_2.C.t0 GND 0.04742f
C5961 D_FlipFlop_3.3-input-nand_2.C.t3 GND 0.04645f
C5962 D_FlipFlop_3.3-input-nand_2.C.n11 GND 0.26418f
C5963 D_FlipFlop_3.3-input-nand_2.C.n12 GND 0.08722f
C5964 D_FlipFlop_3.3-input-nand_2.C.t1 GND 0.04645f
C5965 D_FlipFlop_3.3-input-nand_2.C.n13 GND 0.293f
C5966 D_FlipFlop_3.3-input-nand_2.C.t4 GND 0.17045f
C5967 D_FlipFlop_3.3-input-nand_2.C.n14 GND 0.05129f
C5968 D_FlipFlop_3.3-input-nand_2.Vout.t4 GND 0.35515f
C5969 D_FlipFlop_3.3-input-nand_2.Vout.n0 GND 0.10375f
C5970 D_FlipFlop_3.3-input-nand_2.Vout.n1 GND 0.04502f
C5971 D_FlipFlop_3.3-input-nand_2.Vout.t3 GND 0.04632f
C5972 D_FlipFlop_3.3-input-nand_2.Vout.n2 GND 0.22028f
C5973 D_FlipFlop_3.3-input-nand_2.Vout.n3 GND 0.05002f
C5974 D_FlipFlop_3.3-input-nand_2.Vout.t7 GND 0.35517f
C5975 D_FlipFlop_3.3-input-nand_2.Vout.n4 GND 0.36759f
C5976 D_FlipFlop_3.3-input-nand_2.Vout.t5 GND 0.18465f
C5977 D_FlipFlop_3.3-input-nand_2.Vout.n5 GND 0.18106f
C5978 D_FlipFlop_3.3-input-nand_2.Vout.n6 GND 0.10557f
C5979 D_FlipFlop_3.3-input-nand_2.Vout.n7 GND 0.01331f
C5980 D_FlipFlop_3.3-input-nand_2.Vout.n8 GND 0.01454f
C5981 D_FlipFlop_3.3-input-nand_2.Vout.t0 GND 0.04918f
C5982 D_FlipFlop_3.3-input-nand_2.Vout.t1 GND 0.04817f
C5983 D_FlipFlop_3.3-input-nand_2.Vout.n9 GND 0.27396f
C5984 D_FlipFlop_3.3-input-nand_2.Vout.n10 GND 0.09115f
C5985 D_FlipFlop_3.3-input-nand_2.Vout.t2 GND 0.04817f
C5986 D_FlipFlop_3.3-input-nand_2.Vout.n11 GND 0.30324f
C5987 D_FlipFlop_3.3-input-nand_2.Vout.t6 GND 0.17747f
C5988 D_FlipFlop_3.3-input-nand_2.Vout.n12 GND 0.19793f
C5989 Nand_Gate_4.B.t9 GND 0.65284f
C5990 Nand_Gate_4.B.n0 GND 0.19071f
C5991 Nand_Gate_4.B.n1 GND 0.08275f
C5992 Nand_Gate_4.B.n2 GND 0.36383f
C5993 Nand_Gate_4.B.t17 GND 0.30365f
C5994 Nand_Gate_4.B.n3 GND 0.09526f
C5995 Nand_Gate_4.B.t1 GND 0.08515f
C5996 Nand_Gate_4.B.n4 GND 0.37081f
C5997 Nand_Gate_4.B.n5 GND 0.09194f
C5998 Nand_Gate_4.B.t13 GND 0.65287f
C5999 Nand_Gate_4.B.n6 GND 0.6416f
C6000 Nand_Gate_4.B.n7 GND 0.07013f
C6001 Nand_Gate_4.B.t16 GND 0.33943f
C6002 Nand_Gate_4.B.n8 GND 0.09778f
C6003 Nand_Gate_4.B.n9 GND 0.0419f
C6004 Nand_Gate_4.B.n10 GND 0.07851f
C6005 Nand_Gate_4.B.n11 GND 0.0988f
C6006 Nand_Gate_4.B.t14 GND 0.65287f
C6007 Nand_Gate_4.B.n12 GND 0.6416f
C6008 Nand_Gate_4.B.n13 GND 0.07013f
C6009 Nand_Gate_4.B.t6 GND 0.33943f
C6010 Nand_Gate_4.B.n14 GND 0.09778f
C6011 Nand_Gate_4.B.n15 GND 0.0419f
C6012 Nand_Gate_4.B.n16 GND 0.07851f
C6013 Nand_Gate_4.B.n17 GND 0.01177f
C6014 Nand_Gate_4.B.n18 GND 0.29516f
C6015 Nand_Gate_4.B.n19 GND 0.08068f
C6016 Nand_Gate_4.B.n20 GND 0.21466f
C6017 Nand_Gate_4.B.t5 GND 0.65287f
C6018 Nand_Gate_4.B.n21 GND 0.65747f
C6019 Nand_Gate_4.B.n22 GND 0.07013f
C6020 Nand_Gate_4.B.t11 GND 0.33943f
C6021 Nand_Gate_4.B.n23 GND 0.09778f
C6022 Nand_Gate_4.B.n24 GND 0.02604f
C6023 Nand_Gate_4.B.n25 GND 0.04058f
C6024 Nand_Gate_4.B.n26 GND 0.40488f
C6025 Nand_Gate_4.B.t12 GND 0.65287f
C6026 Nand_Gate_4.B.n27 GND 0.65747f
C6027 Nand_Gate_4.B.n28 GND 0.07013f
C6028 Nand_Gate_4.B.t4 GND 0.33943f
C6029 Nand_Gate_4.B.n29 GND 0.09778f
C6030 Nand_Gate_4.B.n30 GND 0.02604f
C6031 Nand_Gate_4.B.n31 GND 0.04058f
C6032 Nand_Gate_4.B.n32 GND 0.01177f
C6033 Nand_Gate_4.B.n33 GND 1.0513f
C6034 Nand_Gate_4.B.n34 GND 0.45039f
C6035 Nand_Gate_4.B.n35 GND 0.18158f
C6036 Nand_Gate_4.B.t15 GND 0.65284f
C6037 Nand_Gate_4.B.n36 GND 0.19071f
C6038 Nand_Gate_4.B.n37 GND 0.08275f
C6039 Nand_Gate_4.B.n38 GND 0.36383f
C6040 Nand_Gate_4.B.t7 GND 0.30362f
C6041 Nand_Gate_4.B.n39 GND 0.07854f
C6042 Nand_Gate_4.B.n40 GND 0.1833f
C6043 Nand_Gate_4.B.n41 GND 15.2571f
C6044 Nand_Gate_4.B.t10 GND 0.33944f
C6045 Nand_Gate_4.B.n42 GND 0.36264f
C6046 Nand_Gate_4.B.t8 GND 0.65284f
C6047 Nand_Gate_4.B.n43 GND 1.46118f
C6048 Nand_Gate_4.B.n44 GND 17.2191f
C6049 Nand_Gate_4.B.n45 GND 0.11064f
C6050 Nand_Gate_4.B.n46 GND 0.37019f
C6051 Nand_Gate_4.B.n47 GND 0.80036f
C6052 Nand_Gate_4.B.n48 GND 0.01201f
C6053 Nand_Gate_4.B.n49 GND 0.10601f
C6054 Nand_Gate_4.B.n50 GND 0.06083f
C6055 Nand_Gate_4.B.t2 GND 0.0904f
C6056 Nand_Gate_4.B.t3 GND 0.08855f
C6057 Nand_Gate_4.B.n51 GND 0.50358f
C6058 Nand_Gate_4.B.n52 GND 0.16755f
C6059 Nand_Gate_4.B.t0 GND 0.08855f
C6060 Nand_Gate_4.B.n53 GND 0.1364f
C6061 Nand_Gate_4.B.n54 GND 0.24153f
C6062 a_138533_35417.t1 GND 2.87848f
C6063 a_138533_35417.t2 GND 2.70178f
C6064 a_138533_35417.t3 GND 4.49528f
C6065 a_138533_35417.n0 GND 1.98132f
C6066 a_138533_35417.n1 GND 1.65328f
C6067 a_138533_35417.t0 GND 0.88985f
C6068 Nand_Gate_5.A.t16 GND 0.37676f
C6069 Nand_Gate_5.A.n0 GND 0.11006f
C6070 Nand_Gate_5.A.n1 GND 0.04775f
C6071 Nand_Gate_5.A.n2 GND 0.20997f
C6072 Nand_Gate_5.A.t7 GND 0.17524f
C6073 Nand_Gate_5.A.n3 GND 0.05498f
C6074 Nand_Gate_5.A.t2 GND 0.04914f
C6075 Nand_Gate_5.A.n4 GND 0.214f
C6076 Nand_Gate_5.A.n5 GND 0.05306f
C6077 Nand_Gate_5.A.t8 GND 0.37678f
C6078 Nand_Gate_5.A.n6 GND 0.37028f
C6079 Nand_Gate_5.A.n7 GND 0.04047f
C6080 Nand_Gate_5.A.t12 GND 0.19589f
C6081 Nand_Gate_5.A.n8 GND 0.05643f
C6082 Nand_Gate_5.A.n9 GND 0.02418f
C6083 Nand_Gate_5.A.n10 GND 0.04531f
C6084 Nand_Gate_5.A.n11 GND 0.05702f
C6085 Nand_Gate_5.A.t13 GND 0.37678f
C6086 Nand_Gate_5.A.n12 GND 0.37028f
C6087 Nand_Gate_5.A.n13 GND 0.04047f
C6088 Nand_Gate_5.A.t11 GND 0.19589f
C6089 Nand_Gate_5.A.n14 GND 0.05643f
C6090 Nand_Gate_5.A.n15 GND 0.02418f
C6091 Nand_Gate_5.A.n16 GND 0.04531f
C6092 Nand_Gate_5.A.n18 GND 0.17097f
C6093 Nand_Gate_5.A.n19 GND 0.47611f
C6094 Nand_Gate_5.A.n20 GND 0.21364f
C6095 Nand_Gate_5.A.t15 GND 0.37678f
C6096 Nand_Gate_5.A.n21 GND 0.37943f
C6097 Nand_Gate_5.A.n22 GND 0.04047f
C6098 Nand_Gate_5.A.t5 GND 0.19589f
C6099 Nand_Gate_5.A.n23 GND 0.05643f
C6100 Nand_Gate_5.A.n24 GND 0.01503f
C6101 Nand_Gate_5.A.n25 GND 0.02342f
C6102 Nand_Gate_5.A.n26 GND 0.23366f
C6103 Nand_Gate_5.A.t6 GND 0.37678f
C6104 Nand_Gate_5.A.n27 GND 0.37943f
C6105 Nand_Gate_5.A.n28 GND 0.04047f
C6106 Nand_Gate_5.A.t14 GND 0.19589f
C6107 Nand_Gate_5.A.n29 GND 0.05643f
C6108 Nand_Gate_5.A.n30 GND 0.01503f
C6109 Nand_Gate_5.A.n31 GND 0.02342f
C6110 Nand_Gate_5.A.n33 GND 0.60672f
C6111 Nand_Gate_5.A.n34 GND 0.28162f
C6112 Nand_Gate_5.A.n35 GND 0.10479f
C6113 Nand_Gate_5.A.t10 GND 0.37676f
C6114 Nand_Gate_5.A.n36 GND 0.11006f
C6115 Nand_Gate_5.A.n37 GND 0.04775f
C6116 Nand_Gate_5.A.n38 GND 0.20997f
C6117 Nand_Gate_5.A.t17 GND 0.17522f
C6118 Nand_Gate_5.A.n39 GND 0.02363f
C6119 Nand_Gate_5.A.n40 GND 0.05662f
C6120 Nand_Gate_5.A.n41 GND 2.27298f
C6121 Nand_Gate_5.A.t9 GND 0.1959f
C6122 Nand_Gate_5.A.n42 GND 0.19189f
C6123 Nand_Gate_5.A.n43 GND 0.04047f
C6124 Nand_Gate_5.A.t4 GND 0.37676f
C6125 Nand_Gate_5.A.n44 GND 0.11006f
C6126 Nand_Gate_5.A.n45 GND 0.02739f
C6127 Nand_Gate_5.A.n46 GND 0.03984f
C6128 Nand_Gate_5.A.n47 GND 0.05866f
C6129 Nand_Gate_5.A.n48 GND 3.09538f
C6130 Nand_Gate_5.A.n49 GND 0.20732f
C6131 Nand_Gate_5.A.n50 GND 0.0606f
C6132 Nand_Gate_5.A.n51 GND 0.0223f
C6133 Nand_Gate_5.A.n53 GND 0.06118f
C6134 Nand_Gate_5.A.n54 GND 0.0309f
C6135 Nand_Gate_5.A.t1 GND 0.05217f
C6136 Nand_Gate_5.A.t0 GND 0.0511f
C6137 Nand_Gate_5.A.n55 GND 0.29062f
C6138 Nand_Gate_5.A.n56 GND 0.09483f
C6139 Nand_Gate_5.A.t3 GND 0.0511f
C6140 Nand_Gate_5.A.n57 GND 0.07872f
C6141 Nand_Gate_5.A.n58 GND 0.13939f
C6142 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 GND 0.05201f
C6143 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 GND 0.22649f
C6144 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 GND 0.05616f
C6145 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 GND 0.39877f
C6146 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 GND 0.39189f
C6147 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 GND 0.04283f
C6148 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 GND 0.20732f
C6149 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 GND 0.05972f
C6150 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 GND 0.02559f
C6151 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 GND 0.04796f
C6152 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 GND 0.10804f
C6153 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 GND 0.10804f
C6154 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 GND 0.06475f
C6155 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 GND 0.05421f
C6156 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 GND 0.05522f
C6157 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 GND 0.05409f
C6158 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 GND 0.30759f
C6159 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 GND 0.17406f
C6160 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 GND 0.03715f
C6161 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 GND 0.0608f
C6162 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 GND 0.13827f
C6163 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 GND 0.06674f
C6164 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 GND 0.24183f
C6165 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 GND 0.23689f
C6166 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 GND 0.04996f
C6167 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 GND 0.46511f
C6168 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 GND 0.13587f
C6169 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 GND 0.03381f
C6170 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 GND 0.04918f
C6171 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 GND 0.12602f
C6172 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 GND 0.12602f
C6173 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 GND 0.0655f
C6174 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 GND 0.06323f
C6175 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 GND 0.07525f
C6176 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 GND 0.38033f
C6177 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 GND 0.1927f
C6178 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 GND 0.04607f
C6179 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 GND 0.10477f
C6180 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 GND 0.05057f
C6181 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 GND 0.35243f
C6182 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 GND 0.3654f
C6183 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 GND 0.03953f
C6184 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 GND 0.05278f
C6185 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 GND 0.27708f
C6186 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 GND 0.27709f
C6187 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 GND 0.17949f
C6188 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 GND 0.03786f
C6189 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 GND 0.35241f
C6190 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 GND 0.10295f
C6191 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 GND 0.02562f
C6192 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 GND 0.03726f
C6193 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 GND 0.09548f
C6194 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 GND 0.09548f
C6195 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 GND 0.04963f
C6196 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 GND 0.04792f
C6197 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 GND 0.28399f
C6198 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 GND 0.04798f
C6199 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 GND 0.02725f
C6200 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 GND 0.05277f
C6201 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 GND 0.36775f
C6202 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 GND 0.38129f
C6203 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 GND 0.04125f
C6204 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 GND 0.05508f
C6205 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 GND 0.28913f
C6206 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 GND 0.28914f
C6207 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 GND 0.1873f
C6208 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 GND 0.0395f
C6209 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 GND 0.36774f
C6210 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 GND 0.10743f
C6211 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 GND 0.02673f
C6212 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 GND 0.03888f
C6213 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 GND 0.09964f
C6214 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 GND 0.09964f
C6215 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 GND 0.05179f
C6216 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 GND 0.05f
C6217 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 GND 0.29633f
C6218 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 GND 0.06358f
C6219 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 GND 0.03611f
C6220 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 GND 0.06992f
C6221 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 GND 0.25335f
C6222 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 GND 0.24817f
C6223 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 GND 0.05234f
C6224 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 GND 0.48726f
C6225 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 GND 0.14234f
C6226 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 GND 0.03542f
C6227 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 GND 0.05152f
C6228 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 GND 0.13202f
C6229 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 GND 0.13202f
C6230 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 GND 0.06862f
C6231 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 GND 0.06624f
C6232 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 GND 0.07883f
C6233 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 GND 0.39844f
C6234 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 GND 0.20187f
C6235 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 GND 0.05201f
C6236 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 GND 0.22649f
C6237 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 GND 0.05616f
C6238 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 GND 0.39877f
C6239 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 GND 0.39189f
C6240 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 GND 0.04283f
C6241 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 GND 0.20732f
C6242 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 GND 0.05972f
C6243 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 GND 0.02559f
C6244 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 GND 0.04796f
C6245 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 GND 0.10804f
C6246 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 GND 0.10804f
C6247 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 GND 0.06475f
C6248 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 GND 0.05421f
C6249 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 GND 0.05522f
C6250 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 GND 0.05409f
C6251 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 GND 0.30759f
C6252 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 GND 0.17406f
C6253 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 GND 0.03715f
C6254 Nand_Gate_6.B.t16 GND 0.66019f
C6255 Nand_Gate_6.B.n0 GND 0.19286f
C6256 Nand_Gate_6.B.n1 GND 0.08368f
C6257 Nand_Gate_6.B.n2 GND 0.36793f
C6258 Nand_Gate_6.B.t5 GND 0.30707f
C6259 Nand_Gate_6.B.n3 GND 0.09633f
C6260 Nand_Gate_6.B.t2 GND 0.08611f
C6261 Nand_Gate_6.B.n4 GND 0.37499f
C6262 Nand_Gate_6.B.n5 GND 0.09297f
C6263 Nand_Gate_6.B.t10 GND 0.66022f
C6264 Nand_Gate_6.B.n6 GND 0.64883f
C6265 Nand_Gate_6.B.n7 GND 0.07092f
C6266 Nand_Gate_6.B.t17 GND 0.34325f
C6267 Nand_Gate_6.B.n8 GND 0.09888f
C6268 Nand_Gate_6.B.n9 GND 0.04237f
C6269 Nand_Gate_6.B.n10 GND 0.0794f
C6270 Nand_Gate_6.B.n11 GND 0.09991f
C6271 Nand_Gate_6.B.t15 GND 0.66022f
C6272 Nand_Gate_6.B.n12 GND 0.64883f
C6273 Nand_Gate_6.B.n13 GND 0.07092f
C6274 Nand_Gate_6.B.t11 GND 0.34325f
C6275 Nand_Gate_6.B.n14 GND 0.09888f
C6276 Nand_Gate_6.B.n15 GND 0.04237f
C6277 Nand_Gate_6.B.n16 GND 0.0794f
C6278 Nand_Gate_6.B.n17 GND 0.0119f
C6279 Nand_Gate_6.B.n18 GND 0.29848f
C6280 Nand_Gate_6.B.n19 GND 0.08159f
C6281 Nand_Gate_6.B.n20 GND 0.21708f
C6282 Nand_Gate_6.B.t6 GND 0.66022f
C6283 Nand_Gate_6.B.n21 GND 0.66487f
C6284 Nand_Gate_6.B.n22 GND 0.07092f
C6285 Nand_Gate_6.B.t12 GND 0.34325f
C6286 Nand_Gate_6.B.n23 GND 0.09888f
C6287 Nand_Gate_6.B.n24 GND 0.02633f
C6288 Nand_Gate_6.B.n25 GND 0.04104f
C6289 Nand_Gate_6.B.n26 GND 0.40943f
C6290 Nand_Gate_6.B.t13 GND 0.66022f
C6291 Nand_Gate_6.B.n27 GND 0.66487f
C6292 Nand_Gate_6.B.n28 GND 0.07092f
C6293 Nand_Gate_6.B.t7 GND 0.34325f
C6294 Nand_Gate_6.B.n29 GND 0.09888f
C6295 Nand_Gate_6.B.n30 GND 0.02633f
C6296 Nand_Gate_6.B.n31 GND 0.04104f
C6297 Nand_Gate_6.B.n32 GND 0.0119f
C6298 Nand_Gate_6.B.n33 GND 1.06314f
C6299 Nand_Gate_6.B.n34 GND 0.43942f
C6300 Nand_Gate_6.B.n35 GND 0.18362f
C6301 Nand_Gate_6.B.t4 GND 0.66019f
C6302 Nand_Gate_6.B.n36 GND 0.19286f
C6303 Nand_Gate_6.B.n37 GND 0.08368f
C6304 Nand_Gate_6.B.n38 GND 0.36793f
C6305 Nand_Gate_6.B.t9 GND 0.30704f
C6306 Nand_Gate_6.B.n39 GND 0.09546f
C6307 Nand_Gate_6.B.n40 GND 0.22172f
C6308 Nand_Gate_6.B.n41 GND 8.79656f
C6309 Nand_Gate_6.B.t8 GND 0.34326f
C6310 Nand_Gate_6.B.n42 GND 0.36672f
C6311 Nand_Gate_6.B.t14 GND 0.66019f
C6312 Nand_Gate_6.B.n43 GND 1.50275f
C6313 Nand_Gate_6.B.n44 GND 11.1675f
C6314 Nand_Gate_6.B.n45 GND 0.11189f
C6315 Nand_Gate_6.B.n46 GND 0.37436f
C6316 Nand_Gate_6.B.n47 GND 0.80937f
C6317 Nand_Gate_6.B.n48 GND 0.01215f
C6318 Nand_Gate_6.B.n49 GND 0.10721f
C6319 Nand_Gate_6.B.n50 GND 0.06151f
C6320 Nand_Gate_6.B.t0 GND 0.09142f
C6321 Nand_Gate_6.B.t1 GND 0.08955f
C6322 Nand_Gate_6.B.n51 GND 0.50925f
C6323 Nand_Gate_6.B.n52 GND 0.16944f
C6324 Nand_Gate_6.B.t3 GND 0.08955f
C6325 Nand_Gate_6.B.n53 GND 0.13794f
C6326 Nand_Gate_6.B.n54 GND 0.24424f
C6327 Nand_Gate_5.Vout.t1 GND 0.07306f
C6328 Nand_Gate_5.Vout.n0 GND 0.0415f
C6329 Nand_Gate_5.Vout.n1 GND 0.08035f
C6330 Nand_Gate_5.Vout.t3 GND 0.29114f
C6331 Nand_Gate_5.Vout.n2 GND 0.28519f
C6332 Nand_Gate_5.Vout.n3 GND 0.06015f
C6333 Nand_Gate_5.Vout.t4 GND 0.55994f
C6334 Nand_Gate_5.Vout.n4 GND 0.16357f
C6335 Nand_Gate_5.Vout.n5 GND 0.0407f
C6336 Nand_Gate_5.Vout.n6 GND 0.05921f
C6337 Nand_Gate_5.Vout.n7 GND 1.13762f
C6338 Nand_Gate_5.Vout.n8 GND 1.13762f
C6339 Nand_Gate_5.Vout.n9 GND 0.07886f
C6340 Nand_Gate_5.Vout.t2 GND 0.07612f
C6341 Nand_Gate_5.Vout.t0 GND 0.09059f
C6342 Nand_Gate_5.Vout.n10 GND 0.45787f
C6343 Nand_Gate_5.Vout.n11 GND 0.23199f
C6344 CDAC8_0.switch_5.Z.t2 GND 0.03054f
C6345 CDAC8_0.switch_5.Z.t1 GND 0.03054f
C6346 CDAC8_0.switch_5.Z.n0 GND 0.11035f
C6347 CDAC8_0.switch_5.Z.n1 GND 0.254f
C6348 CDAC8_0.switch_5.Z.t3 GND 0.03207f
C6349 CDAC8_0.switch_5.Z.t6 GND 5.60901f
C6350 CDAC8_0.switch_5.Z.n2 GND 1.99837f
C6351 CDAC8_0.switch_5.Z.t5 GND 5.4744f
C6352 CDAC8_0.switch_5.Z.t9 GND 5.4744f
C6353 CDAC8_0.switch_5.Z.t7 GND 5.39614f
C6354 CDAC8_0.switch_5.Z.n3 GND 1.42238f
C6355 CDAC8_0.switch_5.Z.t4 GND 5.39614f
C6356 CDAC8_0.switch_5.Z.n4 GND 1.67019f
C6357 CDAC8_0.switch_5.Z.n5 GND 2.09417f
C6358 CDAC8_0.switch_5.Z.n6 GND 2.09417f
C6359 CDAC8_0.switch_5.Z.t8 GND 5.39614f
C6360 CDAC8_0.switch_5.Z.n7 GND 1.67019f
C6361 CDAC8_0.switch_5.Z.t11 GND 5.39614f
C6362 CDAC8_0.switch_5.Z.n8 GND 1.42238f
C6363 CDAC8_0.switch_5.Z.t10 GND 5.60901f
C6364 CDAC8_0.switch_5.Z.n9 GND 1.95831f
C6365 CDAC8_0.switch_5.Z.n10 GND 0.46579f
C6366 CDAC8_0.switch_5.Z.n11 GND 0.10945f
C6367 CDAC8_0.switch_5.Z.t0 GND 0.03205f
C6368 Q3.t8 GND 0.11803f
C6369 Q3.n0 GND 0.03448f
C6370 Q3.n1 GND 0.01496f
C6371 Q3.n2 GND 0.06578f
C6372 Q3.t5 GND 0.05414f
C6373 Q3.t2 GND 0.0154f
C6374 Q3.n3 GND 0.0755f
C6375 Q3.n4 GND 0.01853f
C6376 Q3.t1 GND 0.01634f
C6377 Q3.t0 GND 0.01601f
C6378 Q3.n5 GND 0.09105f
C6379 Q3.n6 GND 0.03029f
C6380 Q3.t3 GND 0.01601f
C6381 Q3.n7 GND 0.02466f
C6382 Q3.n8 GND 0.04061f
C6383 Q3.n9 GND 0.02001f
C6384 Q3.n11 GND 0.03887f
C6385 Q3.n12 GND 5.74071f
C6386 Q3.t6 GND 0.06147f
C6387 Q3.t4 GND 0.11834f
C6388 Q3.t7 GND 0.06147f
C6389 Q3.n13 GND 0.09574f
C6390 Q3.n14 GND 0.09629f
C6391 Q3.t9 GND 0.1052f
C6392 Q3.n15 GND 1.21087f
C6393 CDAC8_0.switch_2.Z.t3 GND 0.03087f
C6394 CDAC8_0.switch_2.Z.t2 GND 0.02943f
C6395 CDAC8_0.switch_2.Z.t1 GND 0.02943f
C6396 CDAC8_0.switch_2.Z.n0 GND 0.10631f
C6397 CDAC8_0.switch_2.Z.n1 GND 0.24452f
C6398 CDAC8_0.switch_2.Z.n2 GND 0.03182f
C6399 CDAC8_0.switch_2.Z.t5 GND 6.50564f
C6400 CDAC8_0.switch_2.Z.t4 GND 6.4338f
C6401 CDAC8_0.switch_2.Z.n3 GND 1.02469f
C6402 CDAC8_0.switch_2.Z.n4 GND 0.01025f
C6403 CDAC8_0.switch_2.Z.t0 GND 0.03087f
C6404 CDAC8_0.switch_2.Z.n5 GND 0.12722f
C6405 Q6.t3 GND 0.01626f
C6406 Q6.n0 GND 0.07974f
C6407 Q6.n1 GND 0.01957f
C6408 Q6.t0 GND 0.01726f
C6409 Q6.t1 GND 0.01691f
C6410 Q6.n2 GND 0.09616f
C6411 Q6.n3 GND 0.03199f
C6412 Q6.t2 GND 0.01691f
C6413 Q6.n4 GND 0.02605f
C6414 Q6.n5 GND 0.0372f
C6415 Q6.n6 GND 0.0192f
C6416 Q6.t8 GND 0.12466f
C6417 Q6.n7 GND 0.03642f
C6418 Q6.n8 GND 0.0158f
C6419 Q6.n9 GND 0.06947f
C6420 Q6.t6 GND 0.05798f
C6421 Q6.n11 GND 0.01555f
C6422 Q6.n13 GND 3.34141f
C6423 Q6.t4 GND 0.12498f
C6424 Q6.t5 GND 0.12498f
C6425 Q6.t9 GND 0.06492f
C6426 Q6.n14 GND 0.10112f
C6427 Q6.n15 GND 0.1017f
C6428 Q6.t7 GND 0.05702f
C6429 Q6.n16 GND 1.27887f
C6430 D_FlipFlop_5.3-input-nand_2.C.t5 GND 0.3425f
C6431 D_FlipFlop_5.3-input-nand_2.C.n0 GND 0.3551f
C6432 D_FlipFlop_5.3-input-nand_2.C.n1 GND 0.03842f
C6433 D_FlipFlop_5.3-input-nand_2.C.n2 GND 0.05129f
C6434 D_FlipFlop_5.3-input-nand_2.C.t6 GND 0.17045f
C6435 D_FlipFlop_5.3-input-nand_2.C.t2 GND 0.04645f
C6436 D_FlipFlop_5.3-input-nand_2.C.n3 GND 0.293f
C6437 D_FlipFlop_5.3-input-nand_2.C.t1 GND 0.04742f
C6438 D_FlipFlop_5.3-input-nand_2.C.t3 GND 0.04645f
C6439 D_FlipFlop_5.3-input-nand_2.C.n4 GND 0.26418f
C6440 D_FlipFlop_5.3-input-nand_2.C.n5 GND 0.08722f
C6441 D_FlipFlop_5.3-input-nand_2.C.n6 GND 0.124f
C6442 D_FlipFlop_5.3-input-nand_2.C.n7 GND 0.04823f
C6443 D_FlipFlop_5.3-input-nand_2.C.t7 GND 0.17806f
C6444 D_FlipFlop_5.3-input-nand_2.C.t4 GND 0.34248f
C6445 D_FlipFlop_5.3-input-nand_2.C.n8 GND 0.10005f
C6446 D_FlipFlop_5.3-input-nand_2.C.n9 GND 0.04279f
C6447 D_FlipFlop_5.3-input-nand_2.C.n10 GND 0.079f
C6448 D_FlipFlop_5.3-input-nand_2.C.n11 GND 0.13677f
C6449 D_FlipFlop_5.3-input-nand_2.C.n12 GND 0.10181f
C6450 D_FlipFlop_5.3-input-nand_2.C.n13 GND 0.09193f
C6451 D_FlipFlop_5.3-input-nand_2.C.t0 GND 0.04477f
C6452 D_FlipFlop_5.3-input-nand_2.C.n14 GND 0.11971f
C6453 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 GND 0.36784f
C6454 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 GND 0.10746f
C6455 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 GND 0.04662f
C6456 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 GND 0.205f
C6457 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 GND 0.1838f
C6458 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 GND 0.04989f
C6459 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 GND 0.31407f
C6460 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 GND 0.05094f
C6461 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 GND 0.04989f
C6462 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 GND 0.28374f
C6463 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 GND 0.09258f
C6464 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 GND 0.01095f
C6465 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 GND 0.01378f
C6466 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 GND 0.36785f
C6467 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 GND 0.38072f
C6468 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 GND 0.19125f
C6469 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 GND 0.18752f
C6470 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 GND 0.10934f
C6471 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 GND 0.0518f
C6472 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 GND 0.04798f
C6473 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 GND 0.22815f
C6474 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 GND 0.04998f
C6475 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 GND 0.02839f
C6476 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 GND 0.05497f
C6477 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 GND 0.38308f
C6478 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 GND 0.39717f
C6479 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 GND 0.04297f
C6480 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 GND 0.05737f
C6481 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 GND 0.30118f
C6482 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 GND 0.30119f
C6483 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 GND 0.1951f
C6484 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 GND 0.04115f
C6485 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 GND 0.38306f
C6486 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 GND 0.1119f
C6487 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 GND 0.02784f
C6488 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 GND 0.0405f
C6489 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 GND 0.10379f
C6490 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 GND 0.10379f
C6491 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 GND 0.05395f
C6492 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 GND 0.05208f
C6493 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 GND 0.30868f
C6494 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 GND 0.45666f
C6495 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 GND 0.47347f
C6496 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 GND 0.05122f
C6497 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 GND 0.05969f
C6498 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 GND 0.15961f
C6499 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 GND 0.12257f
C6500 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 GND 0.23742f
C6501 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 GND 0.45664f
C6502 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 GND 0.1334f
C6503 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 GND 0.05705f
C6504 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 GND 0.10533f
C6505 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 GND 0.18236f
C6506 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 GND 0.13574f
C6507 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 GND 0.06431f
C6508 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 GND 0.16533f
C6509 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 GND 0.06323f
C6510 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 GND 0.06194f
C6511 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 GND 0.35224f
C6512 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 GND 0.11629f
C6513 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 GND 0.06194f
C6514 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 GND 0.39067f
C6515 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 GND 0.22727f
C6516 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 GND 0.06839f
C6517 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 GND 0.36784f
C6518 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 GND 0.10746f
C6519 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 GND 0.04662f
C6520 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 GND 0.205f
C6521 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 GND 0.1838f
C6522 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 GND 0.04989f
C6523 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 GND 0.31407f
C6524 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 GND 0.05094f
C6525 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 GND 0.04989f
C6526 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 GND 0.28374f
C6527 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 GND 0.09441f
C6528 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 GND 0.01506f
C6529 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 GND 0.01378f
C6530 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 GND 0.36785f
C6531 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 GND 0.38072f
C6532 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 GND 0.19125f
C6533 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 GND 0.18752f
C6534 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 GND 0.10934f
C6535 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 GND 0.0518f
C6536 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 GND 0.04798f
C6537 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 GND 0.22815f
C6538 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 GND 0.05969f
C6539 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 GND 0.15961f
C6540 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 GND 0.12257f
C6541 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 GND 0.23742f
C6542 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 GND 0.45664f
C6543 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 GND 0.1334f
C6544 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 GND 0.05705f
C6545 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 GND 0.10533f
C6546 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 GND 0.18236f
C6547 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 GND 0.13574f
C6548 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 GND 0.06431f
C6549 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 GND 0.45666f
C6550 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 GND 0.47347f
C6551 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 GND 0.05122f
C6552 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 GND 0.06839f
C6553 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 GND 0.22727f
C6554 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 GND 0.06194f
C6555 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 GND 0.39067f
C6556 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 GND 0.06323f
C6557 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 GND 0.06194f
C6558 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 GND 0.35224f
C6559 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 GND 0.11629f
C6560 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 GND 0.16533f
C6561 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 GND 0.36784f
C6562 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 GND 0.10746f
C6563 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 GND 0.04662f
C6564 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 GND 0.04798f
C6565 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 GND 0.22815f
C6566 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 GND 0.0518f
C6567 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 GND 0.36785f
C6568 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 GND 0.38072f
C6569 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 GND 0.19125f
C6570 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 GND 0.18752f
C6571 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 GND 0.10934f
C6572 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 GND 0.01378f
C6573 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 GND 0.01506f
C6574 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 GND 0.05094f
C6575 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 GND 0.04989f
C6576 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 GND 0.28374f
C6577 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 GND 0.09441f
C6578 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 GND 0.04989f
C6579 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 GND 0.31407f
C6580 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 GND 0.1838f
C6581 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 GND 0.205f
C6582 D_FlipFlop_0.3-input-nand_2.Vout.t6 GND 0.35515f
C6583 D_FlipFlop_0.3-input-nand_2.Vout.n0 GND 0.10375f
C6584 D_FlipFlop_0.3-input-nand_2.Vout.n1 GND 0.04502f
C6585 D_FlipFlop_0.3-input-nand_2.Vout.t2 GND 0.04632f
C6586 D_FlipFlop_0.3-input-nand_2.Vout.n2 GND 0.22028f
C6587 D_FlipFlop_0.3-input-nand_2.Vout.n3 GND 0.05002f
C6588 D_FlipFlop_0.3-input-nand_2.Vout.t5 GND 0.35517f
C6589 D_FlipFlop_0.3-input-nand_2.Vout.n4 GND 0.36759f
C6590 D_FlipFlop_0.3-input-nand_2.Vout.t7 GND 0.18465f
C6591 D_FlipFlop_0.3-input-nand_2.Vout.n5 GND 0.18106f
C6592 D_FlipFlop_0.3-input-nand_2.Vout.n6 GND 0.10557f
C6593 D_FlipFlop_0.3-input-nand_2.Vout.n7 GND 0.01331f
C6594 D_FlipFlop_0.3-input-nand_2.Vout.n8 GND 0.01454f
C6595 D_FlipFlop_0.3-input-nand_2.Vout.t1 GND 0.04918f
C6596 D_FlipFlop_0.3-input-nand_2.Vout.t0 GND 0.04817f
C6597 D_FlipFlop_0.3-input-nand_2.Vout.n9 GND 0.27396f
C6598 D_FlipFlop_0.3-input-nand_2.Vout.n10 GND 0.09115f
C6599 D_FlipFlop_0.3-input-nand_2.Vout.t3 GND 0.04817f
C6600 D_FlipFlop_0.3-input-nand_2.Vout.n11 GND 0.30324f
C6601 D_FlipFlop_0.3-input-nand_2.Vout.t4 GND 0.17747f
C6602 D_FlipFlop_0.3-input-nand_2.Vout.n12 GND 0.19793f
C6603 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 GND 0.36784f
C6604 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 GND 0.10746f
C6605 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 GND 0.04662f
C6606 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 GND 0.04798f
C6607 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 GND 0.22815f
C6608 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 GND 0.0518f
C6609 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 GND 0.36785f
C6610 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 GND 0.38072f
C6611 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 GND 0.19125f
C6612 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 GND 0.18752f
C6613 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 GND 0.10934f
C6614 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 GND 0.01378f
C6615 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 GND 0.01506f
C6616 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 GND 0.05094f
C6617 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 GND 0.04989f
C6618 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 GND 0.28374f
C6619 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 GND 0.09441f
C6620 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 GND 0.04989f
C6621 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 GND 0.31407f
C6622 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 GND 0.1838f
C6623 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 GND 0.205f
C6624 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 GND 0.45666f
C6625 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 GND 0.47347f
C6626 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 GND 0.05122f
C6627 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 GND 0.06839f
C6628 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 GND 0.22727f
C6629 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 GND 0.06194f
C6630 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 GND 0.39067f
C6631 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 GND 0.06323f
C6632 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 GND 0.06194f
C6633 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 GND 0.35224f
C6634 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 GND 0.11629f
C6635 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 GND 0.16533f
C6636 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 GND 0.06431f
C6637 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 GND 0.23742f
C6638 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 GND 0.45664f
C6639 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 GND 0.1334f
C6640 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 GND 0.05705f
C6641 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 GND 0.10533f
C6642 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 GND 0.18236f
C6643 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 GND 0.13574f
C6644 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 GND 0.12257f
C6645 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 GND 0.05969f
C6646 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 GND 0.15961f
C6647 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 GND 0.36784f
C6648 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 GND 0.10746f
C6649 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 GND 0.04662f
C6650 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 GND 0.205f
C6651 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 GND 0.1838f
C6652 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 GND 0.04989f
C6653 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 GND 0.31407f
C6654 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 GND 0.05094f
C6655 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 GND 0.04989f
C6656 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 GND 0.28374f
C6657 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 GND 0.09258f
C6658 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 GND 0.01095f
C6659 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 GND 0.01378f
C6660 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 GND 0.36785f
C6661 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 GND 0.38072f
C6662 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 GND 0.19125f
C6663 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 GND 0.18752f
C6664 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 GND 0.10934f
C6665 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 GND 0.0518f
C6666 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 GND 0.04798f
C6667 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 GND 0.22815f
C6668 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 GND 0.38055f
C6669 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 GND 0.39456f
C6670 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 GND 0.04269f
C6671 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 GND 0.04965f
C6672 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 GND 0.04808f
C6673 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 GND 0.10214f
C6674 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 GND 0.19785f
C6675 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 GND 0.38054f
C6676 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 GND 0.11117f
C6677 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 GND 0.04754f
C6678 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 GND 0.08777f
C6679 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 GND 0.15197f
C6680 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 GND 0.11312f
C6681 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 GND 0.05359f
C6682 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 GND 0.13778f
C6683 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 GND 0.05269f
C6684 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 GND 0.05162f
C6685 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 GND 0.29353f
C6686 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 GND 0.09691f
C6687 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 GND 0.05162f
C6688 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 GND 0.32556f
C6689 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 GND 0.18939f
C6690 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 GND 0.05699f
C6691 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 GND 0.05958f
C6692 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 GND 0.0577f
C6693 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 GND 0.12257f
C6694 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 GND 0.23742f
C6695 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 GND 0.45664f
C6696 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 GND 0.1334f
C6697 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 GND 0.05705f
C6698 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 GND 0.10533f
C6699 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 GND 0.18236f
C6700 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 GND 0.13574f
C6701 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 GND 0.06431f
C6702 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 GND 0.45666f
C6703 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 GND 0.47347f
C6704 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 GND 0.05122f
C6705 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 GND 0.06839f
C6706 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 GND 0.22727f
C6707 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 GND 0.06194f
C6708 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 GND 0.39067f
C6709 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 GND 0.06323f
C6710 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 GND 0.06194f
C6711 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 GND 0.35224f
C6712 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 GND 0.11629f
C6713 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 GND 0.16533f
C6714 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 GND 0.36784f
C6715 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 GND 0.10746f
C6716 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 GND 0.04662f
C6717 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 GND 0.04798f
C6718 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 GND 0.22815f
C6719 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 GND 0.0518f
C6720 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 GND 0.36785f
C6721 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 GND 0.38072f
C6722 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 GND 0.19125f
C6723 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 GND 0.18752f
C6724 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 GND 0.10934f
C6725 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 GND 0.01378f
C6726 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 GND 0.01095f
C6727 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 GND 0.05094f
C6728 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 GND 0.04989f
C6729 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 GND 0.28374f
C6730 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 GND 0.09258f
C6731 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 GND 0.04989f
C6732 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 GND 0.31407f
C6733 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 GND 0.1838f
C6734 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 GND 0.205f
C6735 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 GND 0.05958f
C6736 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 GND 0.0577f
C6737 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 GND 0.12257f
C6738 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 GND 0.23742f
C6739 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 GND 0.45664f
C6740 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 GND 0.1334f
C6741 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 GND 0.05705f
C6742 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 GND 0.10533f
C6743 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 GND 0.18236f
C6744 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 GND 0.13574f
C6745 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 GND 0.06431f
C6746 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 GND 0.45666f
C6747 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 GND 0.47347f
C6748 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 GND 0.05122f
C6749 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 GND 0.06839f
C6750 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 GND 0.22727f
C6751 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 GND 0.06194f
C6752 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 GND 0.39067f
C6753 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 GND 0.06323f
C6754 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 GND 0.06194f
C6755 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 GND 0.35224f
C6756 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 GND 0.11629f
C6757 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 GND 0.16533f
C6758 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 GND 0.07037f
C6759 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 GND 0.16004f
C6760 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 GND 0.07725f
C6761 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 GND 0.2799f
C6762 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 GND 0.27418f
C6763 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 GND 0.05783f
C6764 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 GND 0.53832f
C6765 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 GND 0.15726f
C6766 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 GND 0.03913f
C6767 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 GND 0.05692f
C6768 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 GND 0.14585f
C6769 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 GND 0.14585f
C6770 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 GND 0.07581f
C6771 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 GND 0.07318f
C6772 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 GND 0.07454f
C6773 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 GND 0.07302f
C6774 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 GND 0.41525f
C6775 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 GND 0.23391f
C6776 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 GND 0.22303f
C6777 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 GND 0.04607f
C6778 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 GND 0.10477f
C6779 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 GND 0.05057f
C6780 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 GND 0.35243f
C6781 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 GND 0.3654f
C6782 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 GND 0.03953f
C6783 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 GND 0.05278f
C6784 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 GND 0.27708f
C6785 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 GND 0.27709f
C6786 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 GND 0.17949f
C6787 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 GND 0.03786f
C6788 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 GND 0.35241f
C6789 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 GND 0.10295f
C6790 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 GND 0.02562f
C6791 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 GND 0.03726f
C6792 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 GND 0.09548f
C6793 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 GND 0.09548f
C6794 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 GND 0.04963f
C6795 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 GND 0.04792f
C6796 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 GND 0.28399f
C6797 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 GND 0.45666f
C6798 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 GND 0.47347f
C6799 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 GND 0.05122f
C6800 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 GND 0.06839f
C6801 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 GND 0.22727f
C6802 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 GND 0.06194f
C6803 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 GND 0.39067f
C6804 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 GND 0.06323f
C6805 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 GND 0.06194f
C6806 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 GND 0.35224f
C6807 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 GND 0.11629f
C6808 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 GND 0.16533f
C6809 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 GND 0.06431f
C6810 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 GND 0.23742f
C6811 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 GND 0.45664f
C6812 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 GND 0.1334f
C6813 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 GND 0.05705f
C6814 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 GND 0.10533f
C6815 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 GND 0.18236f
C6816 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 GND 0.13574f
C6817 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 GND 0.12257f
C6818 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 GND 0.0577f
C6819 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 GND 0.05958f
C6820 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 GND 0.06323f
C6821 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 GND 0.07525f
C6822 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 GND 0.38033f
C6823 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 GND 0.1927f
C6824 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 GND 0.0655f
C6825 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 GND 0.24183f
C6826 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 GND 0.23689f
C6827 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 GND 0.04996f
C6828 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 GND 0.46511f
C6829 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 GND 0.13587f
C6830 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 GND 0.03381f
C6831 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 GND 0.04918f
C6832 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 GND 0.12602f
C6833 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 GND 0.12602f
C6834 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 GND 0.06674f
C6835 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 GND 0.0608f
C6836 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 GND 0.13827f
C6837 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 GND 0.04607f
C6838 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 GND 0.10477f
C6839 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 GND 0.05057f
C6840 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 GND 0.35243f
C6841 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 GND 0.3654f
C6842 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 GND 0.03953f
C6843 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 GND 0.05278f
C6844 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 GND 0.27708f
C6845 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 GND 0.27709f
C6846 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 GND 0.17949f
C6847 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 GND 0.03786f
C6848 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 GND 0.35241f
C6849 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 GND 0.10295f
C6850 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 GND 0.02562f
C6851 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 GND 0.03726f
C6852 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 GND 0.09548f
C6853 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 GND 0.09548f
C6854 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 GND 0.04963f
C6855 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 GND 0.04792f
C6856 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 GND 0.28399f
C6857 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 GND 0.06358f
C6858 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 GND 0.03611f
C6859 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 GND 0.06992f
C6860 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 GND 0.25335f
C6861 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 GND 0.24817f
C6862 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 GND 0.05234f
C6863 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 GND 0.48726f
C6864 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 GND 0.14234f
C6865 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 GND 0.03542f
C6866 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 GND 0.05152f
C6867 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 GND 0.13202f
C6868 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 GND 0.13202f
C6869 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 GND 0.06862f
C6870 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 GND 0.06624f
C6871 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 GND 0.07883f
C6872 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 GND 0.39844f
C6873 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 GND 0.20187f
C6874 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 GND 0.04998f
C6875 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 GND 0.02839f
C6876 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 GND 0.05497f
C6877 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 GND 0.38308f
C6878 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 GND 0.39717f
C6879 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 GND 0.04297f
C6880 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 GND 0.05737f
C6881 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 GND 0.30118f
C6882 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 GND 0.30119f
C6883 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 GND 0.1951f
C6884 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 GND 0.04115f
C6885 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 GND 0.38306f
C6886 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 GND 0.1119f
C6887 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 GND 0.02784f
C6888 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 GND 0.0405f
C6889 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 GND 0.10379f
C6890 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 GND 0.10379f
C6891 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 GND 0.05395f
C6892 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 GND 0.05208f
C6893 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 GND 0.30868f
C6894 FFCLR.t35 GND 0.57049f
C6895 FFCLR.n0 GND 0.16666f
C6896 FFCLR.n1 GND 0.07231f
C6897 FFCLR.n2 GND 0.31794f
C6898 FFCLR.t6 GND 0.26535f
C6899 FFCLR.n3 GND 0.08324f
C6900 FFCLR.t2 GND 0.07441f
C6901 FFCLR.n4 GND 0.32404f
C6902 FFCLR.n5 GND 0.08034f
C6903 FFCLR.t41 GND 0.57052f
C6904 FFCLR.n6 GND 0.56067f
C6905 FFCLR.n7 GND 0.06128f
C6906 FFCLR.t34 GND 0.29661f
C6907 FFCLR.n8 GND 0.08544f
C6908 FFCLR.n9 GND 0.03662f
C6909 FFCLR.n10 GND 0.06861f
C6910 FFCLR.n11 GND 0.08634f
C6911 FFCLR.t32 GND 0.57052f
C6912 FFCLR.n12 GND 0.56067f
C6913 FFCLR.n13 GND 0.06128f
C6914 FFCLR.t40 GND 0.29661f
C6915 FFCLR.n14 GND 0.08544f
C6916 FFCLR.n15 GND 0.03662f
C6917 FFCLR.n16 GND 0.06861f
C6918 FFCLR.n17 GND 0.01029f
C6919 FFCLR.n18 GND 0.25889f
C6920 FFCLR.n19 GND 0.72092f
C6921 FFCLR.n20 GND 0.32349f
C6922 FFCLR.t39 GND 0.57052f
C6923 FFCLR.n21 GND 0.57454f
C6924 FFCLR.n22 GND 0.06128f
C6925 FFCLR.t11 GND 0.29661f
C6926 FFCLR.n23 GND 0.08544f
C6927 FFCLR.n24 GND 0.02276f
C6928 FFCLR.n25 GND 0.03546f
C6929 FFCLR.n26 GND 0.35381f
C6930 FFCLR.t13 GND 0.57052f
C6931 FFCLR.n27 GND 0.57454f
C6932 FFCLR.n28 GND 0.06128f
C6933 FFCLR.t38 GND 0.29661f
C6934 FFCLR.n29 GND 0.08544f
C6935 FFCLR.n30 GND 0.02276f
C6936 FFCLR.n31 GND 0.03546f
C6937 FFCLR.n32 GND 0.01029f
C6938 FFCLR.n33 GND 0.9187f
C6939 FFCLR.n34 GND 0.43004f
C6940 FFCLR.n35 GND 0.15867f
C6941 FFCLR.t26 GND 0.57049f
C6942 FFCLR.n36 GND 0.16666f
C6943 FFCLR.n37 GND 0.07231f
C6944 FFCLR.n38 GND 0.31794f
C6945 FFCLR.t44 GND 0.26532f
C6946 FFCLR.n39 GND 0.03217f
C6947 FFCLR.n40 GND 0.07753f
C6948 FFCLR.n41 GND 0.0209f
C6949 FFCLR.t19 GND 0.57052f
C6950 FFCLR.n42 GND 0.59152f
C6951 FFCLR.n43 GND 0.06399f
C6952 FFCLR.n44 GND 0.08544f
C6953 FFCLR.t27 GND 0.26647f
C6954 FFCLR.n45 GND 0.53562f
C6955 FFCLR.n46 GND 0.15225f
C6956 FFCLR.t33 GND 0.29663f
C6957 FFCLR.n47 GND 0.2767f
C6958 FFCLR.n48 GND 0.06128f
C6959 FFCLR.t53 GND 0.57049f
C6960 FFCLR.n49 GND 0.16666f
C6961 FFCLR.n50 GND 0.05533f
C6962 FFCLR.n51 GND 0.09347f
C6963 FFCLR.n52 GND 0.35381f
C6964 FFCLR.t8 GND 0.29663f
C6965 FFCLR.n53 GND 0.2767f
C6966 FFCLR.n54 GND 0.06128f
C6967 FFCLR.t23 GND 0.57049f
C6968 FFCLR.n55 GND 0.16666f
C6969 FFCLR.n56 GND 0.05533f
C6970 FFCLR.n57 GND 0.09347f
C6971 FFCLR.n58 GND 0.01029f
C6972 FFCLR.n59 GND 0.89843f
C6973 FFCLR.n60 GND 0.50081f
C6974 FFCLR.t37 GND 0.57052f
C6975 FFCLR.n61 GND 0.59152f
C6976 FFCLR.n62 GND 0.06399f
C6977 FFCLR.n63 GND 0.08544f
C6978 FFCLR.t45 GND 0.26644f
C6979 FFCLR.n64 GND 0.57937f
C6980 FFCLR.n65 GND 0.3227f
C6981 FFCLR.n66 GND 0.15225f
C6982 FFCLR.t50 GND 0.29663f
C6983 FFCLR.n67 GND 0.2767f
C6984 FFCLR.n68 GND 0.06128f
C6985 FFCLR.t12 GND 0.57049f
C6986 FFCLR.n69 GND 0.16666f
C6987 FFCLR.n70 GND 0.05533f
C6988 FFCLR.n71 GND 0.09347f
C6989 FFCLR.n72 GND 0.35381f
C6990 FFCLR.t22 GND 0.29663f
C6991 FFCLR.n73 GND 0.2767f
C6992 FFCLR.n74 GND 0.06128f
C6993 FFCLR.t42 GND 0.57049f
C6994 FFCLR.n75 GND 0.16666f
C6995 FFCLR.n76 GND 0.05533f
C6996 FFCLR.n77 GND 0.09347f
C6997 FFCLR.n78 GND 0.01029f
C6998 FFCLR.n79 GND 0.89843f
C6999 FFCLR.n80 GND 0.50081f
C7000 FFCLR.t14 GND 0.57052f
C7001 FFCLR.n81 GND 0.59152f
C7002 FFCLR.n82 GND 0.06399f
C7003 FFCLR.n83 GND 0.08544f
C7004 FFCLR.t7 GND 0.26644f
C7005 FFCLR.n84 GND 0.57937f
C7006 FFCLR.n85 GND 0.3227f
C7007 FFCLR.n86 GND 0.15225f
C7008 FFCLR.t24 GND 0.29663f
C7009 FFCLR.n87 GND 0.2767f
C7010 FFCLR.n88 GND 0.06128f
C7011 FFCLR.t31 GND 0.57049f
C7012 FFCLR.n89 GND 0.16666f
C7013 FFCLR.n90 GND 0.05533f
C7014 FFCLR.n91 GND 0.09347f
C7015 FFCLR.n92 GND 0.35381f
C7016 FFCLR.t56 GND 0.29663f
C7017 FFCLR.n93 GND 0.2767f
C7018 FFCLR.n94 GND 0.06128f
C7019 FFCLR.t4 GND 0.57049f
C7020 FFCLR.n95 GND 0.16666f
C7021 FFCLR.n96 GND 0.05533f
C7022 FFCLR.n97 GND 0.09347f
C7023 FFCLR.n98 GND 0.01029f
C7024 FFCLR.n99 GND 0.89843f
C7025 FFCLR.n100 GND 0.80733f
C7026 FFCLR.n101 GND 0.10925f
C7027 FFCLR.t54 GND 0.29663f
C7028 FFCLR.n102 GND 0.2767f
C7029 FFCLR.n103 GND 0.06128f
C7030 FFCLR.t17 GND 0.57049f
C7031 FFCLR.n104 GND 0.16666f
C7032 FFCLR.n105 GND 0.05533f
C7033 FFCLR.n106 GND 0.09347f
C7034 FFCLR.n107 GND 0.35381f
C7035 FFCLR.t28 GND 0.29663f
C7036 FFCLR.n108 GND 0.2767f
C7037 FFCLR.n109 GND 0.06128f
C7038 FFCLR.t46 GND 0.57049f
C7039 FFCLR.n110 GND 0.16666f
C7040 FFCLR.n111 GND 0.05533f
C7041 FFCLR.n112 GND 0.09347f
C7042 FFCLR.n113 GND 0.01029f
C7043 FFCLR.n114 GND 0.89843f
C7044 FFCLR.n115 GND 0.12892f
C7045 FFCLR.n116 GND 0.15225f
C7046 FFCLR.n117 GND 0.3227f
C7047 FFCLR.t43 GND 0.57052f
C7048 FFCLR.n118 GND 0.59152f
C7049 FFCLR.n119 GND 0.06399f
C7050 FFCLR.n120 GND 0.08544f
C7051 FFCLR.t49 GND 0.26644f
C7052 FFCLR.n121 GND 0.20748f
C7053 FFCLR.n122 GND 0.59187f
C7054 FFCLR.n123 GND 1.01694f
C7055 FFCLR.t10 GND 0.29663f
C7056 FFCLR.n124 GND 0.2767f
C7057 FFCLR.n125 GND 0.06128f
C7058 FFCLR.t29 GND 0.57049f
C7059 FFCLR.n126 GND 0.16666f
C7060 FFCLR.n127 GND 0.05533f
C7061 FFCLR.n128 GND 0.09347f
C7062 FFCLR.n129 GND 0.35381f
C7063 FFCLR.t36 GND 0.29663f
C7064 FFCLR.n130 GND 0.2767f
C7065 FFCLR.n131 GND 0.06128f
C7066 FFCLR.t59 GND 0.57049f
C7067 FFCLR.n132 GND 0.16666f
C7068 FFCLR.n133 GND 0.05533f
C7069 FFCLR.n134 GND 0.09347f
C7070 FFCLR.n135 GND 0.01029f
C7071 FFCLR.n136 GND 0.89843f
C7072 FFCLR.n137 GND 0.12892f
C7073 FFCLR.n138 GND 0.15225f
C7074 FFCLR.n139 GND 0.3227f
C7075 FFCLR.t15 GND 0.57052f
C7076 FFCLR.n140 GND 0.59152f
C7077 FFCLR.n141 GND 0.06399f
C7078 FFCLR.n142 GND 0.08544f
C7079 FFCLR.t9 GND 0.26644f
C7080 FFCLR.n143 GND 0.20748f
C7081 FFCLR.n144 GND 1.12885f
C7082 FFCLR.n145 GND 1.60761f
C7083 FFCLR.t21 GND 0.29663f
C7084 FFCLR.n146 GND 0.2767f
C7085 FFCLR.n147 GND 0.06128f
C7086 FFCLR.t25 GND 0.57049f
C7087 FFCLR.n148 GND 0.16666f
C7088 FFCLR.n149 GND 0.05533f
C7089 FFCLR.n150 GND 0.09347f
C7090 FFCLR.n151 GND 0.35381f
C7091 FFCLR.t51 GND 0.29663f
C7092 FFCLR.n152 GND 0.2767f
C7093 FFCLR.n153 GND 0.06128f
C7094 FFCLR.t57 GND 0.57049f
C7095 FFCLR.n154 GND 0.16666f
C7096 FFCLR.n155 GND 0.05533f
C7097 FFCLR.n156 GND 0.09347f
C7098 FFCLR.n157 GND 0.01029f
C7099 FFCLR.n158 GND 0.89843f
C7100 FFCLR.n159 GND 0.12892f
C7101 FFCLR.n160 GND 0.15225f
C7102 FFCLR.n161 GND 0.3227f
C7103 FFCLR.t52 GND 0.57052f
C7104 FFCLR.n162 GND 0.59152f
C7105 FFCLR.n163 GND 0.06399f
C7106 FFCLR.n164 GND 0.08544f
C7107 FFCLR.t5 GND 0.26644f
C7108 FFCLR.n165 GND 0.20748f
C7109 FFCLR.n166 GND 1.66583f
C7110 FFCLR.n167 GND 2.19829f
C7111 FFCLR.t58 GND 0.29663f
C7112 FFCLR.n168 GND 0.2767f
C7113 FFCLR.n169 GND 0.06128f
C7114 FFCLR.t18 GND 0.57049f
C7115 FFCLR.n170 GND 0.16666f
C7116 FFCLR.n171 GND 0.05533f
C7117 FFCLR.n172 GND 0.09347f
C7118 FFCLR.n173 GND 0.35381f
C7119 FFCLR.t30 GND 0.29663f
C7120 FFCLR.n174 GND 0.2767f
C7121 FFCLR.n175 GND 0.06128f
C7122 FFCLR.t47 GND 0.57049f
C7123 FFCLR.n176 GND 0.16666f
C7124 FFCLR.n177 GND 0.05533f
C7125 FFCLR.n178 GND 0.09347f
C7126 FFCLR.n179 GND 0.01029f
C7127 FFCLR.n180 GND 0.89843f
C7128 FFCLR.n181 GND 0.12892f
C7129 FFCLR.n182 GND 0.15225f
C7130 FFCLR.n183 GND 0.3227f
C7131 FFCLR.t20 GND 0.57052f
C7132 FFCLR.n184 GND 0.59152f
C7133 FFCLR.n185 GND 0.06399f
C7134 FFCLR.n186 GND 0.08544f
C7135 FFCLR.t55 GND 0.26644f
C7136 FFCLR.n187 GND 0.20748f
C7137 FFCLR.n188 GND 2.27122f
C7138 FFCLR.n189 GND 3.08826f
C7139 FFCLR.n190 GND 0.993f
C7140 FFCLR.n191 GND 15.2532f
C7141 FFCLR.t16 GND 0.29663f
C7142 FFCLR.n192 GND 0.29056f
C7143 FFCLR.n193 GND 0.06128f
C7144 FFCLR.t48 GND 0.57049f
C7145 FFCLR.n194 GND 0.16666f
C7146 FFCLR.n195 GND 0.04147f
C7147 FFCLR.n196 GND 0.06032f
C7148 FFCLR.n197 GND 0.08883f
C7149 FFCLR.n198 GND 16.1053f
C7150 FFCLR.n199 GND 0.31392f
C7151 FFCLR.n200 GND 0.09176f
C7152 FFCLR.n201 GND 0.03377f
C7153 FFCLR.n202 GND 0.01045f
C7154 FFCLR.n203 GND 0.09264f
C7155 FFCLR.n204 GND 0.04678f
C7156 FFCLR.t1 GND 0.079f
C7157 FFCLR.t0 GND 0.07738f
C7158 FFCLR.n205 GND 0.44006f
C7159 FFCLR.n206 GND 0.14359f
C7160 FFCLR.t3 GND 0.07738f
C7161 FFCLR.n207 GND 0.1192f
C7162 FFCLR.n208 GND 0.21106f
C7163 Nand_Gate_6.A.t7 GND 0.27993f
C7164 Nand_Gate_6.A.n0 GND 0.08177f
C7165 Nand_Gate_6.A.n1 GND 0.03548f
C7166 Nand_Gate_6.A.n2 GND 0.15601f
C7167 Nand_Gate_6.A.t11 GND 0.1302f
C7168 Nand_Gate_6.A.n3 GND 0.04085f
C7169 Nand_Gate_6.A.t2 GND 0.03651f
C7170 Nand_Gate_6.A.n4 GND 0.159f
C7171 Nand_Gate_6.A.n5 GND 0.03942f
C7172 Nand_Gate_6.A.t4 GND 0.27994f
C7173 Nand_Gate_6.A.n6 GND 0.27511f
C7174 Nand_Gate_6.A.n7 GND 0.03007f
C7175 Nand_Gate_6.A.t10 GND 0.14554f
C7176 Nand_Gate_6.A.n8 GND 0.04192f
C7177 Nand_Gate_6.A.n9 GND 0.01797f
C7178 Nand_Gate_6.A.n10 GND 0.03367f
C7179 Nand_Gate_6.A.n11 GND 0.04236f
C7180 Nand_Gate_6.A.t6 GND 0.27994f
C7181 Nand_Gate_6.A.n12 GND 0.27511f
C7182 Nand_Gate_6.A.n13 GND 0.03007f
C7183 Nand_Gate_6.A.t8 GND 0.14554f
C7184 Nand_Gate_6.A.n14 GND 0.04192f
C7185 Nand_Gate_6.A.n15 GND 0.01797f
C7186 Nand_Gate_6.A.n16 GND 0.03367f
C7187 Nand_Gate_6.A.n18 GND 0.12656f
C7188 Nand_Gate_6.A.n19 GND 0.03459f
C7189 Nand_Gate_6.A.n20 GND 0.09204f
C7190 Nand_Gate_6.A.t9 GND 0.14555f
C7191 Nand_Gate_6.A.n21 GND 0.14257f
C7192 Nand_Gate_6.A.n22 GND 0.03007f
C7193 Nand_Gate_6.A.t5 GND 0.27993f
C7194 Nand_Gate_6.A.n23 GND 0.08177f
C7195 Nand_Gate_6.A.n24 GND 0.02035f
C7196 Nand_Gate_6.A.n25 GND 0.0296f
C7197 Nand_Gate_6.A.n26 GND 0.14551f
C7198 Nand_Gate_6.A.n27 GND 0.25531f
C7199 Nand_Gate_6.A.n28 GND 0.15873f
C7200 Nand_Gate_6.A.n29 GND 0.34318f
C7201 Nand_Gate_6.A.n31 GND 0.04546f
C7202 Nand_Gate_6.A.n32 GND 0.02608f
C7203 Nand_Gate_6.A.t1 GND 0.03876f
C7204 Nand_Gate_6.A.t0 GND 0.03797f
C7205 Nand_Gate_6.A.n33 GND 0.21593f
C7206 Nand_Gate_6.A.n34 GND 0.07184f
C7207 Nand_Gate_6.A.t3 GND 0.03797f
C7208 Nand_Gate_6.A.n35 GND 0.05849f
C7209 Nand_Gate_6.A.n36 GND 0.10356f
C7210 Nand_Gate_5.B.t9 GND 0.09725f
C7211 Nand_Gate_5.B.n0 GND 0.02801f
C7212 Nand_Gate_5.B.n1 GND 0.01201f
C7213 Nand_Gate_5.B.n2 GND 0.02249f
C7214 Nand_Gate_5.B.t8 GND 0.18705f
C7215 Nand_Gate_5.B.n3 GND 0.18382f
C7216 Nand_Gate_5.B.n4 GND 0.02009f
C7217 Nand_Gate_5.B.t11 GND 0.09725f
C7218 Nand_Gate_5.B.n5 GND 0.02801f
C7219 Nand_Gate_5.B.n6 GND 0.01201f
C7220 Nand_Gate_5.B.n7 GND 0.02249f
C7221 Nand_Gate_5.B.n8 GND 0.05912f
C7222 Nand_Gate_5.B.n9 GND 0.05912f
C7223 Nand_Gate_5.B.n10 GND 0.02009f
C7224 Nand_Gate_5.B.n11 GND 0.18382f
C7225 Nand_Gate_5.B.t10 GND 0.16795f
C7226 Nand_Gate_5.B.n12 GND 1.59684f
C7227 Nand_Gate_5.B.t6 GND 0.09725f
C7228 Nand_Gate_5.B.t4 GND 0.18704f
C7229 Nand_Gate_5.B.n13 GND 0.05464f
C7230 Nand_Gate_5.B.n14 GND 0.02337f
C7231 Nand_Gate_5.B.n15 GND 0.04314f
C7232 Nand_Gate_5.B.n16 GND 0.36438f
C7233 Nand_Gate_5.B.n17 GND 2.13619f
C7234 Nand_Gate_5.B.t5 GND 0.16927f
C7235 Nand_Gate_5.B.n18 GND 0.05464f
C7236 Nand_Gate_5.B.n19 GND 0.02371f
C7237 Nand_Gate_5.B.n20 GND 0.10424f
C7238 Nand_Gate_5.B.t7 GND 0.087f
C7239 Nand_Gate_5.B.n21 GND 0.02729f
C7240 Nand_Gate_5.B.t1 GND 0.0244f
C7241 Nand_Gate_5.B.n22 GND 0.11964f
C7242 Nand_Gate_5.B.n23 GND 0.02727f
C7243 Nand_Gate_5.B.t3 GND 0.0259f
C7244 Nand_Gate_5.B.t0 GND 0.02537f
C7245 Nand_Gate_5.B.n24 GND 0.14428f
C7246 Nand_Gate_5.B.n25 GND 0.04708f
C7247 Nand_Gate_5.B.t2 GND 0.02537f
C7248 Nand_Gate_5.B.n26 GND 0.03908f
C7249 Nand_Gate_5.B.n27 GND 0.0692f
C7250 CDAC8_0.switch_9.Z.t2 GND 0.03608f
C7251 CDAC8_0.switch_9.Z.t1 GND 0.0344f
C7252 CDAC8_0.switch_9.Z.t3 GND 0.0344f
C7253 CDAC8_0.switch_9.Z.n0 GND 0.12427f
C7254 CDAC8_0.switch_9.Z.n1 GND 0.28559f
C7255 CDAC8_0.switch_9.Z.n2 GND 0.0372f
C7256 CDAC8_0.switch_9.Z.t25 GND 6.43398f
C7257 CDAC8_0.switch_9.Z.t23 GND 6.07647f
C7258 CDAC8_0.switch_9.Z.n3 GND 3.42262f
C7259 CDAC8_0.switch_9.Z.t32 GND 6.07647f
C7260 CDAC8_0.switch_9.Z.n4 GND 1.60172f
C7261 CDAC8_0.switch_9.Z.n5 GND 1.3726f
C7262 CDAC8_0.switch_9.Z.t28 GND 6.43398f
C7263 CDAC8_0.switch_9.Z.t27 GND 6.07647f
C7264 CDAC8_0.switch_9.Z.n6 GND 3.42262f
C7265 CDAC8_0.switch_9.Z.t35 GND 6.07647f
C7266 CDAC8_0.switch_9.Z.n7 GND 1.60172f
C7267 CDAC8_0.switch_9.Z.t31 GND 6.44738f
C7268 CDAC8_0.switch_9.Z.t24 GND 6.07647f
C7269 CDAC8_0.switch_9.Z.n8 GND 3.47318f
C7270 CDAC8_0.switch_9.Z.t26 GND 6.07647f
C7271 CDAC8_0.switch_9.Z.n9 GND 1.75389f
C7272 CDAC8_0.switch_9.Z.t30 GND 6.07647f
C7273 CDAC8_0.switch_9.Z.n10 GND 1.88076f
C7274 CDAC8_0.switch_9.Z.t10 GND 6.07647f
C7275 CDAC8_0.switch_9.Z.n11 GND 2.07349f
C7276 CDAC8_0.switch_9.Z.t14 GND 6.07647f
C7277 CDAC8_0.switch_9.Z.n12 GND 2.07349f
C7278 CDAC8_0.switch_9.Z.t13 GND 6.07647f
C7279 CDAC8_0.switch_9.Z.n13 GND 2.07349f
C7280 CDAC8_0.switch_9.Z.t18 GND 6.07647f
C7281 CDAC8_0.switch_9.Z.n14 GND 2.07349f
C7282 CDAC8_0.switch_9.Z.t17 GND 6.07647f
C7283 CDAC8_0.switch_9.Z.n15 GND 2.07349f
C7284 CDAC8_0.switch_9.Z.t34 GND 6.07647f
C7285 CDAC8_0.switch_9.Z.n16 GND 2.07349f
C7286 CDAC8_0.switch_9.Z.t6 GND 6.07647f
C7287 CDAC8_0.switch_9.Z.n17 GND 2.07349f
C7288 CDAC8_0.switch_9.Z.t5 GND 6.07647f
C7289 CDAC8_0.switch_9.Z.n18 GND 2.07349f
C7290 CDAC8_0.switch_9.Z.t9 GND 6.07647f
C7291 CDAC8_0.switch_9.Z.n19 GND 1.72859f
C7292 CDAC8_0.switch_9.Z.t29 GND 6.44738f
C7293 CDAC8_0.switch_9.Z.t20 GND 6.07647f
C7294 CDAC8_0.switch_9.Z.n20 GND 3.47318f
C7295 CDAC8_0.switch_9.Z.t22 GND 6.07647f
C7296 CDAC8_0.switch_9.Z.n21 GND 1.75389f
C7297 CDAC8_0.switch_9.Z.n22 GND 1.99f
C7298 CDAC8_0.switch_9.Z.n23 GND 1.99f
C7299 CDAC8_0.switch_9.Z.t11 GND 6.07647f
C7300 CDAC8_0.switch_9.Z.n24 GND 1.72859f
C7301 CDAC8_0.switch_9.Z.t7 GND 6.07647f
C7302 CDAC8_0.switch_9.Z.n25 GND 2.07349f
C7303 CDAC8_0.switch_9.Z.t8 GND 6.07647f
C7304 CDAC8_0.switch_9.Z.n26 GND 2.07349f
C7305 CDAC8_0.switch_9.Z.t4 GND 6.07647f
C7306 CDAC8_0.switch_9.Z.n27 GND 2.07349f
C7307 CDAC8_0.switch_9.Z.t19 GND 6.07647f
C7308 CDAC8_0.switch_9.Z.n28 GND 2.07349f
C7309 CDAC8_0.switch_9.Z.t21 GND 6.07647f
C7310 CDAC8_0.switch_9.Z.n29 GND 2.07349f
C7311 CDAC8_0.switch_9.Z.t15 GND 6.07647f
C7312 CDAC8_0.switch_9.Z.n30 GND 2.07349f
C7313 CDAC8_0.switch_9.Z.t16 GND 6.07647f
C7314 CDAC8_0.switch_9.Z.n31 GND 2.07349f
C7315 CDAC8_0.switch_9.Z.t12 GND 6.07647f
C7316 CDAC8_0.switch_9.Z.n32 GND 2.07349f
C7317 CDAC8_0.switch_9.Z.t33 GND 6.07647f
C7318 CDAC8_0.switch_9.Z.n33 GND 1.88076f
C7319 CDAC8_0.switch_9.Z.n34 GND 1.32914f
C7320 CDAC8_0.switch_9.Z.n35 GND 1.3012f
C7321 CDAC8_0.switch_9.Z.n36 GND 0.01846f
C7322 CDAC8_0.switch_9.Z.t0 GND 0.03608f
C7323 CDAC8_0.switch_9.Z.n37 GND 0.149f
C7324 D_FlipFlop_2.3-input-nand_2.C.t1 GND 0.04477f
C7325 D_FlipFlop_2.3-input-nand_2.C.n0 GND 0.11971f
C7326 D_FlipFlop_2.3-input-nand_2.C.n1 GND 0.09193f
C7327 D_FlipFlop_2.3-input-nand_2.C.t4 GND 0.17806f
C7328 D_FlipFlop_2.3-input-nand_2.C.t5 GND 0.34248f
C7329 D_FlipFlop_2.3-input-nand_2.C.n2 GND 0.10005f
C7330 D_FlipFlop_2.3-input-nand_2.C.n3 GND 0.04279f
C7331 D_FlipFlop_2.3-input-nand_2.C.n4 GND 0.079f
C7332 D_FlipFlop_2.3-input-nand_2.C.n5 GND 0.13677f
C7333 D_FlipFlop_2.3-input-nand_2.C.n6 GND 0.10181f
C7334 D_FlipFlop_2.3-input-nand_2.C.n7 GND 0.04823f
C7335 D_FlipFlop_2.3-input-nand_2.C.t7 GND 0.3425f
C7336 D_FlipFlop_2.3-input-nand_2.C.n8 GND 0.3551f
C7337 D_FlipFlop_2.3-input-nand_2.C.n9 GND 0.03842f
C7338 D_FlipFlop_2.3-input-nand_2.C.n10 GND 0.05129f
C7339 D_FlipFlop_2.3-input-nand_2.C.t6 GND 0.17045f
C7340 D_FlipFlop_2.3-input-nand_2.C.t0 GND 0.04645f
C7341 D_FlipFlop_2.3-input-nand_2.C.n11 GND 0.293f
C7342 D_FlipFlop_2.3-input-nand_2.C.t3 GND 0.04742f
C7343 D_FlipFlop_2.3-input-nand_2.C.t2 GND 0.04645f
C7344 D_FlipFlop_2.3-input-nand_2.C.n12 GND 0.26418f
C7345 D_FlipFlop_2.3-input-nand_2.C.n13 GND 0.08722f
C7346 D_FlipFlop_2.3-input-nand_2.C.n14 GND 0.124f
C7347 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 GND 0.04607f
C7348 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 GND 0.10477f
C7349 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 GND 0.05057f
C7350 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 GND 0.35243f
C7351 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 GND 0.3654f
C7352 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 GND 0.03953f
C7353 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 GND 0.05278f
C7354 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 GND 0.27708f
C7355 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 GND 0.27709f
C7356 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 GND 0.17949f
C7357 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 GND 0.03786f
C7358 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 GND 0.35241f
C7359 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 GND 0.10295f
C7360 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 GND 0.02562f
C7361 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 GND 0.03726f
C7362 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 GND 0.09548f
C7363 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 GND 0.09548f
C7364 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 GND 0.04963f
C7365 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 GND 0.04792f
C7366 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 GND 0.28399f
C7367 And_Gate_3.Vout.t1 GND 0.08912f
C7368 And_Gate_3.Inverter_0.Vout GND 0.02589f
C7369 And_Gate_3.Vout.n0 GND 0.09833f
C7370 And_Gate_3.Vout.t5 GND 0.68307f
C7371 D_FlipFlop_4.3-input-nand_0.C GND -0.40609f
C7372 And_Gate_3.Vout.n1 GND 0.70821f
C7373 And_Gate_3.Vout.n2 GND 0.07662f
C7374 And_Gate_3.Vout.n3 GND 0.1023f
C7375 And_Gate_3.Vout.t3 GND 0.31442f
C7376 D_FlipFlop_4.CLK GND -0.02336f
C7377 And_Gate_3.Vout.n4 GND 0.2457f
C7378 And_Gate_3.Vout.t2 GND 0.68304f
C7379 D_FlipFlop_4.3-input-nand_1.C GND -0.22831f
C7380 And_Gate_3.Vout.t4 GND 0.35514f
C7381 D_FlipFlop_4.Inverter_1.Vin GND -0.22174f
C7382 And_Gate_3.Vout.n5 GND 0.37451f
C7383 And_Gate_3.Vout.t7 GND 0.68304f
C7384 And_Gate_3.Vout.n6 GND 0.60464f
C7385 And_Gate_3.Vout.n7 GND 0.6063f
C7386 And_Gate_3.Vout.n8 GND 0.37942f
C7387 And_Gate_3.Vout.t6 GND 0.31441f
C7388 And_Gate_3.Vout.n9 GND 0.06377f
C7389 And_Gate_3.Vout.n10 GND 0.15007f
C7390 And_Gate_3.Vout.n11 GND 6.09909f
C7391 And_Gate_3.Vout.t0 GND 0.09306f
C7392 And_Gate_3.Vout.n12 GND 4.81721f
C7393 And_Gate_3.Vout.n13 GND 0.21212f
C7394 D_FlipFlop_0.CLK.t1 GND 0.0601f
C7395 D_FlipFlop_0.CLK.t3 GND 0.46171f
C7396 D_FlipFlop_0.CLK.n0 GND 0.47871f
C7397 D_FlipFlop_0.CLK.n1 GND 0.05179f
C7398 D_FlipFlop_0.CLK.n2 GND 0.06915f
C7399 D_FlipFlop_0.CLK.t6 GND 0.21251f
C7400 D_FlipFlop_0.CLK.n3 GND 0.19074f
C7401 D_FlipFlop_0.CLK.n4 GND 0.06086f
C7402 D_FlipFlop_0.CLK.t5 GND 0.46169f
C7403 D_FlipFlop_0.CLK.t7 GND 0.24006f
C7404 D_FlipFlop_0.CLK.n5 GND 0.25315f
C7405 D_FlipFlop_0.CLK.t4 GND 0.46169f
C7406 D_FlipFlop_0.CLK.n6 GND 0.4087f
C7407 D_FlipFlop_0.CLK.n7 GND 0.40982f
C7408 D_FlipFlop_0.CLK.n8 GND 0.25646f
C7409 D_FlipFlop_0.CLK.t2 GND 0.21252f
C7410 D_FlipFlop_0.CLK.n9 GND 0.01225f
C7411 D_FlipFlop_0.CLK.n10 GND 0.03152f
C7412 D_FlipFlop_0.CLK.n11 GND 1.48264f
C7413 D_FlipFlop_0.CLK.n12 GND 0.85866f
C7414 D_FlipFlop_0.CLK.n13 GND 0.01206f
C7415 D_FlipFlop_0.CLK.n14 GND 0.06203f
C7416 D_FlipFlop_0.CLK.t0 GND 0.06278f
C7417 D_FlipFlop_0.CLK.n15 GND 0.40066f
C7418 And_Gate_4.Vout.t1 GND 0.1132f
C7419 And_Gate_4.Inverter_0.Vout GND -0.36385f
C7420 And_Gate_4.Vout.n0 GND 0.06429f
C7421 And_Gate_4.Vout.n1 GND 0.12449f
C7422 And_Gate_4.Vout.t5 GND 0.86757f
C7423 D_FlipFlop_2.3-input-nand_0.C GND -0.51578f
C7424 And_Gate_4.Vout.n2 GND 0.89951f
C7425 And_Gate_4.Vout.n3 GND 0.09731f
C7426 And_Gate_4.Vout.n4 GND 0.12993f
C7427 And_Gate_4.Vout.t6 GND 0.39932f
C7428 D_FlipFlop_2.CLK GND 0.05804f
C7429 And_Gate_4.Vout.n5 GND 0.3804f
C7430 And_Gate_4.Vout.n6 GND 0.11436f
C7431 And_Gate_4.Vout.t4 GND 0.86753f
C7432 D_FlipFlop_2.3-input-nand_1.C GND -0.28998f
C7433 And_Gate_4.Vout.t7 GND 0.45107f
C7434 D_FlipFlop_2.Inverter_1.Vin GND -0.28164f
C7435 And_Gate_4.Vout.n7 GND 0.47567f
C7436 And_Gate_4.Vout.t3 GND 0.86753f
C7437 And_Gate_4.Vout.n8 GND 0.76796f
C7438 And_Gate_4.Vout.n9 GND 0.77006f
C7439 And_Gate_4.Vout.n10 GND 0.4819f
C7440 And_Gate_4.Vout.t2 GND 0.39933f
C7441 And_Gate_4.Vout.n11 GND 15.5365f
C7442 And_Gate_4.Vout.n12 GND 12.546f
C7443 And_Gate_4.Vout.n13 GND 0.12217f
C7444 And_Gate_4.Vout.t0 GND 0.11796f
C7445 And_Gate_4.Vout.n14 GND 0.69909f
C7446 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 GND 0.0608f
C7447 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 GND 0.13827f
C7448 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 GND 0.06674f
C7449 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 GND 0.24183f
C7450 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 GND 0.23689f
C7451 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 GND 0.04996f
C7452 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 GND 0.46511f
C7453 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 GND 0.13587f
C7454 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 GND 0.03381f
C7455 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 GND 0.04918f
C7456 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 GND 0.12602f
C7457 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 GND 0.12602f
C7458 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 GND 0.0655f
C7459 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 GND 0.06323f
C7460 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 GND 0.07525f
C7461 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 GND 0.38033f
C7462 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 GND 0.1927f
C7463 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 GND 0.04607f
C7464 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 GND 0.10477f
C7465 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 GND 0.05057f
C7466 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 GND 0.35243f
C7467 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 GND 0.3654f
C7468 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 GND 0.03953f
C7469 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 GND 0.05278f
C7470 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 GND 0.27708f
C7471 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 GND 0.27709f
C7472 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 GND 0.17949f
C7473 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 GND 0.03786f
C7474 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 GND 0.35241f
C7475 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 GND 0.10295f
C7476 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 GND 0.02562f
C7477 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 GND 0.03726f
C7478 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 GND 0.09548f
C7479 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 GND 0.09548f
C7480 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 GND 0.04963f
C7481 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 GND 0.04792f
C7482 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 GND 0.28399f
C7483 Nand_Gate_2.B.t10 GND 0.33127f
C7484 Nand_Gate_2.B.n0 GND 0.09677f
C7485 Nand_Gate_2.B.n1 GND 0.04199f
C7486 Nand_Gate_2.B.n2 GND 0.18462f
C7487 Nand_Gate_2.B.t5 GND 0.15408f
C7488 Nand_Gate_2.B.n3 GND 0.04834f
C7489 Nand_Gate_2.B.n4 GND 0.12256f
C7490 Nand_Gate_2.B.t1 GND 0.04493f
C7491 Nand_Gate_2.B.n5 GND 0.06922f
C7492 Nand_Gate_2.B.t2 GND 0.04587f
C7493 Nand_Gate_2.B.t3 GND 0.04493f
C7494 Nand_Gate_2.B.n6 GND 0.25554f
C7495 Nand_Gate_2.B.n7 GND 0.08338f
C7496 Nand_Gate_2.B.n8 GND 0.02717f
C7497 Nand_Gate_2.B.n9 GND 0.05379f
C7498 Nand_Gate_2.B.t7 GND 0.33129f
C7499 Nand_Gate_2.B.n10 GND 0.32557f
C7500 Nand_Gate_2.B.n11 GND 0.03558f
C7501 Nand_Gate_2.B.t4 GND 0.17224f
C7502 Nand_Gate_2.B.n12 GND 0.04961f
C7503 Nand_Gate_2.B.n13 GND 0.02126f
C7504 Nand_Gate_2.B.n14 GND 0.03984f
C7505 Nand_Gate_2.B.n15 GND 0.05014f
C7506 Nand_Gate_2.B.t6 GND 0.33129f
C7507 Nand_Gate_2.B.n16 GND 0.32557f
C7508 Nand_Gate_2.B.n17 GND 0.03558f
C7509 Nand_Gate_2.B.t8 GND 0.17224f
C7510 Nand_Gate_2.B.n18 GND 0.04961f
C7511 Nand_Gate_2.B.n19 GND 0.02126f
C7512 Nand_Gate_2.B.n20 GND 0.03984f
C7513 Nand_Gate_2.B.n22 GND 0.15033f
C7514 Nand_Gate_2.B.n23 GND 0.41862f
C7515 Nand_Gate_2.B.n24 GND 0.18785f
C7516 Nand_Gate_2.B.t11 GND 0.17224f
C7517 Nand_Gate_2.B.t9 GND 0.33127f
C7518 Nand_Gate_2.B.n25 GND 0.09677f
C7519 Nand_Gate_2.B.n26 GND 0.04139f
C7520 Nand_Gate_2.B.n27 GND 0.07641f
C7521 Nand_Gate_2.B.n28 GND 0.87221f
C7522 Nand_Gate_2.B.n29 GND 1.18609f
C7523 Nand_Gate_2.B.n30 GND 0.05328f
C7524 Nand_Gate_2.B.n31 GND 0.01961f
C7525 Nand_Gate_2.B.n33 GND 0.04665f
C7526 Nand_Gate_2.B.t0 GND 0.04321f
C7527 Nand_Gate_2.B.n34 GND 0.18816f
C7528 And_Gate_1.Vout.t1 GND 0.08622f
C7529 And_Gate_1.Inverter_0.Vout GND 0.02505f
C7530 And_Gate_1.Vout.n0 GND 0.09513f
C7531 And_Gate_1.Vout.t6 GND 0.66083f
C7532 D_FlipFlop_7.3-input-nand_0.C GND -0.39286f
C7533 And_Gate_1.Vout.n1 GND 0.68515f
C7534 And_Gate_1.Vout.n2 GND 0.07412f
C7535 And_Gate_1.Vout.n3 GND 0.09897f
C7536 And_Gate_1.Vout.t3 GND 0.30416f
C7537 D_FlipFlop_7.CLK GND -0.06024f
C7538 And_Gate_1.Vout.n4 GND 0.24717f
C7539 And_Gate_1.Vout.n5 GND 0.08711f
C7540 And_Gate_1.Vout.t2 GND 0.6608f
C7541 D_FlipFlop_7.3-input-nand_1.C GND -0.22088f
C7542 And_Gate_1.Vout.t4 GND 0.34358f
C7543 D_FlipFlop_7.Inverter_1.Vin GND -0.21452f
C7544 And_Gate_1.Vout.n6 GND 0.36232f
C7545 And_Gate_1.Vout.t7 GND 0.6608f
C7546 And_Gate_1.Vout.n7 GND 0.58495f
C7547 And_Gate_1.Vout.n8 GND 0.58655f
C7548 And_Gate_1.Vout.n9 GND 0.36707f
C7549 And_Gate_1.Vout.t5 GND 0.30417f
C7550 And_Gate_1.Vout.n10 GND 0.04337f
C7551 And_Gate_1.Vout.n11 GND 0.10365f
C7552 And_Gate_1.Vout.n12 GND 16.2797f
C7553 And_Gate_1.Vout.t0 GND 0.09003f
C7554 And_Gate_1.Vout.n13 GND 13.6324f
C7555 And_Gate_1.Vout.n14 GND 0.20521f
C7556 Nand_Gate_2.A.t8 GND 0.62844f
C7557 Nand_Gate_2.A.n0 GND 0.18359f
C7558 Nand_Gate_2.A.n1 GND 0.07966f
C7559 Nand_Gate_2.A.n2 GND 0.35024f
C7560 Nand_Gate_2.A.t11 GND 0.2923f
C7561 Nand_Gate_2.A.n3 GND 0.0917f
C7562 Nand_Gate_2.A.t1 GND 0.08197f
C7563 Nand_Gate_2.A.n4 GND 0.35696f
C7564 Nand_Gate_2.A.n5 GND 0.0885f
C7565 Nand_Gate_2.A.t16 GND 0.62847f
C7566 Nand_Gate_2.A.n6 GND 0.61763f
C7567 Nand_Gate_2.A.n7 GND 0.06751f
C7568 Nand_Gate_2.A.t17 GND 0.32674f
C7569 Nand_Gate_2.A.n8 GND 0.09412f
C7570 Nand_Gate_2.A.n9 GND 0.04034f
C7571 Nand_Gate_2.A.n10 GND 0.07558f
C7572 Nand_Gate_2.A.n11 GND 0.09511f
C7573 Nand_Gate_2.A.t4 GND 0.62847f
C7574 Nand_Gate_2.A.n12 GND 0.61763f
C7575 Nand_Gate_2.A.n13 GND 0.06751f
C7576 Nand_Gate_2.A.t15 GND 0.32674f
C7577 Nand_Gate_2.A.n14 GND 0.09412f
C7578 Nand_Gate_2.A.n15 GND 0.04034f
C7579 Nand_Gate_2.A.n16 GND 0.07558f
C7580 Nand_Gate_2.A.n17 GND 0.01133f
C7581 Nand_Gate_2.A.n18 GND 0.28519f
C7582 Nand_Gate_2.A.n19 GND 0.79416f
C7583 Nand_Gate_2.A.n20 GND 0.35636f
C7584 Nand_Gate_2.A.t6 GND 0.62847f
C7585 Nand_Gate_2.A.n21 GND 0.6329f
C7586 Nand_Gate_2.A.n22 GND 0.06751f
C7587 Nand_Gate_2.A.t9 GND 0.32674f
C7588 Nand_Gate_2.A.n23 GND 0.09412f
C7589 Nand_Gate_2.A.n24 GND 0.02507f
C7590 Nand_Gate_2.A.n25 GND 0.03906f
C7591 Nand_Gate_2.A.n26 GND 0.38975f
C7592 Nand_Gate_2.A.t10 GND 0.62847f
C7593 Nand_Gate_2.A.n27 GND 0.6329f
C7594 Nand_Gate_2.A.n28 GND 0.06751f
C7595 Nand_Gate_2.A.t5 GND 0.32674f
C7596 Nand_Gate_2.A.n29 GND 0.09412f
C7597 Nand_Gate_2.A.n30 GND 0.02507f
C7598 Nand_Gate_2.A.n31 GND 0.03906f
C7599 Nand_Gate_2.A.n32 GND 0.01133f
C7600 Nand_Gate_2.A.n33 GND 1.01202f
C7601 Nand_Gate_2.A.n34 GND 0.47041f
C7602 Nand_Gate_2.A.n35 GND 0.17479f
C7603 Nand_Gate_2.A.t13 GND 0.62844f
C7604 Nand_Gate_2.A.n36 GND 0.18359f
C7605 Nand_Gate_2.A.n37 GND 0.07966f
C7606 Nand_Gate_2.A.n38 GND 0.35024f
C7607 Nand_Gate_2.A.t7 GND 0.29227f
C7608 Nand_Gate_2.A.n39 GND 0.03875f
C7609 Nand_Gate_2.A.n40 GND 0.09293f
C7610 Nand_Gate_2.A.n41 GND 8.01087f
C7611 Nand_Gate_2.A.t14 GND 0.32676f
C7612 Nand_Gate_2.A.n42 GND 0.32008f
C7613 Nand_Gate_2.A.n43 GND 0.06751f
C7614 Nand_Gate_2.A.t12 GND 0.62844f
C7615 Nand_Gate_2.A.n44 GND 0.18359f
C7616 Nand_Gate_2.A.n45 GND 0.04568f
C7617 Nand_Gate_2.A.n46 GND 0.06645f
C7618 Nand_Gate_2.A.n47 GND 0.09785f
C7619 Nand_Gate_2.A.n48 GND 9.45741f
C7620 Nand_Gate_2.A.n49 GND 0.34581f
C7621 Nand_Gate_2.A.n50 GND 0.10108f
C7622 Nand_Gate_2.A.n51 GND 0.0372f
C7623 Nand_Gate_2.A.n52 GND 0.01151f
C7624 Nand_Gate_2.A.n53 GND 0.10205f
C7625 Nand_Gate_2.A.n54 GND 0.05153f
C7626 Nand_Gate_2.A.t3 GND 0.08702f
C7627 Nand_Gate_2.A.t0 GND 0.08524f
C7628 Nand_Gate_2.A.n55 GND 0.48477f
C7629 Nand_Gate_2.A.n56 GND 0.15818f
C7630 Nand_Gate_2.A.t2 GND 0.08524f
C7631 Nand_Gate_2.A.n57 GND 0.13131f
C7632 Nand_Gate_2.A.n58 GND 0.2325f
C7633 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 GND 0.07024f
C7634 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 GND 0.03989f
C7635 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 GND 0.07725f
C7636 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 GND 0.2799f
C7637 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 GND 0.27418f
C7638 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 GND 0.05783f
C7639 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 GND 0.53832f
C7640 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 GND 0.15726f
C7641 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 GND 0.03913f
C7642 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 GND 0.05692f
C7643 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 GND 0.14585f
C7644 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 GND 0.14585f
C7645 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 GND 0.07581f
C7646 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 GND 0.07318f
C7647 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 GND 0.07454f
C7648 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 GND 0.07302f
C7649 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 GND 0.41525f
C7650 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 GND 0.23391f
C7651 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 GND 0.22303f
C7652 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 GND 0.06624f
C7653 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 GND 0.07883f
C7654 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 GND 0.39844f
C7655 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 GND 0.20187f
C7656 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 GND 0.06862f
C7657 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 GND 0.25335f
C7658 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 GND 0.24817f
C7659 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 GND 0.05234f
C7660 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 GND 0.48726f
C7661 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 GND 0.14234f
C7662 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 GND 0.03542f
C7663 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 GND 0.05152f
C7664 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 GND 0.13202f
C7665 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 GND 0.13202f
C7666 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 GND 0.06992f
C7667 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 GND 0.03611f
C7668 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 GND 0.06358f
C7669 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 GND 0.04998f
C7670 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 GND 0.02839f
C7671 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 GND 0.05497f
C7672 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 GND 0.38308f
C7673 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 GND 0.39717f
C7674 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 GND 0.04297f
C7675 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 GND 0.05737f
C7676 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 GND 0.30118f
C7677 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 GND 0.30119f
C7678 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 GND 0.1951f
C7679 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 GND 0.04115f
C7680 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 GND 0.38306f
C7681 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 GND 0.1119f
C7682 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 GND 0.02784f
C7683 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 GND 0.0405f
C7684 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 GND 0.10379f
C7685 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 GND 0.10379f
C7686 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 GND 0.05395f
C7687 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 GND 0.05208f
C7688 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 GND 0.30868f
C7689 Nand_Gate_0.A.t9 GND 0.75629f
C7690 Nand_Gate_0.A.n0 GND 0.22093f
C7691 Nand_Gate_0.A.n1 GND 0.09586f
C7692 Nand_Gate_0.A.n2 GND 0.42149f
C7693 Nand_Gate_0.A.t13 GND 0.35177f
C7694 Nand_Gate_0.A.n3 GND 0.11036f
C7695 Nand_Gate_0.A.t1 GND 0.09865f
C7696 Nand_Gate_0.A.n4 GND 0.42957f
C7697 Nand_Gate_0.A.n5 GND 0.10651f
C7698 Nand_Gate_0.A.t14 GND 0.75632f
C7699 Nand_Gate_0.A.n6 GND 0.74327f
C7700 Nand_Gate_0.A.n7 GND 0.08124f
C7701 Nand_Gate_0.A.t8 GND 0.39321f
C7702 Nand_Gate_0.A.n8 GND 0.11327f
C7703 Nand_Gate_0.A.n9 GND 0.04854f
C7704 Nand_Gate_0.A.n10 GND 0.09095f
C7705 Nand_Gate_0.A.n11 GND 0.11446f
C7706 Nand_Gate_0.A.t7 GND 0.75632f
C7707 Nand_Gate_0.A.n12 GND 0.74327f
C7708 Nand_Gate_0.A.n13 GND 0.08124f
C7709 Nand_Gate_0.A.t12 GND 0.39321f
C7710 Nand_Gate_0.A.n14 GND 0.11327f
C7711 Nand_Gate_0.A.n15 GND 0.04854f
C7712 Nand_Gate_0.A.n16 GND 0.09095f
C7713 Nand_Gate_0.A.n17 GND 0.01364f
C7714 Nand_Gate_0.A.n18 GND 0.34321f
C7715 Nand_Gate_0.A.n19 GND 0.95571f
C7716 Nand_Gate_0.A.n20 GND 0.42885f
C7717 Nand_Gate_0.A.t15 GND 0.75632f
C7718 Nand_Gate_0.A.n21 GND 0.76165f
C7719 Nand_Gate_0.A.n22 GND 0.08124f
C7720 Nand_Gate_0.A.t17 GND 0.39321f
C7721 Nand_Gate_0.A.n23 GND 0.11327f
C7722 Nand_Gate_0.A.n24 GND 0.03017f
C7723 Nand_Gate_0.A.n25 GND 0.04701f
C7724 Nand_Gate_0.A.n26 GND 0.46904f
C7725 Nand_Gate_0.A.t6 GND 0.75632f
C7726 Nand_Gate_0.A.n27 GND 0.76165f
C7727 Nand_Gate_0.A.n28 GND 0.08124f
C7728 Nand_Gate_0.A.t10 GND 0.39321f
C7729 Nand_Gate_0.A.n29 GND 0.11327f
C7730 Nand_Gate_0.A.n30 GND 0.03017f
C7731 Nand_Gate_0.A.n31 GND 0.04701f
C7732 Nand_Gate_0.A.n32 GND 0.01364f
C7733 Nand_Gate_0.A.n33 GND 1.2179f
C7734 Nand_Gate_0.A.n34 GND 0.5679f
C7735 Nand_Gate_0.A.n35 GND 0.21035f
C7736 Nand_Gate_0.A.t5 GND 0.75629f
C7737 Nand_Gate_0.A.n36 GND 0.22093f
C7738 Nand_Gate_0.A.n37 GND 0.09586f
C7739 Nand_Gate_0.A.n38 GND 0.42149f
C7740 Nand_Gate_0.A.t16 GND 0.35173f
C7741 Nand_Gate_0.A.n39 GND 0.04484f
C7742 Nand_Gate_0.A.n40 GND 0.10776f
C7743 Nand_Gate_0.A.n41 GND 14.747f
C7744 Nand_Gate_0.A.t11 GND 0.39323f
C7745 Nand_Gate_0.A.n42 GND 0.38519f
C7746 Nand_Gate_0.A.n43 GND 0.08124f
C7747 Nand_Gate_0.A.t4 GND 0.75629f
C7748 Nand_Gate_0.A.n44 GND 0.22093f
C7749 Nand_Gate_0.A.n45 GND 0.05497f
C7750 Nand_Gate_0.A.n46 GND 0.07997f
C7751 Nand_Gate_0.A.n47 GND 0.11775f
C7752 Nand_Gate_0.A.n48 GND 16.5226f
C7753 Nand_Gate_0.A.n49 GND 0.41616f
C7754 Nand_Gate_0.A.n50 GND 0.12165f
C7755 Nand_Gate_0.A.n51 GND 0.04477f
C7756 Nand_Gate_0.A.n52 GND 0.01385f
C7757 Nand_Gate_0.A.n53 GND 0.12281f
C7758 Nand_Gate_0.A.n54 GND 0.06202f
C7759 Nand_Gate_0.A.t3 GND 0.10473f
C7760 Nand_Gate_0.A.t0 GND 0.10258f
C7761 Nand_Gate_0.A.n55 GND 0.58338f
C7762 Nand_Gate_0.A.n56 GND 0.19036f
C7763 Nand_Gate_0.A.t2 GND 0.10258f
C7764 Nand_Gate_0.A.n57 GND 0.15802f
C7765 Nand_Gate_0.A.n58 GND 0.2798f
C7766 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 GND 0.05201f
C7767 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 GND 0.22649f
C7768 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 GND 0.05616f
C7769 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 GND 0.39877f
C7770 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 GND 0.39189f
C7771 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 GND 0.04283f
C7772 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 GND 0.20732f
C7773 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 GND 0.05972f
C7774 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 GND 0.02559f
C7775 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 GND 0.04796f
C7776 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 GND 0.10804f
C7777 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 GND 0.10804f
C7778 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 GND 0.06475f
C7779 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 GND 0.05421f
C7780 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 GND 0.05522f
C7781 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 GND 0.05409f
C7782 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 GND 0.30759f
C7783 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 GND 0.17406f
C7784 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 GND 0.03715f
C7785 Comparator_0.Vout GND 0.14103f
C7786 D_FlipFlop_7.D.t33 GND 1.14081f
C7787 D_FlipFlop_7.D.n0 GND 0.33301f
C7788 D_FlipFlop_7.D.t1 GND 4.00728f
C7789 D_FlipFlop_7.D.t2 GND 0.88528f
C7790 D_FlipFlop_7.D.n1 GND 3.0992f
C7791 D_FlipFlop_7.D.t0 GND 1.67549f
C7792 D_FlipFlop_7.D.n2 GND -7.39606f
C7793 D_FlipFlop_7.D.n3 GND 8.35956f
C7794 D_FlipFlop_7.D.n4 GND 2.50292f
C7795 D_FlipFlop_7.D.t20 GND 0.30279f
C7796 D_FlipFlop_0.Inverter_0.Vin GND -0.22043f
C7797 D_FlipFlop_7.D.n5 GND 0.29756f
C7798 D_FlipFlop_7.D.n6 GND 0.03252f
C7799 D_FlipFlop_7.D.t30 GND 0.15742f
C7800 D_FlipFlop_7.D.n7 GND 0.04535f
C7801 D_FlipFlop_7.D.n8 GND 0.01943f
C7802 D_FlipFlop_7.D.n9 GND 0.03641f
C7803 D_FlipFlop_7.D.t27 GND 0.30279f
C7804 D_FlipFlop_0.3-input-nand_0.B GND -0.22043f
C7805 D_FlipFlop_7.D.n11 GND 0.29756f
C7806 D_FlipFlop_7.D.n12 GND 0.03252f
C7807 D_FlipFlop_7.D.t23 GND 0.15742f
C7808 D_FlipFlop_7.D.n13 GND 0.04535f
C7809 D_FlipFlop_7.D.n14 GND 0.01943f
C7810 D_FlipFlop_7.D.n15 GND 0.03641f
C7811 D_FlipFlop_7.D.n16 GND 0.04561f
C7812 D_FlipFlop_7.D.n17 GND 0.27556f
C7813 D_FlipFlop_7.D.t31 GND 0.30279f
C7814 D_FlipFlop_3.Inverter_0.Vin GND -0.22043f
C7815 D_FlipFlop_7.D.n18 GND 0.29756f
C7816 D_FlipFlop_7.D.n19 GND 0.03252f
C7817 D_FlipFlop_7.D.t11 GND 0.15742f
C7818 D_FlipFlop_7.D.n20 GND 0.04535f
C7819 D_FlipFlop_7.D.n21 GND 0.01943f
C7820 D_FlipFlop_7.D.n22 GND 0.03641f
C7821 D_FlipFlop_7.D.t4 GND 0.30279f
C7822 D_FlipFlop_3.3-input-nand_0.B GND -0.22043f
C7823 D_FlipFlop_7.D.n24 GND 0.29756f
C7824 D_FlipFlop_7.D.n25 GND 0.03252f
C7825 D_FlipFlop_7.D.t32 GND 0.15742f
C7826 D_FlipFlop_7.D.n26 GND 0.04535f
C7827 D_FlipFlop_7.D.n27 GND 0.01943f
C7828 D_FlipFlop_7.D.n28 GND 0.03641f
C7829 D_FlipFlop_7.D.n29 GND 0.04561f
C7830 D_FlipFlop_7.D.n30 GND 0.14341f
C7831 D_FlipFlop_7.D.n31 GND 0.73537f
C7832 D_FlipFlop_7.D.t14 GND 0.30279f
C7833 D_FlipFlop_2.Inverter_0.Vin GND -0.22043f
C7834 D_FlipFlop_7.D.n32 GND 0.29756f
C7835 D_FlipFlop_7.D.n33 GND 0.03252f
C7836 D_FlipFlop_7.D.t17 GND 0.15742f
C7837 D_FlipFlop_7.D.n34 GND 0.04535f
C7838 D_FlipFlop_7.D.n35 GND 0.01943f
C7839 D_FlipFlop_7.D.n36 GND 0.03641f
C7840 D_FlipFlop_7.D.t24 GND 0.30279f
C7841 D_FlipFlop_2.3-input-nand_0.B GND -0.22043f
C7842 D_FlipFlop_7.D.n38 GND 0.29756f
C7843 D_FlipFlop_7.D.n39 GND 0.03252f
C7844 D_FlipFlop_7.D.t8 GND 0.15742f
C7845 D_FlipFlop_7.D.n40 GND 0.04535f
C7846 D_FlipFlop_7.D.n41 GND 0.01943f
C7847 D_FlipFlop_7.D.n42 GND 0.03641f
C7848 D_FlipFlop_7.D.n43 GND 0.04561f
C7849 D_FlipFlop_7.D.n44 GND 0.14341f
C7850 D_FlipFlop_7.D.n45 GND 0.57322f
C7851 D_FlipFlop_7.D.t19 GND 0.30279f
C7852 D_FlipFlop_1.Inverter_0.Vin GND -0.22043f
C7853 D_FlipFlop_7.D.n46 GND 0.29756f
C7854 D_FlipFlop_7.D.n47 GND 0.03252f
C7855 D_FlipFlop_7.D.t29 GND 0.15742f
C7856 D_FlipFlop_7.D.n48 GND 0.04535f
C7857 D_FlipFlop_7.D.n49 GND 0.01943f
C7858 D_FlipFlop_7.D.n50 GND 0.03641f
C7859 D_FlipFlop_7.D.t26 GND 0.30279f
C7860 D_FlipFlop_1.3-input-nand_0.B GND -0.22043f
C7861 D_FlipFlop_7.D.n52 GND 0.29756f
C7862 D_FlipFlop_7.D.n53 GND 0.03252f
C7863 D_FlipFlop_7.D.t22 GND 0.15742f
C7864 D_FlipFlop_7.D.n54 GND 0.04535f
C7865 D_FlipFlop_7.D.n55 GND 0.01943f
C7866 D_FlipFlop_7.D.n56 GND 0.03641f
C7867 D_FlipFlop_7.D.n57 GND 0.04561f
C7868 D_FlipFlop_7.D.n58 GND 0.14341f
C7869 D_FlipFlop_7.D.n59 GND 0.74234f
C7870 D_FlipFlop_7.D.t21 GND 0.30279f
C7871 D_FlipFlop_4.Inverter_0.Vin GND -0.22043f
C7872 D_FlipFlop_7.D.n60 GND 0.29756f
C7873 D_FlipFlop_7.D.n61 GND 0.03252f
C7874 D_FlipFlop_7.D.t13 GND 0.15742f
C7875 D_FlipFlop_7.D.n62 GND 0.04535f
C7876 D_FlipFlop_7.D.n63 GND 0.01943f
C7877 D_FlipFlop_7.D.n64 GND 0.03641f
C7878 D_FlipFlop_7.D.t28 GND 0.30279f
C7879 D_FlipFlop_4.3-input-nand_0.B GND -0.22043f
C7880 D_FlipFlop_7.D.n66 GND 0.29756f
C7881 D_FlipFlop_7.D.n67 GND 0.03252f
C7882 D_FlipFlop_7.D.t3 GND 0.15742f
C7883 D_FlipFlop_7.D.n68 GND 0.04535f
C7884 D_FlipFlop_7.D.n69 GND 0.01943f
C7885 D_FlipFlop_7.D.n70 GND 0.03641f
C7886 D_FlipFlop_7.D.n71 GND 0.04561f
C7887 D_FlipFlop_7.D.n72 GND 0.14341f
C7888 D_FlipFlop_7.D.n73 GND 0.74234f
C7889 D_FlipFlop_7.D.t5 GND 0.30279f
C7890 D_FlipFlop_5.Inverter_0.Vin GND -0.22043f
C7891 D_FlipFlop_7.D.n74 GND 0.29756f
C7892 D_FlipFlop_7.D.n75 GND 0.03252f
C7893 D_FlipFlop_7.D.t16 GND 0.15742f
C7894 D_FlipFlop_7.D.n76 GND 0.04535f
C7895 D_FlipFlop_7.D.n77 GND 0.01943f
C7896 D_FlipFlop_7.D.n78 GND 0.03641f
C7897 D_FlipFlop_7.D.t10 GND 0.30279f
C7898 D_FlipFlop_5.3-input-nand_0.B GND -0.22043f
C7899 D_FlipFlop_7.D.n80 GND 0.29756f
C7900 D_FlipFlop_7.D.n81 GND 0.03252f
C7901 D_FlipFlop_7.D.t7 GND 0.15742f
C7902 D_FlipFlop_7.D.n82 GND 0.04535f
C7903 D_FlipFlop_7.D.n83 GND 0.01943f
C7904 D_FlipFlop_7.D.n84 GND 0.03641f
C7905 D_FlipFlop_7.D.n85 GND 0.04561f
C7906 D_FlipFlop_7.D.n86 GND 0.14341f
C7907 D_FlipFlop_7.D.t34 GND 0.30279f
C7908 D_FlipFlop_7.Inverter_0.Vin GND -0.22043f
C7909 D_FlipFlop_7.D.n87 GND 0.29756f
C7910 D_FlipFlop_7.D.n88 GND 0.03252f
C7911 D_FlipFlop_7.D.t12 GND 0.15742f
C7912 D_FlipFlop_7.D.n89 GND 0.04535f
C7913 D_FlipFlop_7.D.n90 GND 0.01943f
C7914 D_FlipFlop_7.D.n91 GND 0.03641f
C7915 D_FlipFlop_7.D.t6 GND 0.30279f
C7916 D_FlipFlop_7.3-input-nand_0.B GND -0.22043f
C7917 D_FlipFlop_7.D.n93 GND 0.29756f
C7918 D_FlipFlop_7.D.n94 GND 0.03252f
C7919 D_FlipFlop_7.D.t35 GND 0.15742f
C7920 D_FlipFlop_7.D.n95 GND 0.04535f
C7921 D_FlipFlop_7.D.n96 GND 0.01943f
C7922 D_FlipFlop_7.D.n97 GND 0.03641f
C7923 D_FlipFlop_7.D.n98 GND 0.04561f
C7924 D_FlipFlop_7.D.n99 GND 0.27556f
C7925 D_FlipFlop_7.D.t15 GND 0.30279f
C7926 D_FlipFlop_6.Inverter_0.Vin GND -0.22043f
C7927 D_FlipFlop_7.D.n100 GND 0.29756f
C7928 D_FlipFlop_7.D.n101 GND 0.03252f
C7929 D_FlipFlop_7.D.t18 GND 0.15742f
C7930 D_FlipFlop_7.D.n102 GND 0.04535f
C7931 D_FlipFlop_7.D.n103 GND 0.01943f
C7932 D_FlipFlop_7.D.n104 GND 0.03641f
C7933 D_FlipFlop_7.D.t25 GND 0.30279f
C7934 D_FlipFlop_6.3-input-nand_0.B GND -0.22043f
C7935 D_FlipFlop_7.D.n106 GND 0.29756f
C7936 D_FlipFlop_7.D.n107 GND 0.03252f
C7937 D_FlipFlop_7.D.t9 GND 0.15742f
C7938 D_FlipFlop_7.D.n108 GND 0.04535f
C7939 D_FlipFlop_7.D.n109 GND 0.01943f
C7940 D_FlipFlop_7.D.n110 GND 0.03641f
C7941 D_FlipFlop_7.D.n111 GND 0.04561f
C7942 D_FlipFlop_7.D.n112 GND 0.14341f
C7943 D_FlipFlop_7.D.n113 GND 0.73537f
C7944 D_FlipFlop_7.D.n114 GND 0.67663f
C7945 D_FlipFlop_7.D.n115 GND 2.25004f
C7946 D_FlipFlop_7.D.n116 GND 1.03924f
C7947 D_FlipFlop_1.3-input-nand_2.C.t1 GND 0.04477f
C7948 D_FlipFlop_1.3-input-nand_2.C.n0 GND 0.11971f
C7949 D_FlipFlop_1.3-input-nand_2.C.n1 GND 0.09193f
C7950 D_FlipFlop_1.3-input-nand_2.C.t4 GND 0.17806f
C7951 D_FlipFlop_1.3-input-nand_2.C.t5 GND 0.34248f
C7952 D_FlipFlop_1.3-input-nand_2.C.n2 GND 0.10005f
C7953 D_FlipFlop_1.3-input-nand_2.C.n3 GND 0.04279f
C7954 D_FlipFlop_1.3-input-nand_2.C.n4 GND 0.079f
C7955 D_FlipFlop_1.3-input-nand_2.C.n5 GND 0.13677f
C7956 D_FlipFlop_1.3-input-nand_2.C.n6 GND 0.10181f
C7957 D_FlipFlop_1.3-input-nand_2.C.n7 GND 0.04823f
C7958 D_FlipFlop_1.3-input-nand_2.C.t6 GND 0.3425f
C7959 D_FlipFlop_1.3-input-nand_2.C.n8 GND 0.3551f
C7960 D_FlipFlop_1.3-input-nand_2.C.n9 GND 0.03842f
C7961 D_FlipFlop_1.3-input-nand_2.C.n10 GND 0.05129f
C7962 D_FlipFlop_1.3-input-nand_2.C.t7 GND 0.17045f
C7963 D_FlipFlop_1.3-input-nand_2.C.t0 GND 0.04645f
C7964 D_FlipFlop_1.3-input-nand_2.C.n11 GND 0.293f
C7965 D_FlipFlop_1.3-input-nand_2.C.t2 GND 0.04742f
C7966 D_FlipFlop_1.3-input-nand_2.C.t3 GND 0.04645f
C7967 D_FlipFlop_1.3-input-nand_2.C.n12 GND 0.26418f
C7968 D_FlipFlop_1.3-input-nand_2.C.n13 GND 0.08722f
C7969 D_FlipFlop_1.3-input-nand_2.C.n14 GND 0.124f
C7970 D_FlipFlop_1.3-input-nand_2.Vout.t6 GND 0.35515f
C7971 D_FlipFlop_1.3-input-nand_2.Vout.n0 GND 0.10375f
C7972 D_FlipFlop_1.3-input-nand_2.Vout.n1 GND 0.04502f
C7973 D_FlipFlop_1.3-input-nand_2.Vout.t1 GND 0.04632f
C7974 D_FlipFlop_1.3-input-nand_2.Vout.n2 GND 0.22028f
C7975 D_FlipFlop_1.3-input-nand_2.Vout.n3 GND 0.05002f
C7976 D_FlipFlop_1.3-input-nand_2.Vout.t5 GND 0.35517f
C7977 D_FlipFlop_1.3-input-nand_2.Vout.n4 GND 0.36759f
C7978 D_FlipFlop_1.3-input-nand_2.Vout.t7 GND 0.18465f
C7979 D_FlipFlop_1.3-input-nand_2.Vout.n5 GND 0.18106f
C7980 D_FlipFlop_1.3-input-nand_2.Vout.n6 GND 0.10557f
C7981 D_FlipFlop_1.3-input-nand_2.Vout.n7 GND 0.01331f
C7982 D_FlipFlop_1.3-input-nand_2.Vout.n8 GND 0.01454f
C7983 D_FlipFlop_1.3-input-nand_2.Vout.t3 GND 0.04918f
C7984 D_FlipFlop_1.3-input-nand_2.Vout.t0 GND 0.04817f
C7985 D_FlipFlop_1.3-input-nand_2.Vout.n9 GND 0.27396f
C7986 D_FlipFlop_1.3-input-nand_2.Vout.n10 GND 0.09115f
C7987 D_FlipFlop_1.3-input-nand_2.Vout.t2 GND 0.04817f
C7988 D_FlipFlop_1.3-input-nand_2.Vout.n11 GND 0.30324f
C7989 D_FlipFlop_1.3-input-nand_2.Vout.t4 GND 0.17747f
C7990 D_FlipFlop_1.3-input-nand_2.Vout.n12 GND 0.19793f
C7991 CDAC8_0.switch_6.Z.t2 GND 0.03493f
C7992 CDAC8_0.switch_6.Z.t3 GND 0.0333f
C7993 CDAC8_0.switch_6.Z.t1 GND 0.0333f
C7994 CDAC8_0.switch_6.Z.n0 GND 0.1203f
C7995 CDAC8_0.switch_6.Z.n1 GND 0.27648f
C7996 CDAC8_0.switch_6.Z.n2 GND 0.03601f
C7997 CDAC8_0.switch_6.Z.n3 GND 1.50056f
C7998 CDAC8_0.switch_6.Z.n4 GND 1.08953f
C7999 CDAC8_0.switch_6.Z.t41 GND 5.88261f
C8000 CDAC8_0.switch_6.Z.n5 GND 1.36404f
C8001 CDAC8_0.switch_6.Z.t10 GND 5.88261f
C8002 CDAC8_0.switch_6.Z.n6 GND 1.36404f
C8003 CDAC8_0.switch_6.Z.t29 GND 5.88261f
C8004 CDAC8_0.switch_6.Z.n7 GND 1.36404f
C8005 CDAC8_0.switch_6.Z.t63 GND 5.96794f
C8006 CDAC8_0.switch_6.Z.t32 GND 5.96794f
C8007 CDAC8_0.switch_6.Z.n8 GND 2.23974f
C8008 CDAC8_0.switch_6.Z.n9 GND 2.23974f
C8009 CDAC8_0.switch_6.Z.t62 GND 5.88261f
C8010 CDAC8_0.switch_6.Z.n10 GND 1.36404f
C8011 CDAC8_0.switch_6.Z.n11 GND 1.12959f
C8012 CDAC8_0.switch_6.Z.n12 GND 1.12959f
C8013 CDAC8_0.switch_6.Z.t45 GND 5.88261f
C8014 CDAC8_0.switch_6.Z.n13 GND 1.36404f
C8015 CDAC8_0.switch_6.Z.n14 GND 1.12959f
C8016 CDAC8_0.switch_6.Z.n15 GND 1.12959f
C8017 CDAC8_0.switch_6.Z.t7 GND 5.88261f
C8018 CDAC8_0.switch_6.Z.n16 GND 1.36404f
C8019 CDAC8_0.switch_6.Z.t34 GND 5.88261f
C8020 CDAC8_0.switch_6.Z.n17 GND 1.36404f
C8021 CDAC8_0.switch_6.Z.n18 GND 1.12959f
C8022 CDAC8_0.switch_6.Z.n19 GND 1.12959f
C8023 CDAC8_0.switch_6.Z.t67 GND 5.88261f
C8024 CDAC8_0.switch_6.Z.n20 GND 1.36404f
C8025 CDAC8_0.switch_6.Z.t9 GND 5.88261f
C8026 CDAC8_0.switch_6.Z.n21 GND 1.36404f
C8027 CDAC8_0.switch_6.Z.t46 GND 5.88261f
C8028 CDAC8_0.switch_6.Z.n22 GND 1.36404f
C8029 CDAC8_0.switch_6.Z.t53 GND 5.88261f
C8030 CDAC8_0.switch_6.Z.n23 GND 1.36404f
C8031 CDAC8_0.switch_6.Z.t17 GND 5.88261f
C8032 CDAC8_0.switch_6.Z.n24 GND 1.36404f
C8033 CDAC8_0.switch_6.Z.t15 GND 5.88261f
C8034 CDAC8_0.switch_6.Z.n25 GND 1.36404f
C8035 CDAC8_0.switch_6.Z.t58 GND 5.88261f
C8036 CDAC8_0.switch_6.Z.n26 GND 1.36404f
C8037 CDAC8_0.switch_6.Z.t22 GND 5.88261f
C8038 CDAC8_0.switch_6.Z.n27 GND 1.36404f
C8039 CDAC8_0.switch_6.Z.t65 GND 5.88261f
C8040 CDAC8_0.switch_6.Z.n28 GND 1.36404f
C8041 CDAC8_0.switch_6.Z.t61 GND 5.88261f
C8042 CDAC8_0.switch_6.Z.n29 GND 1.36404f
C8043 CDAC8_0.switch_6.Z.t25 GND 5.88261f
C8044 CDAC8_0.switch_6.Z.n30 GND 1.36404f
C8045 CDAC8_0.switch_6.Z.t5 GND 6.12449f
C8046 CDAC8_0.switch_6.Z.t37 GND 6.12449f
C8047 CDAC8_0.switch_6.Z.n31 GND 2.41525f
C8048 CDAC8_0.switch_6.Z.n32 GND 2.41525f
C8049 CDAC8_0.switch_6.Z.t59 GND 5.88261f
C8050 CDAC8_0.switch_6.Z.n33 GND 1.36404f
C8051 CDAC8_0.switch_6.Z.n34 GND 1.12959f
C8052 CDAC8_0.switch_6.Z.n35 GND 1.12959f
C8053 CDAC8_0.switch_6.Z.t27 GND 5.88261f
C8054 CDAC8_0.switch_6.Z.n36 GND 1.36404f
C8055 CDAC8_0.switch_6.Z.n37 GND 1.12959f
C8056 CDAC8_0.switch_6.Z.n38 GND 1.12959f
C8057 CDAC8_0.switch_6.Z.t33 GND 5.88261f
C8058 CDAC8_0.switch_6.Z.n39 GND 1.36404f
C8059 CDAC8_0.switch_6.Z.n40 GND 1.12959f
C8060 CDAC8_0.switch_6.Z.n41 GND 1.12959f
C8061 CDAC8_0.switch_6.Z.t56 GND 5.88261f
C8062 CDAC8_0.switch_6.Z.n42 GND 1.24121f
C8063 CDAC8_0.switch_6.Z.n43 GND 0.7957f
C8064 CDAC8_0.switch_6.Z.t13 GND 5.88261f
C8065 CDAC8_0.switch_6.Z.n44 GND 1.36404f
C8066 CDAC8_0.switch_6.Z.t48 GND 5.88261f
C8067 CDAC8_0.switch_6.Z.n45 GND 1.36404f
C8068 CDAC8_0.switch_6.Z.t30 GND 5.88261f
C8069 CDAC8_0.switch_6.Z.n46 GND 1.36404f
C8070 CDAC8_0.switch_6.Z.t19 GND 5.88261f
C8071 CDAC8_0.switch_6.Z.n47 GND 1.36404f
C8072 CDAC8_0.switch_6.Z.t18 GND 5.88261f
C8073 CDAC8_0.switch_6.Z.n48 GND 1.36404f
C8074 CDAC8_0.switch_6.Z.t11 GND 5.88261f
C8075 CDAC8_0.switch_6.Z.n49 GND 1.36404f
C8076 CDAC8_0.switch_6.Z.t52 GND 5.88261f
C8077 CDAC8_0.switch_6.Z.n50 GND 1.36404f
C8078 CDAC8_0.switch_6.Z.t44 GND 5.88261f
C8079 CDAC8_0.switch_6.Z.n51 GND 1.36404f
C8080 CDAC8_0.switch_6.Z.t43 GND 5.88261f
C8081 CDAC8_0.switch_6.Z.n52 GND 1.36404f
C8082 CDAC8_0.switch_6.Z.t31 GND 5.96794f
C8083 CDAC8_0.switch_6.Z.t47 GND 5.96794f
C8084 CDAC8_0.switch_6.Z.n53 GND 2.23974f
C8085 CDAC8_0.switch_6.Z.n54 GND 2.23974f
C8086 CDAC8_0.switch_6.Z.t28 GND 5.88261f
C8087 CDAC8_0.switch_6.Z.n55 GND 1.36404f
C8088 CDAC8_0.switch_6.Z.n56 GND 1.12959f
C8089 CDAC8_0.switch_6.Z.n57 GND 1.12959f
C8090 CDAC8_0.switch_6.Z.t54 GND 5.88261f
C8091 CDAC8_0.switch_6.Z.n58 GND 1.36404f
C8092 CDAC8_0.switch_6.Z.n59 GND 1.24989f
C8093 CDAC8_0.switch_6.Z.n60 GND 1.24989f
C8094 CDAC8_0.switch_6.Z.t40 GND 5.88261f
C8095 CDAC8_0.switch_6.Z.n61 GND 1.36404f
C8096 CDAC8_0.switch_6.Z.n62 GND 1.08953f
C8097 CDAC8_0.switch_6.Z.t66 GND 5.88261f
C8098 CDAC8_0.switch_6.Z.n63 GND 1.36404f
C8099 CDAC8_0.switch_6.Z.n64 GND 1.12959f
C8100 CDAC8_0.switch_6.Z.n65 GND 1.12959f
C8101 CDAC8_0.switch_6.Z.t14 GND 5.88261f
C8102 CDAC8_0.switch_6.Z.n66 GND 1.36404f
C8103 CDAC8_0.switch_6.Z.n67 GND 0.6433f
C8104 CDAC8_0.switch_6.Z.t21 GND 5.88261f
C8105 CDAC8_0.switch_6.Z.n68 GND 1.36404f
C8106 CDAC8_0.switch_6.Z.n69 GND 1.12959f
C8107 CDAC8_0.switch_6.Z.n70 GND 1.12959f
C8108 CDAC8_0.switch_6.Z.t8 GND 5.88261f
C8109 CDAC8_0.switch_6.Z.n71 GND 1.36404f
C8110 CDAC8_0.switch_6.Z.n72 GND 1.12959f
C8111 CDAC8_0.switch_6.Z.n73 GND 1.12959f
C8112 CDAC8_0.switch_6.Z.t35 GND 5.88261f
C8113 CDAC8_0.switch_6.Z.n74 GND 1.36404f
C8114 CDAC8_0.switch_6.Z.n75 GND 1.12959f
C8115 CDAC8_0.switch_6.Z.n76 GND 1.12959f
C8116 CDAC8_0.switch_6.Z.t16 GND 5.88261f
C8117 CDAC8_0.switch_6.Z.n77 GND 1.36404f
C8118 CDAC8_0.switch_6.Z.n78 GND 1.12959f
C8119 CDAC8_0.switch_6.Z.n79 GND 1.12959f
C8120 CDAC8_0.switch_6.Z.t60 GND 5.88261f
C8121 CDAC8_0.switch_6.Z.n80 GND 1.36404f
C8122 CDAC8_0.switch_6.Z.t6 GND 5.88261f
C8123 CDAC8_0.switch_6.Z.n81 GND 1.36404f
C8124 CDAC8_0.switch_6.Z.n82 GND 1.12959f
C8125 CDAC8_0.switch_6.Z.n83 GND 1.12959f
C8126 CDAC8_0.switch_6.Z.t57 GND 5.88261f
C8127 CDAC8_0.switch_6.Z.n84 GND 1.36404f
C8128 CDAC8_0.switch_6.Z.n85 GND 1.12959f
C8129 CDAC8_0.switch_6.Z.t55 GND 5.88261f
C8130 CDAC8_0.switch_6.Z.n86 GND 1.36404f
C8131 CDAC8_0.switch_6.Z.t26 GND 5.88261f
C8132 CDAC8_0.switch_6.Z.n87 GND 1.36404f
C8133 CDAC8_0.switch_6.Z.t38 GND 5.88261f
C8134 CDAC8_0.switch_6.Z.n88 GND 1.36404f
C8135 CDAC8_0.switch_6.Z.t36 GND 6.12449f
C8136 CDAC8_0.switch_6.Z.t50 GND 6.12449f
C8137 CDAC8_0.switch_6.Z.n89 GND 2.41525f
C8138 CDAC8_0.switch_6.Z.n90 GND 2.41525f
C8139 CDAC8_0.switch_6.Z.t24 GND 5.88261f
C8140 CDAC8_0.switch_6.Z.n91 GND 1.36404f
C8141 CDAC8_0.switch_6.Z.n92 GND 1.12959f
C8142 CDAC8_0.switch_6.Z.n93 GND 1.12959f
C8143 CDAC8_0.switch_6.Z.t39 GND 5.88261f
C8144 CDAC8_0.switch_6.Z.n94 GND 1.36404f
C8145 CDAC8_0.switch_6.Z.n95 GND 1.12959f
C8146 CDAC8_0.switch_6.Z.n96 GND 1.12959f
C8147 CDAC8_0.switch_6.Z.t64 GND 5.88261f
C8148 CDAC8_0.switch_6.Z.n97 GND 1.36404f
C8149 CDAC8_0.switch_6.Z.n98 GND 1.12959f
C8150 CDAC8_0.switch_6.Z.n99 GND 1.12959f
C8151 CDAC8_0.switch_6.Z.t4 GND 5.88261f
C8152 CDAC8_0.switch_6.Z.n100 GND 1.24121f
C8153 CDAC8_0.switch_6.Z.n101 GND 2.49363f
C8154 CDAC8_0.switch_6.Z.n102 GND 2.49363f
C8155 CDAC8_0.switch_6.Z.n103 GND 0.7957f
C8156 CDAC8_0.switch_6.Z.n104 GND 1.12959f
C8157 CDAC8_0.switch_6.Z.t23 GND 5.88261f
C8158 CDAC8_0.switch_6.Z.n105 GND 1.36404f
C8159 CDAC8_0.switch_6.Z.n106 GND 1.12959f
C8160 CDAC8_0.switch_6.Z.n107 GND 1.12959f
C8161 CDAC8_0.switch_6.Z.t49 GND 5.88261f
C8162 CDAC8_0.switch_6.Z.n108 GND 1.36404f
C8163 CDAC8_0.switch_6.Z.n109 GND 1.12959f
C8164 CDAC8_0.switch_6.Z.n110 GND 1.12959f
C8165 CDAC8_0.switch_6.Z.t51 GND 5.88261f
C8166 CDAC8_0.switch_6.Z.n111 GND 1.36404f
C8167 CDAC8_0.switch_6.Z.n112 GND 1.12959f
C8168 CDAC8_0.switch_6.Z.n113 GND 1.12959f
C8169 CDAC8_0.switch_6.Z.t20 GND 5.88261f
C8170 CDAC8_0.switch_6.Z.n114 GND 1.36404f
C8171 CDAC8_0.switch_6.Z.n115 GND 1.12959f
C8172 CDAC8_0.switch_6.Z.n116 GND 1.12959f
C8173 CDAC8_0.switch_6.Z.t42 GND 5.88261f
C8174 CDAC8_0.switch_6.Z.n117 GND 1.36404f
C8175 CDAC8_0.switch_6.Z.n118 GND 1.12959f
C8176 CDAC8_0.switch_6.Z.n119 GND 1.12959f
C8177 CDAC8_0.switch_6.Z.t12 GND 5.88261f
C8178 CDAC8_0.switch_6.Z.n120 GND 1.36404f
C8179 CDAC8_0.switch_6.Z.n121 GND 0.6433f
C8180 CDAC8_0.switch_6.Z.n122 GND 1.45909f
C8181 CDAC8_0.switch_6.Z.n123 GND 1.93832f
C8182 CDAC8_0.switch_6.Z.n124 GND 0.01787f
C8183 CDAC8_0.switch_6.Z.t0 GND 0.03493f
C8184 CDAC8_0.switch_6.Z.n125 GND 0.14424f
C8185 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 GND 0.06323f
C8186 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 GND 0.07525f
C8187 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 GND 0.38033f
C8188 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 GND 0.1927f
C8189 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 GND 0.0655f
C8190 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 GND 0.24183f
C8191 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 GND 0.23689f
C8192 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 GND 0.04996f
C8193 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 GND 0.46511f
C8194 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 GND 0.13587f
C8195 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 GND 0.03381f
C8196 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 GND 0.04918f
C8197 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 GND 0.12602f
C8198 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 GND 0.12602f
C8199 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 GND 0.06674f
C8200 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 GND 0.0608f
C8201 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 GND 0.13827f
C8202 CDAC8_0.switch_8.Z.t2 GND 0.03182f
C8203 CDAC8_0.switch_8.Z.t1 GND 0.03182f
C8204 CDAC8_0.switch_8.Z.n0 GND 0.11498f
C8205 CDAC8_0.switch_8.Z.n1 GND 0.24282f
C8206 CDAC8_0.switch_8.Z.n2 GND 0.03442f
C8207 CDAC8_0.switch_8.Z.t14 GND 5.70386f
C8208 CDAC8_0.switch_8.Z.n3 GND 1.9642f
C8209 CDAC8_0.switch_8.Z.t6 GND 5.70386f
C8210 CDAC8_0.switch_8.Z.t4 GND 5.9531f
C8211 CDAC8_0.switch_8.Z.t17 GND 5.62231f
C8212 CDAC8_0.switch_8.Z.n4 GND 3.16681f
C8213 CDAC8_0.switch_8.Z.t19 GND 5.62231f
C8214 CDAC8_0.switch_8.Z.n5 GND 1.91851f
C8215 CDAC8_0.switch_8.Z.t15 GND 5.62231f
C8216 CDAC8_0.switch_8.Z.n6 GND 1.91851f
C8217 CDAC8_0.switch_8.Z.t9 GND 5.62231f
C8218 CDAC8_0.switch_8.Z.n7 GND 1.6228f
C8219 CDAC8_0.switch_8.Z.t13 GND 5.62231f
C8220 CDAC8_0.switch_8.Z.n8 GND 1.74019f
C8221 CDAC8_0.switch_8.Z.t18 GND 5.62231f
C8222 CDAC8_0.switch_8.Z.n9 GND 1.59939f
C8223 CDAC8_0.switch_8.Z.t12 GND 5.9531f
C8224 CDAC8_0.switch_8.Z.t8 GND 5.62231f
C8225 CDAC8_0.switch_8.Z.n10 GND 3.16681f
C8226 CDAC8_0.switch_8.Z.t10 GND 5.62231f
C8227 CDAC8_0.switch_8.Z.n11 GND 1.91851f
C8228 CDAC8_0.switch_8.Z.t7 GND 5.62231f
C8229 CDAC8_0.switch_8.Z.n12 GND 1.91851f
C8230 CDAC8_0.switch_8.Z.t16 GND 5.62231f
C8231 CDAC8_0.switch_8.Z.n13 GND 1.6228f
C8232 CDAC8_0.switch_8.Z.n14 GND 1.12092f
C8233 CDAC8_0.switch_8.Z.n15 GND 1.12092f
C8234 CDAC8_0.switch_8.Z.t11 GND 5.62231f
C8235 CDAC8_0.switch_8.Z.n16 GND 1.59939f
C8236 CDAC8_0.switch_8.Z.t5 GND 5.62231f
C8237 CDAC8_0.switch_8.Z.n17 GND 1.74019f
C8238 CDAC8_0.switch_8.Z.n18 GND 1.92246f
C8239 CDAC8_0.switch_8.Z.n19 GND 0.48531f
C8240 CDAC8_0.switch_8.Z.n20 GND 0.01245f
C8241 CDAC8_0.switch_8.Z.n21 GND 0.0507f
C8242 CDAC8_0.switch_8.Z.t3 GND 0.03342f
C8243 CDAC8_0.switch_8.Z.n22 GND 0.09316f
C8244 CDAC8_0.switch_8.Z.t0 GND 0.0334f
C8245 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 GND 0.07037f
C8246 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 GND 0.16004f
C8247 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 GND 0.07725f
C8248 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 GND 0.2799f
C8249 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 GND 0.27418f
C8250 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 GND 0.05783f
C8251 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 GND 0.53832f
C8252 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 GND 0.15726f
C8253 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 GND 0.03913f
C8254 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 GND 0.05692f
C8255 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 GND 0.14585f
C8256 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 GND 0.14585f
C8257 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 GND 0.07581f
C8258 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 GND 0.07318f
C8259 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 GND 0.07454f
C8260 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 GND 0.07302f
C8261 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 GND 0.41525f
C8262 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 GND 0.23391f
C8263 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 GND 0.22303f
C8264 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 GND 0.45666f
C8265 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 GND 0.47347f
C8266 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 GND 0.05122f
C8267 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 GND 0.05958f
C8268 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 GND 0.0577f
C8269 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 GND 0.12257f
C8270 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 GND 0.23742f
C8271 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 GND 0.45664f
C8272 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 GND 0.1334f
C8273 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 GND 0.05705f
C8274 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 GND 0.10533f
C8275 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 GND 0.18236f
C8276 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 GND 0.13574f
C8277 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 GND 0.06431f
C8278 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 GND 0.16533f
C8279 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 GND 0.06323f
C8280 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 GND 0.06194f
C8281 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 GND 0.35224f
C8282 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 GND 0.11629f
C8283 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 GND 0.06194f
C8284 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 GND 0.39067f
C8285 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 GND 0.22727f
C8286 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 GND 0.06839f
C8287 D_FlipFlop_6.3-input-nand_2.C.t6 GND 0.3425f
C8288 D_FlipFlop_6.3-input-nand_2.C.n0 GND 0.3551f
C8289 D_FlipFlop_6.3-input-nand_2.C.n1 GND 0.03842f
C8290 D_FlipFlop_6.3-input-nand_2.C.t2 GND 0.04477f
C8291 D_FlipFlop_6.3-input-nand_2.C.n2 GND 0.11971f
C8292 D_FlipFlop_6.3-input-nand_2.C.n3 GND 0.09193f
C8293 D_FlipFlop_6.3-input-nand_2.C.t7 GND 0.17806f
C8294 D_FlipFlop_6.3-input-nand_2.C.t4 GND 0.34248f
C8295 D_FlipFlop_6.3-input-nand_2.C.n4 GND 0.10005f
C8296 D_FlipFlop_6.3-input-nand_2.C.n5 GND 0.04279f
C8297 D_FlipFlop_6.3-input-nand_2.C.n6 GND 0.079f
C8298 D_FlipFlop_6.3-input-nand_2.C.n7 GND 0.13677f
C8299 D_FlipFlop_6.3-input-nand_2.C.n8 GND 0.10181f
C8300 D_FlipFlop_6.3-input-nand_2.C.n9 GND 0.04823f
C8301 D_FlipFlop_6.3-input-nand_2.C.n10 GND 0.124f
C8302 D_FlipFlop_6.3-input-nand_2.C.t1 GND 0.04742f
C8303 D_FlipFlop_6.3-input-nand_2.C.t0 GND 0.04645f
C8304 D_FlipFlop_6.3-input-nand_2.C.n11 GND 0.26418f
C8305 D_FlipFlop_6.3-input-nand_2.C.n12 GND 0.08722f
C8306 D_FlipFlop_6.3-input-nand_2.C.t3 GND 0.04645f
C8307 D_FlipFlop_6.3-input-nand_2.C.n13 GND 0.293f
C8308 D_FlipFlop_6.3-input-nand_2.C.t5 GND 0.17045f
C8309 D_FlipFlop_6.3-input-nand_2.C.n14 GND 0.05129f
C8310 VDD.n0 GND 0.02334f
C8311 VDD.t240 GND 0.02334f
C8312 VDD.t343 GND 0.02334f
C8313 VDD.n1 GND 0.03166f
C8314 VDD.n2 GND 0.0536f
C8315 VDD.n3 GND 0.05074f
C8316 VDD.n4 GND 0.0536f
C8317 VDD.n5 GND 0.04999f
C8318 VDD.n6 GND 0.04999f
C8319 VDD.t830 GND 0.63568f
C8320 VDD.n7 GND 0.04999f
C8321 VDD.n8 GND 0.05074f
C8322 VDD.n9 GND 0.05074f
C8323 VDD.n10 GND 0.02967f
C8324 VDD.n11 GND 0.02522f
C8325 VDD.n12 GND 0.0536f
C8326 VDD.n13 GND 0.05074f
C8327 VDD.n14 GND 0.02967f
C8328 VDD.n15 GND 0.02522f
C8329 VDD.t603 GND 0.63568f
C8330 VDD.n16 GND 0.04999f
C8331 VDD.n17 GND 0.05074f
C8332 VDD.n18 GND 0.05074f
C8333 VDD.n19 GND 0.02967f
C8334 VDD.n20 GND 0.02522f
C8335 VDD.n21 GND 0.0536f
C8336 VDD.t604 GND 0.02321f
C8337 VDD.t831 GND 0.02321f
C8338 VDD.n22 GND 0.10855f
C8339 VDD.t852 GND 0.02321f
C8340 VDD.t834 GND 0.02321f
C8341 VDD.n23 GND 0.10855f
C8342 VDD.n24 GND 0.04152f
C8343 VDD.n25 GND 0.03166f
C8344 VDD.n26 GND 0.05074f
C8345 VDD.n27 GND 0.02967f
C8346 VDD.n28 GND 0.02522f
C8347 VDD.t241 GND 0.63568f
C8348 VDD.n29 GND 0.04999f
C8349 VDD.n30 GND 0.05074f
C8350 VDD.n31 GND 0.05074f
C8351 VDD.n32 GND 0.02967f
C8352 VDD.n33 GND 0.02522f
C8353 VDD.n34 GND 0.0536f
C8354 VDD.n35 GND 0.0263f
C8355 VDD.n36 GND 0.05074f
C8356 VDD.n37 GND 0.02967f
C8357 VDD.n38 GND 0.02522f
C8358 VDD.t867 GND 0.74438f
C8359 VDD.n39 GND 0.05074f
C8360 VDD.n40 GND 0.05074f
C8361 VDD.n41 GND 0.02967f
C8362 VDD.n43 GND 0.62973f
C8363 VDD.n44 GND 0.02746f
C8364 VDD.t868 GND 0.02334f
C8365 VDD.t630 GND 0.02334f
C8366 VDD.n45 GND 0.0731f
C8367 VDD.n46 GND 0.02746f
C8368 VDD.n47 GND 0.05074f
C8369 VDD.n48 GND 0.02967f
C8370 VDD.n49 GND 0.05074f
C8371 VDD.n50 GND 0.35737f
C8372 VDD.t629 GND 0.33785f
C8373 VDD.t1089 GND 0.30977f
C8374 VDD.n52 GND 0.05074f
C8375 VDD.n53 GND 0.05074f
C8376 VDD.n54 GND 0.09132f
C8377 VDD.t77 GND 0.33785f
C8378 VDD.n55 GND 0.05074f
C8379 VDD.n56 GND 0.05074f
C8380 VDD.t1090 GND 0.02321f
C8381 VDD.t78 GND 0.02321f
C8382 VDD.n57 GND 0.10855f
C8383 VDD.n58 GND 0.02334f
C8384 VDD.n59 GND 0.03131f
C8385 VDD.t647 GND 0.02321f
C8386 VDD.t352 GND 0.02321f
C8387 VDD.n60 GND 0.10855f
C8388 VDD.n61 GND 0.03131f
C8389 VDD.n62 GND 0.02746f
C8390 VDD.n63 GND 0.05074f
C8391 VDD.n64 GND 0.02967f
C8392 VDD.n65 GND 0.05074f
C8393 VDD.n66 GND 0.35737f
C8394 VDD.t646 GND 0.33785f
C8395 VDD.t351 GND 0.33785f
C8396 VDD.n68 GND 0.05074f
C8397 VDD.n69 GND 0.05074f
C8398 VDD.t879 GND 0.02334f
C8399 VDD.n70 GND 0.0731f
C8400 VDD.n71 GND 0.02746f
C8401 VDD.n72 GND 0.05074f
C8402 VDD.n73 GND 0.02967f
C8403 VDD.n74 GND 0.05074f
C8404 VDD.n75 GND 0.35737f
C8405 VDD.t878 GND 0.33785f
C8406 VDD.t1065 GND 0.30977f
C8407 VDD.n77 GND 0.05074f
C8408 VDD.n78 GND 0.05074f
C8409 VDD.n79 GND 0.09132f
C8410 VDD.t957 GND 0.33785f
C8411 VDD.n80 GND 0.05074f
C8412 VDD.n81 GND 0.05074f
C8413 VDD.t1066 GND 0.02321f
C8414 VDD.t958 GND 0.02321f
C8415 VDD.n82 GND 0.10855f
C8416 VDD.n83 GND 0.02334f
C8417 VDD.n84 GND 0.03131f
C8418 VDD.t922 GND 0.02321f
C8419 VDD.t839 GND 0.02321f
C8420 VDD.n85 GND 0.10855f
C8421 VDD.n86 GND 0.03131f
C8422 VDD.n87 GND 0.02746f
C8423 VDD.n88 GND 0.05074f
C8424 VDD.n89 GND 0.02967f
C8425 VDD.n90 GND 0.05074f
C8426 VDD.n91 GND 0.35737f
C8427 VDD.t921 GND 0.33785f
C8428 VDD.t838 GND 0.33785f
C8429 VDD.n93 GND 0.05074f
C8430 VDD.n94 GND 0.05074f
C8431 VDD.t171 GND 0.02334f
C8432 VDD.n95 GND 0.0731f
C8433 VDD.n96 GND 0.02746f
C8434 VDD.n97 GND 0.05074f
C8435 VDD.n98 GND 0.02967f
C8436 VDD.n99 GND 0.05074f
C8437 VDD.n100 GND 0.35737f
C8438 VDD.t170 GND 0.33785f
C8439 VDD.t1026 GND 0.30977f
C8440 VDD.n102 GND 0.05074f
C8441 VDD.n103 GND 0.05074f
C8442 VDD.n104 GND 0.09132f
C8443 VDD.t976 GND 0.33785f
C8444 VDD.n105 GND 0.05074f
C8445 VDD.n106 GND 0.05074f
C8446 VDD.t1027 GND 0.02321f
C8447 VDD.t977 GND 0.02321f
C8448 VDD.n107 GND 0.10855f
C8449 VDD.n108 GND 0.02334f
C8450 VDD.n109 GND 0.03131f
C8451 VDD.t129 GND 0.02321f
C8452 VDD.t620 GND 0.02321f
C8453 VDD.n110 GND 0.10855f
C8454 VDD.n111 GND 0.03131f
C8455 VDD.n112 GND 0.02746f
C8456 VDD.n113 GND 0.05074f
C8457 VDD.n114 GND 0.02967f
C8458 VDD.n115 GND 0.05074f
C8459 VDD.n116 GND 0.35737f
C8460 VDD.t128 GND 0.33785f
C8461 VDD.t619 GND 0.33785f
C8462 VDD.n118 GND 0.05074f
C8463 VDD.n119 GND 0.05074f
C8464 VDD.t847 GND 0.02334f
C8465 VDD.n120 GND 0.0731f
C8466 VDD.n121 GND 0.02746f
C8467 VDD.n122 GND 0.05074f
C8468 VDD.n123 GND 0.02967f
C8469 VDD.n124 GND 0.05074f
C8470 VDD.n125 GND 0.35737f
C8471 VDD.t846 GND 0.33785f
C8472 VDD.t1072 GND 0.30977f
C8473 VDD.n127 GND 0.05074f
C8474 VDD.n128 GND 0.05074f
C8475 VDD.n129 GND 0.09132f
C8476 VDD.t654 GND 0.33785f
C8477 VDD.n130 GND 0.05074f
C8478 VDD.n131 GND 0.05074f
C8479 VDD.t1073 GND 0.02321f
C8480 VDD.t655 GND 0.02321f
C8481 VDD.n132 GND 0.10855f
C8482 VDD.n133 GND 0.02334f
C8483 VDD.n134 GND 0.03131f
C8484 VDD.t371 GND 0.02321f
C8485 VDD.t214 GND 0.02321f
C8486 VDD.n135 GND 0.10855f
C8487 VDD.n136 GND 0.03131f
C8488 VDD.n137 GND 0.02746f
C8489 VDD.n138 GND 0.05074f
C8490 VDD.n139 GND 0.02967f
C8491 VDD.n140 GND 0.05074f
C8492 VDD.n141 GND 0.35737f
C8493 VDD.t370 GND 0.33785f
C8494 VDD.t213 GND 0.33785f
C8495 VDD.n143 GND 0.05074f
C8496 VDD.n144 GND 0.05074f
C8497 VDD.n145 GND 0.02334f
C8498 VDD.n146 GND 0.09132f
C8499 VDD.n148 GND 0.35737f
C8500 VDD.n149 GND 0.02746f
C8501 VDD.n150 GND 0.02967f
C8502 VDD.n151 GND 0.02746f
C8503 VDD.n152 GND 0.04999f
C8504 VDD.n153 GND 0.24979f
C8505 VDD.n154 GND 0.24979f
C8506 VDD.n155 GND 0.04999f
C8507 VDD.n156 GND 0.02746f
C8508 VDD.n157 GND 0.09132f
C8509 VDD.n158 GND 0.34336f
C8510 VDD.n159 GND 0.02334f
C8511 VDD.n160 GND 0.09132f
C8512 VDD.n162 GND 0.35737f
C8513 VDD.n163 GND 0.02746f
C8514 VDD.n164 GND 0.02967f
C8515 VDD.n165 GND 0.02746f
C8516 VDD.n166 GND 0.04999f
C8517 VDD.n167 GND 0.24979f
C8518 VDD.n168 GND 0.24979f
C8519 VDD.n169 GND 0.04999f
C8520 VDD.n170 GND 0.02746f
C8521 VDD.n171 GND 0.02967f
C8522 VDD.n172 GND 0.02746f
C8523 VDD.n173 GND 0.04999f
C8524 VDD.n174 GND 0.33547f
C8525 VDD.n175 GND 0.33547f
C8526 VDD.n176 GND 0.04999f
C8527 VDD.n177 GND 0.02746f
C8528 VDD.n178 GND 0.09132f
C8529 VDD.n179 GND 0.33799f
C8530 VDD.n180 GND 0.02334f
C8531 VDD.n181 GND 0.09132f
C8532 VDD.n183 GND 0.35737f
C8533 VDD.n184 GND 0.02746f
C8534 VDD.n185 GND 0.02967f
C8535 VDD.n186 GND 0.02746f
C8536 VDD.n187 GND 0.04999f
C8537 VDD.n188 GND 0.24979f
C8538 VDD.n189 GND 0.24979f
C8539 VDD.n190 GND 0.04999f
C8540 VDD.n191 GND 0.02746f
C8541 VDD.n192 GND 0.09132f
C8542 VDD.n193 GND 0.34336f
C8543 VDD.n194 GND 0.02334f
C8544 VDD.n195 GND 0.09132f
C8545 VDD.n197 GND 0.35737f
C8546 VDD.n198 GND 0.02746f
C8547 VDD.n199 GND 0.02967f
C8548 VDD.n200 GND 0.02746f
C8549 VDD.n201 GND 0.04999f
C8550 VDD.n202 GND 0.24979f
C8551 VDD.n203 GND 0.24979f
C8552 VDD.n204 GND 0.04999f
C8553 VDD.n205 GND 0.02746f
C8554 VDD.n206 GND 0.02967f
C8555 VDD.n207 GND 0.02746f
C8556 VDD.n208 GND 0.04999f
C8557 VDD.n209 GND 0.33547f
C8558 VDD.n210 GND 0.33547f
C8559 VDD.n211 GND 0.04999f
C8560 VDD.n212 GND 0.02746f
C8561 VDD.n213 GND 0.09132f
C8562 VDD.n214 GND 0.33799f
C8563 VDD.n215 GND 0.02334f
C8564 VDD.n216 GND 0.09132f
C8565 VDD.n218 GND 0.35737f
C8566 VDD.n219 GND 0.02746f
C8567 VDD.n220 GND 0.02967f
C8568 VDD.n221 GND 0.02746f
C8569 VDD.n222 GND 0.04999f
C8570 VDD.n223 GND 0.24979f
C8571 VDD.n224 GND 0.24979f
C8572 VDD.n225 GND 0.04999f
C8573 VDD.n226 GND 0.02746f
C8574 VDD.n227 GND 0.09132f
C8575 VDD.n228 GND 0.34336f
C8576 VDD.n229 GND 0.02334f
C8577 VDD.n230 GND 0.09132f
C8578 VDD.n232 GND 0.35737f
C8579 VDD.n233 GND 0.02746f
C8580 VDD.n234 GND 0.02967f
C8581 VDD.n235 GND 0.02746f
C8582 VDD.n236 GND 0.04999f
C8583 VDD.n237 GND 0.24979f
C8584 VDD.n238 GND 0.24979f
C8585 VDD.n239 GND 0.04999f
C8586 VDD.n240 GND 0.02746f
C8587 VDD.n241 GND 0.02967f
C8588 VDD.n242 GND 0.02746f
C8589 VDD.n243 GND 0.04999f
C8590 VDD.n244 GND 0.33547f
C8591 VDD.n245 GND 0.33547f
C8592 VDD.n246 GND 0.04999f
C8593 VDD.n247 GND 0.02746f
C8594 VDD.n248 GND 0.09132f
C8595 VDD.n249 GND 0.33799f
C8596 VDD.n250 GND 0.02334f
C8597 VDD.n251 GND 0.09132f
C8598 VDD.n253 GND 0.35737f
C8599 VDD.n254 GND 0.02746f
C8600 VDD.n255 GND 0.02967f
C8601 VDD.n256 GND 0.02746f
C8602 VDD.n257 GND 0.04999f
C8603 VDD.n258 GND 0.24979f
C8604 VDD.n259 GND 0.24979f
C8605 VDD.n260 GND 0.04999f
C8606 VDD.n261 GND 0.02746f
C8607 VDD.n262 GND 0.09132f
C8608 VDD.n263 GND 0.34336f
C8609 VDD.n264 GND 0.02334f
C8610 VDD.n265 GND 0.09132f
C8611 VDD.n267 GND 0.35737f
C8612 VDD.n268 GND 0.02746f
C8613 VDD.n269 GND 0.02967f
C8614 VDD.n270 GND 0.02746f
C8615 VDD.n271 GND 0.04999f
C8616 VDD.n272 GND 0.24979f
C8617 VDD.n273 GND 0.24979f
C8618 VDD.n274 GND 0.04999f
C8619 VDD.n275 GND 0.02746f
C8620 VDD.n276 GND 0.02967f
C8621 VDD.n277 GND 0.02746f
C8622 VDD.n278 GND 0.04999f
C8623 VDD.n279 GND 0.33547f
C8624 VDD.n280 GND 0.33547f
C8625 VDD.n281 GND 0.04999f
C8626 VDD.n282 GND 0.02746f
C8627 VDD.n283 GND 0.09132f
C8628 VDD.n284 GND 0.01588f
C8629 VDD.n285 GND 0.37306f
C8630 VDD.t402 GND 2.03691f
C8631 VDD.n286 GND 0.51013f
C8632 VDD.n287 GND 0.32274f
C8633 VDD.n288 GND 0.32274f
C8634 VDD.n289 GND 0.55808f
C8635 VDD.n290 GND 3.99444f
C8636 VDD.n291 GND 0.3293f
C8637 VDD.n292 GND 1.66742f
C8638 VDD.t786 GND 4.164f
C8639 VDD.n294 GND 0.24939f
C8640 VDD.n295 GND 0.24939f
C8641 VDD.n296 GND 0.2271f
C8642 VDD.n297 GND 0.26346f
C8643 VDD.n298 GND 0.27199f
C8644 VDD.n299 GND 3.88046f
C8645 VDD.n300 GND 0.247f
C8646 VDD.n301 GND 4.164f
C8647 VDD.n302 GND 0.4484f
C8648 VDD.n303 GND 0.247f
C8649 VDD.t90 GND 1.61986f
C8650 VDD.t787 GND 1.61986f
C8651 VDD.n304 GND 0.91137f
C8652 VDD.t566 GND 0.2545f
C8653 VDD.n305 GND 1.05193f
C8654 VDD.n306 GND 1.48433f
C8655 VDD.n307 GND 0.51021f
C8656 VDD.n308 GND 1.11174f
C8657 VDD.n309 GND 6.13237f
C8658 VDD.n310 GND 7.25759f
C8659 VDD.n311 GND 8.5293f
C8660 VDD.n312 GND 2.14681f
C8661 VDD.n313 GND 1.79532f
C8662 VDD.n314 GND 0.88826f
C8663 VDD.n315 GND 0.54045f
C8664 VDD.n316 GND 1.18129f
C8665 VDD.n317 GND 4.98286f
C8666 VDD.n318 GND 4.78027f
C8667 VDD.n319 GND 4.33377f
C8668 VDD.n320 GND 1.02378f
C8669 VDD.n321 GND 0.45423f
C8670 VDD.n322 GND 1.14224f
C8671 VDD.n323 GND 3.01256f
C8672 VDD.n324 GND 0.14878f
C8673 VDD.n325 GND 0.0704f
C8674 VDD.n326 GND 0.19384f
C8675 VDD.n327 GND 0.2271f
C8676 VDD.n328 GND 0.24939f
C8677 VDD.t89 GND 4.3411f
C8678 VDD.n330 GND 0.24939f
C8679 VDD.n331 GND 0.14592f
C8680 VDD.n332 GND 0.1451f
C8681 VDD.n333 GND 0.14592f
C8682 VDD.n334 GND 0.27199f
C8683 VDD.n335 GND 0.47144f
C8684 VDD.n336 GND 6.86348f
C8685 VDD.n337 GND 6.86348f
C8686 VDD.t401 GND 5.34916f
C8687 VDD.n338 GND 0.5627f
C8688 VDD.n339 GND 0.44303f
C8689 VDD.n340 GND 0.08304f
C8690 VDD.n341 GND 0.61662f
C8691 VDD.t964 GND 0.02334f
C8692 VDD.n342 GND 0.02746f
C8693 VDD.n343 GND 0.05074f
C8694 VDD.n344 GND 0.02967f
C8695 VDD.n345 GND 0.05074f
C8696 VDD.n346 GND 0.62973f
C8697 VDD.t963 GND 0.74438f
C8698 VDD.n348 GND 0.04999f
C8699 VDD.t11 GND 0.63568f
C8700 VDD.n349 GND 0.05074f
C8701 VDD.n350 GND 0.05074f
C8702 VDD.n351 GND 0.02967f
C8703 VDD.n352 GND 0.02522f
C8704 VDD.t12 GND 0.02334f
C8705 VDD.t79 GND 0.02334f
C8706 VDD.n353 GND 0.13341f
C8707 VDD.n354 GND 0.0263f
C8708 VDD.n355 GND 0.0536f
C8709 VDD.n356 GND 0.05074f
C8710 VDD.n357 GND 0.02967f
C8711 VDD.n358 GND 0.02522f
C8712 VDD.n359 GND 0.04999f
C8713 VDD.t333 GND 0.63568f
C8714 VDD.n360 GND 0.05074f
C8715 VDD.n361 GND 0.05074f
C8716 VDD.n362 GND 0.02967f
C8717 VDD.n363 GND 0.02522f
C8718 VDD.n364 GND 0.03166f
C8719 VDD.n365 GND 0.0536f
C8720 VDD.n366 GND 0.05074f
C8721 VDD.n367 GND 0.02967f
C8722 VDD.n368 GND 0.02522f
C8723 VDD.n369 GND 0.04999f
C8724 VDD.t555 GND 0.63568f
C8725 VDD.n370 GND 0.05074f
C8726 VDD.n371 GND 0.05074f
C8727 VDD.n372 GND 0.02967f
C8728 VDD.n373 GND 0.02522f
C8729 VDD.t395 GND 0.02321f
C8730 VDD.t557 GND 0.02321f
C8731 VDD.n374 GND 0.10855f
C8732 VDD.t334 GND 0.02321f
C8733 VDD.t556 GND 0.02321f
C8734 VDD.n375 GND 0.10855f
C8735 VDD.n376 GND 0.04152f
C8736 VDD.n377 GND 0.02334f
C8737 VDD.n378 GND 0.0536f
C8738 VDD.n379 GND 0.05074f
C8739 VDD.n380 GND 0.02967f
C8740 VDD.n381 GND 0.02522f
C8741 VDD.n382 GND 0.04999f
C8742 VDD.t249 GND 0.63568f
C8743 VDD.n383 GND 0.05074f
C8744 VDD.n384 GND 0.05074f
C8745 VDD.n385 GND 0.02967f
C8746 VDD.n386 GND 0.02522f
C8747 VDD.t577 GND 0.02334f
C8748 VDD.t250 GND 0.02334f
C8749 VDD.n387 GND 0.13341f
C8750 VDD.n388 GND 0.0263f
C8751 VDD.n389 GND 0.0536f
C8752 VDD.n390 GND 0.05074f
C8753 VDD.n391 GND 0.02967f
C8754 VDD.n392 GND 0.02522f
C8755 VDD.n393 GND 0.04999f
C8756 VDD.t75 GND 0.63568f
C8757 VDD.n394 GND 0.05074f
C8758 VDD.n395 GND 0.05074f
C8759 VDD.n396 GND 0.02967f
C8760 VDD.n397 GND 0.02522f
C8761 VDD.n398 GND 0.03166f
C8762 VDD.n399 GND 0.0536f
C8763 VDD.n400 GND 0.05074f
C8764 VDD.n401 GND 0.02967f
C8765 VDD.n402 GND 0.02522f
C8766 VDD.n403 GND 0.04999f
C8767 VDD.t233 GND 0.63568f
C8768 VDD.n404 GND 0.05074f
C8769 VDD.n405 GND 0.05074f
C8770 VDD.n406 GND 0.02967f
C8771 VDD.n407 GND 0.02522f
C8772 VDD.t76 GND 0.02321f
C8773 VDD.t975 GND 0.02321f
C8774 VDD.n408 GND 0.10855f
C8775 VDD.t108 GND 0.02321f
C8776 VDD.t234 GND 0.02321f
C8777 VDD.n409 GND 0.10855f
C8778 VDD.n410 GND 0.04152f
C8779 VDD.n411 GND 0.02334f
C8780 VDD.n412 GND 0.0536f
C8781 VDD.n413 GND 0.05074f
C8782 VDD.n414 GND 0.02967f
C8783 VDD.n415 GND 0.02522f
C8784 VDD.t58 GND 0.63568f
C8785 VDD.n416 GND 0.05074f
C8786 VDD.n417 GND 0.05074f
C8787 VDD.n418 GND 0.09132f
C8788 VDD.n419 GND 0.04999f
C8789 VDD.t204 GND 0.63568f
C8790 VDD.n420 GND 0.05074f
C8791 VDD.n421 GND 0.05074f
C8792 VDD.n422 GND 0.02967f
C8793 VDD.n423 GND 0.02522f
C8794 VDD.t59 GND 0.02334f
C8795 VDD.n424 GND 0.0731f
C8796 VDD.n425 GND 0.01798f
C8797 VDD.n426 GND 0.02334f
C8798 VDD.n427 GND 0.0536f
C8799 VDD.n428 GND 0.05074f
C8800 VDD.n429 GND 0.02967f
C8801 VDD.n430 GND 0.02522f
C8802 VDD.n431 GND 0.04999f
C8803 VDD.t988 GND 0.63568f
C8804 VDD.n432 GND 0.05074f
C8805 VDD.n433 GND 0.05074f
C8806 VDD.n434 GND 0.02967f
C8807 VDD.n435 GND 0.02522f
C8808 VDD.t205 GND 0.02321f
C8809 VDD.t990 GND 0.02321f
C8810 VDD.n436 GND 0.10855f
C8811 VDD.t273 GND 0.02321f
C8812 VDD.t989 GND 0.02321f
C8813 VDD.n437 GND 0.10855f
C8814 VDD.n438 GND 0.04152f
C8815 VDD.n439 GND 0.02334f
C8816 VDD.n440 GND 0.0536f
C8817 VDD.n441 GND 0.05074f
C8818 VDD.n442 GND 0.02967f
C8819 VDD.n443 GND 0.02522f
C8820 VDD.n444 GND 0.04999f
C8821 VDD.t339 GND 0.63568f
C8822 VDD.n445 GND 0.05074f
C8823 VDD.n446 GND 0.05074f
C8824 VDD.n447 GND 0.02967f
C8825 VDD.n448 GND 0.02522f
C8826 VDD.t959 GND 0.02334f
C8827 VDD.t340 GND 0.02334f
C8828 VDD.n449 GND 0.13341f
C8829 VDD.n450 GND 0.0263f
C8830 VDD.n451 GND 0.0536f
C8831 VDD.n452 GND 0.05074f
C8832 VDD.n453 GND 0.02967f
C8833 VDD.n454 GND 0.02522f
C8834 VDD.n455 GND 0.04999f
C8835 VDD.t335 GND 0.63568f
C8836 VDD.n456 GND 0.05074f
C8837 VDD.n457 GND 0.05074f
C8838 VDD.n458 GND 0.02967f
C8839 VDD.n459 GND 0.02522f
C8840 VDD.n460 GND 0.03166f
C8841 VDD.n461 GND 0.0536f
C8842 VDD.n462 GND 0.05074f
C8843 VDD.n463 GND 0.02967f
C8844 VDD.n464 GND 0.02522f
C8845 VDD.n465 GND 0.04999f
C8846 VDD.t362 GND 0.63568f
C8847 VDD.n466 GND 0.05074f
C8848 VDD.n467 GND 0.05074f
C8849 VDD.n468 GND 0.02967f
C8850 VDD.n469 GND 0.02522f
C8851 VDD.t398 GND 0.02321f
C8852 VDD.t363 GND 0.02321f
C8853 VDD.n470 GND 0.10855f
C8854 VDD.t336 GND 0.02321f
C8855 VDD.t785 GND 0.02321f
C8856 VDD.n471 GND 0.10855f
C8857 VDD.n472 GND 0.04152f
C8858 VDD.n473 GND 0.02334f
C8859 VDD.n474 GND 0.0536f
C8860 VDD.n475 GND 0.05074f
C8861 VDD.n476 GND 0.02967f
C8862 VDD.n477 GND 0.02522f
C8863 VDD.n478 GND 0.02522f
C8864 VDD.n479 GND 0.04999f
C8865 VDD.n480 GND 0.68843f
C8866 VDD.n481 GND 0.04999f
C8867 VDD.n482 GND 0.05074f
C8868 VDD.n483 GND 0.06295f
C8869 VDD.n484 GND 0.0536f
C8870 VDD.n485 GND 0.02522f
C8871 VDD.n486 GND 0.04999f
C8872 VDD.n487 GND 0.5126f
C8873 VDD.n488 GND 0.02522f
C8874 VDD.n489 GND 0.04999f
C8875 VDD.n490 GND 0.5126f
C8876 VDD.n491 GND 0.04999f
C8877 VDD.n492 GND 0.05074f
C8878 VDD.n493 GND 0.06295f
C8879 VDD.n494 GND 0.0536f
C8880 VDD.n495 GND 0.02522f
C8881 VDD.n496 GND 0.04999f
C8882 VDD.n497 GND 0.5126f
C8883 VDD.n498 GND 0.02522f
C8884 VDD.n499 GND 0.04999f
C8885 VDD.n500 GND 0.5126f
C8886 VDD.n501 GND 0.04999f
C8887 VDD.n502 GND 0.05074f
C8888 VDD.n503 GND 0.06295f
C8889 VDD.n504 GND 0.0536f
C8890 VDD.n505 GND 0.02522f
C8891 VDD.n506 GND 0.04999f
C8892 VDD.n507 GND 0.68843f
C8893 VDD.n508 GND 0.02522f
C8894 VDD.n509 GND 0.04999f
C8895 VDD.n510 GND 0.68843f
C8896 VDD.n511 GND 0.04999f
C8897 VDD.n512 GND 0.05074f
C8898 VDD.n513 GND 0.06295f
C8899 VDD.n514 GND 0.0536f
C8900 VDD.n515 GND 0.02522f
C8901 VDD.n516 GND 0.04999f
C8902 VDD.n517 GND 0.5126f
C8903 VDD.n518 GND 0.02522f
C8904 VDD.n519 GND 0.04999f
C8905 VDD.n520 GND 0.5126f
C8906 VDD.n521 GND 0.04999f
C8907 VDD.n522 GND 0.05074f
C8908 VDD.n523 GND 0.06295f
C8909 VDD.n524 GND 0.0536f
C8910 VDD.n525 GND 0.02522f
C8911 VDD.n526 GND 0.04999f
C8912 VDD.n527 GND 0.68843f
C8913 VDD.n528 GND 0.68843f
C8914 VDD.n529 GND 0.04999f
C8915 VDD.n530 GND 0.02746f
C8916 VDD.n531 GND 0.02967f
C8917 VDD.n532 GND 0.02746f
C8918 VDD.n533 GND 0.04999f
C8919 VDD.n534 GND 0.68843f
C8920 VDD.n535 GND 0.02522f
C8921 VDD.n536 GND 0.04999f
C8922 VDD.n537 GND 0.68843f
C8923 VDD.n538 GND 0.04999f
C8924 VDD.n539 GND 0.05074f
C8925 VDD.n540 GND 0.06295f
C8926 VDD.n541 GND 0.0536f
C8927 VDD.n542 GND 0.02522f
C8928 VDD.n543 GND 0.04999f
C8929 VDD.n544 GND 0.5126f
C8930 VDD.n545 GND 0.02522f
C8931 VDD.n546 GND 0.04999f
C8932 VDD.n547 GND 0.5126f
C8933 VDD.n548 GND 0.04999f
C8934 VDD.n549 GND 0.05074f
C8935 VDD.n550 GND 0.06295f
C8936 VDD.n551 GND 0.0536f
C8937 VDD.n552 GND 0.02522f
C8938 VDD.n553 GND 0.04999f
C8939 VDD.n554 GND 0.5126f
C8940 VDD.n555 GND 0.02522f
C8941 VDD.n556 GND 0.04999f
C8942 VDD.n557 GND 0.5126f
C8943 VDD.n558 GND 0.04999f
C8944 VDD.n559 GND 0.05074f
C8945 VDD.n560 GND 0.06295f
C8946 VDD.n561 GND 0.0536f
C8947 VDD.n562 GND 0.02522f
C8948 VDD.n563 GND 0.04999f
C8949 VDD.n564 GND 0.68843f
C8950 VDD.n565 GND 0.02522f
C8951 VDD.n566 GND 0.04999f
C8952 VDD.n567 GND 0.68843f
C8953 VDD.n568 GND 0.04999f
C8954 VDD.n569 GND 0.05074f
C8955 VDD.n570 GND 0.06295f
C8956 VDD.n571 GND 0.0536f
C8957 VDD.n572 GND 0.02522f
C8958 VDD.n573 GND 0.04999f
C8959 VDD.n574 GND 0.5126f
C8960 VDD.n575 GND 0.02522f
C8961 VDD.n576 GND 0.04999f
C8962 VDD.n577 GND 0.5126f
C8963 VDD.n578 GND 0.04999f
C8964 VDD.n579 GND 0.05074f
C8965 VDD.n580 GND 0.06295f
C8966 VDD.n581 GND 0.0536f
C8967 VDD.n582 GND 0.02522f
C8968 VDD.n583 GND 0.04999f
C8969 VDD.n584 GND 0.5126f
C8970 VDD.n585 GND 0.02522f
C8971 VDD.n586 GND 0.04999f
C8972 VDD.n587 GND 0.5126f
C8973 VDD.n588 GND 0.04999f
C8974 VDD.n589 GND 0.05074f
C8975 VDD.n590 GND 0.06295f
C8976 VDD.n591 GND 0.0536f
C8977 VDD.n592 GND 0.02522f
C8978 VDD.n593 GND 0.04999f
C8979 VDD.n594 GND 0.68843f
C8980 VDD.n595 GND 0.68843f
C8981 VDD.n596 GND 0.04999f
C8982 VDD.n597 GND 0.02746f
C8983 VDD.n598 GND 0.09132f
C8984 VDD.n599 GND 0.01798f
C8985 VDD.n600 GND 0.09868f
C8986 VDD.n601 GND 0.26626f
C8987 VDD.t606 GND 0.02334f
C8988 VDD.n602 GND 0.02746f
C8989 VDD.n603 GND 0.05074f
C8990 VDD.n604 GND 0.02967f
C8991 VDD.n605 GND 0.05074f
C8992 VDD.n606 GND 0.62973f
C8993 VDD.t605 GND 0.74438f
C8994 VDD.n608 GND 0.04999f
C8995 VDD.t353 GND 0.63568f
C8996 VDD.n609 GND 0.05074f
C8997 VDD.n610 GND 0.05074f
C8998 VDD.n611 GND 0.02967f
C8999 VDD.n612 GND 0.02522f
C9000 VDD.t354 GND 0.02334f
C9001 VDD.t843 GND 0.02334f
C9002 VDD.n613 GND 0.13341f
C9003 VDD.n614 GND 0.0263f
C9004 VDD.n615 GND 0.0536f
C9005 VDD.n616 GND 0.05074f
C9006 VDD.n617 GND 0.02967f
C9007 VDD.n618 GND 0.02522f
C9008 VDD.n619 GND 0.04999f
C9009 VDD.t120 GND 0.63568f
C9010 VDD.n620 GND 0.05074f
C9011 VDD.n621 GND 0.05074f
C9012 VDD.n622 GND 0.02967f
C9013 VDD.n623 GND 0.02522f
C9014 VDD.n624 GND 0.03166f
C9015 VDD.n625 GND 0.0536f
C9016 VDD.n626 GND 0.05074f
C9017 VDD.n627 GND 0.02967f
C9018 VDD.n628 GND 0.02522f
C9019 VDD.n629 GND 0.04999f
C9020 VDD.t41 GND 0.63568f
C9021 VDD.n630 GND 0.05074f
C9022 VDD.n631 GND 0.05074f
C9023 VDD.n632 GND 0.02967f
C9024 VDD.n633 GND 0.02522f
C9025 VDD.t965 GND 0.02321f
C9026 VDD.t42 GND 0.02321f
C9027 VDD.n634 GND 0.10855f
C9028 VDD.t121 GND 0.02321f
C9029 VDD.t45 GND 0.02321f
C9030 VDD.n635 GND 0.10855f
C9031 VDD.n636 GND 0.04152f
C9032 VDD.n637 GND 0.02334f
C9033 VDD.n638 GND 0.0536f
C9034 VDD.n639 GND 0.05074f
C9035 VDD.n640 GND 0.02967f
C9036 VDD.n641 GND 0.02522f
C9037 VDD.n642 GND 0.04999f
C9038 VDD.t384 GND 0.63568f
C9039 VDD.n643 GND 0.05074f
C9040 VDD.n644 GND 0.05074f
C9041 VDD.n645 GND 0.02967f
C9042 VDD.n646 GND 0.02522f
C9043 VDD.t842 GND 0.02334f
C9044 VDD.t385 GND 0.02334f
C9045 VDD.n647 GND 0.13341f
C9046 VDD.n648 GND 0.0263f
C9047 VDD.n649 GND 0.0536f
C9048 VDD.n650 GND 0.05074f
C9049 VDD.n651 GND 0.02967f
C9050 VDD.n652 GND 0.02522f
C9051 VDD.n653 GND 0.04999f
C9052 VDD.t220 GND 0.63568f
C9053 VDD.n654 GND 0.05074f
C9054 VDD.n655 GND 0.05074f
C9055 VDD.n656 GND 0.02967f
C9056 VDD.n657 GND 0.02522f
C9057 VDD.n658 GND 0.03166f
C9058 VDD.n659 GND 0.0536f
C9059 VDD.n660 GND 0.05074f
C9060 VDD.n661 GND 0.02967f
C9061 VDD.n662 GND 0.02522f
C9062 VDD.n663 GND 0.04999f
C9063 VDD.t166 GND 0.63568f
C9064 VDD.n664 GND 0.05074f
C9065 VDD.n665 GND 0.05074f
C9066 VDD.n666 GND 0.02967f
C9067 VDD.n667 GND 0.02522f
C9068 VDD.t221 GND 0.02321f
C9069 VDD.t613 GND 0.02321f
C9070 VDD.n668 GND 0.10855f
C9071 VDD.t853 GND 0.02321f
C9072 VDD.t167 GND 0.02321f
C9073 VDD.n669 GND 0.10855f
C9074 VDD.n670 GND 0.04152f
C9075 VDD.n671 GND 0.02334f
C9076 VDD.n672 GND 0.0536f
C9077 VDD.n673 GND 0.05074f
C9078 VDD.n674 GND 0.02967f
C9079 VDD.n675 GND 0.02522f
C9080 VDD.t43 GND 0.63568f
C9081 VDD.n676 GND 0.05074f
C9082 VDD.n677 GND 0.05074f
C9083 VDD.n678 GND 0.09132f
C9084 VDD.n679 GND 0.04999f
C9085 VDD.t164 GND 0.63568f
C9086 VDD.n680 GND 0.05074f
C9087 VDD.n681 GND 0.05074f
C9088 VDD.n682 GND 0.02967f
C9089 VDD.n683 GND 0.02522f
C9090 VDD.t44 GND 0.02334f
C9091 VDD.n684 GND 0.0731f
C9092 VDD.n685 GND 0.01798f
C9093 VDD.n686 GND 0.02334f
C9094 VDD.n687 GND 0.0536f
C9095 VDD.n688 GND 0.05074f
C9096 VDD.n689 GND 0.02967f
C9097 VDD.n690 GND 0.02522f
C9098 VDD.n691 GND 0.04999f
C9099 VDD.t60 GND 0.63568f
C9100 VDD.n692 GND 0.05074f
C9101 VDD.n693 GND 0.05074f
C9102 VDD.n694 GND 0.02967f
C9103 VDD.n695 GND 0.02522f
C9104 VDD.t165 GND 0.02321f
C9105 VDD.t62 GND 0.02321f
C9106 VDD.n696 GND 0.10855f
C9107 VDD.t614 GND 0.02321f
C9108 VDD.t61 GND 0.02321f
C9109 VDD.n697 GND 0.10855f
C9110 VDD.n698 GND 0.04152f
C9111 VDD.n699 GND 0.02334f
C9112 VDD.n700 GND 0.0536f
C9113 VDD.n701 GND 0.05074f
C9114 VDD.n702 GND 0.02967f
C9115 VDD.n703 GND 0.02522f
C9116 VDD.n704 GND 0.04999f
C9117 VDD.t356 GND 0.63568f
C9118 VDD.n705 GND 0.05074f
C9119 VDD.n706 GND 0.05074f
C9120 VDD.n707 GND 0.02967f
C9121 VDD.n708 GND 0.02522f
C9122 VDD.t844 GND 0.02334f
C9123 VDD.t357 GND 0.02334f
C9124 VDD.n709 GND 0.13341f
C9125 VDD.n710 GND 0.0263f
C9126 VDD.n711 GND 0.0536f
C9127 VDD.n712 GND 0.05074f
C9128 VDD.n713 GND 0.02967f
C9129 VDD.n714 GND 0.02522f
C9130 VDD.n715 GND 0.04999f
C9131 VDD.t63 GND 0.63568f
C9132 VDD.n716 GND 0.05074f
C9133 VDD.n717 GND 0.05074f
C9134 VDD.n718 GND 0.02967f
C9135 VDD.n719 GND 0.02522f
C9136 VDD.n720 GND 0.03166f
C9137 VDD.n721 GND 0.0536f
C9138 VDD.n722 GND 0.05074f
C9139 VDD.n723 GND 0.02967f
C9140 VDD.n724 GND 0.02522f
C9141 VDD.n725 GND 0.04999f
C9142 VDD.t278 GND 0.63568f
C9143 VDD.n726 GND 0.05074f
C9144 VDD.n727 GND 0.05074f
C9145 VDD.n728 GND 0.02967f
C9146 VDD.n729 GND 0.02522f
C9147 VDD.t64 GND 0.02321f
C9148 VDD.t560 GND 0.02321f
C9149 VDD.n730 GND 0.10855f
C9150 VDD.t294 GND 0.02321f
C9151 VDD.t279 GND 0.02321f
C9152 VDD.n731 GND 0.10855f
C9153 VDD.n732 GND 0.04152f
C9154 VDD.n733 GND 0.02334f
C9155 VDD.n734 GND 0.0536f
C9156 VDD.n735 GND 0.05074f
C9157 VDD.n736 GND 0.02967f
C9158 VDD.n737 GND 0.02522f
C9159 VDD.n738 GND 0.02522f
C9160 VDD.n739 GND 0.04999f
C9161 VDD.n740 GND 0.68843f
C9162 VDD.n741 GND 0.04999f
C9163 VDD.n742 GND 0.05074f
C9164 VDD.n743 GND 0.06295f
C9165 VDD.n744 GND 0.0536f
C9166 VDD.n745 GND 0.02522f
C9167 VDD.n746 GND 0.04999f
C9168 VDD.n747 GND 0.5126f
C9169 VDD.n748 GND 0.02522f
C9170 VDD.n749 GND 0.04999f
C9171 VDD.n750 GND 0.5126f
C9172 VDD.n751 GND 0.04999f
C9173 VDD.n752 GND 0.05074f
C9174 VDD.n753 GND 0.06295f
C9175 VDD.n754 GND 0.0536f
C9176 VDD.n755 GND 0.02522f
C9177 VDD.n756 GND 0.04999f
C9178 VDD.n757 GND 0.5126f
C9179 VDD.n758 GND 0.02522f
C9180 VDD.n759 GND 0.04999f
C9181 VDD.n760 GND 0.5126f
C9182 VDD.n761 GND 0.04999f
C9183 VDD.n762 GND 0.05074f
C9184 VDD.n763 GND 0.06295f
C9185 VDD.n764 GND 0.0536f
C9186 VDD.n765 GND 0.02522f
C9187 VDD.n766 GND 0.04999f
C9188 VDD.n767 GND 0.68843f
C9189 VDD.n768 GND 0.02522f
C9190 VDD.n769 GND 0.04999f
C9191 VDD.n770 GND 0.68843f
C9192 VDD.n771 GND 0.04999f
C9193 VDD.n772 GND 0.05074f
C9194 VDD.n773 GND 0.06295f
C9195 VDD.n774 GND 0.0536f
C9196 VDD.n775 GND 0.02522f
C9197 VDD.n776 GND 0.04999f
C9198 VDD.n777 GND 0.5126f
C9199 VDD.n778 GND 0.02522f
C9200 VDD.n779 GND 0.04999f
C9201 VDD.n780 GND 0.5126f
C9202 VDD.n781 GND 0.04999f
C9203 VDD.n782 GND 0.05074f
C9204 VDD.n783 GND 0.06295f
C9205 VDD.n784 GND 0.0536f
C9206 VDD.n785 GND 0.02522f
C9207 VDD.n786 GND 0.04999f
C9208 VDD.n787 GND 0.68843f
C9209 VDD.n788 GND 0.68843f
C9210 VDD.n789 GND 0.04999f
C9211 VDD.n790 GND 0.02746f
C9212 VDD.n791 GND 0.02967f
C9213 VDD.n792 GND 0.02746f
C9214 VDD.n793 GND 0.04999f
C9215 VDD.n794 GND 0.68843f
C9216 VDD.n795 GND 0.02522f
C9217 VDD.n796 GND 0.04999f
C9218 VDD.n797 GND 0.68843f
C9219 VDD.n798 GND 0.04999f
C9220 VDD.n799 GND 0.05074f
C9221 VDD.n800 GND 0.06295f
C9222 VDD.n801 GND 0.0536f
C9223 VDD.n802 GND 0.02522f
C9224 VDD.n803 GND 0.04999f
C9225 VDD.n804 GND 0.5126f
C9226 VDD.n805 GND 0.02522f
C9227 VDD.n806 GND 0.04999f
C9228 VDD.n807 GND 0.5126f
C9229 VDD.n808 GND 0.04999f
C9230 VDD.n809 GND 0.05074f
C9231 VDD.n810 GND 0.06295f
C9232 VDD.n811 GND 0.0536f
C9233 VDD.n812 GND 0.02522f
C9234 VDD.n813 GND 0.04999f
C9235 VDD.n814 GND 0.5126f
C9236 VDD.n815 GND 0.02522f
C9237 VDD.n816 GND 0.04999f
C9238 VDD.n817 GND 0.5126f
C9239 VDD.n818 GND 0.04999f
C9240 VDD.n819 GND 0.05074f
C9241 VDD.n820 GND 0.06295f
C9242 VDD.n821 GND 0.0536f
C9243 VDD.n822 GND 0.02522f
C9244 VDD.n823 GND 0.04999f
C9245 VDD.n824 GND 0.68843f
C9246 VDD.n825 GND 0.02522f
C9247 VDD.n826 GND 0.04999f
C9248 VDD.n827 GND 0.68843f
C9249 VDD.n828 GND 0.04999f
C9250 VDD.n829 GND 0.05074f
C9251 VDD.n830 GND 0.06295f
C9252 VDD.n831 GND 0.0536f
C9253 VDD.n832 GND 0.02522f
C9254 VDD.n833 GND 0.04999f
C9255 VDD.n834 GND 0.5126f
C9256 VDD.n835 GND 0.02522f
C9257 VDD.n836 GND 0.04999f
C9258 VDD.n837 GND 0.5126f
C9259 VDD.n838 GND 0.04999f
C9260 VDD.n839 GND 0.05074f
C9261 VDD.n840 GND 0.06295f
C9262 VDD.n841 GND 0.0536f
C9263 VDD.n842 GND 0.02522f
C9264 VDD.n843 GND 0.04999f
C9265 VDD.n844 GND 0.5126f
C9266 VDD.n845 GND 0.02522f
C9267 VDD.n846 GND 0.04999f
C9268 VDD.n847 GND 0.5126f
C9269 VDD.n848 GND 0.04999f
C9270 VDD.n849 GND 0.05074f
C9271 VDD.n850 GND 0.06295f
C9272 VDD.n851 GND 0.0536f
C9273 VDD.n852 GND 0.02522f
C9274 VDD.n853 GND 0.04999f
C9275 VDD.n854 GND 0.68843f
C9276 VDD.n855 GND 0.68843f
C9277 VDD.n856 GND 0.04999f
C9278 VDD.n857 GND 0.02746f
C9279 VDD.n858 GND 0.09132f
C9280 VDD.n859 GND 0.01798f
C9281 VDD.n860 GND 0.09868f
C9282 VDD.n861 GND 0.3275f
C9283 VDD.t866 GND 0.02334f
C9284 VDD.n862 GND 0.02746f
C9285 VDD.n863 GND 0.05074f
C9286 VDD.n864 GND 0.02967f
C9287 VDD.n865 GND 0.05074f
C9288 VDD.n866 GND 0.62973f
C9289 VDD.t865 GND 0.74438f
C9290 VDD.n868 GND 0.04999f
C9291 VDD.t247 GND 0.63568f
C9292 VDD.n869 GND 0.05074f
C9293 VDD.n870 GND 0.05074f
C9294 VDD.n871 GND 0.02967f
C9295 VDD.n872 GND 0.02522f
C9296 VDD.t248 GND 0.02334f
C9297 VDD.t624 GND 0.02334f
C9298 VDD.n873 GND 0.13341f
C9299 VDD.n874 GND 0.0263f
C9300 VDD.n875 GND 0.0536f
C9301 VDD.n876 GND 0.05074f
C9302 VDD.n877 GND 0.02967f
C9303 VDD.n878 GND 0.02522f
C9304 VDD.n879 GND 0.04999f
C9305 VDD.t601 GND 0.63568f
C9306 VDD.n880 GND 0.05074f
C9307 VDD.n881 GND 0.05074f
C9308 VDD.n882 GND 0.02967f
C9309 VDD.n883 GND 0.02522f
C9310 VDD.n884 GND 0.03166f
C9311 VDD.n885 GND 0.0536f
C9312 VDD.n886 GND 0.05074f
C9313 VDD.n887 GND 0.02967f
C9314 VDD.n888 GND 0.02522f
C9315 VDD.n889 GND 0.04999f
C9316 VDD.t657 GND 0.63568f
C9317 VDD.n890 GND 0.05074f
C9318 VDD.n891 GND 0.05074f
C9319 VDD.n892 GND 0.02967f
C9320 VDD.n893 GND 0.02522f
C9321 VDD.t602 GND 0.02321f
C9322 VDD.t658 GND 0.02321f
C9323 VDD.n894 GND 0.10855f
C9324 VDD.t631 GND 0.02321f
C9325 VDD.t766 GND 0.02321f
C9326 VDD.n895 GND 0.10855f
C9327 VDD.n896 GND 0.04152f
C9328 VDD.n897 GND 0.02334f
C9329 VDD.n898 GND 0.0536f
C9330 VDD.n899 GND 0.05074f
C9331 VDD.n900 GND 0.02967f
C9332 VDD.n901 GND 0.02522f
C9333 VDD.n902 GND 0.04999f
C9334 VDD.t642 GND 0.63568f
C9335 VDD.n903 GND 0.05074f
C9336 VDD.n904 GND 0.05074f
C9337 VDD.n905 GND 0.02967f
C9338 VDD.n906 GND 0.02522f
C9339 VDD.t873 GND 0.02334f
C9340 VDD.t643 GND 0.02334f
C9341 VDD.n907 GND 0.13341f
C9342 VDD.n908 GND 0.0263f
C9343 VDD.n909 GND 0.0536f
C9344 VDD.n910 GND 0.05074f
C9345 VDD.n911 GND 0.02967f
C9346 VDD.n912 GND 0.02522f
C9347 VDD.n913 GND 0.04999f
C9348 VDD.t429 GND 0.63568f
C9349 VDD.n914 GND 0.05074f
C9350 VDD.n915 GND 0.05074f
C9351 VDD.n916 GND 0.02967f
C9352 VDD.n917 GND 0.02522f
C9353 VDD.n918 GND 0.03166f
C9354 VDD.n919 GND 0.0536f
C9355 VDD.n920 GND 0.05074f
C9356 VDD.n921 GND 0.02967f
C9357 VDD.n922 GND 0.02522f
C9358 VDD.n923 GND 0.04999f
C9359 VDD.t174 GND 0.63568f
C9360 VDD.n924 GND 0.05074f
C9361 VDD.n925 GND 0.05074f
C9362 VDD.n926 GND 0.02967f
C9363 VDD.n927 GND 0.02522f
C9364 VDD.t824 GND 0.02321f
C9365 VDD.t910 GND 0.02321f
C9366 VDD.n928 GND 0.10855f
C9367 VDD.t430 GND 0.02321f
C9368 VDD.t175 GND 0.02321f
C9369 VDD.n929 GND 0.10855f
C9370 VDD.n930 GND 0.04152f
C9371 VDD.n931 GND 0.02334f
C9372 VDD.n932 GND 0.0536f
C9373 VDD.n933 GND 0.05074f
C9374 VDD.n934 GND 0.02967f
C9375 VDD.n935 GND 0.02522f
C9376 VDD.t659 GND 0.63568f
C9377 VDD.n936 GND 0.05074f
C9378 VDD.n937 GND 0.05074f
C9379 VDD.n938 GND 0.09132f
C9380 VDD.n939 GND 0.04999f
C9381 VDD.t172 GND 0.63568f
C9382 VDD.n940 GND 0.05074f
C9383 VDD.n941 GND 0.05074f
C9384 VDD.n942 GND 0.02967f
C9385 VDD.n943 GND 0.02522f
C9386 VDD.t660 GND 0.02334f
C9387 VDD.n944 GND 0.0731f
C9388 VDD.n945 GND 0.01798f
C9389 VDD.n946 GND 0.02334f
C9390 VDD.n947 GND 0.0536f
C9391 VDD.n948 GND 0.05074f
C9392 VDD.n949 GND 0.02967f
C9393 VDD.n950 GND 0.02522f
C9394 VDD.n951 GND 0.04999f
C9395 VDD.t346 GND 0.63568f
C9396 VDD.n952 GND 0.05074f
C9397 VDD.n953 GND 0.05074f
C9398 VDD.n954 GND 0.02967f
C9399 VDD.n955 GND 0.02522f
C9400 VDD.t173 GND 0.02321f
C9401 VDD.t347 GND 0.02321f
C9402 VDD.n956 GND 0.10855f
C9403 VDD.t909 GND 0.02321f
C9404 VDD.t348 GND 0.02321f
C9405 VDD.n957 GND 0.10855f
C9406 VDD.n958 GND 0.04152f
C9407 VDD.n959 GND 0.02334f
C9408 VDD.n960 GND 0.0536f
C9409 VDD.n961 GND 0.05074f
C9410 VDD.n962 GND 0.02967f
C9411 VDD.n963 GND 0.02522f
C9412 VDD.n964 GND 0.04999f
C9413 VDD.t9 GND 0.63568f
C9414 VDD.n965 GND 0.05074f
C9415 VDD.n966 GND 0.05074f
C9416 VDD.n967 GND 0.02967f
C9417 VDD.n968 GND 0.02522f
C9418 VDD.t625 GND 0.02334f
C9419 VDD.t10 GND 0.02334f
C9420 VDD.n969 GND 0.13341f
C9421 VDD.n970 GND 0.0263f
C9422 VDD.n971 GND 0.0536f
C9423 VDD.n972 GND 0.05074f
C9424 VDD.n973 GND 0.02967f
C9425 VDD.n974 GND 0.02522f
C9426 VDD.n975 GND 0.04999f
C9427 VDD.t318 GND 0.63568f
C9428 VDD.n976 GND 0.05074f
C9429 VDD.n977 GND 0.05074f
C9430 VDD.n978 GND 0.02967f
C9431 VDD.n979 GND 0.02522f
C9432 VDD.n980 GND 0.03166f
C9433 VDD.n981 GND 0.0536f
C9434 VDD.n982 GND 0.05074f
C9435 VDD.n983 GND 0.02967f
C9436 VDD.n984 GND 0.02522f
C9437 VDD.n985 GND 0.04999f
C9438 VDD.t808 GND 0.63568f
C9439 VDD.n986 GND 0.05074f
C9440 VDD.n987 GND 0.05074f
C9441 VDD.n988 GND 0.02967f
C9442 VDD.n989 GND 0.02522f
C9443 VDD.t540 GND 0.02321f
C9444 VDD.t825 GND 0.02321f
C9445 VDD.n990 GND 0.10855f
C9446 VDD.t319 GND 0.02321f
C9447 VDD.t809 GND 0.02321f
C9448 VDD.n991 GND 0.10855f
C9449 VDD.n992 GND 0.04152f
C9450 VDD.n993 GND 0.02334f
C9451 VDD.n994 GND 0.0536f
C9452 VDD.n995 GND 0.05074f
C9453 VDD.n996 GND 0.02967f
C9454 VDD.n997 GND 0.02522f
C9455 VDD.n998 GND 0.02522f
C9456 VDD.n999 GND 0.04999f
C9457 VDD.n1000 GND 0.68843f
C9458 VDD.n1001 GND 0.04999f
C9459 VDD.n1002 GND 0.05074f
C9460 VDD.n1003 GND 0.06295f
C9461 VDD.n1004 GND 0.0536f
C9462 VDD.n1005 GND 0.02522f
C9463 VDD.n1006 GND 0.04999f
C9464 VDD.n1007 GND 0.5126f
C9465 VDD.n1008 GND 0.02522f
C9466 VDD.n1009 GND 0.04999f
C9467 VDD.n1010 GND 0.5126f
C9468 VDD.n1011 GND 0.04999f
C9469 VDD.n1012 GND 0.05074f
C9470 VDD.n1013 GND 0.06295f
C9471 VDD.n1014 GND 0.0536f
C9472 VDD.n1015 GND 0.02522f
C9473 VDD.n1016 GND 0.04999f
C9474 VDD.n1017 GND 0.5126f
C9475 VDD.n1018 GND 0.02522f
C9476 VDD.n1019 GND 0.04999f
C9477 VDD.n1020 GND 0.5126f
C9478 VDD.n1021 GND 0.04999f
C9479 VDD.n1022 GND 0.05074f
C9480 VDD.n1023 GND 0.06295f
C9481 VDD.n1024 GND 0.0536f
C9482 VDD.n1025 GND 0.02522f
C9483 VDD.n1026 GND 0.04999f
C9484 VDD.n1027 GND 0.68843f
C9485 VDD.n1028 GND 0.02522f
C9486 VDD.n1029 GND 0.04999f
C9487 VDD.n1030 GND 0.68843f
C9488 VDD.n1031 GND 0.04999f
C9489 VDD.n1032 GND 0.05074f
C9490 VDD.n1033 GND 0.06295f
C9491 VDD.n1034 GND 0.0536f
C9492 VDD.n1035 GND 0.02522f
C9493 VDD.n1036 GND 0.04999f
C9494 VDD.n1037 GND 0.5126f
C9495 VDD.n1038 GND 0.02522f
C9496 VDD.n1039 GND 0.04999f
C9497 VDD.n1040 GND 0.5126f
C9498 VDD.n1041 GND 0.04999f
C9499 VDD.n1042 GND 0.05074f
C9500 VDD.n1043 GND 0.06295f
C9501 VDD.n1044 GND 0.0536f
C9502 VDD.n1045 GND 0.02522f
C9503 VDD.n1046 GND 0.04999f
C9504 VDD.n1047 GND 0.68843f
C9505 VDD.n1048 GND 0.68843f
C9506 VDD.n1049 GND 0.04999f
C9507 VDD.n1050 GND 0.02746f
C9508 VDD.n1051 GND 0.02967f
C9509 VDD.n1052 GND 0.02746f
C9510 VDD.n1053 GND 0.04999f
C9511 VDD.n1054 GND 0.68843f
C9512 VDD.n1055 GND 0.02522f
C9513 VDD.n1056 GND 0.04999f
C9514 VDD.n1057 GND 0.68843f
C9515 VDD.n1058 GND 0.04999f
C9516 VDD.n1059 GND 0.05074f
C9517 VDD.n1060 GND 0.06295f
C9518 VDD.n1061 GND 0.0536f
C9519 VDD.n1062 GND 0.02522f
C9520 VDD.n1063 GND 0.04999f
C9521 VDD.n1064 GND 0.5126f
C9522 VDD.n1065 GND 0.02522f
C9523 VDD.n1066 GND 0.04999f
C9524 VDD.n1067 GND 0.5126f
C9525 VDD.n1068 GND 0.04999f
C9526 VDD.n1069 GND 0.05074f
C9527 VDD.n1070 GND 0.06295f
C9528 VDD.n1071 GND 0.0536f
C9529 VDD.n1072 GND 0.02522f
C9530 VDD.n1073 GND 0.04999f
C9531 VDD.n1074 GND 0.5126f
C9532 VDD.n1075 GND 0.02522f
C9533 VDD.n1076 GND 0.04999f
C9534 VDD.n1077 GND 0.5126f
C9535 VDD.n1078 GND 0.04999f
C9536 VDD.n1079 GND 0.05074f
C9537 VDD.n1080 GND 0.06295f
C9538 VDD.n1081 GND 0.0536f
C9539 VDD.n1082 GND 0.02522f
C9540 VDD.n1083 GND 0.04999f
C9541 VDD.n1084 GND 0.68843f
C9542 VDD.n1085 GND 0.02522f
C9543 VDD.n1086 GND 0.04999f
C9544 VDD.n1087 GND 0.68843f
C9545 VDD.n1088 GND 0.04999f
C9546 VDD.n1089 GND 0.05074f
C9547 VDD.n1090 GND 0.06295f
C9548 VDD.n1091 GND 0.0536f
C9549 VDD.n1092 GND 0.02522f
C9550 VDD.n1093 GND 0.04999f
C9551 VDD.n1094 GND 0.5126f
C9552 VDD.n1095 GND 0.02522f
C9553 VDD.n1096 GND 0.04999f
C9554 VDD.n1097 GND 0.5126f
C9555 VDD.n1098 GND 0.04999f
C9556 VDD.n1099 GND 0.05074f
C9557 VDD.n1100 GND 0.06295f
C9558 VDD.n1101 GND 0.0536f
C9559 VDD.n1102 GND 0.02522f
C9560 VDD.n1103 GND 0.04999f
C9561 VDD.n1104 GND 0.5126f
C9562 VDD.n1105 GND 0.02522f
C9563 VDD.n1106 GND 0.04999f
C9564 VDD.n1107 GND 0.5126f
C9565 VDD.n1108 GND 0.04999f
C9566 VDD.n1109 GND 0.05074f
C9567 VDD.n1110 GND 0.06295f
C9568 VDD.n1111 GND 0.0536f
C9569 VDD.n1112 GND 0.02522f
C9570 VDD.n1113 GND 0.04999f
C9571 VDD.n1114 GND 0.68843f
C9572 VDD.n1115 GND 0.68843f
C9573 VDD.n1116 GND 0.04999f
C9574 VDD.n1117 GND 0.02746f
C9575 VDD.n1118 GND 0.09132f
C9576 VDD.n1119 GND 0.01798f
C9577 VDD.n1120 GND 0.09868f
C9578 VDD.n1121 GND 0.3275f
C9579 VDD.t962 GND 0.02334f
C9580 VDD.n1122 GND 0.02746f
C9581 VDD.n1123 GND 0.05074f
C9582 VDD.n1124 GND 0.02967f
C9583 VDD.n1125 GND 0.05074f
C9584 VDD.n1126 GND 0.62973f
C9585 VDD.t961 GND 0.74438f
C9586 VDD.n1128 GND 0.04999f
C9587 VDD.t480 GND 0.63568f
C9588 VDD.n1129 GND 0.05074f
C9589 VDD.n1130 GND 0.05074f
C9590 VDD.n1131 GND 0.02967f
C9591 VDD.n1132 GND 0.02522f
C9592 VDD.t481 GND 0.02334f
C9593 VDD.t883 GND 0.02334f
C9594 VDD.n1133 GND 0.13341f
C9595 VDD.n1134 GND 0.0263f
C9596 VDD.n1135 GND 0.0536f
C9597 VDD.n1136 GND 0.05074f
C9598 VDD.n1137 GND 0.02967f
C9599 VDD.n1138 GND 0.02522f
C9600 VDD.n1139 GND 0.04999f
C9601 VDD.t393 GND 0.63568f
C9602 VDD.n1140 GND 0.05074f
C9603 VDD.n1141 GND 0.05074f
C9604 VDD.n1142 GND 0.02967f
C9605 VDD.n1143 GND 0.02522f
C9606 VDD.n1144 GND 0.03166f
C9607 VDD.n1145 GND 0.0536f
C9608 VDD.n1146 GND 0.05074f
C9609 VDD.n1147 GND 0.02967f
C9610 VDD.n1148 GND 0.02522f
C9611 VDD.n1149 GND 0.04999f
C9612 VDD.t101 GND 0.63568f
C9613 VDD.n1150 GND 0.05074f
C9614 VDD.n1151 GND 0.05074f
C9615 VDD.n1152 GND 0.02967f
C9616 VDD.n1153 GND 0.02522f
C9617 VDD.t394 GND 0.02321f
C9618 VDD.t102 GND 0.02321f
C9619 VDD.n1154 GND 0.10855f
C9620 VDD.t638 GND 0.02321f
C9621 VDD.t275 GND 0.02321f
C9622 VDD.n1155 GND 0.10855f
C9623 VDD.n1156 GND 0.04152f
C9624 VDD.n1157 GND 0.02334f
C9625 VDD.n1158 GND 0.0536f
C9626 VDD.n1159 GND 0.05074f
C9627 VDD.n1160 GND 0.02967f
C9628 VDD.n1161 GND 0.02522f
C9629 VDD.n1162 GND 0.04999f
C9630 VDD.t538 GND 0.63568f
C9631 VDD.n1163 GND 0.05074f
C9632 VDD.n1164 GND 0.05074f
C9633 VDD.n1165 GND 0.02967f
C9634 VDD.n1166 GND 0.02522f
C9635 VDD.t880 GND 0.02334f
C9636 VDD.t539 GND 0.02334f
C9637 VDD.n1167 GND 0.13341f
C9638 VDD.n1168 GND 0.0263f
C9639 VDD.n1169 GND 0.0536f
C9640 VDD.n1170 GND 0.05074f
C9641 VDD.n1171 GND 0.02967f
C9642 VDD.n1172 GND 0.02522f
C9643 VDD.n1173 GND 0.04999f
C9644 VDD.t412 GND 0.63568f
C9645 VDD.n1174 GND 0.05074f
C9646 VDD.n1175 GND 0.05074f
C9647 VDD.n1176 GND 0.02967f
C9648 VDD.n1177 GND 0.02522f
C9649 VDD.n1178 GND 0.03166f
C9650 VDD.n1179 GND 0.0536f
C9651 VDD.n1180 GND 0.05074f
C9652 VDD.n1181 GND 0.02967f
C9653 VDD.n1182 GND 0.02522f
C9654 VDD.n1183 GND 0.04999f
C9655 VDD.t778 GND 0.63568f
C9656 VDD.n1184 GND 0.05074f
C9657 VDD.n1185 GND 0.05074f
C9658 VDD.n1186 GND 0.02967f
C9659 VDD.n1187 GND 0.02522f
C9660 VDD.t413 GND 0.02321f
C9661 VDD.t779 GND 0.02321f
C9662 VDD.n1188 GND 0.10855f
C9663 VDD.t550 GND 0.02321f
C9664 VDD.t966 GND 0.02321f
C9665 VDD.n1189 GND 0.10855f
C9666 VDD.n1190 GND 0.04152f
C9667 VDD.n1191 GND 0.02334f
C9668 VDD.n1192 GND 0.0536f
C9669 VDD.n1193 GND 0.05074f
C9670 VDD.n1194 GND 0.02967f
C9671 VDD.n1195 GND 0.02522f
C9672 VDD.t103 GND 0.63568f
C9673 VDD.n1196 GND 0.05074f
C9674 VDD.n1197 GND 0.05074f
C9675 VDD.n1198 GND 0.09132f
C9676 VDD.n1199 GND 0.04999f
C9677 VDD.t191 GND 0.63568f
C9678 VDD.n1200 GND 0.05074f
C9679 VDD.n1201 GND 0.05074f
C9680 VDD.n1202 GND 0.02967f
C9681 VDD.n1203 GND 0.02522f
C9682 VDD.t104 GND 0.02334f
C9683 VDD.n1204 GND 0.0731f
C9684 VDD.n1205 GND 0.01798f
C9685 VDD.n1206 GND 0.02334f
C9686 VDD.n1207 GND 0.0536f
C9687 VDD.n1208 GND 0.05074f
C9688 VDD.n1209 GND 0.02967f
C9689 VDD.n1210 GND 0.02522f
C9690 VDD.n1211 GND 0.04999f
C9691 VDD.t178 GND 0.63568f
C9692 VDD.n1212 GND 0.05074f
C9693 VDD.n1213 GND 0.05074f
C9694 VDD.n1214 GND 0.02967f
C9695 VDD.n1215 GND 0.02522f
C9696 VDD.t192 GND 0.02321f
C9697 VDD.t180 GND 0.02321f
C9698 VDD.n1216 GND 0.10855f
C9699 VDD.t777 GND 0.02321f
C9700 VDD.t179 GND 0.02321f
C9701 VDD.n1217 GND 0.10855f
C9702 VDD.n1218 GND 0.04152f
C9703 VDD.n1219 GND 0.02334f
C9704 VDD.n1220 GND 0.0536f
C9705 VDD.n1221 GND 0.05074f
C9706 VDD.n1222 GND 0.02967f
C9707 VDD.n1223 GND 0.02522f
C9708 VDD.n1224 GND 0.04999f
C9709 VDD.t211 GND 0.63568f
C9710 VDD.n1225 GND 0.05074f
C9711 VDD.n1226 GND 0.05074f
C9712 VDD.n1227 GND 0.02967f
C9713 VDD.n1228 GND 0.02522f
C9714 VDD.t212 GND 0.02334f
C9715 VDD.t477 GND 0.02334f
C9716 VDD.n1229 GND 0.13341f
C9717 VDD.n1230 GND 0.0263f
C9718 VDD.n1231 GND 0.0536f
C9719 VDD.n1232 GND 0.05074f
C9720 VDD.n1233 GND 0.02967f
C9721 VDD.n1234 GND 0.02522f
C9722 VDD.n1235 GND 0.04999f
C9723 VDD.t360 GND 0.63568f
C9724 VDD.n1236 GND 0.05074f
C9725 VDD.n1237 GND 0.05074f
C9726 VDD.n1238 GND 0.02967f
C9727 VDD.n1239 GND 0.02522f
C9728 VDD.n1240 GND 0.03166f
C9729 VDD.n1241 GND 0.0536f
C9730 VDD.n1242 GND 0.05074f
C9731 VDD.n1243 GND 0.02967f
C9732 VDD.n1244 GND 0.02522f
C9733 VDD.n1245 GND 0.04999f
C9734 VDD.t114 GND 0.63568f
C9735 VDD.n1246 GND 0.05074f
C9736 VDD.n1247 GND 0.05074f
C9737 VDD.n1248 GND 0.02967f
C9738 VDD.n1249 GND 0.02522f
C9739 VDD.t615 GND 0.02321f
C9740 VDD.t115 GND 0.02321f
C9741 VDD.n1250 GND 0.10855f
C9742 VDD.t361 GND 0.02321f
C9743 VDD.t269 GND 0.02321f
C9744 VDD.n1251 GND 0.10855f
C9745 VDD.n1252 GND 0.04152f
C9746 VDD.n1253 GND 0.02334f
C9747 VDD.n1254 GND 0.0536f
C9748 VDD.n1255 GND 0.05074f
C9749 VDD.n1256 GND 0.02967f
C9750 VDD.n1257 GND 0.02522f
C9751 VDD.n1258 GND 0.02522f
C9752 VDD.n1259 GND 0.04999f
C9753 VDD.n1260 GND 0.68843f
C9754 VDD.n1261 GND 0.04999f
C9755 VDD.n1262 GND 0.05074f
C9756 VDD.n1263 GND 0.06295f
C9757 VDD.n1264 GND 0.0536f
C9758 VDD.n1265 GND 0.02522f
C9759 VDD.n1266 GND 0.04999f
C9760 VDD.n1267 GND 0.5126f
C9761 VDD.n1268 GND 0.02522f
C9762 VDD.n1269 GND 0.04999f
C9763 VDD.n1270 GND 0.5126f
C9764 VDD.n1271 GND 0.04999f
C9765 VDD.n1272 GND 0.05074f
C9766 VDD.n1273 GND 0.06295f
C9767 VDD.n1274 GND 0.0536f
C9768 VDD.n1275 GND 0.02522f
C9769 VDD.n1276 GND 0.04999f
C9770 VDD.n1277 GND 0.5126f
C9771 VDD.n1278 GND 0.02522f
C9772 VDD.n1279 GND 0.04999f
C9773 VDD.n1280 GND 0.5126f
C9774 VDD.n1281 GND 0.04999f
C9775 VDD.n1282 GND 0.05074f
C9776 VDD.n1283 GND 0.06295f
C9777 VDD.n1284 GND 0.0536f
C9778 VDD.n1285 GND 0.02522f
C9779 VDD.n1286 GND 0.04999f
C9780 VDD.n1287 GND 0.68843f
C9781 VDD.n1288 GND 0.02522f
C9782 VDD.n1289 GND 0.04999f
C9783 VDD.n1290 GND 0.68843f
C9784 VDD.n1291 GND 0.04999f
C9785 VDD.n1292 GND 0.05074f
C9786 VDD.n1293 GND 0.06295f
C9787 VDD.n1294 GND 0.0536f
C9788 VDD.n1295 GND 0.02522f
C9789 VDD.n1296 GND 0.04999f
C9790 VDD.n1297 GND 0.5126f
C9791 VDD.n1298 GND 0.02522f
C9792 VDD.n1299 GND 0.04999f
C9793 VDD.n1300 GND 0.5126f
C9794 VDD.n1301 GND 0.04999f
C9795 VDD.n1302 GND 0.05074f
C9796 VDD.n1303 GND 0.06295f
C9797 VDD.n1304 GND 0.0536f
C9798 VDD.n1305 GND 0.02522f
C9799 VDD.n1306 GND 0.04999f
C9800 VDD.n1307 GND 0.68843f
C9801 VDD.n1308 GND 0.68843f
C9802 VDD.n1309 GND 0.04999f
C9803 VDD.n1310 GND 0.02746f
C9804 VDD.n1311 GND 0.02967f
C9805 VDD.n1312 GND 0.02746f
C9806 VDD.n1313 GND 0.04999f
C9807 VDD.n1314 GND 0.68843f
C9808 VDD.n1315 GND 0.02522f
C9809 VDD.n1316 GND 0.04999f
C9810 VDD.n1317 GND 0.68843f
C9811 VDD.n1318 GND 0.04999f
C9812 VDD.n1319 GND 0.05074f
C9813 VDD.n1320 GND 0.06295f
C9814 VDD.n1321 GND 0.0536f
C9815 VDD.n1322 GND 0.02522f
C9816 VDD.n1323 GND 0.04999f
C9817 VDD.n1324 GND 0.5126f
C9818 VDD.n1325 GND 0.02522f
C9819 VDD.n1326 GND 0.04999f
C9820 VDD.n1327 GND 0.5126f
C9821 VDD.n1328 GND 0.04999f
C9822 VDD.n1329 GND 0.05074f
C9823 VDD.n1330 GND 0.06295f
C9824 VDD.n1331 GND 0.0536f
C9825 VDD.n1332 GND 0.02522f
C9826 VDD.n1333 GND 0.04999f
C9827 VDD.n1334 GND 0.5126f
C9828 VDD.n1335 GND 0.02522f
C9829 VDD.n1336 GND 0.04999f
C9830 VDD.n1337 GND 0.5126f
C9831 VDD.n1338 GND 0.04999f
C9832 VDD.n1339 GND 0.05074f
C9833 VDD.n1340 GND 0.06295f
C9834 VDD.n1341 GND 0.0536f
C9835 VDD.n1342 GND 0.02522f
C9836 VDD.n1343 GND 0.04999f
C9837 VDD.n1344 GND 0.68843f
C9838 VDD.n1345 GND 0.02522f
C9839 VDD.n1346 GND 0.04999f
C9840 VDD.n1347 GND 0.68843f
C9841 VDD.n1348 GND 0.04999f
C9842 VDD.n1349 GND 0.05074f
C9843 VDD.n1350 GND 0.06295f
C9844 VDD.n1351 GND 0.0536f
C9845 VDD.n1352 GND 0.02522f
C9846 VDD.n1353 GND 0.04999f
C9847 VDD.n1354 GND 0.5126f
C9848 VDD.n1355 GND 0.02522f
C9849 VDD.n1356 GND 0.04999f
C9850 VDD.n1357 GND 0.5126f
C9851 VDD.n1358 GND 0.04999f
C9852 VDD.n1359 GND 0.05074f
C9853 VDD.n1360 GND 0.06295f
C9854 VDD.n1361 GND 0.0536f
C9855 VDD.n1362 GND 0.02522f
C9856 VDD.n1363 GND 0.04999f
C9857 VDD.n1364 GND 0.5126f
C9858 VDD.n1365 GND 0.02522f
C9859 VDD.n1366 GND 0.04999f
C9860 VDD.n1367 GND 0.5126f
C9861 VDD.n1368 GND 0.04999f
C9862 VDD.n1369 GND 0.05074f
C9863 VDD.n1370 GND 0.06295f
C9864 VDD.n1371 GND 0.0536f
C9865 VDD.n1372 GND 0.02522f
C9866 VDD.n1373 GND 0.04999f
C9867 VDD.n1374 GND 0.68843f
C9868 VDD.n1375 GND 0.68843f
C9869 VDD.n1376 GND 0.04999f
C9870 VDD.n1377 GND 0.02746f
C9871 VDD.n1378 GND 0.09132f
C9872 VDD.n1379 GND 0.01798f
C9873 VDD.n1380 GND 0.09868f
C9874 VDD.n1381 GND 0.42233f
C9875 VDD.t610 GND 0.02334f
C9876 VDD.n1382 GND 0.02746f
C9877 VDD.n1383 GND 0.05074f
C9878 VDD.n1384 GND 0.02967f
C9879 VDD.n1385 GND 0.05074f
C9880 VDD.n1386 GND 0.62973f
C9881 VDD.t609 GND 0.74438f
C9882 VDD.n1388 GND 0.04999f
C9883 VDD.t418 GND 0.63568f
C9884 VDD.n1389 GND 0.05074f
C9885 VDD.n1390 GND 0.05074f
C9886 VDD.n1391 GND 0.02967f
C9887 VDD.n1392 GND 0.02522f
C9888 VDD.t641 GND 0.02334f
C9889 VDD.t419 GND 0.02334f
C9890 VDD.n1393 GND 0.13341f
C9891 VDD.n1394 GND 0.0263f
C9892 VDD.n1395 GND 0.0536f
C9893 VDD.n1396 GND 0.05074f
C9894 VDD.n1397 GND 0.02967f
C9895 VDD.n1398 GND 0.02522f
C9896 VDD.n1399 GND 0.04999f
C9897 VDD.t806 GND 0.63568f
C9898 VDD.n1400 GND 0.05074f
C9899 VDD.n1401 GND 0.05074f
C9900 VDD.n1402 GND 0.02967f
C9901 VDD.n1403 GND 0.02522f
C9902 VDD.n1404 GND 0.03166f
C9903 VDD.n1405 GND 0.0536f
C9904 VDD.n1406 GND 0.05074f
C9905 VDD.n1407 GND 0.02967f
C9906 VDD.n1408 GND 0.02522f
C9907 VDD.n1409 GND 0.04999f
C9908 VDD.t4 GND 0.63568f
C9909 VDD.n1410 GND 0.05074f
C9910 VDD.n1411 GND 0.05074f
C9911 VDD.n1412 GND 0.02967f
C9912 VDD.n1413 GND 0.02522f
C9913 VDD.t807 GND 0.02321f
C9914 VDD.t5 GND 0.02321f
C9915 VDD.n1414 GND 0.10855f
C9916 VDD.t982 GND 0.02321f
C9917 VDD.t8 GND 0.02321f
C9918 VDD.n1415 GND 0.10855f
C9919 VDD.n1416 GND 0.04152f
C9920 VDD.n1417 GND 0.02334f
C9921 VDD.n1418 GND 0.0536f
C9922 VDD.n1419 GND 0.05074f
C9923 VDD.n1420 GND 0.02967f
C9924 VDD.n1421 GND 0.02522f
C9925 VDD.n1422 GND 0.04999f
C9926 VDD.t15 GND 0.63568f
C9927 VDD.n1423 GND 0.05074f
C9928 VDD.n1424 GND 0.05074f
C9929 VDD.n1425 GND 0.02967f
C9930 VDD.n1426 GND 0.02522f
C9931 VDD.t417 GND 0.02334f
C9932 VDD.t16 GND 0.02334f
C9933 VDD.n1427 GND 0.13341f
C9934 VDD.n1428 GND 0.0263f
C9935 VDD.n1429 GND 0.0536f
C9936 VDD.n1430 GND 0.05074f
C9937 VDD.n1431 GND 0.02967f
C9938 VDD.n1432 GND 0.02522f
C9939 VDD.n1433 GND 0.04999f
C9940 VDD.t93 GND 0.63568f
C9941 VDD.n1434 GND 0.05074f
C9942 VDD.n1435 GND 0.05074f
C9943 VDD.n1436 GND 0.02967f
C9944 VDD.n1437 GND 0.02522f
C9945 VDD.n1438 GND 0.03166f
C9946 VDD.n1439 GND 0.0536f
C9947 VDD.n1440 GND 0.05074f
C9948 VDD.n1441 GND 0.02967f
C9949 VDD.n1442 GND 0.02522f
C9950 VDD.n1443 GND 0.04999f
C9951 VDD.t769 GND 0.63568f
C9952 VDD.n1444 GND 0.05074f
C9953 VDD.n1445 GND 0.05074f
C9954 VDD.n1446 GND 0.02967f
C9955 VDD.n1447 GND 0.02522f
C9956 VDD.t392 GND 0.02321f
C9957 VDD.t770 GND 0.02321f
C9958 VDD.n1448 GND 0.10855f
C9959 VDD.t94 GND 0.02321f
C9960 VDD.t929 GND 0.02321f
C9961 VDD.n1449 GND 0.10855f
C9962 VDD.n1450 GND 0.04152f
C9963 VDD.n1451 GND 0.02334f
C9964 VDD.n1452 GND 0.0536f
C9965 VDD.n1453 GND 0.05074f
C9966 VDD.n1454 GND 0.02967f
C9967 VDD.n1455 GND 0.02522f
C9968 VDD.t6 GND 0.63568f
C9969 VDD.n1456 GND 0.05074f
C9970 VDD.n1457 GND 0.05074f
C9971 VDD.n1458 GND 0.09132f
C9972 VDD.n1459 GND 0.04999f
C9973 VDD.t771 GND 0.63568f
C9974 VDD.n1460 GND 0.05074f
C9975 VDD.n1461 GND 0.05074f
C9976 VDD.n1462 GND 0.02967f
C9977 VDD.n1463 GND 0.02522f
C9978 VDD.t7 GND 0.02334f
C9979 VDD.n1464 GND 0.0731f
C9980 VDD.n1465 GND 0.01798f
C9981 VDD.n1466 GND 0.02334f
C9982 VDD.n1467 GND 0.0536f
C9983 VDD.n1468 GND 0.05074f
C9984 VDD.n1469 GND 0.02967f
C9985 VDD.n1470 GND 0.02522f
C9986 VDD.n1471 GND 0.04999f
C9987 VDD.t815 GND 0.63568f
C9988 VDD.n1472 GND 0.05074f
C9989 VDD.n1473 GND 0.05074f
C9990 VDD.n1474 GND 0.02967f
C9991 VDD.n1475 GND 0.02522f
C9992 VDD.t928 GND 0.02321f
C9993 VDD.t817 GND 0.02321f
C9994 VDD.n1476 GND 0.10855f
C9995 VDD.t772 GND 0.02321f
C9996 VDD.t816 GND 0.02321f
C9997 VDD.n1477 GND 0.10855f
C9998 VDD.n1478 GND 0.04152f
C9999 VDD.n1479 GND 0.02334f
C10000 VDD.n1480 GND 0.0536f
C10001 VDD.n1481 GND 0.05074f
C10002 VDD.n1482 GND 0.02967f
C10003 VDD.n1483 GND 0.02522f
C10004 VDD.n1484 GND 0.04999f
C10005 VDD.t644 GND 0.63568f
C10006 VDD.n1485 GND 0.05074f
C10007 VDD.n1486 GND 0.05074f
C10008 VDD.n1487 GND 0.02967f
C10009 VDD.n1488 GND 0.02522f
C10010 VDD.t895 GND 0.02334f
C10011 VDD.t645 GND 0.02334f
C10012 VDD.n1489 GND 0.13341f
C10013 VDD.n1490 GND 0.0263f
C10014 VDD.n1491 GND 0.0536f
C10015 VDD.n1492 GND 0.05074f
C10016 VDD.n1493 GND 0.02967f
C10017 VDD.n1494 GND 0.02522f
C10018 VDD.n1495 GND 0.04999f
C10019 VDD.t298 GND 0.63568f
C10020 VDD.n1496 GND 0.05074f
C10021 VDD.n1497 GND 0.05074f
C10022 VDD.n1498 GND 0.02967f
C10023 VDD.n1499 GND 0.02522f
C10024 VDD.n1500 GND 0.03166f
C10025 VDD.n1501 GND 0.0536f
C10026 VDD.n1502 GND 0.05074f
C10027 VDD.n1503 GND 0.02967f
C10028 VDD.n1504 GND 0.02522f
C10029 VDD.n1505 GND 0.04999f
C10030 VDD.t994 GND 0.63568f
C10031 VDD.n1506 GND 0.05074f
C10032 VDD.n1507 GND 0.05074f
C10033 VDD.n1508 GND 0.02967f
C10034 VDD.n1509 GND 0.02522f
C10035 VDD.t299 GND 0.02321f
C10036 VDD.t1107 GND 0.02321f
C10037 VDD.n1510 GND 0.10855f
C10038 VDD.t826 GND 0.02321f
C10039 VDD.t995 GND 0.02321f
C10040 VDD.n1511 GND 0.10855f
C10041 VDD.n1512 GND 0.04152f
C10042 VDD.n1513 GND 0.02334f
C10043 VDD.n1514 GND 0.0536f
C10044 VDD.n1515 GND 0.05074f
C10045 VDD.n1516 GND 0.02967f
C10046 VDD.n1517 GND 0.02522f
C10047 VDD.n1518 GND 0.02522f
C10048 VDD.n1519 GND 0.04999f
C10049 VDD.n1520 GND 0.68843f
C10050 VDD.n1521 GND 0.04999f
C10051 VDD.n1522 GND 0.05074f
C10052 VDD.n1523 GND 0.06295f
C10053 VDD.n1524 GND 0.0536f
C10054 VDD.n1525 GND 0.02522f
C10055 VDD.n1526 GND 0.04999f
C10056 VDD.n1527 GND 0.5126f
C10057 VDD.n1528 GND 0.02522f
C10058 VDD.n1529 GND 0.04999f
C10059 VDD.n1530 GND 0.5126f
C10060 VDD.n1531 GND 0.04999f
C10061 VDD.n1532 GND 0.05074f
C10062 VDD.n1533 GND 0.06295f
C10063 VDD.n1534 GND 0.0536f
C10064 VDD.n1535 GND 0.02522f
C10065 VDD.n1536 GND 0.04999f
C10066 VDD.n1537 GND 0.5126f
C10067 VDD.n1538 GND 0.02522f
C10068 VDD.n1539 GND 0.04999f
C10069 VDD.n1540 GND 0.5126f
C10070 VDD.n1541 GND 0.04999f
C10071 VDD.n1542 GND 0.05074f
C10072 VDD.n1543 GND 0.06295f
C10073 VDD.n1544 GND 0.0536f
C10074 VDD.n1545 GND 0.02522f
C10075 VDD.n1546 GND 0.04999f
C10076 VDD.n1547 GND 0.68843f
C10077 VDD.n1548 GND 0.02522f
C10078 VDD.n1549 GND 0.04999f
C10079 VDD.n1550 GND 0.68843f
C10080 VDD.n1551 GND 0.04999f
C10081 VDD.n1552 GND 0.05074f
C10082 VDD.n1553 GND 0.06295f
C10083 VDD.n1554 GND 0.0536f
C10084 VDD.n1555 GND 0.02522f
C10085 VDD.n1556 GND 0.04999f
C10086 VDD.n1557 GND 0.5126f
C10087 VDD.n1558 GND 0.02522f
C10088 VDD.n1559 GND 0.04999f
C10089 VDD.n1560 GND 0.5126f
C10090 VDD.n1561 GND 0.04999f
C10091 VDD.n1562 GND 0.05074f
C10092 VDD.n1563 GND 0.06295f
C10093 VDD.n1564 GND 0.0536f
C10094 VDD.n1565 GND 0.02522f
C10095 VDD.n1566 GND 0.04999f
C10096 VDD.n1567 GND 0.68843f
C10097 VDD.n1568 GND 0.68843f
C10098 VDD.n1569 GND 0.04999f
C10099 VDD.n1570 GND 0.02746f
C10100 VDD.n1571 GND 0.02967f
C10101 VDD.n1572 GND 0.02746f
C10102 VDD.n1573 GND 0.04999f
C10103 VDD.n1574 GND 0.68843f
C10104 VDD.n1575 GND 0.02522f
C10105 VDD.n1576 GND 0.04999f
C10106 VDD.n1577 GND 0.68843f
C10107 VDD.n1578 GND 0.04999f
C10108 VDD.n1579 GND 0.05074f
C10109 VDD.n1580 GND 0.06295f
C10110 VDD.n1581 GND 0.0536f
C10111 VDD.n1582 GND 0.02522f
C10112 VDD.n1583 GND 0.04999f
C10113 VDD.n1584 GND 0.5126f
C10114 VDD.n1585 GND 0.02522f
C10115 VDD.n1586 GND 0.04999f
C10116 VDD.n1587 GND 0.5126f
C10117 VDD.n1588 GND 0.04999f
C10118 VDD.n1589 GND 0.05074f
C10119 VDD.n1590 GND 0.06295f
C10120 VDD.n1591 GND 0.0536f
C10121 VDD.n1592 GND 0.02522f
C10122 VDD.n1593 GND 0.04999f
C10123 VDD.n1594 GND 0.5126f
C10124 VDD.n1595 GND 0.02522f
C10125 VDD.n1596 GND 0.04999f
C10126 VDD.n1597 GND 0.5126f
C10127 VDD.n1598 GND 0.04999f
C10128 VDD.n1599 GND 0.05074f
C10129 VDD.n1600 GND 0.06295f
C10130 VDD.n1601 GND 0.0536f
C10131 VDD.n1602 GND 0.02522f
C10132 VDD.n1603 GND 0.04999f
C10133 VDD.n1604 GND 0.68843f
C10134 VDD.n1605 GND 0.02522f
C10135 VDD.n1606 GND 0.04999f
C10136 VDD.n1607 GND 0.68843f
C10137 VDD.n1608 GND 0.04999f
C10138 VDD.n1609 GND 0.05074f
C10139 VDD.n1610 GND 0.06295f
C10140 VDD.n1611 GND 0.0536f
C10141 VDD.n1612 GND 0.02522f
C10142 VDD.n1613 GND 0.04999f
C10143 VDD.n1614 GND 0.5126f
C10144 VDD.n1615 GND 0.02522f
C10145 VDD.n1616 GND 0.04999f
C10146 VDD.n1617 GND 0.5126f
C10147 VDD.n1618 GND 0.04999f
C10148 VDD.n1619 GND 0.05074f
C10149 VDD.n1620 GND 0.06295f
C10150 VDD.n1621 GND 0.0536f
C10151 VDD.n1622 GND 0.02522f
C10152 VDD.n1623 GND 0.04999f
C10153 VDD.n1624 GND 0.5126f
C10154 VDD.n1625 GND 0.02522f
C10155 VDD.n1626 GND 0.04999f
C10156 VDD.n1627 GND 0.5126f
C10157 VDD.n1628 GND 0.04999f
C10158 VDD.n1629 GND 0.05074f
C10159 VDD.n1630 GND 0.06295f
C10160 VDD.n1631 GND 0.0536f
C10161 VDD.n1632 GND 0.02522f
C10162 VDD.n1633 GND 0.04999f
C10163 VDD.n1634 GND 0.68843f
C10164 VDD.n1635 GND 0.68843f
C10165 VDD.n1636 GND 0.04999f
C10166 VDD.n1637 GND 0.02746f
C10167 VDD.n1638 GND 0.09132f
C10168 VDD.n1639 GND 0.01798f
C10169 VDD.n1640 GND 0.09868f
C10170 VDD.n1641 GND 0.42233f
C10171 VDD.t864 GND 0.02334f
C10172 VDD.n1642 GND 0.02746f
C10173 VDD.n1643 GND 0.05074f
C10174 VDD.n1644 GND 0.02967f
C10175 VDD.n1645 GND 0.05074f
C10176 VDD.n1646 GND 0.62973f
C10177 VDD.t863 GND 0.74438f
C10178 VDD.n1648 GND 0.04999f
C10179 VDD.t243 GND 0.63568f
C10180 VDD.n1649 GND 0.05074f
C10181 VDD.n1650 GND 0.05074f
C10182 VDD.n1651 GND 0.02967f
C10183 VDD.n1652 GND 0.02522f
C10184 VDD.t244 GND 0.02334f
C10185 VDD.t793 GND 0.02334f
C10186 VDD.n1653 GND 0.13341f
C10187 VDD.n1654 GND 0.0263f
C10188 VDD.n1655 GND 0.0536f
C10189 VDD.n1656 GND 0.05074f
C10190 VDD.n1657 GND 0.02967f
C10191 VDD.n1658 GND 0.02522f
C10192 VDD.n1659 GND 0.04999f
C10193 VDD.t599 GND 0.63568f
C10194 VDD.n1660 GND 0.05074f
C10195 VDD.n1661 GND 0.05074f
C10196 VDD.n1662 GND 0.02967f
C10197 VDD.n1663 GND 0.02522f
C10198 VDD.n1664 GND 0.03166f
C10199 VDD.n1665 GND 0.0536f
C10200 VDD.n1666 GND 0.05074f
C10201 VDD.n1667 GND 0.02967f
C10202 VDD.n1668 GND 0.02522f
C10203 VDD.n1669 GND 0.04999f
C10204 VDD.t923 GND 0.63568f
C10205 VDD.n1670 GND 0.05074f
C10206 VDD.n1671 GND 0.05074f
C10207 VDD.n1672 GND 0.02967f
C10208 VDD.n1673 GND 0.02522f
C10209 VDD.t600 GND 0.02321f
C10210 VDD.t924 GND 0.02321f
C10211 VDD.n1674 GND 0.10855f
C10212 VDD.t875 GND 0.02321f
C10213 VDD.t927 GND 0.02321f
C10214 VDD.n1675 GND 0.10855f
C10215 VDD.n1676 GND 0.04152f
C10216 VDD.n1677 GND 0.02334f
C10217 VDD.n1678 GND 0.0536f
C10218 VDD.n1679 GND 0.05074f
C10219 VDD.n1680 GND 0.02967f
C10220 VDD.n1681 GND 0.02522f
C10221 VDD.n1682 GND 0.04999f
C10222 VDD.t358 GND 0.63568f
C10223 VDD.n1683 GND 0.05074f
C10224 VDD.n1684 GND 0.05074f
C10225 VDD.n1685 GND 0.02967f
C10226 VDD.n1686 GND 0.02522f
C10227 VDD.t790 GND 0.02334f
C10228 VDD.t359 GND 0.02334f
C10229 VDD.n1687 GND 0.13341f
C10230 VDD.n1688 GND 0.0263f
C10231 VDD.n1689 GND 0.0536f
C10232 VDD.n1690 GND 0.05074f
C10233 VDD.n1691 GND 0.02967f
C10234 VDD.n1692 GND 0.02522f
C10235 VDD.n1693 GND 0.04999f
C10236 VDD.t567 GND 0.63568f
C10237 VDD.n1694 GND 0.05074f
C10238 VDD.n1695 GND 0.05074f
C10239 VDD.n1696 GND 0.02967f
C10240 VDD.n1697 GND 0.02522f
C10241 VDD.n1698 GND 0.03166f
C10242 VDD.n1699 GND 0.0536f
C10243 VDD.n1700 GND 0.05074f
C10244 VDD.n1701 GND 0.02967f
C10245 VDD.n1702 GND 0.02522f
C10246 VDD.n1703 GND 0.04999f
C10247 VDD.t597 GND 0.63568f
C10248 VDD.n1704 GND 0.05074f
C10249 VDD.n1705 GND 0.05074f
C10250 VDD.n1706 GND 0.02967f
C10251 VDD.n1707 GND 0.02522f
C10252 VDD.t568 GND 0.02321f
C10253 VDD.t991 GND 0.02321f
C10254 VDD.n1708 GND 0.10855f
C10255 VDD.t979 GND 0.02321f
C10256 VDD.t598 GND 0.02321f
C10257 VDD.n1709 GND 0.10855f
C10258 VDD.n1710 GND 0.04152f
C10259 VDD.n1711 GND 0.02334f
C10260 VDD.n1712 GND 0.0536f
C10261 VDD.n1713 GND 0.05074f
C10262 VDD.n1714 GND 0.02967f
C10263 VDD.n1715 GND 0.02522f
C10264 VDD.t925 GND 0.63568f
C10265 VDD.n1716 GND 0.05074f
C10266 VDD.n1717 GND 0.05074f
C10267 VDD.n1718 GND 0.09132f
C10268 VDD.n1719 GND 0.04999f
C10269 VDD.t595 GND 0.63568f
C10270 VDD.n1720 GND 0.05074f
C10271 VDD.n1721 GND 0.05074f
C10272 VDD.n1722 GND 0.02967f
C10273 VDD.n1723 GND 0.02522f
C10274 VDD.t926 GND 0.02334f
C10275 VDD.n1724 GND 0.0731f
C10276 VDD.n1725 GND 0.01798f
C10277 VDD.n1726 GND 0.02334f
C10278 VDD.n1727 GND 0.0536f
C10279 VDD.n1728 GND 0.05074f
C10280 VDD.n1729 GND 0.02967f
C10281 VDD.n1730 GND 0.02522f
C10282 VDD.n1731 GND 0.04999f
C10283 VDD.t157 GND 0.63568f
C10284 VDD.n1732 GND 0.05074f
C10285 VDD.n1733 GND 0.05074f
C10286 VDD.n1734 GND 0.02967f
C10287 VDD.n1735 GND 0.02522f
C10288 VDD.t596 GND 0.02321f
C10289 VDD.t158 GND 0.02321f
C10290 VDD.n1736 GND 0.10855f
C10291 VDD.t992 GND 0.02321f
C10292 VDD.t159 GND 0.02321f
C10293 VDD.n1737 GND 0.10855f
C10294 VDD.n1738 GND 0.04152f
C10295 VDD.n1739 GND 0.02334f
C10296 VDD.n1740 GND 0.0536f
C10297 VDD.n1741 GND 0.05074f
C10298 VDD.n1742 GND 0.02967f
C10299 VDD.n1743 GND 0.02522f
C10300 VDD.n1744 GND 0.04999f
C10301 VDD.t27 GND 0.63568f
C10302 VDD.n1745 GND 0.05074f
C10303 VDD.n1746 GND 0.05074f
C10304 VDD.n1747 GND 0.02967f
C10305 VDD.n1748 GND 0.02522f
C10306 VDD.t28 GND 0.02334f
C10307 VDD.t383 GND 0.02334f
C10308 VDD.n1749 GND 0.13341f
C10309 VDD.n1750 GND 0.0263f
C10310 VDD.n1751 GND 0.0536f
C10311 VDD.n1752 GND 0.05074f
C10312 VDD.n1753 GND 0.02967f
C10313 VDD.n1754 GND 0.02522f
C10314 VDD.n1755 GND 0.04999f
C10315 VDD.t422 GND 0.63568f
C10316 VDD.n1756 GND 0.05074f
C10317 VDD.n1757 GND 0.05074f
C10318 VDD.n1758 GND 0.02967f
C10319 VDD.n1759 GND 0.02522f
C10320 VDD.n1760 GND 0.03166f
C10321 VDD.n1761 GND 0.0536f
C10322 VDD.n1762 GND 0.05074f
C10323 VDD.n1763 GND 0.02967f
C10324 VDD.n1764 GND 0.02522f
C10325 VDD.n1765 GND 0.04999f
C10326 VDD.t54 GND 0.63568f
C10327 VDD.n1766 GND 0.05074f
C10328 VDD.n1767 GND 0.05074f
C10329 VDD.n1768 GND 0.02967f
C10330 VDD.n1769 GND 0.02522f
C10331 VDD.t423 GND 0.02321f
C10332 VDD.t265 GND 0.02321f
C10333 VDD.n1770 GND 0.10855f
C10334 VDD.t936 GND 0.02321f
C10335 VDD.t55 GND 0.02321f
C10336 VDD.n1771 GND 0.10855f
C10337 VDD.n1772 GND 0.04152f
C10338 VDD.n1773 GND 0.02334f
C10339 VDD.n1774 GND 0.0536f
C10340 VDD.n1775 GND 0.05074f
C10341 VDD.n1776 GND 0.02967f
C10342 VDD.n1777 GND 0.02522f
C10343 VDD.n1778 GND 0.02522f
C10344 VDD.n1779 GND 0.04999f
C10345 VDD.n1780 GND 0.68843f
C10346 VDD.n1781 GND 0.04999f
C10347 VDD.n1782 GND 0.05074f
C10348 VDD.n1783 GND 0.06295f
C10349 VDD.n1784 GND 0.0536f
C10350 VDD.n1785 GND 0.02522f
C10351 VDD.n1786 GND 0.04999f
C10352 VDD.n1787 GND 0.5126f
C10353 VDD.n1788 GND 0.02522f
C10354 VDD.n1789 GND 0.04999f
C10355 VDD.n1790 GND 0.5126f
C10356 VDD.n1791 GND 0.04999f
C10357 VDD.n1792 GND 0.05074f
C10358 VDD.n1793 GND 0.06295f
C10359 VDD.n1794 GND 0.0536f
C10360 VDD.n1795 GND 0.02522f
C10361 VDD.n1796 GND 0.04999f
C10362 VDD.n1797 GND 0.5126f
C10363 VDD.n1798 GND 0.02522f
C10364 VDD.n1799 GND 0.04999f
C10365 VDD.n1800 GND 0.5126f
C10366 VDD.n1801 GND 0.04999f
C10367 VDD.n1802 GND 0.05074f
C10368 VDD.n1803 GND 0.06295f
C10369 VDD.n1804 GND 0.0536f
C10370 VDD.n1805 GND 0.02522f
C10371 VDD.n1806 GND 0.04999f
C10372 VDD.n1807 GND 0.68843f
C10373 VDD.n1808 GND 0.02522f
C10374 VDD.n1809 GND 0.04999f
C10375 VDD.n1810 GND 0.68843f
C10376 VDD.n1811 GND 0.04999f
C10377 VDD.n1812 GND 0.05074f
C10378 VDD.n1813 GND 0.06295f
C10379 VDD.n1814 GND 0.0536f
C10380 VDD.n1815 GND 0.02522f
C10381 VDD.n1816 GND 0.04999f
C10382 VDD.n1817 GND 0.5126f
C10383 VDD.n1818 GND 0.02522f
C10384 VDD.n1819 GND 0.04999f
C10385 VDD.n1820 GND 0.5126f
C10386 VDD.n1821 GND 0.04999f
C10387 VDD.n1822 GND 0.05074f
C10388 VDD.n1823 GND 0.06295f
C10389 VDD.n1824 GND 0.0536f
C10390 VDD.n1825 GND 0.02522f
C10391 VDD.n1826 GND 0.04999f
C10392 VDD.n1827 GND 0.68843f
C10393 VDD.n1828 GND 0.68843f
C10394 VDD.n1829 GND 0.04999f
C10395 VDD.n1830 GND 0.02746f
C10396 VDD.n1831 GND 0.02967f
C10397 VDD.n1832 GND 0.02746f
C10398 VDD.n1833 GND 0.04999f
C10399 VDD.n1834 GND 0.68843f
C10400 VDD.n1835 GND 0.02522f
C10401 VDD.n1836 GND 0.04999f
C10402 VDD.n1837 GND 0.68843f
C10403 VDD.n1838 GND 0.04999f
C10404 VDD.n1839 GND 0.05074f
C10405 VDD.n1840 GND 0.06295f
C10406 VDD.n1841 GND 0.0536f
C10407 VDD.n1842 GND 0.02522f
C10408 VDD.n1843 GND 0.04999f
C10409 VDD.n1844 GND 0.5126f
C10410 VDD.n1845 GND 0.02522f
C10411 VDD.n1846 GND 0.04999f
C10412 VDD.n1847 GND 0.5126f
C10413 VDD.n1848 GND 0.04999f
C10414 VDD.n1849 GND 0.05074f
C10415 VDD.n1850 GND 0.06295f
C10416 VDD.n1851 GND 0.0536f
C10417 VDD.n1852 GND 0.02522f
C10418 VDD.n1853 GND 0.04999f
C10419 VDD.n1854 GND 0.5126f
C10420 VDD.n1855 GND 0.02522f
C10421 VDD.n1856 GND 0.04999f
C10422 VDD.n1857 GND 0.5126f
C10423 VDD.n1858 GND 0.04999f
C10424 VDD.n1859 GND 0.05074f
C10425 VDD.n1860 GND 0.06295f
C10426 VDD.n1861 GND 0.0536f
C10427 VDD.n1862 GND 0.02522f
C10428 VDD.n1863 GND 0.04999f
C10429 VDD.n1864 GND 0.68843f
C10430 VDD.n1865 GND 0.02522f
C10431 VDD.n1866 GND 0.04999f
C10432 VDD.n1867 GND 0.68843f
C10433 VDD.n1868 GND 0.04999f
C10434 VDD.n1869 GND 0.05074f
C10435 VDD.n1870 GND 0.06295f
C10436 VDD.n1871 GND 0.0536f
C10437 VDD.n1872 GND 0.02522f
C10438 VDD.n1873 GND 0.04999f
C10439 VDD.n1874 GND 0.5126f
C10440 VDD.n1875 GND 0.02522f
C10441 VDD.n1876 GND 0.04999f
C10442 VDD.n1877 GND 0.5126f
C10443 VDD.n1878 GND 0.04999f
C10444 VDD.n1879 GND 0.05074f
C10445 VDD.n1880 GND 0.06295f
C10446 VDD.n1881 GND 0.0536f
C10447 VDD.n1882 GND 0.02522f
C10448 VDD.n1883 GND 0.04999f
C10449 VDD.n1884 GND 0.5126f
C10450 VDD.n1885 GND 0.02522f
C10451 VDD.n1886 GND 0.04999f
C10452 VDD.n1887 GND 0.5126f
C10453 VDD.n1888 GND 0.04999f
C10454 VDD.n1889 GND 0.05074f
C10455 VDD.n1890 GND 0.06295f
C10456 VDD.n1891 GND 0.0536f
C10457 VDD.n1892 GND 0.02522f
C10458 VDD.n1893 GND 0.04999f
C10459 VDD.n1894 GND 0.68843f
C10460 VDD.n1895 GND 0.68843f
C10461 VDD.n1896 GND 0.04999f
C10462 VDD.n1897 GND 0.02746f
C10463 VDD.n1898 GND 0.09132f
C10464 VDD.n1899 GND 0.01798f
C10465 VDD.n1900 GND 0.09868f
C10466 VDD.n1901 GND 0.3275f
C10467 VDD.t650 GND 0.02334f
C10468 VDD.n1902 GND 0.02746f
C10469 VDD.n1903 GND 0.05074f
C10470 VDD.n1904 GND 0.02967f
C10471 VDD.n1905 GND 0.05074f
C10472 VDD.n1906 GND 0.62973f
C10473 VDD.t649 GND 0.74438f
C10474 VDD.n1908 GND 0.04999f
C10475 VDD.t439 GND 0.63568f
C10476 VDD.n1909 GND 0.05074f
C10477 VDD.n1910 GND 0.05074f
C10478 VDD.n1911 GND 0.02967f
C10479 VDD.n1912 GND 0.02522f
C10480 VDD.t733 GND 0.02334f
C10481 VDD.t440 GND 0.02334f
C10482 VDD.n1913 GND 0.13341f
C10483 VDD.n1914 GND 0.0263f
C10484 VDD.n1915 GND 0.0536f
C10485 VDD.n1916 GND 0.05074f
C10486 VDD.n1917 GND 0.02967f
C10487 VDD.n1918 GND 0.02522f
C10488 VDD.n1919 GND 0.04999f
C10489 VDD.t572 GND 0.63568f
C10490 VDD.n1920 GND 0.05074f
C10491 VDD.n1921 GND 0.05074f
C10492 VDD.n1922 GND 0.02967f
C10493 VDD.n1923 GND 0.02522f
C10494 VDD.n1924 GND 0.03166f
C10495 VDD.n1925 GND 0.0536f
C10496 VDD.n1926 GND 0.05074f
C10497 VDD.n1927 GND 0.02967f
C10498 VDD.n1928 GND 0.02522f
C10499 VDD.n1929 GND 0.04999f
C10500 VDD.t1020 GND 0.63568f
C10501 VDD.n1930 GND 0.05074f
C10502 VDD.n1931 GND 0.05074f
C10503 VDD.n1932 GND 0.02967f
C10504 VDD.n1933 GND 0.02522f
C10505 VDD.t651 GND 0.02321f
C10506 VDD.t1021 GND 0.02321f
C10507 VDD.n1934 GND 0.10855f
C10508 VDD.t573 GND 0.02321f
C10509 VDD.t1067 GND 0.02321f
C10510 VDD.n1935 GND 0.10855f
C10511 VDD.n1936 GND 0.04152f
C10512 VDD.n1937 GND 0.02334f
C10513 VDD.n1938 GND 0.0536f
C10514 VDD.n1939 GND 0.05074f
C10515 VDD.n1940 GND 0.02967f
C10516 VDD.n1941 GND 0.02522f
C10517 VDD.n1942 GND 0.04999f
C10518 VDD.t500 GND 0.63568f
C10519 VDD.n1943 GND 0.05074f
C10520 VDD.n1944 GND 0.05074f
C10521 VDD.n1945 GND 0.02967f
C10522 VDD.n1946 GND 0.02522f
C10523 VDD.t501 GND 0.02334f
C10524 VDD.t671 GND 0.02334f
C10525 VDD.n1947 GND 0.13232f
C10526 VDD.n1948 GND 0.06172f
C10527 VDD.n1950 GND 0.0536f
C10528 VDD.n1951 GND 0.05074f
C10529 VDD.n1952 GND 0.02967f
C10530 VDD.n1953 GND 0.02522f
C10531 VDD.n1954 GND 0.04999f
C10532 VDD.t149 GND 0.63568f
C10533 VDD.n1955 GND 0.05074f
C10534 VDD.n1956 GND 0.05074f
C10535 VDD.n1957 GND 0.02967f
C10536 VDD.n1958 GND 0.02522f
C10537 VDD.n1959 GND 0.0536f
C10538 VDD.n1960 GND 0.05074f
C10539 VDD.n1961 GND 0.09652f
C10540 VDD.t571 GND 0.02321f
C10541 VDD.t36 GND 0.02321f
C10542 VDD.n1962 GND 0.10855f
C10543 VDD.t150 GND 0.02321f
C10544 VDD.t105 GND 0.02321f
C10545 VDD.n1963 GND 0.10855f
C10546 VDD.n1964 GND 0.0536f
C10547 VDD.n1965 GND 0.05074f
C10548 VDD.n1966 GND 0.0536f
C10549 VDD.n1967 GND 0.04999f
C10550 VDD.n1968 GND 0.04999f
C10551 VDD.n1969 GND 0.05074f
C10552 VDD.n1970 GND 0.02967f
C10553 VDD.n1971 GND 0.02522f
C10554 VDD.n1972 GND 0.04999f
C10555 VDD.n1973 GND 0.02522f
C10556 VDD.n1974 GND 0.04999f
C10557 VDD.n1975 GND 0.5126f
C10558 VDD.n1976 GND 0.5126f
C10559 VDD.n1977 GND 0.02522f
C10560 VDD.n1978 GND 0.02522f
C10561 VDD.n1979 GND 0.02967f
C10562 VDD.n1980 GND 0.05074f
C10563 VDD.t1074 GND 0.63568f
C10564 VDD.n1981 GND 0.05074f
C10565 VDD.n1982 GND 0.05074f
C10566 VDD.n1983 GND 0.09132f
C10567 VDD.n1984 GND 0.04999f
C10568 VDD.t106 GND 0.63568f
C10569 VDD.n1985 GND 0.05074f
C10570 VDD.n1986 GND 0.05074f
C10571 VDD.n1987 GND 0.02967f
C10572 VDD.n1988 GND 0.02522f
C10573 VDD.t1075 GND 0.02334f
C10574 VDD.n1989 GND 0.0731f
C10575 VDD.n1990 GND 0.01798f
C10576 VDD.n1991 GND 0.02334f
C10577 VDD.n1992 GND 0.0536f
C10578 VDD.n1993 GND 0.05074f
C10579 VDD.n1994 GND 0.02967f
C10580 VDD.n1995 GND 0.02522f
C10581 VDD.n1996 GND 0.04999f
C10582 VDD.t29 GND 0.63568f
C10583 VDD.n1997 GND 0.05074f
C10584 VDD.n1998 GND 0.05074f
C10585 VDD.n1999 GND 0.02967f
C10586 VDD.n2000 GND 0.02522f
C10587 VDD.t768 GND 0.02321f
C10588 VDD.t30 GND 0.02321f
C10589 VDD.n2001 GND 0.10855f
C10590 VDD.t107 GND 0.02321f
C10591 VDD.t999 GND 0.02321f
C10592 VDD.n2002 GND 0.10855f
C10593 VDD.n2003 GND 0.04152f
C10594 VDD.n2004 GND 0.02334f
C10595 VDD.n2005 GND 0.0536f
C10596 VDD.n2006 GND 0.05074f
C10597 VDD.n2007 GND 0.02967f
C10598 VDD.n2008 GND 0.02522f
C10599 VDD.n2009 GND 0.04999f
C10600 VDD.t522 GND 0.63568f
C10601 VDD.n2010 GND 0.05074f
C10602 VDD.n2011 GND 0.05074f
C10603 VDD.n2012 GND 0.02967f
C10604 VDD.n2013 GND 0.02522f
C10605 VDD.t523 GND 0.02334f
C10606 VDD.t695 GND 0.02334f
C10607 VDD.n2014 GND 0.13341f
C10608 VDD.n2015 GND 0.0263f
C10609 VDD.n2016 GND 0.0536f
C10610 VDD.n2017 GND 0.05074f
C10611 VDD.n2018 GND 0.02967f
C10612 VDD.n2019 GND 0.02522f
C10613 VDD.n2020 GND 0.04999f
C10614 VDD.t193 GND 0.63568f
C10615 VDD.n2021 GND 0.05074f
C10616 VDD.n2022 GND 0.05074f
C10617 VDD.n2023 GND 0.02967f
C10618 VDD.n2024 GND 0.02522f
C10619 VDD.n2025 GND 0.03166f
C10620 VDD.n2026 GND 0.0536f
C10621 VDD.n2027 GND 0.05074f
C10622 VDD.n2028 GND 0.02967f
C10623 VDD.n2029 GND 0.02522f
C10624 VDD.n2030 GND 0.04999f
C10625 VDD.t546 GND 0.63568f
C10626 VDD.n2031 GND 0.05074f
C10627 VDD.n2032 GND 0.05074f
C10628 VDD.n2033 GND 0.02967f
C10629 VDD.n2034 GND 0.02522f
C10630 VDD.t307 GND 0.02321f
C10631 VDD.t547 GND 0.02321f
C10632 VDD.n2035 GND 0.10855f
C10633 VDD.t194 GND 0.02321f
C10634 VDD.t896 GND 0.02321f
C10635 VDD.n2036 GND 0.10855f
C10636 VDD.n2037 GND 0.04152f
C10637 VDD.t304 GND 0.02334f
C10638 VDD.n2038 GND 0.02746f
C10639 VDD.n2039 GND 0.05074f
C10640 VDD.n2040 GND 0.02967f
C10641 VDD.n2041 GND 0.05074f
C10642 VDD.n2042 GND 0.62973f
C10643 VDD.t303 GND 0.74438f
C10644 VDD.n2044 GND 0.04999f
C10645 VDD.t461 GND 0.63568f
C10646 VDD.n2045 GND 0.05074f
C10647 VDD.n2046 GND 0.05074f
C10648 VDD.n2047 GND 0.02967f
C10649 VDD.n2048 GND 0.02522f
C10650 VDD.t749 GND 0.02334f
C10651 VDD.t462 GND 0.02334f
C10652 VDD.n2049 GND 0.13341f
C10653 VDD.n2050 GND 0.0263f
C10654 VDD.n2051 GND 0.0536f
C10655 VDD.n2052 GND 0.05074f
C10656 VDD.n2053 GND 0.02967f
C10657 VDD.n2054 GND 0.02522f
C10658 VDD.n2055 GND 0.04999f
C10659 VDD.t415 GND 0.63568f
C10660 VDD.n2056 GND 0.05074f
C10661 VDD.n2057 GND 0.05074f
C10662 VDD.n2058 GND 0.02967f
C10663 VDD.n2059 GND 0.02522f
C10664 VDD.n2060 GND 0.03166f
C10665 VDD.n2061 GND 0.0536f
C10666 VDD.n2062 GND 0.05074f
C10667 VDD.n2063 GND 0.02967f
C10668 VDD.n2064 GND 0.02522f
C10669 VDD.n2065 GND 0.04999f
C10670 VDD.t1016 GND 0.63568f
C10671 VDD.n2066 GND 0.05074f
C10672 VDD.n2067 GND 0.05074f
C10673 VDD.n2068 GND 0.02967f
C10674 VDD.n2069 GND 0.02522f
C10675 VDD.t416 GND 0.02321f
C10676 VDD.t1086 GND 0.02321f
C10677 VDD.n2070 GND 0.10855f
C10678 VDD.t984 GND 0.02321f
C10679 VDD.t1017 GND 0.02321f
C10680 VDD.n2071 GND 0.10855f
C10681 VDD.n2072 GND 0.04152f
C10682 VDD.n2073 GND 0.02334f
C10683 VDD.n2074 GND 0.0536f
C10684 VDD.n2075 GND 0.05074f
C10685 VDD.n2076 GND 0.02967f
C10686 VDD.n2077 GND 0.02522f
C10687 VDD.n2078 GND 0.04999f
C10688 VDD.t526 GND 0.63568f
C10689 VDD.n2079 GND 0.05074f
C10690 VDD.n2080 GND 0.05074f
C10691 VDD.n2081 GND 0.02967f
C10692 VDD.n2082 GND 0.02522f
C10693 VDD.t527 GND 0.02334f
C10694 VDD.t701 GND 0.02334f
C10695 VDD.n2083 GND 0.13232f
C10696 VDD.n2084 GND 0.06172f
C10697 VDD.n2086 GND 0.0536f
C10698 VDD.n2087 GND 0.05074f
C10699 VDD.n2088 GND 0.02967f
C10700 VDD.n2089 GND 0.02522f
C10701 VDD.n2090 GND 0.04999f
C10702 VDD.t261 GND 0.63568f
C10703 VDD.n2091 GND 0.05074f
C10704 VDD.n2092 GND 0.05074f
C10705 VDD.n2093 GND 0.02967f
C10706 VDD.n2094 GND 0.02522f
C10707 VDD.n2095 GND 0.0536f
C10708 VDD.n2096 GND 0.05074f
C10709 VDD.n2097 GND 0.09652f
C10710 VDD.t877 GND 0.02321f
C10711 VDD.t563 GND 0.02321f
C10712 VDD.n2098 GND 0.10855f
C10713 VDD.t262 GND 0.02321f
C10714 VDD.t906 GND 0.02321f
C10715 VDD.n2099 GND 0.10855f
C10716 VDD.n2100 GND 0.0536f
C10717 VDD.n2101 GND 0.05074f
C10718 VDD.n2102 GND 0.0536f
C10719 VDD.n2103 GND 0.04999f
C10720 VDD.n2104 GND 0.04999f
C10721 VDD.n2105 GND 0.05074f
C10722 VDD.n2106 GND 0.02967f
C10723 VDD.n2107 GND 0.02522f
C10724 VDD.n2108 GND 0.04999f
C10725 VDD.n2109 GND 0.02522f
C10726 VDD.n2110 GND 0.04999f
C10727 VDD.n2111 GND 0.5126f
C10728 VDD.n2112 GND 0.5126f
C10729 VDD.n2113 GND 0.02522f
C10730 VDD.n2114 GND 0.02522f
C10731 VDD.n2115 GND 0.02967f
C10732 VDD.n2116 GND 0.05074f
C10733 VDD.t1068 GND 0.63568f
C10734 VDD.n2117 GND 0.05074f
C10735 VDD.n2118 GND 0.05074f
C10736 VDD.n2119 GND 0.09132f
C10737 VDD.n2120 GND 0.04999f
C10738 VDD.t564 GND 0.63568f
C10739 VDD.n2121 GND 0.05074f
C10740 VDD.n2122 GND 0.05074f
C10741 VDD.n2123 GND 0.02967f
C10742 VDD.n2124 GND 0.02522f
C10743 VDD.t1069 GND 0.02334f
C10744 VDD.n2125 GND 0.0731f
C10745 VDD.n2126 GND 0.01798f
C10746 VDD.n2127 GND 0.02334f
C10747 VDD.n2128 GND 0.0536f
C10748 VDD.n2129 GND 0.05074f
C10749 VDD.n2130 GND 0.02967f
C10750 VDD.n2131 GND 0.02522f
C10751 VDD.n2132 GND 0.04999f
C10752 VDD.t848 GND 0.63568f
C10753 VDD.n2133 GND 0.05074f
C10754 VDD.n2134 GND 0.05074f
C10755 VDD.n2135 GND 0.02967f
C10756 VDD.n2136 GND 0.02522f
C10757 VDD.t907 GND 0.02321f
C10758 VDD.t849 GND 0.02321f
C10759 VDD.n2137 GND 0.10855f
C10760 VDD.t565 GND 0.02321f
C10761 VDD.t1106 GND 0.02321f
C10762 VDD.n2138 GND 0.10855f
C10763 VDD.n2139 GND 0.04152f
C10764 VDD.n2140 GND 0.02334f
C10765 VDD.n2141 GND 0.0536f
C10766 VDD.n2142 GND 0.05074f
C10767 VDD.n2143 GND 0.02967f
C10768 VDD.n2144 GND 0.02522f
C10769 VDD.n2145 GND 0.04999f
C10770 VDD.t467 GND 0.63568f
C10771 VDD.n2146 GND 0.05074f
C10772 VDD.n2147 GND 0.05074f
C10773 VDD.n2148 GND 0.02967f
C10774 VDD.n2149 GND 0.02522f
C10775 VDD.t468 GND 0.02334f
C10776 VDD.t743 GND 0.02334f
C10777 VDD.n2150 GND 0.13341f
C10778 VDD.n2151 GND 0.0263f
C10779 VDD.n2152 GND 0.0536f
C10780 VDD.n2153 GND 0.05074f
C10781 VDD.n2154 GND 0.02967f
C10782 VDD.n2155 GND 0.02522f
C10783 VDD.n2156 GND 0.04999f
C10784 VDD.t634 GND 0.63568f
C10785 VDD.n2157 GND 0.05074f
C10786 VDD.n2158 GND 0.05074f
C10787 VDD.n2159 GND 0.02967f
C10788 VDD.n2160 GND 0.02522f
C10789 VDD.n2161 GND 0.03166f
C10790 VDD.n2162 GND 0.0536f
C10791 VDD.n2163 GND 0.05074f
C10792 VDD.n2164 GND 0.02967f
C10793 VDD.n2165 GND 0.02522f
C10794 VDD.n2166 GND 0.04999f
C10795 VDD.t548 GND 0.63568f
C10796 VDD.n2167 GND 0.05074f
C10797 VDD.n2168 GND 0.05074f
C10798 VDD.n2169 GND 0.02967f
C10799 VDD.n2170 GND 0.02522f
C10800 VDD.t818 GND 0.02321f
C10801 VDD.t549 GND 0.02321f
C10802 VDD.n2171 GND 0.10855f
C10803 VDD.t635 GND 0.02321f
C10804 VDD.t775 GND 0.02321f
C10805 VDD.n2172 GND 0.10855f
C10806 VDD.n2173 GND 0.04152f
C10807 VDD.t66 GND 0.02334f
C10808 VDD.n2174 GND 0.02746f
C10809 VDD.n2175 GND 0.05074f
C10810 VDD.n2176 GND 0.02967f
C10811 VDD.n2177 GND 0.05074f
C10812 VDD.n2178 GND 0.62973f
C10813 VDD.t65 GND 0.74438f
C10814 VDD.n2180 GND 0.04999f
C10815 VDD.t498 GND 0.63568f
C10816 VDD.n2181 GND 0.05074f
C10817 VDD.n2182 GND 0.05074f
C10818 VDD.n2183 GND 0.02967f
C10819 VDD.n2184 GND 0.02522f
C10820 VDD.t685 GND 0.02334f
C10821 VDD.t499 GND 0.02334f
C10822 VDD.n2185 GND 0.13341f
C10823 VDD.n2186 GND 0.0263f
C10824 VDD.n2187 GND 0.0536f
C10825 VDD.n2188 GND 0.05074f
C10826 VDD.n2189 GND 0.02967f
C10827 VDD.n2190 GND 0.02522f
C10828 VDD.n2191 GND 0.04999f
C10829 VDD.t396 GND 0.63568f
C10830 VDD.n2192 GND 0.05074f
C10831 VDD.n2193 GND 0.05074f
C10832 VDD.n2194 GND 0.02967f
C10833 VDD.n2195 GND 0.02522f
C10834 VDD.n2196 GND 0.03166f
C10835 VDD.n2197 GND 0.0536f
C10836 VDD.n2198 GND 0.05074f
C10837 VDD.n2199 GND 0.02967f
C10838 VDD.n2200 GND 0.02522f
C10839 VDD.n2201 GND 0.04999f
C10840 VDD.t1042 GND 0.63568f
C10841 VDD.n2202 GND 0.05074f
C10842 VDD.n2203 GND 0.05074f
C10843 VDD.n2204 GND 0.02967f
C10844 VDD.n2205 GND 0.02522f
C10845 VDD.t814 GND 0.02321f
C10846 VDD.t1098 GND 0.02321f
C10847 VDD.n2206 GND 0.10855f
C10848 VDD.t397 GND 0.02321f
C10849 VDD.t1043 GND 0.02321f
C10850 VDD.n2207 GND 0.10855f
C10851 VDD.n2208 GND 0.04152f
C10852 VDD.n2209 GND 0.02334f
C10853 VDD.n2210 GND 0.0536f
C10854 VDD.n2211 GND 0.05074f
C10855 VDD.n2212 GND 0.02967f
C10856 VDD.n2213 GND 0.02522f
C10857 VDD.n2214 GND 0.04999f
C10858 VDD.t449 GND 0.63568f
C10859 VDD.n2215 GND 0.05074f
C10860 VDD.n2216 GND 0.05074f
C10861 VDD.n2217 GND 0.02967f
C10862 VDD.n2218 GND 0.02522f
C10863 VDD.t450 GND 0.02334f
C10864 VDD.t723 GND 0.02334f
C10865 VDD.n2219 GND 0.13232f
C10866 VDD.n2220 GND 0.06172f
C10867 VDD.n2222 GND 0.0536f
C10868 VDD.n2223 GND 0.05074f
C10869 VDD.n2224 GND 0.02967f
C10870 VDD.n2225 GND 0.02522f
C10871 VDD.n2226 GND 0.04999f
C10872 VDD.t133 GND 0.63568f
C10873 VDD.n2227 GND 0.05074f
C10874 VDD.n2228 GND 0.05074f
C10875 VDD.n2229 GND 0.02967f
C10876 VDD.n2230 GND 0.02522f
C10877 VDD.n2231 GND 0.0536f
C10878 VDD.n2232 GND 0.05074f
C10879 VDD.n2233 GND 0.09652f
C10880 VDD.t300 GND 0.02321f
C10881 VDD.t255 GND 0.02321f
C10882 VDD.n2234 GND 0.10855f
C10883 VDD.t134 GND 0.02321f
C10884 VDD.t96 GND 0.02321f
C10885 VDD.n2235 GND 0.10855f
C10886 VDD.n2236 GND 0.0536f
C10887 VDD.n2237 GND 0.05074f
C10888 VDD.n2238 GND 0.0536f
C10889 VDD.n2239 GND 0.04999f
C10890 VDD.n2240 GND 0.04999f
C10891 VDD.n2241 GND 0.05074f
C10892 VDD.n2242 GND 0.02967f
C10893 VDD.n2243 GND 0.02522f
C10894 VDD.n2244 GND 0.04999f
C10895 VDD.n2245 GND 0.02522f
C10896 VDD.n2246 GND 0.04999f
C10897 VDD.n2247 GND 0.5126f
C10898 VDD.n2248 GND 0.5126f
C10899 VDD.n2249 GND 0.02522f
C10900 VDD.n2250 GND 0.02522f
C10901 VDD.n2251 GND 0.02967f
C10902 VDD.n2252 GND 0.05074f
C10903 VDD.t1082 GND 0.63568f
C10904 VDD.n2253 GND 0.05074f
C10905 VDD.n2254 GND 0.05074f
C10906 VDD.n2255 GND 0.09132f
C10907 VDD.n2256 GND 0.04999f
C10908 VDD.t97 GND 0.63568f
C10909 VDD.n2257 GND 0.05074f
C10910 VDD.n2258 GND 0.05074f
C10911 VDD.n2259 GND 0.02967f
C10912 VDD.n2260 GND 0.02522f
C10913 VDD.t1083 GND 0.02334f
C10914 VDD.n2261 GND 0.0731f
C10915 VDD.n2262 GND 0.01798f
C10916 VDD.n2263 GND 0.02334f
C10917 VDD.n2264 GND 0.0536f
C10918 VDD.n2265 GND 0.05074f
C10919 VDD.n2266 GND 0.02967f
C10920 VDD.n2267 GND 0.02522f
C10921 VDD.n2268 GND 0.04999f
C10922 VDD.t143 GND 0.63568f
C10923 VDD.n2269 GND 0.05074f
C10924 VDD.n2270 GND 0.05074f
C10925 VDD.n2271 GND 0.02967f
C10926 VDD.n2272 GND 0.02522f
C10927 VDD.t98 GND 0.02321f
C10928 VDD.t144 GND 0.02321f
C10929 VDD.n2273 GND 0.10855f
C10930 VDD.t776 GND 0.02321f
C10931 VDD.t933 GND 0.02321f
C10932 VDD.n2274 GND 0.10855f
C10933 VDD.n2275 GND 0.04152f
C10934 VDD.n2276 GND 0.02334f
C10935 VDD.n2277 GND 0.0536f
C10936 VDD.n2278 GND 0.05074f
C10937 VDD.n2279 GND 0.02967f
C10938 VDD.n2280 GND 0.02522f
C10939 VDD.n2281 GND 0.04999f
C10940 VDD.t473 GND 0.63568f
C10941 VDD.n2282 GND 0.05074f
C10942 VDD.n2283 GND 0.05074f
C10943 VDD.n2284 GND 0.02967f
C10944 VDD.n2285 GND 0.02522f
C10945 VDD.t474 GND 0.02334f
C10946 VDD.t751 GND 0.02334f
C10947 VDD.n2286 GND 0.13341f
C10948 VDD.n2287 GND 0.0263f
C10949 VDD.n2288 GND 0.0536f
C10950 VDD.n2289 GND 0.05074f
C10951 VDD.n2290 GND 0.02967f
C10952 VDD.n2291 GND 0.02522f
C10953 VDD.n2292 GND 0.04999f
C10954 VDD.t541 GND 0.63568f
C10955 VDD.n2293 GND 0.05074f
C10956 VDD.n2294 GND 0.05074f
C10957 VDD.n2295 GND 0.02967f
C10958 VDD.n2296 GND 0.02522f
C10959 VDD.n2297 GND 0.03166f
C10960 VDD.n2298 GND 0.0536f
C10961 VDD.n2299 GND 0.05074f
C10962 VDD.n2300 GND 0.02967f
C10963 VDD.n2301 GND 0.02522f
C10964 VDD.n2302 GND 0.04999f
C10965 VDD.t788 GND 0.63568f
C10966 VDD.n2303 GND 0.05074f
C10967 VDD.n2304 GND 0.05074f
C10968 VDD.n2305 GND 0.02967f
C10969 VDD.n2306 GND 0.02522f
C10970 VDD.t542 GND 0.02321f
C10971 VDD.t897 GND 0.02321f
C10972 VDD.n2307 GND 0.10855f
C10973 VDD.t870 GND 0.02321f
C10974 VDD.t789 GND 0.02321f
C10975 VDD.n2308 GND 0.10855f
C10976 VDD.n2309 GND 0.04152f
C10977 VDD.t26 GND 0.02334f
C10978 VDD.n2310 GND 0.02746f
C10979 VDD.n2311 GND 0.05074f
C10980 VDD.n2312 GND 0.02967f
C10981 VDD.n2313 GND 0.05074f
C10982 VDD.n2314 GND 0.62973f
C10983 VDD.t25 GND 0.74438f
C10984 VDD.n2316 GND 0.04999f
C10985 VDD.t508 GND 0.63568f
C10986 VDD.n2317 GND 0.05074f
C10987 VDD.n2318 GND 0.05074f
C10988 VDD.n2319 GND 0.02967f
C10989 VDD.n2320 GND 0.02522f
C10990 VDD.t697 GND 0.02334f
C10991 VDD.t509 GND 0.02334f
C10992 VDD.n2321 GND 0.13341f
C10993 VDD.n2322 GND 0.0263f
C10994 VDD.n2323 GND 0.0536f
C10995 VDD.n2324 GND 0.05074f
C10996 VDD.n2325 GND 0.02967f
C10997 VDD.n2326 GND 0.02522f
C10998 VDD.n2327 GND 0.04999f
C10999 VDD.t858 GND 0.63568f
C11000 VDD.n2328 GND 0.05074f
C11001 VDD.n2329 GND 0.05074f
C11002 VDD.n2330 GND 0.02967f
C11003 VDD.n2331 GND 0.02522f
C11004 VDD.n2332 GND 0.03166f
C11005 VDD.n2333 GND 0.0536f
C11006 VDD.n2334 GND 0.05074f
C11007 VDD.n2335 GND 0.02967f
C11008 VDD.n2336 GND 0.02522f
C11009 VDD.n2337 GND 0.04999f
C11010 VDD.t1050 GND 0.63568f
C11011 VDD.n2338 GND 0.05074f
C11012 VDD.n2339 GND 0.05074f
C11013 VDD.n2340 GND 0.02967f
C11014 VDD.n2341 GND 0.02522f
C11015 VDD.t937 GND 0.02321f
C11016 VDD.t1051 GND 0.02321f
C11017 VDD.n2342 GND 0.10855f
C11018 VDD.t859 GND 0.02321f
C11019 VDD.t1094 GND 0.02321f
C11020 VDD.n2343 GND 0.10855f
C11021 VDD.n2344 GND 0.04152f
C11022 VDD.n2345 GND 0.02334f
C11023 VDD.n2346 GND 0.0536f
C11024 VDD.n2347 GND 0.05074f
C11025 VDD.n2348 GND 0.02967f
C11026 VDD.n2349 GND 0.02522f
C11027 VDD.n2350 GND 0.04999f
C11028 VDD.t518 GND 0.63568f
C11029 VDD.n2351 GND 0.05074f
C11030 VDD.n2352 GND 0.05074f
C11031 VDD.n2353 GND 0.02967f
C11032 VDD.n2354 GND 0.02522f
C11033 VDD.t519 GND 0.02334f
C11034 VDD.t689 GND 0.02334f
C11035 VDD.n2355 GND 0.13232f
C11036 VDD.n2356 GND 0.06172f
C11037 VDD.n2358 GND 0.0536f
C11038 VDD.n2359 GND 0.05074f
C11039 VDD.n2360 GND 0.02967f
C11040 VDD.n2361 GND 0.02522f
C11041 VDD.n2362 GND 0.04999f
C11042 VDD.t266 GND 0.63568f
C11043 VDD.n2363 GND 0.05074f
C11044 VDD.n2364 GND 0.05074f
C11045 VDD.n2365 GND 0.02967f
C11046 VDD.n2366 GND 0.02522f
C11047 VDD.n2367 GND 0.0536f
C11048 VDD.n2368 GND 0.05074f
C11049 VDD.n2369 GND 0.09652f
C11050 VDD.t582 GND 0.02321f
C11051 VDD.t219 GND 0.02321f
C11052 VDD.n2370 GND 0.10855f
C11053 VDD.t267 GND 0.02321f
C11054 VDD.t216 GND 0.02321f
C11055 VDD.n2371 GND 0.10855f
C11056 VDD.n2372 GND 0.0536f
C11057 VDD.n2373 GND 0.05074f
C11058 VDD.n2374 GND 0.0536f
C11059 VDD.n2375 GND 0.04999f
C11060 VDD.n2376 GND 0.04999f
C11061 VDD.n2377 GND 0.05074f
C11062 VDD.n2378 GND 0.02967f
C11063 VDD.n2379 GND 0.02522f
C11064 VDD.n2380 GND 0.04999f
C11065 VDD.n2381 GND 0.02522f
C11066 VDD.n2382 GND 0.04999f
C11067 VDD.n2383 GND 0.5126f
C11068 VDD.n2384 GND 0.5126f
C11069 VDD.n2385 GND 0.02522f
C11070 VDD.n2386 GND 0.02522f
C11071 VDD.n2387 GND 0.02967f
C11072 VDD.n2388 GND 0.05074f
C11073 VDD.t1010 GND 0.63568f
C11074 VDD.n2389 GND 0.05074f
C11075 VDD.n2390 GND 0.05074f
C11076 VDD.n2391 GND 0.09132f
C11077 VDD.n2392 GND 0.04999f
C11078 VDD.t217 GND 0.63568f
C11079 VDD.n2393 GND 0.05074f
C11080 VDD.n2394 GND 0.05074f
C11081 VDD.n2395 GND 0.02967f
C11082 VDD.n2396 GND 0.02522f
C11083 VDD.t1011 GND 0.02334f
C11084 VDD.n2397 GND 0.0731f
C11085 VDD.n2398 GND 0.01798f
C11086 VDD.n2399 GND 0.02334f
C11087 VDD.n2400 GND 0.0536f
C11088 VDD.n2401 GND 0.05074f
C11089 VDD.n2402 GND 0.02967f
C11090 VDD.n2403 GND 0.02522f
C11091 VDD.n2404 GND 0.04999f
C11092 VDD.t91 GND 0.63568f
C11093 VDD.n2405 GND 0.05074f
C11094 VDD.n2406 GND 0.05074f
C11095 VDD.n2407 GND 0.02967f
C11096 VDD.n2408 GND 0.02522f
C11097 VDD.t218 GND 0.02321f
C11098 VDD.t92 GND 0.02321f
C11099 VDD.n2409 GND 0.10855f
C11100 VDD.t589 GND 0.02321f
C11101 VDD.t616 GND 0.02321f
C11102 VDD.n2410 GND 0.10855f
C11103 VDD.n2411 GND 0.04152f
C11104 VDD.n2412 GND 0.02334f
C11105 VDD.n2413 GND 0.0536f
C11106 VDD.n2414 GND 0.05074f
C11107 VDD.n2415 GND 0.02967f
C11108 VDD.n2416 GND 0.02522f
C11109 VDD.n2417 GND 0.04999f
C11110 VDD.t532 GND 0.63568f
C11111 VDD.n2418 GND 0.05074f
C11112 VDD.n2419 GND 0.05074f
C11113 VDD.n2420 GND 0.02967f
C11114 VDD.n2421 GND 0.02522f
C11115 VDD.t533 GND 0.02334f
C11116 VDD.t703 GND 0.02334f
C11117 VDD.n2422 GND 0.13341f
C11118 VDD.n2423 GND 0.0263f
C11119 VDD.n2424 GND 0.0536f
C11120 VDD.n2425 GND 0.05074f
C11121 VDD.n2426 GND 0.02967f
C11122 VDD.n2427 GND 0.02522f
C11123 VDD.n2428 GND 0.04999f
C11124 VDD.t160 GND 0.63568f
C11125 VDD.n2429 GND 0.05074f
C11126 VDD.n2430 GND 0.05074f
C11127 VDD.n2431 GND 0.02967f
C11128 VDD.n2432 GND 0.02522f
C11129 VDD.n2433 GND 0.03166f
C11130 VDD.n2434 GND 0.0536f
C11131 VDD.n2435 GND 0.05074f
C11132 VDD.n2436 GND 0.02967f
C11133 VDD.n2437 GND 0.02522f
C11134 VDD.n2438 GND 0.04999f
C11135 VDD.t590 GND 0.63568f
C11136 VDD.n2439 GND 0.05074f
C11137 VDD.n2440 GND 0.05074f
C11138 VDD.n2441 GND 0.02967f
C11139 VDD.n2442 GND 0.02522f
C11140 VDD.t161 GND 0.02321f
C11141 VDD.t591 GND 0.02321f
C11142 VDD.n2443 GND 0.10855f
C11143 VDD.t899 GND 0.02321f
C11144 VDD.t802 GND 0.02321f
C11145 VDD.n2444 GND 0.10855f
C11146 VDD.n2445 GND 0.04152f
C11147 VDD.t797 GND 0.02334f
C11148 VDD.n2446 GND 0.02746f
C11149 VDD.n2447 GND 0.05074f
C11150 VDD.n2448 GND 0.02967f
C11151 VDD.n2449 GND 0.05074f
C11152 VDD.n2450 GND 0.62973f
C11153 VDD.t796 GND 0.74438f
C11154 VDD.n2452 GND 0.04999f
C11155 VDD.t504 GND 0.63568f
C11156 VDD.n2453 GND 0.05074f
C11157 VDD.n2454 GND 0.05074f
C11158 VDD.n2455 GND 0.02967f
C11159 VDD.n2456 GND 0.02522f
C11160 VDD.t691 GND 0.02334f
C11161 VDD.t505 GND 0.02334f
C11162 VDD.n2457 GND 0.13341f
C11163 VDD.n2458 GND 0.0263f
C11164 VDD.n2459 GND 0.0536f
C11165 VDD.n2460 GND 0.05074f
C11166 VDD.n2461 GND 0.02967f
C11167 VDD.n2462 GND 0.02522f
C11168 VDD.n2463 GND 0.04999f
C11169 VDD.t800 GND 0.63568f
C11170 VDD.n2464 GND 0.05074f
C11171 VDD.n2465 GND 0.05074f
C11172 VDD.n2466 GND 0.02967f
C11173 VDD.n2467 GND 0.02522f
C11174 VDD.n2468 GND 0.03166f
C11175 VDD.n2469 GND 0.0536f
C11176 VDD.n2470 GND 0.05074f
C11177 VDD.n2471 GND 0.02967f
C11178 VDD.n2472 GND 0.02522f
C11179 VDD.n2473 GND 0.04999f
C11180 VDD.t1048 GND 0.63568f
C11181 VDD.n2474 GND 0.05074f
C11182 VDD.n2475 GND 0.05074f
C11183 VDD.n2476 GND 0.02967f
C11184 VDD.n2477 GND 0.02522f
C11185 VDD.t801 GND 0.02321f
C11186 VDD.t1100 GND 0.02321f
C11187 VDD.n2478 GND 0.10855f
C11188 VDD.t876 GND 0.02321f
C11189 VDD.t1049 GND 0.02321f
C11190 VDD.n2479 GND 0.10855f
C11191 VDD.n2480 GND 0.04152f
C11192 VDD.n2481 GND 0.02334f
C11193 VDD.n2482 GND 0.0536f
C11194 VDD.n2483 GND 0.05074f
C11195 VDD.n2484 GND 0.02967f
C11196 VDD.n2485 GND 0.02522f
C11197 VDD.n2486 GND 0.04999f
C11198 VDD.t441 GND 0.63568f
C11199 VDD.n2487 GND 0.05074f
C11200 VDD.n2488 GND 0.05074f
C11201 VDD.n2489 GND 0.02967f
C11202 VDD.n2490 GND 0.02522f
C11203 VDD.t442 GND 0.02334f
C11204 VDD.t715 GND 0.02334f
C11205 VDD.n2491 GND 0.13232f
C11206 VDD.n2492 GND 0.06172f
C11207 VDD.n2494 GND 0.0536f
C11208 VDD.n2495 GND 0.05074f
C11209 VDD.n2496 GND 0.02967f
C11210 VDD.n2497 GND 0.02522f
C11211 VDD.n2498 GND 0.04999f
C11212 VDD.t328 GND 0.63568f
C11213 VDD.n2499 GND 0.05074f
C11214 VDD.n2500 GND 0.05074f
C11215 VDD.n2501 GND 0.02967f
C11216 VDD.n2502 GND 0.02522f
C11217 VDD.n2503 GND 0.0536f
C11218 VDD.n2504 GND 0.05074f
C11219 VDD.n2505 GND 0.09652f
C11220 VDD.t329 GND 0.02321f
C11221 VDD.t20 GND 0.02321f
C11222 VDD.n2506 GND 0.10855f
C11223 VDD.t1102 GND 0.02321f
C11224 VDD.t592 GND 0.02321f
C11225 VDD.n2507 GND 0.10855f
C11226 VDD.n2508 GND 0.0536f
C11227 VDD.n2509 GND 0.05074f
C11228 VDD.n2510 GND 0.0536f
C11229 VDD.n2511 GND 0.04999f
C11230 VDD.n2512 GND 0.04999f
C11231 VDD.n2513 GND 0.05074f
C11232 VDD.n2514 GND 0.02967f
C11233 VDD.n2515 GND 0.02522f
C11234 VDD.n2516 GND 0.04999f
C11235 VDD.n2517 GND 0.02522f
C11236 VDD.n2518 GND 0.04999f
C11237 VDD.n2519 GND 0.5126f
C11238 VDD.n2520 GND 0.5126f
C11239 VDD.n2521 GND 0.02522f
C11240 VDD.n2522 GND 0.02522f
C11241 VDD.n2523 GND 0.02967f
C11242 VDD.n2524 GND 0.05074f
C11243 VDD.t1038 GND 0.63568f
C11244 VDD.n2525 GND 0.05074f
C11245 VDD.n2526 GND 0.05074f
C11246 VDD.n2527 GND 0.09132f
C11247 VDD.n2528 GND 0.04999f
C11248 VDD.t593 GND 0.63568f
C11249 VDD.n2529 GND 0.05074f
C11250 VDD.n2530 GND 0.05074f
C11251 VDD.n2531 GND 0.02967f
C11252 VDD.n2532 GND 0.02522f
C11253 VDD.t1039 GND 0.02334f
C11254 VDD.n2533 GND 0.0731f
C11255 VDD.n2534 GND 0.01798f
C11256 VDD.n2535 GND 0.02334f
C11257 VDD.n2536 GND 0.0536f
C11258 VDD.n2537 GND 0.05074f
C11259 VDD.n2538 GND 0.02967f
C11260 VDD.n2539 GND 0.02522f
C11261 VDD.n2540 GND 0.04999f
C11262 VDD.t199 GND 0.63568f
C11263 VDD.n2541 GND 0.05074f
C11264 VDD.n2542 GND 0.05074f
C11265 VDD.n2543 GND 0.02967f
C11266 VDD.n2544 GND 0.02522f
C11267 VDD.t594 GND 0.02321f
C11268 VDD.t767 GND 0.02321f
C11269 VDD.n2545 GND 0.10855f
C11270 VDD.t905 GND 0.02321f
C11271 VDD.t200 GND 0.02321f
C11272 VDD.n2546 GND 0.10855f
C11273 VDD.n2547 GND 0.04152f
C11274 VDD.n2548 GND 0.02334f
C11275 VDD.n2549 GND 0.0536f
C11276 VDD.n2550 GND 0.05074f
C11277 VDD.n2551 GND 0.02967f
C11278 VDD.n2552 GND 0.02522f
C11279 VDD.n2553 GND 0.04999f
C11280 VDD.t451 GND 0.63568f
C11281 VDD.n2554 GND 0.05074f
C11282 VDD.n2555 GND 0.05074f
C11283 VDD.n2556 GND 0.02967f
C11284 VDD.n2557 GND 0.02522f
C11285 VDD.t452 GND 0.02334f
C11286 VDD.t731 GND 0.02334f
C11287 VDD.n2558 GND 0.13341f
C11288 VDD.n2559 GND 0.0263f
C11289 VDD.n2560 GND 0.0536f
C11290 VDD.n2561 GND 0.05074f
C11291 VDD.n2562 GND 0.02967f
C11292 VDD.n2563 GND 0.02522f
C11293 VDD.n2564 GND 0.04999f
C11294 VDD.t39 GND 0.63568f
C11295 VDD.n2565 GND 0.05074f
C11296 VDD.n2566 GND 0.05074f
C11297 VDD.n2567 GND 0.02967f
C11298 VDD.n2568 GND 0.02522f
C11299 VDD.n2569 GND 0.03166f
C11300 VDD.n2570 GND 0.0536f
C11301 VDD.n2571 GND 0.05074f
C11302 VDD.n2572 GND 0.02967f
C11303 VDD.n2573 GND 0.02522f
C11304 VDD.n2574 GND 0.04999f
C11305 VDD.t69 GND 0.63568f
C11306 VDD.n2575 GND 0.05074f
C11307 VDD.n2576 GND 0.05074f
C11308 VDD.n2577 GND 0.02967f
C11309 VDD.n2578 GND 0.02522f
C11310 VDD.t628 GND 0.02321f
C11311 VDD.t375 GND 0.02321f
C11312 VDD.n2579 GND 0.10855f
C11313 VDD.t40 GND 0.02321f
C11314 VDD.t70 GND 0.02321f
C11315 VDD.n2580 GND 0.10855f
C11316 VDD.n2581 GND 0.04152f
C11317 VDD.t765 GND 0.02334f
C11318 VDD.n2582 GND 0.02746f
C11319 VDD.n2583 GND 0.05074f
C11320 VDD.n2584 GND 0.02967f
C11321 VDD.n2585 GND 0.05074f
C11322 VDD.n2586 GND 0.62973f
C11323 VDD.t764 GND 0.74438f
C11324 VDD.n2588 GND 0.04999f
C11325 VDD.t536 GND 0.63568f
C11326 VDD.n2589 GND 0.05074f
C11327 VDD.n2590 GND 0.05074f
C11328 VDD.n2591 GND 0.02967f
C11329 VDD.n2592 GND 0.02522f
C11330 VDD.t717 GND 0.02334f
C11331 VDD.t537 GND 0.02334f
C11332 VDD.n2593 GND 0.13341f
C11333 VDD.n2594 GND 0.0263f
C11334 VDD.n2595 GND 0.0536f
C11335 VDD.n2596 GND 0.05074f
C11336 VDD.n2597 GND 0.02967f
C11337 VDD.n2598 GND 0.02522f
C11338 VDD.n2599 GND 0.04999f
C11339 VDD.t67 GND 0.63568f
C11340 VDD.n2600 GND 0.05074f
C11341 VDD.n2601 GND 0.05074f
C11342 VDD.n2602 GND 0.02967f
C11343 VDD.n2603 GND 0.02522f
C11344 VDD.n2604 GND 0.03166f
C11345 VDD.n2605 GND 0.0536f
C11346 VDD.n2606 GND 0.05074f
C11347 VDD.n2607 GND 0.02967f
C11348 VDD.n2608 GND 0.02522f
C11349 VDD.n2609 GND 0.04999f
C11350 VDD.t1022 GND 0.63568f
C11351 VDD.n2610 GND 0.05074f
C11352 VDD.n2611 GND 0.05074f
C11353 VDD.n2612 GND 0.02967f
C11354 VDD.n2613 GND 0.02522f
C11355 VDD.t68 GND 0.02321f
C11356 VDD.t1023 GND 0.02321f
C11357 VDD.n2614 GND 0.10855f
C11358 VDD.t586 GND 0.02321f
C11359 VDD.t1071 GND 0.02321f
C11360 VDD.n2615 GND 0.10855f
C11361 VDD.n2616 GND 0.04152f
C11362 VDD.n2617 GND 0.02334f
C11363 VDD.n2618 GND 0.0536f
C11364 VDD.n2619 GND 0.05074f
C11365 VDD.n2620 GND 0.02967f
C11366 VDD.n2621 GND 0.02522f
C11367 VDD.n2622 GND 0.04999f
C11368 VDD.t488 GND 0.63568f
C11369 VDD.n2623 GND 0.05074f
C11370 VDD.n2624 GND 0.05074f
C11371 VDD.n2625 GND 0.02967f
C11372 VDD.n2626 GND 0.02522f
C11373 VDD.t489 GND 0.02334f
C11374 VDD.t669 GND 0.02334f
C11375 VDD.n2627 GND 0.13232f
C11376 VDD.n2628 GND 0.06172f
C11377 VDD.n2630 GND 0.0536f
C11378 VDD.n2631 GND 0.05074f
C11379 VDD.n2632 GND 0.02967f
C11380 VDD.n2633 GND 0.02522f
C11381 VDD.n2634 GND 0.04999f
C11382 VDD.t31 GND 0.63568f
C11383 VDD.n2635 GND 0.05074f
C11384 VDD.n2636 GND 0.05074f
C11385 VDD.n2637 GND 0.02967f
C11386 VDD.n2638 GND 0.02522f
C11387 VDD.n2639 GND 0.0536f
C11388 VDD.n2640 GND 0.05074f
C11389 VDD.n2641 GND 0.09652f
C11390 VDD.t32 GND 0.02321f
C11391 VDD.t617 GND 0.02321f
C11392 VDD.n2642 GND 0.10855f
C11393 VDD.t894 GND 0.02321f
C11394 VDD.t387 GND 0.02321f
C11395 VDD.n2643 GND 0.10855f
C11396 VDD.n2644 GND 0.0536f
C11397 VDD.n2645 GND 0.05074f
C11398 VDD.n2646 GND 0.0536f
C11399 VDD.n2647 GND 0.04999f
C11400 VDD.n2648 GND 0.04999f
C11401 VDD.n2649 GND 0.05074f
C11402 VDD.n2650 GND 0.02967f
C11403 VDD.n2651 GND 0.02522f
C11404 VDD.n2652 GND 0.04999f
C11405 VDD.n2653 GND 0.02522f
C11406 VDD.n2654 GND 0.04999f
C11407 VDD.n2655 GND 0.5126f
C11408 VDD.n2656 GND 0.5126f
C11409 VDD.n2657 GND 0.02522f
C11410 VDD.n2658 GND 0.02522f
C11411 VDD.n2659 GND 0.02967f
C11412 VDD.n2660 GND 0.05074f
C11413 VDD.t1062 GND 0.63568f
C11414 VDD.n2661 GND 0.05074f
C11415 VDD.n2662 GND 0.05074f
C11416 VDD.n2663 GND 0.09132f
C11417 VDD.n2664 GND 0.04999f
C11418 VDD.t388 GND 0.63568f
C11419 VDD.n2665 GND 0.05074f
C11420 VDD.n2666 GND 0.05074f
C11421 VDD.n2667 GND 0.02967f
C11422 VDD.n2668 GND 0.02522f
C11423 VDD.t1063 GND 0.02334f
C11424 VDD.n2669 GND 0.0731f
C11425 VDD.n2670 GND 0.01798f
C11426 VDD.n2671 GND 0.02334f
C11427 VDD.n2672 GND 0.0536f
C11428 VDD.n2673 GND 0.05074f
C11429 VDD.n2674 GND 0.02967f
C11430 VDD.n2675 GND 0.02522f
C11431 VDD.n2676 GND 0.04999f
C11432 VDD.t344 GND 0.63568f
C11433 VDD.n2677 GND 0.05074f
C11434 VDD.n2678 GND 0.05074f
C11435 VDD.n2679 GND 0.02967f
C11436 VDD.n2680 GND 0.02522f
C11437 VDD.t389 GND 0.02321f
C11438 VDD.t345 GND 0.02321f
C11439 VDD.n2681 GND 0.10855f
C11440 VDD.t618 GND 0.02321f
C11441 VDD.t1103 GND 0.02321f
C11442 VDD.n2682 GND 0.10855f
C11443 VDD.n2683 GND 0.04152f
C11444 VDD.n2684 GND 0.02334f
C11445 VDD.n2685 GND 0.0536f
C11446 VDD.n2686 GND 0.05074f
C11447 VDD.n2687 GND 0.02967f
C11448 VDD.n2688 GND 0.02522f
C11449 VDD.n2689 GND 0.04999f
C11450 VDD.t469 GND 0.63568f
C11451 VDD.n2690 GND 0.05074f
C11452 VDD.n2691 GND 0.05074f
C11453 VDD.n2692 GND 0.02967f
C11454 VDD.n2693 GND 0.02522f
C11455 VDD.t470 GND 0.02334f
C11456 VDD.t747 GND 0.02334f
C11457 VDD.n2694 GND 0.13341f
C11458 VDD.n2695 GND 0.0263f
C11459 VDD.n2696 GND 0.0536f
C11460 VDD.n2697 GND 0.05074f
C11461 VDD.n2698 GND 0.02967f
C11462 VDD.n2699 GND 0.02522f
C11463 VDD.n2700 GND 0.04999f
C11464 VDD.t892 GND 0.63568f
C11465 VDD.n2701 GND 0.05074f
C11466 VDD.n2702 GND 0.05074f
C11467 VDD.n2703 GND 0.02967f
C11468 VDD.n2704 GND 0.02522f
C11469 VDD.n2705 GND 0.03166f
C11470 VDD.n2706 GND 0.0536f
C11471 VDD.n2707 GND 0.05074f
C11472 VDD.n2708 GND 0.02967f
C11473 VDD.n2709 GND 0.02522f
C11474 VDD.n2710 GND 0.04999f
C11475 VDD.t2 GND 0.63568f
C11476 VDD.n2711 GND 0.05074f
C11477 VDD.n2712 GND 0.05074f
C11478 VDD.n2713 GND 0.02967f
C11479 VDD.n2714 GND 0.02522f
C11480 VDD.t1101 GND 0.02321f
C11481 VDD.t900 GND 0.02321f
C11482 VDD.n2715 GND 0.10855f
C11483 VDD.t893 GND 0.02321f
C11484 VDD.t3 GND 0.02321f
C11485 VDD.n2716 GND 0.10855f
C11486 VDD.n2717 GND 0.04152f
C11487 VDD.t125 GND 0.02334f
C11488 VDD.n2718 GND 0.02746f
C11489 VDD.n2719 GND 0.05074f
C11490 VDD.n2720 GND 0.02967f
C11491 VDD.n2721 GND 0.05074f
C11492 VDD.n2722 GND 0.62973f
C11493 VDD.t124 GND 0.74438f
C11494 VDD.n2724 GND 0.04999f
C11495 VDD.t455 GND 0.63568f
C11496 VDD.n2725 GND 0.05074f
C11497 VDD.n2726 GND 0.05074f
C11498 VDD.n2727 GND 0.02967f
C11499 VDD.n2728 GND 0.02522f
C11500 VDD.t739 GND 0.02334f
C11501 VDD.t456 GND 0.02334f
C11502 VDD.n2729 GND 0.13341f
C11503 VDD.n2730 GND 0.0263f
C11504 VDD.n2731 GND 0.0536f
C11505 VDD.n2732 GND 0.05074f
C11506 VDD.n2733 GND 0.02967f
C11507 VDD.n2734 GND 0.02522f
C11508 VDD.n2735 GND 0.04999f
C11509 VDD.t0 GND 0.63568f
C11510 VDD.n2736 GND 0.05074f
C11511 VDD.n2737 GND 0.05074f
C11512 VDD.n2738 GND 0.02967f
C11513 VDD.n2739 GND 0.02522f
C11514 VDD.n2740 GND 0.03166f
C11515 VDD.n2741 GND 0.0536f
C11516 VDD.n2742 GND 0.05074f
C11517 VDD.n2743 GND 0.02967f
C11518 VDD.n2744 GND 0.02522f
C11519 VDD.n2745 GND 0.04999f
C11520 VDD.t1018 GND 0.63568f
C11521 VDD.n2746 GND 0.05074f
C11522 VDD.n2747 GND 0.05074f
C11523 VDD.n2748 GND 0.02967f
C11524 VDD.n2749 GND 0.02522f
C11525 VDD.t1 GND 0.02321f
C11526 VDD.t1087 GND 0.02321f
C11527 VDD.n2750 GND 0.10855f
C11528 VDD.t230 GND 0.02321f
C11529 VDD.t1019 GND 0.02321f
C11530 VDD.n2751 GND 0.10855f
C11531 VDD.n2752 GND 0.04152f
C11532 VDD.n2753 GND 0.02334f
C11533 VDD.n2754 GND 0.0536f
C11534 VDD.n2755 GND 0.05074f
C11535 VDD.n2756 GND 0.02967f
C11536 VDD.n2757 GND 0.02522f
C11537 VDD.n2758 GND 0.04999f
C11538 VDD.t514 GND 0.63568f
C11539 VDD.n2759 GND 0.05074f
C11540 VDD.n2760 GND 0.05074f
C11541 VDD.n2761 GND 0.02967f
C11542 VDD.n2762 GND 0.02522f
C11543 VDD.t515 GND 0.02334f
C11544 VDD.t683 GND 0.02334f
C11545 VDD.n2763 GND 0.13232f
C11546 VDD.n2764 GND 0.06172f
C11547 VDD.n2766 GND 0.0536f
C11548 VDD.n2767 GND 0.05074f
C11549 VDD.n2768 GND 0.02967f
C11550 VDD.n2769 GND 0.02522f
C11551 VDD.n2770 GND 0.04999f
C11552 VDD.t373 GND 0.63568f
C11553 VDD.n2771 GND 0.05074f
C11554 VDD.n2772 GND 0.05074f
C11555 VDD.n2773 GND 0.02967f
C11556 VDD.n2774 GND 0.02522f
C11557 VDD.n2775 GND 0.0536f
C11558 VDD.n2776 GND 0.05074f
C11559 VDD.n2777 GND 0.09652f
C11560 VDD.t374 GND 0.02321f
C11561 VDD.t201 GND 0.02321f
C11562 VDD.n2778 GND 0.10855f
C11563 VDD.t611 GND 0.02321f
C11564 VDD.t81 GND 0.02321f
C11565 VDD.n2779 GND 0.10855f
C11566 VDD.n2780 GND 0.0536f
C11567 VDD.n2781 GND 0.05074f
C11568 VDD.n2782 GND 0.0536f
C11569 VDD.n2783 GND 0.04999f
C11570 VDD.n2784 GND 0.04999f
C11571 VDD.n2785 GND 0.05074f
C11572 VDD.n2786 GND 0.02967f
C11573 VDD.n2787 GND 0.02522f
C11574 VDD.n2788 GND 0.04999f
C11575 VDD.n2789 GND 0.02522f
C11576 VDD.n2790 GND 0.04999f
C11577 VDD.n2791 GND 0.5126f
C11578 VDD.n2792 GND 0.5126f
C11579 VDD.n2793 GND 0.02522f
C11580 VDD.n2794 GND 0.02522f
C11581 VDD.n2795 GND 0.02967f
C11582 VDD.n2796 GND 0.05074f
C11583 VDD.t1006 GND 0.63568f
C11584 VDD.n2797 GND 0.05074f
C11585 VDD.n2798 GND 0.05074f
C11586 VDD.n2799 GND 0.09132f
C11587 VDD.n2800 GND 0.04999f
C11588 VDD.t82 GND 0.63568f
C11589 VDD.n2801 GND 0.05074f
C11590 VDD.n2802 GND 0.05074f
C11591 VDD.n2803 GND 0.02967f
C11592 VDD.n2804 GND 0.02522f
C11593 VDD.t1007 GND 0.02334f
C11594 VDD.n2805 GND 0.0731f
C11595 VDD.n2806 GND 0.01798f
C11596 VDD.n2807 GND 0.02334f
C11597 VDD.n2808 GND 0.0536f
C11598 VDD.n2809 GND 0.05074f
C11599 VDD.n2810 GND 0.02967f
C11600 VDD.n2811 GND 0.02522f
C11601 VDD.n2812 GND 0.04999f
C11602 VDD.t168 GND 0.63568f
C11603 VDD.n2813 GND 0.05074f
C11604 VDD.n2814 GND 0.05074f
C11605 VDD.n2815 GND 0.02967f
C11606 VDD.n2816 GND 0.02522f
C11607 VDD.t83 GND 0.02321f
C11608 VDD.t169 GND 0.02321f
C11609 VDD.n2817 GND 0.10855f
C11610 VDD.t588 GND 0.02321f
C11611 VDD.t326 GND 0.02321f
C11612 VDD.n2818 GND 0.10855f
C11613 VDD.n2819 GND 0.04152f
C11614 VDD.n2820 GND 0.02334f
C11615 VDD.n2821 GND 0.0536f
C11616 VDD.n2822 GND 0.05074f
C11617 VDD.n2823 GND 0.02967f
C11618 VDD.n2824 GND 0.02522f
C11619 VDD.n2825 GND 0.04999f
C11620 VDD.t524 GND 0.63568f
C11621 VDD.n2826 GND 0.05074f
C11622 VDD.n2827 GND 0.05074f
C11623 VDD.n2828 GND 0.02967f
C11624 VDD.n2829 GND 0.02522f
C11625 VDD.t525 GND 0.02334f
C11626 VDD.t699 GND 0.02334f
C11627 VDD.n2830 GND 0.13341f
C11628 VDD.n2831 GND 0.0263f
C11629 VDD.n2832 GND 0.0536f
C11630 VDD.n2833 GND 0.05074f
C11631 VDD.n2834 GND 0.02967f
C11632 VDD.n2835 GND 0.02522f
C11633 VDD.n2836 GND 0.04999f
C11634 VDD.t99 GND 0.63568f
C11635 VDD.n2837 GND 0.05074f
C11636 VDD.n2838 GND 0.05074f
C11637 VDD.n2839 GND 0.02967f
C11638 VDD.n2840 GND 0.02522f
C11639 VDD.n2841 GND 0.03166f
C11640 VDD.n2842 GND 0.0536f
C11641 VDD.n2843 GND 0.05074f
C11642 VDD.n2844 GND 0.02967f
C11643 VDD.n2845 GND 0.02522f
C11644 VDD.n2846 GND 0.04999f
C11645 VDD.t292 GND 0.63568f
C11646 VDD.n2847 GND 0.05074f
C11647 VDD.n2848 GND 0.05074f
C11648 VDD.n2849 GND 0.02967f
C11649 VDD.n2850 GND 0.02522f
C11650 VDD.t861 GND 0.02321f
C11651 VDD.t293 GND 0.02321f
C11652 VDD.n2851 GND 0.10855f
C11653 VDD.t100 GND 0.02321f
C11654 VDD.t953 GND 0.02321f
C11655 VDD.n2852 GND 0.10855f
C11656 VDD.n2853 GND 0.04152f
C11657 VDD.t154 GND 0.02334f
C11658 VDD.n2854 GND 0.02746f
C11659 VDD.n2855 GND 0.05074f
C11660 VDD.n2856 GND 0.02967f
C11661 VDD.n2857 GND 0.05074f
C11662 VDD.n2858 GND 0.62973f
C11663 VDD.t153 GND 0.74438f
C11664 VDD.n2860 GND 0.04999f
C11665 VDD.t502 GND 0.63568f
C11666 VDD.n2861 GND 0.05074f
C11667 VDD.n2862 GND 0.05074f
C11668 VDD.n2863 GND 0.02967f
C11669 VDD.n2864 GND 0.02522f
C11670 VDD.t687 GND 0.02334f
C11671 VDD.t503 GND 0.02334f
C11672 VDD.n2865 GND 0.13341f
C11673 VDD.n2866 GND 0.0263f
C11674 VDD.n2867 GND 0.0536f
C11675 VDD.n2868 GND 0.05074f
C11676 VDD.n2869 GND 0.02967f
C11677 VDD.n2870 GND 0.02522f
C11678 VDD.n2871 GND 0.04999f
C11679 VDD.t934 GND 0.63568f
C11680 VDD.n2872 GND 0.05074f
C11681 VDD.n2873 GND 0.05074f
C11682 VDD.n2874 GND 0.02967f
C11683 VDD.n2875 GND 0.02522f
C11684 VDD.n2876 GND 0.03166f
C11685 VDD.n2877 GND 0.0536f
C11686 VDD.n2878 GND 0.05074f
C11687 VDD.n2879 GND 0.02967f
C11688 VDD.n2880 GND 0.02522f
C11689 VDD.n2881 GND 0.04999f
C11690 VDD.t1045 GND 0.63568f
C11691 VDD.n2882 GND 0.05074f
C11692 VDD.n2883 GND 0.05074f
C11693 VDD.n2884 GND 0.02967f
C11694 VDD.n2885 GND 0.02522f
C11695 VDD.t952 GND 0.02321f
C11696 VDD.t1099 GND 0.02321f
C11697 VDD.n2886 GND 0.10855f
C11698 VDD.t935 GND 0.02321f
C11699 VDD.t1046 GND 0.02321f
C11700 VDD.n2887 GND 0.10855f
C11701 VDD.n2888 GND 0.04152f
C11702 VDD.n2889 GND 0.02334f
C11703 VDD.n2890 GND 0.0536f
C11704 VDD.n2891 GND 0.05074f
C11705 VDD.n2892 GND 0.02967f
C11706 VDD.n2893 GND 0.02522f
C11707 VDD.n2894 GND 0.04999f
C11708 VDD.t437 GND 0.63568f
C11709 VDD.n2895 GND 0.05074f
C11710 VDD.n2896 GND 0.05074f
C11711 VDD.n2897 GND 0.02967f
C11712 VDD.n2898 GND 0.02522f
C11713 VDD.t438 GND 0.02334f
C11714 VDD.t711 GND 0.02334f
C11715 VDD.n2899 GND 0.13232f
C11716 VDD.n2900 GND 0.06172f
C11717 VDD.n2902 GND 0.0536f
C11718 VDD.n2903 GND 0.05074f
C11719 VDD.n2904 GND 0.02967f
C11720 VDD.n2905 GND 0.02522f
C11721 VDD.n2906 GND 0.04999f
C11722 VDD.t821 GND 0.63568f
C11723 VDD.n2907 GND 0.05074f
C11724 VDD.n2908 GND 0.05074f
C11725 VDD.n2909 GND 0.02967f
C11726 VDD.n2910 GND 0.02522f
C11727 VDD.n2911 GND 0.0536f
C11728 VDD.n2912 GND 0.05074f
C11729 VDD.n2913 GND 0.09652f
C11730 VDD.t956 GND 0.02321f
C11731 VDD.t311 GND 0.02321f
C11732 VDD.n2914 GND 0.10855f
C11733 VDD.t822 GND 0.02321f
C11734 VDD.t1104 GND 0.02321f
C11735 VDD.n2915 GND 0.10855f
C11736 VDD.n2916 GND 0.0536f
C11737 VDD.n2917 GND 0.05074f
C11738 VDD.n2918 GND 0.0536f
C11739 VDD.n2919 GND 0.04999f
C11740 VDD.n2920 GND 0.04999f
C11741 VDD.n2921 GND 0.05074f
C11742 VDD.n2922 GND 0.02967f
C11743 VDD.n2923 GND 0.02522f
C11744 VDD.n2924 GND 0.04999f
C11745 VDD.n2925 GND 0.02522f
C11746 VDD.n2926 GND 0.04999f
C11747 VDD.n2927 GND 0.5126f
C11748 VDD.n2928 GND 0.5126f
C11749 VDD.n2929 GND 0.02522f
C11750 VDD.n2930 GND 0.02522f
C11751 VDD.n2931 GND 0.02967f
C11752 VDD.n2932 GND 0.05074f
C11753 VDD.t1034 GND 0.63568f
C11754 VDD.n2933 GND 0.05074f
C11755 VDD.n2934 GND 0.05074f
C11756 VDD.n2935 GND 0.09132f
C11757 VDD.n2936 GND 0.04999f
C11758 VDD.t308 GND 0.63568f
C11759 VDD.n2937 GND 0.05074f
C11760 VDD.n2938 GND 0.05074f
C11761 VDD.n2939 GND 0.02967f
C11762 VDD.n2940 GND 0.02522f
C11763 VDD.t1035 GND 0.02334f
C11764 VDD.n2941 GND 0.0731f
C11765 VDD.n2942 GND 0.01798f
C11766 VDD.n2943 GND 0.02334f
C11767 VDD.n2944 GND 0.0536f
C11768 VDD.n2945 GND 0.05074f
C11769 VDD.n2946 GND 0.02967f
C11770 VDD.n2947 GND 0.02522f
C11771 VDD.n2948 GND 0.04999f
C11772 VDD.t196 GND 0.63568f
C11773 VDD.n2949 GND 0.05074f
C11774 VDD.n2950 GND 0.05074f
C11775 VDD.n2951 GND 0.02967f
C11776 VDD.n2952 GND 0.02522f
C11777 VDD.t1105 GND 0.02321f
C11778 VDD.t198 GND 0.02321f
C11779 VDD.n2953 GND 0.10855f
C11780 VDD.t309 GND 0.02321f
C11781 VDD.t197 GND 0.02321f
C11782 VDD.n2954 GND 0.10855f
C11783 VDD.n2955 GND 0.04152f
C11784 VDD.n2956 GND 0.02334f
C11785 VDD.n2957 GND 0.0536f
C11786 VDD.n2958 GND 0.05074f
C11787 VDD.n2959 GND 0.02967f
C11788 VDD.n2960 GND 0.02522f
C11789 VDD.n2961 GND 0.04999f
C11790 VDD.t447 GND 0.63568f
C11791 VDD.n2962 GND 0.05074f
C11792 VDD.n2963 GND 0.05074f
C11793 VDD.n2964 GND 0.02967f
C11794 VDD.n2965 GND 0.02522f
C11795 VDD.t448 GND 0.02334f
C11796 VDD.t725 GND 0.02334f
C11797 VDD.n2966 GND 0.13341f
C11798 VDD.n2967 GND 0.0263f
C11799 VDD.n2968 GND 0.0536f
C11800 VDD.n2969 GND 0.05074f
C11801 VDD.n2970 GND 0.02967f
C11802 VDD.n2971 GND 0.02522f
C11803 VDD.n2972 GND 0.04999f
C11804 VDD.t296 GND 0.63568f
C11805 VDD.n2973 GND 0.05074f
C11806 VDD.n2974 GND 0.05074f
C11807 VDD.n2975 GND 0.02967f
C11808 VDD.n2976 GND 0.02522f
C11809 VDD.n2977 GND 0.03166f
C11810 VDD.n2978 GND 0.0536f
C11811 VDD.n2979 GND 0.05074f
C11812 VDD.n2980 GND 0.02967f
C11813 VDD.n2981 GND 0.02522f
C11814 VDD.n2982 GND 0.04999f
C11815 VDD.t626 GND 0.63568f
C11816 VDD.n2983 GND 0.05074f
C11817 VDD.n2984 GND 0.05074f
C11818 VDD.n2985 GND 0.02967f
C11819 VDD.n2986 GND 0.02522f
C11820 VDD.t297 GND 0.02321f
C11821 VDD.t627 GND 0.02321f
C11822 VDD.n2987 GND 0.10855f
C11823 VDD.t327 GND 0.02321f
C11824 VDD.t943 GND 0.02321f
C11825 VDD.n2988 GND 0.10855f
C11826 VDD.n2989 GND 0.04152f
C11827 VDD.t942 GND 0.02334f
C11828 VDD.n2990 GND 0.02746f
C11829 VDD.n2991 GND 0.05074f
C11830 VDD.n2992 GND 0.02967f
C11831 VDD.n2993 GND 0.05074f
C11832 VDD.n2994 GND 0.62973f
C11833 VDD.t941 GND 0.74438f
C11834 VDD.n2996 GND 0.04999f
C11835 VDD.t528 GND 0.63568f
C11836 VDD.n2997 GND 0.05074f
C11837 VDD.n2998 GND 0.05074f
C11838 VDD.n2999 GND 0.02967f
C11839 VDD.n3000 GND 0.02522f
C11840 VDD.t713 GND 0.02334f
C11841 VDD.t529 GND 0.02334f
C11842 VDD.n3001 GND 0.13341f
C11843 VDD.n3002 GND 0.0263f
C11844 VDD.n3003 GND 0.0536f
C11845 VDD.n3004 GND 0.05074f
C11846 VDD.n3005 GND 0.02967f
C11847 VDD.n3006 GND 0.02522f
C11848 VDD.n3007 GND 0.04999f
C11849 VDD.t151 GND 0.63568f
C11850 VDD.n3008 GND 0.05074f
C11851 VDD.n3009 GND 0.05074f
C11852 VDD.n3010 GND 0.02967f
C11853 VDD.n3011 GND 0.02522f
C11854 VDD.n3012 GND 0.03166f
C11855 VDD.n3013 GND 0.0536f
C11856 VDD.n3014 GND 0.05074f
C11857 VDD.n3015 GND 0.02967f
C11858 VDD.n3016 GND 0.02522f
C11859 VDD.n3017 GND 0.04999f
C11860 VDD.t1014 GND 0.63568f
C11861 VDD.n3018 GND 0.05074f
C11862 VDD.n3019 GND 0.05074f
C11863 VDD.n3020 GND 0.02967f
C11864 VDD.n3021 GND 0.02522f
C11865 VDD.t938 GND 0.02321f
C11866 VDD.t1015 GND 0.02321f
C11867 VDD.n3022 GND 0.10855f
C11868 VDD.t152 GND 0.02321f
C11869 VDD.t1064 GND 0.02321f
C11870 VDD.n3023 GND 0.10855f
C11871 VDD.n3024 GND 0.04152f
C11872 VDD.n3025 GND 0.02334f
C11873 VDD.n3026 GND 0.0536f
C11874 VDD.n3027 GND 0.05074f
C11875 VDD.n3028 GND 0.02967f
C11876 VDD.n3029 GND 0.02522f
C11877 VDD.n3030 GND 0.04999f
C11878 VDD.t484 GND 0.63568f
C11879 VDD.n3031 GND 0.05074f
C11880 VDD.n3032 GND 0.05074f
C11881 VDD.n3033 GND 0.02967f
C11882 VDD.n3034 GND 0.02522f
C11883 VDD.t485 GND 0.02334f
C11884 VDD.t665 GND 0.02334f
C11885 VDD.n3035 GND 0.13232f
C11886 VDD.n3036 GND 0.06172f
C11887 VDD.n3037 GND 0.76206f
C11888 VDD.t1140 GND 0.16977f
C11889 VDD.n3038 GND 0.17097f
C11890 VDD.n3039 GND 0.01824f
C11891 VDD.t726 GND 0.08826f
C11892 VDD.n3040 GND 0.02543f
C11893 VDD.n3042 GND 0.01055f
C11894 VDD.n3043 GND 0.02883f
C11895 VDD.t1134 GND 0.16976f
C11896 VDD.n3044 GND 0.04959f
C11897 VDD.n3045 GND 0.02152f
C11898 VDD.n3046 GND 0.09461f
C11899 VDD.t666 GND 0.07895f
C11900 VDD.n3047 GND 0.04531f
C11901 VDD.n3048 GND 0.14048f
C11902 VDD.t1120 GND 0.16977f
C11903 VDD.n3049 GND 0.17097f
C11904 VDD.n3050 GND 0.01824f
C11905 VDD.t728 GND 0.08826f
C11906 VDD.n3051 GND 0.02543f
C11907 VDD.n3053 GND 0.01055f
C11908 VDD.n3055 GND 0.18033f
C11909 VDD.n3056 GND 0.21978f
C11910 VDD.n3057 GND 0.76206f
C11911 VDD.t678 GND 0.08827f
C11912 VDD.n3058 GND 0.08234f
C11913 VDD.n3059 GND 0.01824f
C11914 VDD.t1126 GND 0.16976f
C11915 VDD.n3060 GND 0.04959f
C11916 VDD.n3061 GND 0.01646f
C11917 VDD.n3062 GND 0.02781f
C11918 VDD.n3063 GND 0.02883f
C11919 VDD.t1157 GND 0.16977f
C11920 VDD.n3064 GND 0.17602f
C11921 VDD.n3065 GND 0.01904f
C11922 VDD.n3066 GND 0.02543f
C11923 VDD.t754 GND 0.07929f
C11924 VDD.n3067 GND 0.15939f
C11925 VDD.n3068 GND 0.04531f
C11926 VDD.t720 GND 0.08827f
C11927 VDD.n3069 GND 0.08234f
C11928 VDD.n3070 GND 0.01824f
C11929 VDD.t1125 GND 0.16976f
C11930 VDD.n3071 GND 0.04959f
C11931 VDD.n3072 GND 0.01646f
C11932 VDD.n3073 GND 0.02781f
C11933 VDD.n3075 GND 0.1744f
C11934 VDD.n3076 GND 0.18262f
C11935 VDD.t1158 GND 0.16976f
C11936 VDD.n3077 GND 0.04959f
C11937 VDD.n3078 GND 0.01646f
C11938 VDD.n3079 GND 0.02781f
C11939 VDD.t1119 GND 0.16977f
C11940 VDD.n3080 GND 0.17602f
C11941 VDD.n3081 GND 0.01904f
C11942 VDD.n3082 GND 0.02543f
C11943 VDD.t716 GND 0.07929f
C11944 VDD.n3083 GND 0.15939f
C11945 VDD.n3084 GND 0.04531f
C11946 VDD.t746 GND 0.08827f
C11947 VDD.n3085 GND 0.08234f
C11948 VDD.n3086 GND 0.01824f
C11949 VDD.t1139 GND 0.16976f
C11950 VDD.n3087 GND 0.04959f
C11951 VDD.n3088 GND 0.01646f
C11952 VDD.n3089 GND 0.02781f
C11953 VDD.n3090 GND 0.10528f
C11954 VDD.n3091 GND 0.26745f
C11955 VDD.n3093 GND 0.01824f
C11956 VDD.n3094 GND 0.08234f
C11957 VDD.t668 GND 0.07819f
C11958 VDD.n3095 GND 0.14455f
C11959 VDD.n3096 GND 0.76206f
C11960 VDD.t662 GND 0.08827f
C11961 VDD.n3097 GND 0.08234f
C11962 VDD.n3098 GND 0.01824f
C11963 VDD.t1135 GND 0.16976f
C11964 VDD.n3099 GND 0.04959f
C11965 VDD.n3100 GND 0.01646f
C11966 VDD.n3101 GND 0.02781f
C11967 VDD.n3102 GND 0.02883f
C11968 VDD.t1143 GND 0.16977f
C11969 VDD.n3103 GND 0.17602f
C11970 VDD.n3104 GND 0.01904f
C11971 VDD.n3105 GND 0.02543f
C11972 VDD.t672 GND 0.07929f
C11973 VDD.n3106 GND 0.15939f
C11974 VDD.n3107 GND 0.04531f
C11975 VDD.t744 GND 0.08827f
C11976 VDD.n3108 GND 0.08234f
C11977 VDD.n3109 GND 0.01824f
C11978 VDD.t1111 GND 0.16976f
C11979 VDD.n3110 GND 0.04959f
C11980 VDD.n3111 GND 0.01646f
C11981 VDD.n3112 GND 0.02781f
C11982 VDD.n3114 GND 0.1744f
C11983 VDD.n3115 GND 0.18262f
C11984 VDD.t676 GND 0.08827f
C11985 VDD.n3116 GND 0.08234f
C11986 VDD.n3117 GND 0.01824f
C11987 VDD.t1127 GND 0.16976f
C11988 VDD.n3118 GND 0.04959f
C11989 VDD.n3119 GND 0.01646f
C11990 VDD.n3120 GND 0.02781f
C11991 VDD.n3121 GND 0.02883f
C11992 VDD.t1136 GND 0.16977f
C11993 VDD.n3122 GND 0.17602f
C11994 VDD.n3123 GND 0.01904f
C11995 VDD.n3124 GND 0.02543f
C11996 VDD.t692 GND 0.07929f
C11997 VDD.n3125 GND 0.15939f
C11998 VDD.n3126 GND 0.04531f
C11999 VDD.t760 GND 0.08827f
C12000 VDD.n3127 GND 0.08234f
C12001 VDD.n3128 GND 0.01824f
C12002 VDD.t1153 GND 0.16976f
C12003 VDD.n3129 GND 0.04959f
C12004 VDD.n3130 GND 0.01646f
C12005 VDD.n3131 GND 0.02781f
C12006 VDD.n3133 GND 0.1744f
C12007 VDD.n3134 GND 0.18262f
C12008 VDD.n3135 GND 1.91602f
C12009 VDD.t706 GND 0.08827f
C12010 VDD.n3136 GND 0.08234f
C12011 VDD.n3137 GND 0.01824f
C12012 VDD.t1113 GND 0.16976f
C12013 VDD.n3138 GND 0.04959f
C12014 VDD.n3139 GND 0.01646f
C12015 VDD.n3140 GND 0.02781f
C12016 VDD.n3141 GND 0.02883f
C12017 VDD.t1124 GND 0.16977f
C12018 VDD.n3142 GND 0.17602f
C12019 VDD.n3143 GND 0.01904f
C12020 VDD.n3144 GND 0.02543f
C12021 VDD.t752 GND 0.07929f
C12022 VDD.n3145 GND 0.15939f
C12023 VDD.n3146 GND 0.04531f
C12024 VDD.t674 GND 0.08827f
C12025 VDD.n3147 GND 0.08234f
C12026 VDD.n3148 GND 0.01824f
C12027 VDD.t1128 GND 0.16976f
C12028 VDD.n3149 GND 0.04959f
C12029 VDD.n3150 GND 0.01646f
C12030 VDD.n3151 GND 0.02781f
C12031 VDD.n3153 GND 0.1744f
C12032 VDD.n3154 GND 0.18262f
C12033 VDD.t1132 GND 0.16976f
C12034 VDD.n3155 GND 0.04959f
C12035 VDD.n3156 GND 0.01646f
C12036 VDD.n3157 GND 0.02781f
C12037 VDD.t1110 GND 0.16977f
C12038 VDD.n3158 GND 0.17602f
C12039 VDD.n3159 GND 0.01904f
C12040 VDD.n3160 GND 0.02543f
C12041 VDD.t748 GND 0.07929f
C12042 VDD.n3161 GND 0.15939f
C12043 VDD.n3162 GND 0.04531f
C12044 VDD.t742 GND 0.08827f
C12045 VDD.n3163 GND 0.08234f
C12046 VDD.n3164 GND 0.01824f
C12047 VDD.t1141 GND 0.16976f
C12048 VDD.n3165 GND 0.04959f
C12049 VDD.n3166 GND 0.01646f
C12050 VDD.n3167 GND 0.02781f
C12051 VDD.n3168 GND 0.10528f
C12052 VDD.n3169 GND 0.26745f
C12053 VDD.n3171 GND 0.01824f
C12054 VDD.n3172 GND 0.08234f
C12055 VDD.t700 GND 0.07819f
C12056 VDD.n3173 GND 0.14455f
C12057 VDD.t1149 GND 0.16976f
C12058 VDD.n3174 GND 0.04959f
C12059 VDD.n3175 GND 0.01646f
C12060 VDD.n3176 GND 0.02781f
C12061 VDD.t1121 GND 0.16977f
C12062 VDD.n3177 GND 0.17602f
C12063 VDD.n3178 GND 0.01904f
C12064 VDD.n3179 GND 0.02543f
C12065 VDD.t732 GND 0.07929f
C12066 VDD.n3180 GND 0.15939f
C12067 VDD.n3181 GND 0.04531f
C12068 VDD.t694 GND 0.08827f
C12069 VDD.n3182 GND 0.08234f
C12070 VDD.n3183 GND 0.01824f
C12071 VDD.t1116 GND 0.16976f
C12072 VDD.n3184 GND 0.04959f
C12073 VDD.n3185 GND 0.01646f
C12074 VDD.n3186 GND 0.02781f
C12075 VDD.n3187 GND 0.10528f
C12076 VDD.n3188 GND 0.26745f
C12077 VDD.n3190 GND 0.01824f
C12078 VDD.n3191 GND 0.08234f
C12079 VDD.t670 GND 0.07819f
C12080 VDD.n3192 GND 0.14455f
C12081 VDD.n3193 GND 1.56549f
C12082 VDD.n3194 GND 0.99189f
C12083 VDD.n3195 GND 0.37775f
C12084 VDD.n3196 GND 0.38258f
C12085 VDD.n3197 GND 1.56538f
C12086 VDD.n3198 GND 1.57029f
C12087 VDD.n3199 GND 0.80146f
C12088 VDD.t756 GND 0.08827f
C12089 VDD.n3200 GND 0.08234f
C12090 VDD.n3201 GND 0.01824f
C12091 VDD.t1156 GND 0.16976f
C12092 VDD.n3202 GND 0.04959f
C12093 VDD.n3203 GND 0.01646f
C12094 VDD.n3204 GND 0.02781f
C12095 VDD.n3205 GND 0.02883f
C12096 VDD.t1154 GND 0.16977f
C12097 VDD.n3206 GND 0.17602f
C12098 VDD.n3207 GND 0.01904f
C12099 VDD.n3208 GND 0.02543f
C12100 VDD.t758 GND 0.07929f
C12101 VDD.n3209 GND 0.15939f
C12102 VDD.n3210 GND 0.04531f
C12103 VDD.t680 GND 0.08827f
C12104 VDD.n3211 GND 0.08234f
C12105 VDD.n3212 GND 0.01824f
C12106 VDD.t1122 GND 0.16976f
C12107 VDD.n3213 GND 0.04959f
C12108 VDD.n3214 GND 0.01646f
C12109 VDD.n3215 GND 0.02781f
C12110 VDD.n3217 GND 0.1744f
C12111 VDD.n3218 GND 0.18262f
C12112 VDD.t1155 GND 0.16976f
C12113 VDD.n3219 GND 0.04959f
C12114 VDD.n3220 GND 0.01646f
C12115 VDD.n3221 GND 0.02781f
C12116 VDD.t1151 GND 0.16977f
C12117 VDD.n3222 GND 0.17602f
C12118 VDD.n3223 GND 0.01904f
C12119 VDD.n3224 GND 0.02543f
C12120 VDD.t684 GND 0.07929f
C12121 VDD.n3225 GND 0.15939f
C12122 VDD.n3226 GND 0.04531f
C12123 VDD.t750 GND 0.08827f
C12124 VDD.n3227 GND 0.08234f
C12125 VDD.n3228 GND 0.01824f
C12126 VDD.t1138 GND 0.16976f
C12127 VDD.n3229 GND 0.04959f
C12128 VDD.n3230 GND 0.01646f
C12129 VDD.n3231 GND 0.02781f
C12130 VDD.n3232 GND 0.10528f
C12131 VDD.n3233 GND 0.26745f
C12132 VDD.n3235 GND 0.01824f
C12133 VDD.n3236 GND 0.08234f
C12134 VDD.t722 GND 0.07819f
C12135 VDD.n3237 GND 0.14455f
C12136 VDD.n3238 GND 1.56538f
C12137 VDD.n3239 GND 1.57029f
C12138 VDD.n3240 GND 0.76206f
C12139 VDD.n3241 GND 0.76206f
C12140 VDD.n3242 GND 1.57029f
C12141 VDD.t1130 GND 0.16976f
C12142 VDD.n3243 GND 0.04959f
C12143 VDD.n3244 GND 0.01646f
C12144 VDD.n3245 GND 0.02781f
C12145 VDD.t1133 GND 0.16977f
C12146 VDD.n3246 GND 0.17602f
C12147 VDD.n3247 GND 0.01904f
C12148 VDD.n3248 GND 0.02543f
C12149 VDD.t696 GND 0.07929f
C12150 VDD.n3249 GND 0.15939f
C12151 VDD.n3250 GND 0.04531f
C12152 VDD.t702 GND 0.08827f
C12153 VDD.n3251 GND 0.08234f
C12154 VDD.n3252 GND 0.01824f
C12155 VDD.t1129 GND 0.16976f
C12156 VDD.n3253 GND 0.04959f
C12157 VDD.n3254 GND 0.01646f
C12158 VDD.n3255 GND 0.02781f
C12159 VDD.n3256 GND 0.10528f
C12160 VDD.n3257 GND 0.26745f
C12161 VDD.n3259 GND 0.01824f
C12162 VDD.n3260 GND 0.08234f
C12163 VDD.t688 GND 0.07819f
C12164 VDD.n3261 GND 0.14455f
C12165 VDD.n3262 GND 1.56538f
C12166 VDD.n3263 GND 0.76206f
C12167 VDD.n3264 GND 0.34136f
C12168 VDD.t903 GND 0.02334f
C12169 VDD.t87 GND 0.02334f
C12170 VDD.n3265 GND 0.14146f
C12171 VDD.n3266 GND 0.0536f
C12172 VDD.n3267 GND 0.05074f
C12173 VDD.n3268 GND 0.0536f
C12174 VDD.n3269 GND 0.04999f
C12175 VDD.n3270 GND 0.04999f
C12176 VDD.n3271 GND 0.68843f
C12177 VDD.n3272 GND 0.02522f
C12178 VDD.n3273 GND 0.02522f
C12179 VDD.n3274 GND 0.02967f
C12180 VDD.n3275 GND 0.05074f
C12181 VDD.n3276 GND 0.04999f
C12182 VDD.t88 GND 0.63568f
C12183 VDD.n3277 GND 0.05074f
C12184 VDD.n3278 GND 0.05074f
C12185 VDD.n3279 GND 0.02967f
C12186 VDD.n3280 GND 0.02522f
C12187 VDD.n3281 GND 0.03042f
C12188 VDD.n3282 GND 0.0536f
C12189 VDD.n3283 GND 0.05074f
C12190 VDD.n3284 GND 0.02967f
C12191 VDD.n3285 GND 0.02522f
C12192 VDD.n3286 GND 0.04999f
C12193 VDD.t21 GND 0.63568f
C12194 VDD.n3287 GND 0.05074f
C12195 VDD.n3288 GND 0.05074f
C12196 VDD.n3289 GND 0.02967f
C12197 VDD.n3290 GND 0.02522f
C12198 VDD.n3291 GND 0.0536f
C12199 VDD.n3292 GND 0.05074f
C12200 VDD.n3293 GND 0.02967f
C12201 VDD.n3294 GND 0.02522f
C12202 VDD.n3295 GND 0.02522f
C12203 VDD.n3296 GND 0.04999f
C12204 VDD.n3297 GND 0.68843f
C12205 VDD.n3298 GND 0.04999f
C12206 VDD.n3299 GND 0.05074f
C12207 VDD.n3300 GND 0.19438f
C12208 VDD.n3301 GND 0.03542f
C12209 VDD.t138 GND 0.02552f
C12210 VDD.n3302 GND 0.09114f
C12211 VDD.n3303 GND 0.03545f
C12212 VDD.n3305 GND 0.56273f
C12213 VDD.n3306 GND 0.02746f
C12214 VDD.n3307 GND 0.05074f
C12215 VDD.n3308 GND 0.02967f
C12216 VDD.n3309 GND 0.05074f
C12217 VDD.t998 GND 0.30977f
C12218 VDD.n3310 GND 0.05074f
C12219 VDD.n3311 GND 0.05074f
C12220 VDD.n3312 GND 0.02967f
C12221 VDD.n3313 GND 0.02746f
C12222 VDD.t997 GND 0.02334f
C12223 VDD.n3314 GND 0.34117f
C12224 VDD.t272 GND 0.02334f
C12225 VDD.n3315 GND 0.08128f
C12226 VDD.n3316 GND 0.02746f
C12227 VDD.n3317 GND 0.05074f
C12228 VDD.n3318 GND 0.02967f
C12229 VDD.n3319 GND 0.05074f
C12230 VDD.n3320 GND 0.35737f
C12231 VDD.t271 GND 0.33785f
C12232 VDD.t256 GND 0.30977f
C12233 VDD.n3322 GND 0.05074f
C12234 VDD.n3323 GND 0.05074f
C12235 VDD.n3324 GND 0.02967f
C12236 VDD.n3325 GND 0.02746f
C12237 VDD.n3326 GND 0.02746f
C12238 VDD.n3327 GND 0.05074f
C12239 VDD.n3328 GND 0.02967f
C12240 VDD.n3329 GND 0.05074f
C12241 VDD.n3330 GND 0.04999f
C12242 VDD.n3331 GND 0.24979f
C12243 VDD.n3332 GND 0.04999f
C12244 VDD.n3333 GND 0.24979f
C12245 VDD.t884 GND 0.33785f
C12246 VDD.n3335 GND 0.35737f
C12247 VDD.n3336 GND 0.02746f
C12248 VDD.n3337 GND 0.09132f
C12249 VDD.n3338 GND 0.04596f
C12250 VDD.t132 GND 0.02552f
C12251 VDD.n3339 GND 0.09115f
C12252 VDD.n3340 GND 0.03542f
C12253 VDD.n3342 GND 0.91591f
C12254 VDD.n3343 GND 0.02746f
C12255 VDD.n3344 GND 0.05074f
C12256 VDD.n3345 GND 0.02967f
C12257 VDD.n3346 GND 0.05074f
C12258 VDD.t176 GND 0.30977f
C12259 VDD.n3347 GND 0.05074f
C12260 VDD.n3348 GND 0.05074f
C12261 VDD.n3349 GND 0.02967f
C12262 VDD.n3350 GND 0.02746f
C12263 VDD.t855 GND 0.02334f
C12264 VDD.t734 GND 0.08827f
C12265 VDD.n3351 GND 0.08234f
C12266 VDD.n3352 GND 0.01824f
C12267 VDD.t1152 GND 0.16976f
C12268 VDD.n3353 GND 0.04959f
C12269 VDD.n3354 GND 0.01646f
C12270 VDD.n3355 GND 0.02781f
C12271 VDD.n3356 GND 0.02883f
C12272 VDD.t1114 GND 0.16977f
C12273 VDD.n3357 GND 0.17602f
C12274 VDD.n3358 GND 0.01904f
C12275 VDD.n3359 GND 0.02543f
C12276 VDD.t736 GND 0.07929f
C12277 VDD.n3360 GND 0.15939f
C12278 VDD.n3361 GND 0.04531f
C12279 VDD.t762 GND 0.08827f
C12280 VDD.n3362 GND 0.08234f
C12281 VDD.n3363 GND 0.01824f
C12282 VDD.t1137 GND 0.16976f
C12283 VDD.n3364 GND 0.04959f
C12284 VDD.n3365 GND 0.01646f
C12285 VDD.n3366 GND 0.02781f
C12286 VDD.n3368 GND 0.1744f
C12287 VDD.n3369 GND 0.18262f
C12288 VDD.n3370 GND 0.29196f
C12289 VDD.t783 GND 0.02334f
C12290 VDD.n3371 GND 0.08128f
C12291 VDD.n3372 GND 0.02746f
C12292 VDD.n3373 GND 0.05074f
C12293 VDD.n3374 GND 0.02967f
C12294 VDD.n3375 GND 0.05074f
C12295 VDD.n3376 GND 0.35737f
C12296 VDD.t782 GND 0.33785f
C12297 VDD.t784 GND 0.30977f
C12298 VDD.n3378 GND 0.05074f
C12299 VDD.n3379 GND 0.05074f
C12300 VDD.n3380 GND 0.02967f
C12301 VDD.n3381 GND 0.02746f
C12302 VDD.n3382 GND 0.02746f
C12303 VDD.n3383 GND 0.05074f
C12304 VDD.n3384 GND 0.02967f
C12305 VDD.n3385 GND 0.05074f
C12306 VDD.n3386 GND 0.04999f
C12307 VDD.n3387 GND 0.24979f
C12308 VDD.n3388 GND 0.04999f
C12309 VDD.n3389 GND 0.24979f
C12310 VDD.t206 GND 0.33785f
C12311 VDD.n3391 GND 0.35737f
C12312 VDD.n3392 GND 0.02746f
C12313 VDD.n3393 GND 0.09132f
C12314 VDD.n3394 GND 1.08589f
C12315 VDD.t781 GND 0.03067f
C12316 VDD.n3395 GND 0.14083f
C12317 VDD.n3396 GND 0.03755f
C12318 VDD.t207 GND 0.02552f
C12319 VDD.n3397 GND 0.09115f
C12320 VDD.n3398 GND 0.03755f
C12321 VDD.n3399 GND 0.07974f
C12322 VDD.t813 GND 0.03065f
C12323 VDD.n3400 GND 0.17961f
C12324 VDD.n3401 GND 0.12536f
C12325 VDD.t986 GND 0.02552f
C12326 VDD.n3402 GND 0.09115f
C12327 VDD.n3403 GND 0.03755f
C12328 VDD.n3404 GND 0.07974f
C12329 VDD.t177 GND 0.03065f
C12330 VDD.n3405 GND 0.15984f
C12331 VDD.n3406 GND 0.10559f
C12332 VDD.n3408 GND 0.03542f
C12333 VDD.n3409 GND 0.03042f
C12334 VDD.n3410 GND 0.09132f
C12335 VDD.n3411 GND 0.02746f
C12336 VDD.n3412 GND 0.04999f
C12337 VDD.n3413 GND 0.24979f
C12338 VDD.n3414 GND 0.24979f
C12339 VDD.n3415 GND 0.04999f
C12340 VDD.n3416 GND 0.02746f
C12341 VDD.n3417 GND 0.09132f
C12342 VDD.n3418 GND 0.01581f
C12343 VDD.n3419 GND 0.12361f
C12344 VDD.n3420 GND 0.36368f
C12345 VDD.n3421 GND 0.3214f
C12346 VDD.n3422 GND 0.12361f
C12347 VDD.n3423 GND 0.02746f
C12348 VDD.n3424 GND 0.05074f
C12349 VDD.n3425 GND 0.02967f
C12350 VDD.n3426 GND 0.05074f
C12351 VDD.n3427 GND 0.35737f
C12352 VDD.t854 GND 0.33785f
C12353 VDD.n3429 GND 0.04999f
C12354 VDD.n3430 GND 0.24979f
C12355 VDD.n3431 GND 0.24979f
C12356 VDD.n3432 GND 0.04999f
C12357 VDD.n3433 GND 0.02746f
C12358 VDD.n3434 GND 0.09132f
C12359 VDD.n3435 GND 0.01581f
C12360 VDD.n3436 GND 0.08128f
C12361 VDD.n3437 GND 0.03542f
C12362 VDD.n3438 GND 0.03042f
C12363 VDD.n3439 GND 0.09132f
C12364 VDD.n3440 GND 0.02746f
C12365 VDD.n3441 GND 0.04999f
C12366 VDD.n3442 GND 0.24979f
C12367 VDD.n3443 GND 0.04999f
C12368 VDD.n3444 GND 0.24979f
C12369 VDD.t985 GND 0.33785f
C12370 VDD.n3446 GND 0.35737f
C12371 VDD.n3447 GND 0.02746f
C12372 VDD.n3448 GND 0.09132f
C12373 VDD.n3449 GND 0.04596f
C12374 VDD.n3450 GND 0.80829f
C12375 VDD.n3451 GND 0.68551f
C12376 VDD.n3452 GND 0.02746f
C12377 VDD.n3453 GND 0.05074f
C12378 VDD.n3454 GND 0.02967f
C12379 VDD.n3455 GND 0.05074f
C12380 VDD.t812 GND 0.30977f
C12381 VDD.n3456 GND 0.05074f
C12382 VDD.n3457 GND 0.05074f
C12383 VDD.n3458 GND 0.02967f
C12384 VDD.n3459 GND 0.02746f
C12385 VDD.t811 GND 0.02334f
C12386 VDD.n3460 GND 0.12361f
C12387 VDD.n3461 GND 0.02746f
C12388 VDD.n3462 GND 0.05074f
C12389 VDD.n3463 GND 0.02967f
C12390 VDD.n3464 GND 0.05074f
C12391 VDD.n3465 GND 0.35737f
C12392 VDD.t810 GND 0.33785f
C12393 VDD.n3467 GND 0.04999f
C12394 VDD.n3468 GND 0.24979f
C12395 VDD.n3469 GND 0.24979f
C12396 VDD.n3470 GND 0.04999f
C12397 VDD.n3471 GND 0.02746f
C12398 VDD.n3472 GND 0.09132f
C12399 VDD.n3473 GND 0.01581f
C12400 VDD.n3474 GND 0.08128f
C12401 VDD.n3475 GND 0.03042f
C12402 VDD.n3476 GND 0.09132f
C12403 VDD.n3477 GND 0.02746f
C12404 VDD.n3478 GND 0.04999f
C12405 VDD.n3479 GND 0.24979f
C12406 VDD.n3480 GND 0.04999f
C12407 VDD.n3481 GND 0.24979f
C12408 VDD.t131 GND 0.33785f
C12409 VDD.n3483 GND 0.35737f
C12410 VDD.n3484 GND 0.02746f
C12411 VDD.n3485 GND 0.09132f
C12412 VDD.n3486 GND 0.04596f
C12413 VDD.n3488 GND 0.12536f
C12414 VDD.t270 GND 0.03065f
C12415 VDD.n3489 GND 0.17961f
C12416 VDD.n3490 GND 0.07974f
C12417 VDD.n3491 GND 0.03755f
C12418 VDD.t885 GND 0.02552f
C12419 VDD.n3492 GND 0.09115f
C12420 VDD.n3493 GND 0.03755f
C12421 VDD.n3494 GND 0.07974f
C12422 VDD.t53 GND 0.03065f
C12423 VDD.n3495 GND 0.17961f
C12424 VDD.n3496 GND 0.12536f
C12425 VDD.t123 GND 0.02552f
C12426 VDD.n3497 GND 0.09115f
C12427 VDD.n3498 GND 0.03755f
C12428 VDD.n3499 GND 0.07974f
C12429 VDD.t993 GND 0.03065f
C12430 VDD.n3500 GND 0.33976f
C12431 VDD.n3501 GND 0.28551f
C12432 VDD.n3503 GND 0.03542f
C12433 VDD.n3504 GND 0.03042f
C12434 VDD.n3505 GND 0.09132f
C12435 VDD.n3506 GND 0.02746f
C12436 VDD.n3507 GND 0.04999f
C12437 VDD.n3508 GND 0.24979f
C12438 VDD.n3509 GND 0.24979f
C12439 VDD.n3510 GND 0.04999f
C12440 VDD.n3511 GND 0.02746f
C12441 VDD.n3512 GND 0.09132f
C12442 VDD.n3513 GND 0.01581f
C12443 VDD.n3514 GND 0.12361f
C12444 VDD.n3515 GND 0.50133f
C12445 VDD.n3516 GND 0.50133f
C12446 VDD.n3517 GND 0.12361f
C12447 VDD.n3518 GND 0.02746f
C12448 VDD.n3519 GND 0.05074f
C12449 VDD.n3520 GND 0.02967f
C12450 VDD.n3521 GND 0.05074f
C12451 VDD.n3522 GND 0.35737f
C12452 VDD.t996 GND 0.33785f
C12453 VDD.n3524 GND 0.04999f
C12454 VDD.n3525 GND 0.24979f
C12455 VDD.n3526 GND 0.24979f
C12456 VDD.n3527 GND 0.04999f
C12457 VDD.n3528 GND 0.02746f
C12458 VDD.n3529 GND 0.09132f
C12459 VDD.n3530 GND 0.01581f
C12460 VDD.n3531 GND 0.08128f
C12461 VDD.n3532 GND 0.03542f
C12462 VDD.n3533 GND 0.03042f
C12463 VDD.n3534 GND 0.09132f
C12464 VDD.n3535 GND 0.02746f
C12465 VDD.n3536 GND 0.04999f
C12466 VDD.n3537 GND 0.24979f
C12467 VDD.n3538 GND 0.04999f
C12468 VDD.n3539 GND 0.24979f
C12469 VDD.t122 GND 0.33785f
C12470 VDD.n3541 GND 0.35737f
C12471 VDD.n3542 GND 0.02746f
C12472 VDD.n3543 GND 0.09132f
C12473 VDD.n3544 GND 0.04596f
C12474 VDD.n3545 GND 0.31716f
C12475 VDD.n3546 GND 0.02746f
C12476 VDD.n3547 GND 0.05074f
C12477 VDD.n3548 GND 0.02967f
C12478 VDD.n3549 GND 0.05074f
C12479 VDD.t410 GND 0.30977f
C12480 VDD.n3550 GND 0.05074f
C12481 VDD.n3551 GND 0.05074f
C12482 VDD.n3552 GND 0.02967f
C12483 VDD.n3553 GND 0.02746f
C12484 VDD.t409 GND 0.02334f
C12485 VDD.n3554 GND 0.12361f
C12486 VDD.n3555 GND 0.02746f
C12487 VDD.n3556 GND 0.05074f
C12488 VDD.n3557 GND 0.02967f
C12489 VDD.n3558 GND 0.05074f
C12490 VDD.n3559 GND 0.35737f
C12491 VDD.t408 GND 0.33785f
C12492 VDD.n3561 GND 0.04999f
C12493 VDD.n3562 GND 0.24979f
C12494 VDD.n3563 GND 0.24979f
C12495 VDD.n3564 GND 0.04999f
C12496 VDD.n3565 GND 0.02746f
C12497 VDD.n3566 GND 0.09132f
C12498 VDD.n3567 GND 0.01581f
C12499 VDD.n3568 GND 0.08128f
C12500 VDD.n3569 GND 0.03042f
C12501 VDD.n3570 GND 0.09132f
C12502 VDD.n3571 GND 0.02746f
C12503 VDD.n3572 GND 0.04999f
C12504 VDD.n3573 GND 0.24979f
C12505 VDD.n3574 GND 0.04999f
C12506 VDD.n3575 GND 0.24979f
C12507 VDD.t137 GND 0.33785f
C12508 VDD.n3577 GND 0.35737f
C12509 VDD.n3578 GND 0.02746f
C12510 VDD.n3579 GND 0.09132f
C12511 VDD.n3580 GND 0.04635f
C12512 VDD.n3582 GND 0.12555f
C12513 VDD.t902 GND 0.03065f
C12514 VDD.n3583 GND 0.17979f
C12515 VDD.n3584 GND 0.07974f
C12516 VDD.n3585 GND 0.03755f
C12517 VDD.t569 GND 0.02552f
C12518 VDD.n3586 GND 0.09115f
C12519 VDD.t805 GND 0.03067f
C12520 VDD.n3587 GND 0.03755f
C12521 VDD.n3588 GND 0.07974f
C12522 VDD.t22 GND 0.02552f
C12523 VDD.n3589 GND 0.09139f
C12524 VDD.n3590 GND 0.0569f
C12525 VDD.n3592 GND 0.04596f
C12526 VDD.n3593 GND 0.06295f
C12527 VDD.n3594 GND 0.0536f
C12528 VDD.n3595 GND 0.02522f
C12529 VDD.n3596 GND 0.04999f
C12530 VDD.n3597 GND 0.5126f
C12531 VDD.n3598 GND 0.02522f
C12532 VDD.n3599 GND 0.04999f
C12533 VDD.n3600 GND 0.5126f
C12534 VDD.n3601 GND 0.04999f
C12535 VDD.n3602 GND 0.05074f
C12536 VDD.n3603 GND 0.06295f
C12537 VDD.n3604 GND 0.0536f
C12538 VDD.n3605 GND 0.02522f
C12539 VDD.n3606 GND 0.04999f
C12540 VDD.n3607 GND 0.5126f
C12541 VDD.n3608 GND 0.5126f
C12542 VDD.n3609 GND 0.04999f
C12543 VDD.n3610 GND 0.04999f
C12544 VDD.n3611 GND 0.02522f
C12545 VDD.n3612 GND 0.02522f
C12546 VDD.n3613 GND 0.02967f
C12547 VDD.n3614 GND 0.05074f
C12548 VDD.t86 GND 0.63568f
C12549 VDD.n3615 GND 0.05074f
C12550 VDD.n3616 GND 0.06295f
C12551 VDD.n3617 GND 0.01581f
C12552 VDD.n3618 GND 0.12361f
C12553 VDD.n3619 GND 0.35808f
C12554 VDD.t1115 GND 0.16976f
C12555 VDD.n3620 GND 0.04959f
C12556 VDD.n3621 GND 0.01646f
C12557 VDD.n3622 GND 0.02781f
C12558 VDD.t1147 GND 0.16977f
C12559 VDD.n3623 GND 0.17602f
C12560 VDD.n3624 GND 0.01904f
C12561 VDD.n3625 GND 0.02543f
C12562 VDD.t690 GND 0.07929f
C12563 VDD.n3626 GND 0.15939f
C12564 VDD.n3627 GND 0.04531f
C12565 VDD.t730 GND 0.08827f
C12566 VDD.n3628 GND 0.08234f
C12567 VDD.n3629 GND 0.01824f
C12568 VDD.t1146 GND 0.16976f
C12569 VDD.n3630 GND 0.04959f
C12570 VDD.n3631 GND 0.01646f
C12571 VDD.n3632 GND 0.02781f
C12572 VDD.n3633 GND 0.10528f
C12573 VDD.n3634 GND 0.26745f
C12574 VDD.n3636 GND 0.01824f
C12575 VDD.n3637 GND 0.08234f
C12576 VDD.t714 GND 0.07819f
C12577 VDD.n3638 GND 0.14455f
C12578 VDD.n3639 GND 0.26149f
C12579 VDD.n3640 GND 0.76206f
C12580 VDD.n3641 GND 0.76206f
C12581 VDD.n3642 GND 1.56538f
C12582 VDD.n3643 GND 1.57029f
C12583 VDD.n3644 GND 0.76206f
C12584 VDD.t704 GND 0.08827f
C12585 VDD.n3645 GND 0.08234f
C12586 VDD.n3646 GND 0.01824f
C12587 VDD.t1112 GND 0.16976f
C12588 VDD.n3647 GND 0.04959f
C12589 VDD.n3648 GND 0.01646f
C12590 VDD.n3649 GND 0.02781f
C12591 VDD.n3650 GND 0.02883f
C12592 VDD.t1144 GND 0.16977f
C12593 VDD.n3651 GND 0.17602f
C12594 VDD.n3652 GND 0.01904f
C12595 VDD.n3653 GND 0.02543f
C12596 VDD.t708 GND 0.07929f
C12597 VDD.n3654 GND 0.15939f
C12598 VDD.n3655 GND 0.04531f
C12599 VDD.t740 GND 0.08827f
C12600 VDD.n3656 GND 0.08234f
C12601 VDD.n3657 GND 0.01824f
C12602 VDD.t1145 GND 0.16976f
C12603 VDD.n3658 GND 0.04959f
C12604 VDD.n3659 GND 0.01646f
C12605 VDD.n3660 GND 0.02781f
C12606 VDD.n3662 GND 0.1744f
C12607 VDD.n3663 GND 0.18262f
C12608 VDD.t1131 GND 0.16976f
C12609 VDD.n3664 GND 0.04959f
C12610 VDD.n3665 GND 0.01646f
C12611 VDD.n3666 GND 0.02781f
C12612 VDD.t1109 GND 0.16977f
C12613 VDD.n3667 GND 0.17602f
C12614 VDD.n3668 GND 0.01904f
C12615 VDD.n3669 GND 0.02543f
C12616 VDD.t738 GND 0.07929f
C12617 VDD.n3670 GND 0.15939f
C12618 VDD.n3671 GND 0.04531f
C12619 VDD.t698 GND 0.08827f
C12620 VDD.n3672 GND 0.08234f
C12621 VDD.n3673 GND 0.01824f
C12622 VDD.t1108 GND 0.16976f
C12623 VDD.n3674 GND 0.04959f
C12624 VDD.n3675 GND 0.01646f
C12625 VDD.n3676 GND 0.02781f
C12626 VDD.n3677 GND 0.10528f
C12627 VDD.n3678 GND 0.26745f
C12628 VDD.n3680 GND 0.01824f
C12629 VDD.n3681 GND 0.08234f
C12630 VDD.t682 GND 0.07819f
C12631 VDD.n3682 GND 0.14455f
C12632 VDD.n3683 GND 1.56538f
C12633 VDD.n3684 GND 1.57029f
C12634 VDD.n3685 GND 0.80146f
C12635 VDD.n3686 GND 2.02412f
C12636 VDD.t1117 GND 0.16976f
C12637 VDD.n3687 GND 0.04959f
C12638 VDD.n3688 GND 0.01646f
C12639 VDD.n3689 GND 0.02781f
C12640 VDD.t1150 GND 0.16977f
C12641 VDD.n3690 GND 0.17602f
C12642 VDD.n3691 GND 0.01904f
C12643 VDD.n3692 GND 0.02543f
C12644 VDD.t686 GND 0.07929f
C12645 VDD.n3693 GND 0.15939f
C12646 VDD.n3694 GND 0.04531f
C12647 VDD.t724 GND 0.08827f
C12648 VDD.n3695 GND 0.08234f
C12649 VDD.n3696 GND 0.01824f
C12650 VDD.t1148 GND 0.16976f
C12651 VDD.n3697 GND 0.04959f
C12652 VDD.n3698 GND 0.01646f
C12653 VDD.n3699 GND 0.02781f
C12654 VDD.n3700 GND 0.10528f
C12655 VDD.n3701 GND 0.26745f
C12656 VDD.n3703 GND 0.01824f
C12657 VDD.n3704 GND 0.08234f
C12658 VDD.t710 GND 0.07819f
C12659 VDD.n3705 GND 0.14455f
C12660 VDD.n3706 GND 1.56538f
C12661 VDD.n3707 GND 0.81968f
C12662 VDD.t1142 GND 0.16976f
C12663 VDD.n3708 GND 0.04959f
C12664 VDD.n3709 GND 0.01646f
C12665 VDD.n3710 GND 0.02781f
C12666 VDD.t1123 GND 0.16977f
C12667 VDD.n3711 GND 0.17602f
C12668 VDD.n3712 GND 0.01904f
C12669 VDD.n3713 GND 0.02543f
C12670 VDD.t712 GND 0.07929f
C12671 VDD.n3714 GND 0.15939f
C12672 VDD.n3715 GND 0.04531f
C12673 VDD.t718 GND 0.08827f
C12674 VDD.n3716 GND 0.08234f
C12675 VDD.n3717 GND 0.01824f
C12676 VDD.t1118 GND 0.16976f
C12677 VDD.n3718 GND 0.04959f
C12678 VDD.n3719 GND 0.01646f
C12679 VDD.n3720 GND 0.02781f
C12680 VDD.n3721 GND 0.10528f
C12681 VDD.n3722 GND 0.26745f
C12682 VDD.n3724 GND 0.01824f
C12683 VDD.n3725 GND 0.08234f
C12684 VDD.t664 GND 0.07819f
C12685 VDD.n3726 GND 0.55963f
C12686 VDD.n3728 GND 0.0536f
C12687 VDD.n3729 GND 0.05074f
C12688 VDD.n3730 GND 0.02967f
C12689 VDD.n3731 GND 0.02522f
C12690 VDD.n3732 GND 0.04999f
C12691 VDD.t51 GND 0.63568f
C12692 VDD.n3733 GND 0.05074f
C12693 VDD.n3734 GND 0.05074f
C12694 VDD.n3735 GND 0.02967f
C12695 VDD.n3736 GND 0.02522f
C12696 VDD.n3737 GND 0.0536f
C12697 VDD.n3738 GND 0.05074f
C12698 VDD.n3739 GND 0.09652f
C12699 VDD.t52 GND 0.02321f
C12700 VDD.t283 GND 0.02321f
C12701 VDD.n3740 GND 0.10855f
C12702 VDD.t111 GND 0.02321f
C12703 VDD.t232 GND 0.02321f
C12704 VDD.n3741 GND 0.10855f
C12705 VDD.n3742 GND 0.0536f
C12706 VDD.n3743 GND 0.05074f
C12707 VDD.n3744 GND 0.0536f
C12708 VDD.n3745 GND 0.04999f
C12709 VDD.n3746 GND 0.04999f
C12710 VDD.n3747 GND 0.05074f
C12711 VDD.n3748 GND 0.02967f
C12712 VDD.n3749 GND 0.02522f
C12713 VDD.n3750 GND 0.04999f
C12714 VDD.n3751 GND 0.02522f
C12715 VDD.n3752 GND 0.04999f
C12716 VDD.n3753 GND 0.5126f
C12717 VDD.n3754 GND 0.5126f
C12718 VDD.n3755 GND 0.02522f
C12719 VDD.n3756 GND 0.02522f
C12720 VDD.n3757 GND 0.02967f
C12721 VDD.n3758 GND 0.05074f
C12722 VDD.t1091 GND 0.63568f
C12723 VDD.n3759 GND 0.05074f
C12724 VDD.n3760 GND 0.05074f
C12725 VDD.n3761 GND 0.09132f
C12726 VDD.n3762 GND 0.04999f
C12727 VDD.t284 GND 0.63568f
C12728 VDD.n3763 GND 0.05074f
C12729 VDD.n3764 GND 0.05074f
C12730 VDD.n3765 GND 0.02967f
C12731 VDD.n3766 GND 0.02522f
C12732 VDD.t1092 GND 0.02334f
C12733 VDD.n3767 GND 0.0731f
C12734 VDD.n3768 GND 0.01798f
C12735 VDD.n3769 GND 0.02334f
C12736 VDD.n3770 GND 0.0536f
C12737 VDD.n3771 GND 0.05074f
C12738 VDD.n3772 GND 0.02967f
C12739 VDD.n3773 GND 0.02522f
C12740 VDD.n3774 GND 0.04999f
C12741 VDD.t558 GND 0.63568f
C12742 VDD.n3775 GND 0.05074f
C12743 VDD.n3776 GND 0.05074f
C12744 VDD.n3777 GND 0.02967f
C12745 VDD.n3778 GND 0.02522f
C12746 VDD.t570 GND 0.02321f
C12747 VDD.t559 GND 0.02321f
C12748 VDD.n3779 GND 0.10855f
C12749 VDD.t285 GND 0.02321f
C12750 VDD.t967 GND 0.02321f
C12751 VDD.n3780 GND 0.10855f
C12752 VDD.n3781 GND 0.04152f
C12753 VDD.n3782 GND 0.02334f
C12754 VDD.n3783 GND 0.0536f
C12755 VDD.n3784 GND 0.05074f
C12756 VDD.n3785 GND 0.02967f
C12757 VDD.n3786 GND 0.02522f
C12758 VDD.n3787 GND 0.04999f
C12759 VDD.t445 GND 0.63568f
C12760 VDD.n3788 GND 0.05074f
C12761 VDD.n3789 GND 0.05074f
C12762 VDD.n3790 GND 0.02967f
C12763 VDD.n3791 GND 0.02522f
C12764 VDD.t446 GND 0.02334f
C12765 VDD.t719 GND 0.02334f
C12766 VDD.n3792 GND 0.13341f
C12767 VDD.n3793 GND 0.0263f
C12768 VDD.n3794 GND 0.0536f
C12769 VDD.n3795 GND 0.05074f
C12770 VDD.n3796 GND 0.02967f
C12771 VDD.n3797 GND 0.02522f
C12772 VDD.n3798 GND 0.04999f
C12773 VDD.t427 GND 0.63568f
C12774 VDD.n3799 GND 0.05074f
C12775 VDD.n3800 GND 0.05074f
C12776 VDD.n3801 GND 0.02967f
C12777 VDD.n3802 GND 0.02522f
C12778 VDD.n3803 GND 0.03166f
C12779 VDD.n3804 GND 0.0536f
C12780 VDD.n3805 GND 0.05074f
C12781 VDD.n3806 GND 0.02967f
C12782 VDD.n3807 GND 0.02522f
C12783 VDD.n3808 GND 0.04999f
C12784 VDD.t235 GND 0.63568f
C12785 VDD.n3809 GND 0.05074f
C12786 VDD.n3810 GND 0.05074f
C12787 VDD.n3811 GND 0.02967f
C12788 VDD.n3812 GND 0.02522f
C12789 VDD.t428 GND 0.02321f
C12790 VDD.t236 GND 0.02321f
C12791 VDD.n3813 GND 0.10855f
C12792 VDD.t862 GND 0.02321f
C12793 VDD.t890 GND 0.02321f
C12794 VDD.n3814 GND 0.10855f
C12795 VDD.n3815 GND 0.04152f
C12796 VDD.n3816 GND 0.02334f
C12797 VDD.n3817 GND 0.0536f
C12798 VDD.n3818 GND 0.05074f
C12799 VDD.n3819 GND 0.02967f
C12800 VDD.n3820 GND 0.02522f
C12801 VDD.n3821 GND 0.02522f
C12802 VDD.n3822 GND 0.04999f
C12803 VDD.n3823 GND 0.68843f
C12804 VDD.n3824 GND 0.04999f
C12805 VDD.n3825 GND 0.05074f
C12806 VDD.n3826 GND 0.06295f
C12807 VDD.n3827 GND 0.0536f
C12808 VDD.n3828 GND 0.02522f
C12809 VDD.n3829 GND 0.04999f
C12810 VDD.n3830 GND 0.5126f
C12811 VDD.n3831 GND 0.02522f
C12812 VDD.n3832 GND 0.04999f
C12813 VDD.n3833 GND 0.5126f
C12814 VDD.n3834 GND 0.04999f
C12815 VDD.n3835 GND 0.05074f
C12816 VDD.n3836 GND 0.06295f
C12817 VDD.n3837 GND 0.0536f
C12818 VDD.n3838 GND 0.02522f
C12819 VDD.n3839 GND 0.04999f
C12820 VDD.n3840 GND 0.5126f
C12821 VDD.n3841 GND 0.02522f
C12822 VDD.n3842 GND 0.04999f
C12823 VDD.n3843 GND 0.5126f
C12824 VDD.n3844 GND 0.04999f
C12825 VDD.n3845 GND 0.05074f
C12826 VDD.n3846 GND 0.06295f
C12827 VDD.n3847 GND 0.0536f
C12828 VDD.n3848 GND 0.02522f
C12829 VDD.n3849 GND 0.04999f
C12830 VDD.n3850 GND 0.68843f
C12831 VDD.n3851 GND 0.02522f
C12832 VDD.n3852 GND 0.04999f
C12833 VDD.n3853 GND 0.68843f
C12834 VDD.n3854 GND 0.04999f
C12835 VDD.n3855 GND 0.05074f
C12836 VDD.n3856 GND 0.06295f
C12837 VDD.n3857 GND 0.0536f
C12838 VDD.n3858 GND 0.02522f
C12839 VDD.n3859 GND 0.04999f
C12840 VDD.n3860 GND 0.5126f
C12841 VDD.n3861 GND 0.02522f
C12842 VDD.n3862 GND 0.04999f
C12843 VDD.n3863 GND 0.5126f
C12844 VDD.n3864 GND 0.04999f
C12845 VDD.n3865 GND 0.05074f
C12846 VDD.n3866 GND 0.06295f
C12847 VDD.n3867 GND 0.0536f
C12848 VDD.n3868 GND 0.02522f
C12849 VDD.n3869 GND 0.04999f
C12850 VDD.n3870 GND 0.68843f
C12851 VDD.n3871 GND 0.68843f
C12852 VDD.n3872 GND 0.04999f
C12853 VDD.n3873 GND 0.02746f
C12854 VDD.n3874 GND 0.02967f
C12855 VDD.n3875 GND 0.02746f
C12856 VDD.n3876 GND 0.04999f
C12857 VDD.n3877 GND 0.68843f
C12858 VDD.n3878 GND 0.68843f
C12859 VDD.n3879 GND 0.04999f
C12860 VDD.n3880 GND 0.04999f
C12861 VDD.n3881 GND 0.02522f
C12862 VDD.n3882 GND 0.02522f
C12863 VDD.n3883 GND 0.02967f
C12864 VDD.n3884 GND 0.05074f
C12865 VDD.t231 GND 0.63568f
C12866 VDD.n3885 GND 0.05074f
C12867 VDD.n3886 GND 0.06295f
C12868 VDD.n3887 GND 0.02334f
C12869 VDD.n3888 GND 0.04152f
C12870 VDD.n3889 GND 0.03056f
C12871 VDD.n3890 GND 0.06295f
C12872 VDD.n3891 GND 0.0536f
C12873 VDD.n3892 GND 0.02522f
C12874 VDD.n3893 GND 0.04999f
C12875 VDD.n3894 GND 0.5126f
C12876 VDD.n3895 GND 0.02522f
C12877 VDD.n3896 GND 0.04999f
C12878 VDD.n3897 GND 0.5126f
C12879 VDD.n3898 GND 0.04999f
C12880 VDD.n3899 GND 0.05074f
C12881 VDD.n3900 GND 0.06295f
C12882 VDD.n3901 GND 0.0536f
C12883 VDD.n3902 GND 0.02522f
C12884 VDD.n3903 GND 0.04999f
C12885 VDD.n3904 GND 0.68843f
C12886 VDD.n3905 GND 0.02522f
C12887 VDD.n3906 GND 0.04999f
C12888 VDD.n3907 GND 0.68843f
C12889 VDD.n3908 GND 0.04999f
C12890 VDD.n3909 GND 0.05074f
C12891 VDD.n3910 GND 0.06295f
C12892 VDD.n3911 GND 0.0536f
C12893 VDD.n3912 GND 0.02522f
C12894 VDD.n3913 GND 0.04999f
C12895 VDD.n3914 GND 0.5126f
C12896 VDD.n3915 GND 0.02522f
C12897 VDD.n3916 GND 0.04999f
C12898 VDD.n3917 GND 0.5126f
C12899 VDD.n3918 GND 0.04999f
C12900 VDD.n3919 GND 0.05074f
C12901 VDD.n3920 GND 0.06295f
C12902 VDD.n3921 GND 0.0536f
C12903 VDD.n3922 GND 0.02522f
C12904 VDD.n3923 GND 0.04999f
C12905 VDD.n3924 GND 0.5126f
C12906 VDD.n3925 GND 0.02522f
C12907 VDD.n3926 GND 0.04999f
C12908 VDD.n3927 GND 0.5126f
C12909 VDD.n3928 GND 0.04999f
C12910 VDD.n3929 GND 0.05074f
C12911 VDD.n3930 GND 0.06295f
C12912 VDD.n3931 GND 0.0536f
C12913 VDD.n3932 GND 0.02522f
C12914 VDD.n3933 GND 0.04999f
C12915 VDD.n3934 GND 0.68843f
C12916 VDD.n3935 GND 0.68843f
C12917 VDD.n3936 GND 0.04999f
C12918 VDD.n3937 GND 0.02746f
C12919 VDD.n3938 GND 0.09132f
C12920 VDD.n3939 GND 0.01798f
C12921 VDD.n3940 GND 0.1514f
C12922 VDD.n3941 GND 0.02334f
C12923 VDD.n3942 GND 0.0536f
C12924 VDD.n3943 GND 0.05074f
C12925 VDD.n3944 GND 0.02967f
C12926 VDD.n3945 GND 0.02522f
C12927 VDD.n3946 GND 0.02522f
C12928 VDD.n3947 GND 0.04999f
C12929 VDD.n3948 GND 0.68843f
C12930 VDD.n3949 GND 0.04999f
C12931 VDD.n3950 GND 0.05074f
C12932 VDD.n3951 GND 0.06295f
C12933 VDD.n3952 GND 0.0536f
C12934 VDD.n3953 GND 0.02522f
C12935 VDD.n3954 GND 0.04999f
C12936 VDD.n3955 GND 0.5126f
C12937 VDD.n3956 GND 0.02522f
C12938 VDD.n3957 GND 0.04999f
C12939 VDD.n3958 GND 0.5126f
C12940 VDD.n3959 GND 0.04999f
C12941 VDD.n3960 GND 0.05074f
C12942 VDD.n3961 GND 0.06295f
C12943 VDD.n3962 GND 0.0536f
C12944 VDD.n3963 GND 0.02522f
C12945 VDD.n3964 GND 0.04999f
C12946 VDD.n3965 GND 0.5126f
C12947 VDD.n3966 GND 0.02522f
C12948 VDD.n3967 GND 0.04999f
C12949 VDD.n3968 GND 0.5126f
C12950 VDD.n3969 GND 0.04999f
C12951 VDD.n3970 GND 0.05074f
C12952 VDD.n3971 GND 0.06295f
C12953 VDD.n3972 GND 0.0536f
C12954 VDD.n3973 GND 0.02522f
C12955 VDD.n3974 GND 0.04999f
C12956 VDD.n3975 GND 0.68843f
C12957 VDD.n3976 GND 0.02522f
C12958 VDD.n3977 GND 0.04999f
C12959 VDD.n3978 GND 0.68843f
C12960 VDD.n3979 GND 0.04999f
C12961 VDD.n3980 GND 0.05074f
C12962 VDD.n3981 GND 0.06295f
C12963 VDD.n3982 GND 0.0536f
C12964 VDD.n3983 GND 0.02522f
C12965 VDD.n3984 GND 0.04999f
C12966 VDD.n3985 GND 0.5126f
C12967 VDD.n3986 GND 0.02522f
C12968 VDD.n3987 GND 0.04999f
C12969 VDD.n3988 GND 0.5126f
C12970 VDD.n3989 GND 0.04999f
C12971 VDD.n3990 GND 0.05074f
C12972 VDD.n3991 GND 0.06295f
C12973 VDD.n3992 GND 0.0536f
C12974 VDD.n3993 GND 0.02522f
C12975 VDD.n3994 GND 0.04999f
C12976 VDD.n3995 GND 0.68843f
C12977 VDD.n3996 GND 0.68843f
C12978 VDD.n3997 GND 0.04999f
C12979 VDD.n3998 GND 0.02746f
C12980 VDD.n3999 GND 0.02967f
C12981 VDD.n4000 GND 0.02746f
C12982 VDD.n4001 GND 0.04999f
C12983 VDD.n4002 GND 0.68843f
C12984 VDD.n4003 GND 0.68843f
C12985 VDD.n4004 GND 0.04999f
C12986 VDD.n4005 GND 0.04999f
C12987 VDD.n4006 GND 0.02522f
C12988 VDD.n4007 GND 0.02522f
C12989 VDD.n4008 GND 0.02967f
C12990 VDD.n4009 GND 0.05074f
C12991 VDD.t310 GND 0.63568f
C12992 VDD.n4010 GND 0.05074f
C12993 VDD.n4011 GND 0.06295f
C12994 VDD.n4012 GND 0.02334f
C12995 VDD.n4013 GND 0.04152f
C12996 VDD.n4014 GND 0.03056f
C12997 VDD.n4015 GND 0.06295f
C12998 VDD.n4016 GND 0.0536f
C12999 VDD.n4017 GND 0.02522f
C13000 VDD.n4018 GND 0.04999f
C13001 VDD.n4019 GND 0.5126f
C13002 VDD.n4020 GND 0.02522f
C13003 VDD.n4021 GND 0.04999f
C13004 VDD.n4022 GND 0.5126f
C13005 VDD.n4023 GND 0.04999f
C13006 VDD.n4024 GND 0.05074f
C13007 VDD.n4025 GND 0.06295f
C13008 VDD.n4026 GND 0.0536f
C13009 VDD.n4027 GND 0.02522f
C13010 VDD.n4028 GND 0.04999f
C13011 VDD.n4029 GND 0.68843f
C13012 VDD.n4030 GND 0.02522f
C13013 VDD.n4031 GND 0.04999f
C13014 VDD.n4032 GND 0.68843f
C13015 VDD.n4033 GND 0.04999f
C13016 VDD.n4034 GND 0.05074f
C13017 VDD.n4035 GND 0.06295f
C13018 VDD.n4036 GND 0.0536f
C13019 VDD.n4037 GND 0.02522f
C13020 VDD.n4038 GND 0.04999f
C13021 VDD.n4039 GND 0.5126f
C13022 VDD.n4040 GND 0.02522f
C13023 VDD.n4041 GND 0.04999f
C13024 VDD.n4042 GND 0.5126f
C13025 VDD.n4043 GND 0.04999f
C13026 VDD.n4044 GND 0.05074f
C13027 VDD.n4045 GND 0.06295f
C13028 VDD.n4046 GND 0.0536f
C13029 VDD.n4047 GND 0.02522f
C13030 VDD.n4048 GND 0.04999f
C13031 VDD.n4049 GND 0.5126f
C13032 VDD.n4050 GND 0.02522f
C13033 VDD.n4051 GND 0.04999f
C13034 VDD.n4052 GND 0.5126f
C13035 VDD.n4053 GND 0.04999f
C13036 VDD.n4054 GND 0.05074f
C13037 VDD.n4055 GND 0.06295f
C13038 VDD.n4056 GND 0.0536f
C13039 VDD.n4057 GND 0.02522f
C13040 VDD.n4058 GND 0.04999f
C13041 VDD.n4059 GND 0.68843f
C13042 VDD.n4060 GND 0.68843f
C13043 VDD.n4061 GND 0.04999f
C13044 VDD.n4062 GND 0.02746f
C13045 VDD.n4063 GND 0.09132f
C13046 VDD.n4064 GND 0.01798f
C13047 VDD.n4065 GND 0.1514f
C13048 VDD.n4066 GND 0.02334f
C13049 VDD.n4067 GND 0.0536f
C13050 VDD.n4068 GND 0.05074f
C13051 VDD.n4069 GND 0.02967f
C13052 VDD.n4070 GND 0.02522f
C13053 VDD.n4071 GND 0.02522f
C13054 VDD.n4072 GND 0.04999f
C13055 VDD.n4073 GND 0.68843f
C13056 VDD.n4074 GND 0.04999f
C13057 VDD.n4075 GND 0.05074f
C13058 VDD.n4076 GND 0.06295f
C13059 VDD.n4077 GND 0.0536f
C13060 VDD.n4078 GND 0.02522f
C13061 VDD.n4079 GND 0.04999f
C13062 VDD.n4080 GND 0.5126f
C13063 VDD.n4081 GND 0.02522f
C13064 VDD.n4082 GND 0.04999f
C13065 VDD.n4083 GND 0.5126f
C13066 VDD.n4084 GND 0.04999f
C13067 VDD.n4085 GND 0.05074f
C13068 VDD.n4086 GND 0.06295f
C13069 VDD.n4087 GND 0.0536f
C13070 VDD.n4088 GND 0.02522f
C13071 VDD.n4089 GND 0.04999f
C13072 VDD.n4090 GND 0.5126f
C13073 VDD.n4091 GND 0.02522f
C13074 VDD.n4092 GND 0.04999f
C13075 VDD.n4093 GND 0.5126f
C13076 VDD.n4094 GND 0.04999f
C13077 VDD.n4095 GND 0.05074f
C13078 VDD.n4096 GND 0.06295f
C13079 VDD.n4097 GND 0.0536f
C13080 VDD.n4098 GND 0.02522f
C13081 VDD.n4099 GND 0.04999f
C13082 VDD.n4100 GND 0.68843f
C13083 VDD.n4101 GND 0.02522f
C13084 VDD.n4102 GND 0.04999f
C13085 VDD.n4103 GND 0.68843f
C13086 VDD.n4104 GND 0.04999f
C13087 VDD.n4105 GND 0.05074f
C13088 VDD.n4106 GND 0.06295f
C13089 VDD.n4107 GND 0.0536f
C13090 VDD.n4108 GND 0.02522f
C13091 VDD.n4109 GND 0.04999f
C13092 VDD.n4110 GND 0.5126f
C13093 VDD.n4111 GND 0.02522f
C13094 VDD.n4112 GND 0.04999f
C13095 VDD.n4113 GND 0.5126f
C13096 VDD.n4114 GND 0.04999f
C13097 VDD.n4115 GND 0.05074f
C13098 VDD.n4116 GND 0.06295f
C13099 VDD.n4117 GND 0.0536f
C13100 VDD.n4118 GND 0.02522f
C13101 VDD.n4119 GND 0.04999f
C13102 VDD.n4120 GND 0.68843f
C13103 VDD.n4121 GND 0.68843f
C13104 VDD.n4122 GND 0.04999f
C13105 VDD.n4123 GND 0.02746f
C13106 VDD.n4124 GND 0.02967f
C13107 VDD.n4125 GND 0.02746f
C13108 VDD.n4126 GND 0.04999f
C13109 VDD.n4127 GND 0.68843f
C13110 VDD.n4128 GND 0.68843f
C13111 VDD.n4129 GND 0.04999f
C13112 VDD.n4130 GND 0.04999f
C13113 VDD.n4131 GND 0.02522f
C13114 VDD.n4132 GND 0.02522f
C13115 VDD.n4133 GND 0.02967f
C13116 VDD.n4134 GND 0.05074f
C13117 VDD.t80 GND 0.63568f
C13118 VDD.n4135 GND 0.05074f
C13119 VDD.n4136 GND 0.06295f
C13120 VDD.n4137 GND 0.02334f
C13121 VDD.n4138 GND 0.04152f
C13122 VDD.n4139 GND 0.03056f
C13123 VDD.n4140 GND 0.06295f
C13124 VDD.n4141 GND 0.0536f
C13125 VDD.n4142 GND 0.02522f
C13126 VDD.n4143 GND 0.04999f
C13127 VDD.n4144 GND 0.5126f
C13128 VDD.n4145 GND 0.02522f
C13129 VDD.n4146 GND 0.04999f
C13130 VDD.n4147 GND 0.5126f
C13131 VDD.n4148 GND 0.04999f
C13132 VDD.n4149 GND 0.05074f
C13133 VDD.n4150 GND 0.06295f
C13134 VDD.n4151 GND 0.0536f
C13135 VDD.n4152 GND 0.02522f
C13136 VDD.n4153 GND 0.04999f
C13137 VDD.n4154 GND 0.68843f
C13138 VDD.n4155 GND 0.02522f
C13139 VDD.n4156 GND 0.04999f
C13140 VDD.n4157 GND 0.68843f
C13141 VDD.n4158 GND 0.04999f
C13142 VDD.n4159 GND 0.05074f
C13143 VDD.n4160 GND 0.06295f
C13144 VDD.n4161 GND 0.0536f
C13145 VDD.n4162 GND 0.02522f
C13146 VDD.n4163 GND 0.04999f
C13147 VDD.n4164 GND 0.5126f
C13148 VDD.n4165 GND 0.02522f
C13149 VDD.n4166 GND 0.04999f
C13150 VDD.n4167 GND 0.5126f
C13151 VDD.n4168 GND 0.04999f
C13152 VDD.n4169 GND 0.05074f
C13153 VDD.n4170 GND 0.06295f
C13154 VDD.n4171 GND 0.0536f
C13155 VDD.n4172 GND 0.02522f
C13156 VDD.n4173 GND 0.04999f
C13157 VDD.n4174 GND 0.5126f
C13158 VDD.n4175 GND 0.02522f
C13159 VDD.n4176 GND 0.04999f
C13160 VDD.n4177 GND 0.5126f
C13161 VDD.n4178 GND 0.04999f
C13162 VDD.n4179 GND 0.05074f
C13163 VDD.n4180 GND 0.06295f
C13164 VDD.n4181 GND 0.0536f
C13165 VDD.n4182 GND 0.02522f
C13166 VDD.n4183 GND 0.04999f
C13167 VDD.n4184 GND 0.68843f
C13168 VDD.n4185 GND 0.68843f
C13169 VDD.n4186 GND 0.04999f
C13170 VDD.n4187 GND 0.02746f
C13171 VDD.n4188 GND 0.09132f
C13172 VDD.n4189 GND 0.01798f
C13173 VDD.n4190 GND 0.1514f
C13174 VDD.n4191 GND 0.02334f
C13175 VDD.n4192 GND 0.0536f
C13176 VDD.n4193 GND 0.05074f
C13177 VDD.n4194 GND 0.02967f
C13178 VDD.n4195 GND 0.02522f
C13179 VDD.n4196 GND 0.02522f
C13180 VDD.n4197 GND 0.04999f
C13181 VDD.n4198 GND 0.68843f
C13182 VDD.n4199 GND 0.04999f
C13183 VDD.n4200 GND 0.05074f
C13184 VDD.n4201 GND 0.06295f
C13185 VDD.n4202 GND 0.0536f
C13186 VDD.n4203 GND 0.02522f
C13187 VDD.n4204 GND 0.04999f
C13188 VDD.n4205 GND 0.5126f
C13189 VDD.n4206 GND 0.02522f
C13190 VDD.n4207 GND 0.04999f
C13191 VDD.n4208 GND 0.5126f
C13192 VDD.n4209 GND 0.04999f
C13193 VDD.n4210 GND 0.05074f
C13194 VDD.n4211 GND 0.06295f
C13195 VDD.n4212 GND 0.0536f
C13196 VDD.n4213 GND 0.02522f
C13197 VDD.n4214 GND 0.04999f
C13198 VDD.n4215 GND 0.5126f
C13199 VDD.n4216 GND 0.02522f
C13200 VDD.n4217 GND 0.04999f
C13201 VDD.n4218 GND 0.5126f
C13202 VDD.n4219 GND 0.04999f
C13203 VDD.n4220 GND 0.05074f
C13204 VDD.n4221 GND 0.06295f
C13205 VDD.n4222 GND 0.0536f
C13206 VDD.n4223 GND 0.02522f
C13207 VDD.n4224 GND 0.04999f
C13208 VDD.n4225 GND 0.68843f
C13209 VDD.n4226 GND 0.02522f
C13210 VDD.n4227 GND 0.04999f
C13211 VDD.n4228 GND 0.68843f
C13212 VDD.n4229 GND 0.04999f
C13213 VDD.n4230 GND 0.05074f
C13214 VDD.n4231 GND 0.06295f
C13215 VDD.n4232 GND 0.0536f
C13216 VDD.n4233 GND 0.02522f
C13217 VDD.n4234 GND 0.04999f
C13218 VDD.n4235 GND 0.5126f
C13219 VDD.n4236 GND 0.02522f
C13220 VDD.n4237 GND 0.04999f
C13221 VDD.n4238 GND 0.5126f
C13222 VDD.n4239 GND 0.04999f
C13223 VDD.n4240 GND 0.05074f
C13224 VDD.n4241 GND 0.06295f
C13225 VDD.n4242 GND 0.0536f
C13226 VDD.n4243 GND 0.02522f
C13227 VDD.n4244 GND 0.04999f
C13228 VDD.n4245 GND 0.68843f
C13229 VDD.n4246 GND 0.68843f
C13230 VDD.n4247 GND 0.04999f
C13231 VDD.n4248 GND 0.02746f
C13232 VDD.n4249 GND 0.02967f
C13233 VDD.n4250 GND 0.02746f
C13234 VDD.n4251 GND 0.04999f
C13235 VDD.n4252 GND 0.68843f
C13236 VDD.n4253 GND 0.68843f
C13237 VDD.n4254 GND 0.04999f
C13238 VDD.n4255 GND 0.04999f
C13239 VDD.n4256 GND 0.02522f
C13240 VDD.n4257 GND 0.02522f
C13241 VDD.n4258 GND 0.02967f
C13242 VDD.n4259 GND 0.05074f
C13243 VDD.t386 GND 0.63568f
C13244 VDD.n4260 GND 0.05074f
C13245 VDD.n4261 GND 0.06295f
C13246 VDD.n4262 GND 0.02334f
C13247 VDD.n4263 GND 0.04152f
C13248 VDD.n4264 GND 0.03056f
C13249 VDD.n4265 GND 0.06295f
C13250 VDD.n4266 GND 0.0536f
C13251 VDD.n4267 GND 0.02522f
C13252 VDD.n4268 GND 0.04999f
C13253 VDD.n4269 GND 0.5126f
C13254 VDD.n4270 GND 0.02522f
C13255 VDD.n4271 GND 0.04999f
C13256 VDD.n4272 GND 0.5126f
C13257 VDD.n4273 GND 0.04999f
C13258 VDD.n4274 GND 0.05074f
C13259 VDD.n4275 GND 0.06295f
C13260 VDD.n4276 GND 0.0536f
C13261 VDD.n4277 GND 0.02522f
C13262 VDD.n4278 GND 0.04999f
C13263 VDD.n4279 GND 0.68843f
C13264 VDD.n4280 GND 0.02522f
C13265 VDD.n4281 GND 0.04999f
C13266 VDD.n4282 GND 0.68843f
C13267 VDD.n4283 GND 0.04999f
C13268 VDD.n4284 GND 0.05074f
C13269 VDD.n4285 GND 0.06295f
C13270 VDD.n4286 GND 0.0536f
C13271 VDD.n4287 GND 0.02522f
C13272 VDD.n4288 GND 0.04999f
C13273 VDD.n4289 GND 0.5126f
C13274 VDD.n4290 GND 0.02522f
C13275 VDD.n4291 GND 0.04999f
C13276 VDD.n4292 GND 0.5126f
C13277 VDD.n4293 GND 0.04999f
C13278 VDD.n4294 GND 0.05074f
C13279 VDD.n4295 GND 0.06295f
C13280 VDD.n4296 GND 0.0536f
C13281 VDD.n4297 GND 0.02522f
C13282 VDD.n4298 GND 0.04999f
C13283 VDD.n4299 GND 0.5126f
C13284 VDD.n4300 GND 0.02522f
C13285 VDD.n4301 GND 0.04999f
C13286 VDD.n4302 GND 0.5126f
C13287 VDD.n4303 GND 0.04999f
C13288 VDD.n4304 GND 0.05074f
C13289 VDD.n4305 GND 0.06295f
C13290 VDD.n4306 GND 0.0536f
C13291 VDD.n4307 GND 0.02522f
C13292 VDD.n4308 GND 0.04999f
C13293 VDD.n4309 GND 0.68843f
C13294 VDD.n4310 GND 0.68843f
C13295 VDD.n4311 GND 0.04999f
C13296 VDD.n4312 GND 0.02746f
C13297 VDD.n4313 GND 0.09132f
C13298 VDD.n4314 GND 0.01798f
C13299 VDD.n4315 GND 0.1514f
C13300 VDD.n4316 GND 0.02334f
C13301 VDD.n4317 GND 0.0536f
C13302 VDD.n4318 GND 0.05074f
C13303 VDD.n4319 GND 0.02967f
C13304 VDD.n4320 GND 0.02522f
C13305 VDD.n4321 GND 0.02522f
C13306 VDD.n4322 GND 0.04999f
C13307 VDD.n4323 GND 0.68843f
C13308 VDD.n4324 GND 0.04999f
C13309 VDD.n4325 GND 0.05074f
C13310 VDD.n4326 GND 0.06295f
C13311 VDD.n4327 GND 0.0536f
C13312 VDD.n4328 GND 0.02522f
C13313 VDD.n4329 GND 0.04999f
C13314 VDD.n4330 GND 0.5126f
C13315 VDD.n4331 GND 0.02522f
C13316 VDD.n4332 GND 0.04999f
C13317 VDD.n4333 GND 0.5126f
C13318 VDD.n4334 GND 0.04999f
C13319 VDD.n4335 GND 0.05074f
C13320 VDD.n4336 GND 0.06295f
C13321 VDD.n4337 GND 0.0536f
C13322 VDD.n4338 GND 0.02522f
C13323 VDD.n4339 GND 0.04999f
C13324 VDD.n4340 GND 0.5126f
C13325 VDD.n4341 GND 0.02522f
C13326 VDD.n4342 GND 0.04999f
C13327 VDD.n4343 GND 0.5126f
C13328 VDD.n4344 GND 0.04999f
C13329 VDD.n4345 GND 0.05074f
C13330 VDD.n4346 GND 0.06295f
C13331 VDD.n4347 GND 0.0536f
C13332 VDD.n4348 GND 0.02522f
C13333 VDD.n4349 GND 0.04999f
C13334 VDD.n4350 GND 0.68843f
C13335 VDD.n4351 GND 0.02522f
C13336 VDD.n4352 GND 0.04999f
C13337 VDD.n4353 GND 0.68843f
C13338 VDD.n4354 GND 0.04999f
C13339 VDD.n4355 GND 0.05074f
C13340 VDD.n4356 GND 0.06295f
C13341 VDD.n4357 GND 0.0536f
C13342 VDD.n4358 GND 0.02522f
C13343 VDD.n4359 GND 0.04999f
C13344 VDD.n4360 GND 0.5126f
C13345 VDD.n4361 GND 0.02522f
C13346 VDD.n4362 GND 0.04999f
C13347 VDD.n4363 GND 0.5126f
C13348 VDD.n4364 GND 0.04999f
C13349 VDD.n4365 GND 0.05074f
C13350 VDD.n4366 GND 0.06295f
C13351 VDD.n4367 GND 0.0536f
C13352 VDD.n4368 GND 0.02522f
C13353 VDD.n4369 GND 0.04999f
C13354 VDD.n4370 GND 0.68843f
C13355 VDD.n4371 GND 0.68843f
C13356 VDD.n4372 GND 0.04999f
C13357 VDD.n4373 GND 0.02746f
C13358 VDD.n4374 GND 0.02967f
C13359 VDD.n4375 GND 0.02746f
C13360 VDD.n4376 GND 0.04999f
C13361 VDD.n4377 GND 0.68843f
C13362 VDD.n4378 GND 0.68843f
C13363 VDD.n4379 GND 0.04999f
C13364 VDD.n4380 GND 0.04999f
C13365 VDD.n4381 GND 0.02522f
C13366 VDD.n4382 GND 0.02522f
C13367 VDD.n4383 GND 0.02967f
C13368 VDD.n4384 GND 0.05074f
C13369 VDD.t19 GND 0.63568f
C13370 VDD.n4385 GND 0.05074f
C13371 VDD.n4386 GND 0.06295f
C13372 VDD.n4387 GND 0.02334f
C13373 VDD.n4388 GND 0.04152f
C13374 VDD.n4389 GND 0.03056f
C13375 VDD.n4390 GND 0.06295f
C13376 VDD.n4391 GND 0.0536f
C13377 VDD.n4392 GND 0.02522f
C13378 VDD.n4393 GND 0.04999f
C13379 VDD.n4394 GND 0.5126f
C13380 VDD.n4395 GND 0.02522f
C13381 VDD.n4396 GND 0.04999f
C13382 VDD.n4397 GND 0.5126f
C13383 VDD.n4398 GND 0.04999f
C13384 VDD.n4399 GND 0.05074f
C13385 VDD.n4400 GND 0.06295f
C13386 VDD.n4401 GND 0.0536f
C13387 VDD.n4402 GND 0.02522f
C13388 VDD.n4403 GND 0.04999f
C13389 VDD.n4404 GND 0.68843f
C13390 VDD.n4405 GND 0.02522f
C13391 VDD.n4406 GND 0.04999f
C13392 VDD.n4407 GND 0.68843f
C13393 VDD.n4408 GND 0.04999f
C13394 VDD.n4409 GND 0.05074f
C13395 VDD.n4410 GND 0.06295f
C13396 VDD.n4411 GND 0.0536f
C13397 VDD.n4412 GND 0.02522f
C13398 VDD.n4413 GND 0.04999f
C13399 VDD.n4414 GND 0.5126f
C13400 VDD.n4415 GND 0.02522f
C13401 VDD.n4416 GND 0.04999f
C13402 VDD.n4417 GND 0.5126f
C13403 VDD.n4418 GND 0.04999f
C13404 VDD.n4419 GND 0.05074f
C13405 VDD.n4420 GND 0.06295f
C13406 VDD.n4421 GND 0.0536f
C13407 VDD.n4422 GND 0.02522f
C13408 VDD.n4423 GND 0.04999f
C13409 VDD.n4424 GND 0.5126f
C13410 VDD.n4425 GND 0.02522f
C13411 VDD.n4426 GND 0.04999f
C13412 VDD.n4427 GND 0.5126f
C13413 VDD.n4428 GND 0.04999f
C13414 VDD.n4429 GND 0.05074f
C13415 VDD.n4430 GND 0.06295f
C13416 VDD.n4431 GND 0.0536f
C13417 VDD.n4432 GND 0.02522f
C13418 VDD.n4433 GND 0.04999f
C13419 VDD.n4434 GND 0.68843f
C13420 VDD.n4435 GND 0.68843f
C13421 VDD.n4436 GND 0.04999f
C13422 VDD.n4437 GND 0.02746f
C13423 VDD.n4438 GND 0.09132f
C13424 VDD.n4439 GND 0.01798f
C13425 VDD.n4440 GND 0.1514f
C13426 VDD.n4441 GND 0.02334f
C13427 VDD.n4442 GND 0.0536f
C13428 VDD.n4443 GND 0.05074f
C13429 VDD.n4444 GND 0.02967f
C13430 VDD.n4445 GND 0.02522f
C13431 VDD.n4446 GND 0.02522f
C13432 VDD.n4447 GND 0.04999f
C13433 VDD.n4448 GND 0.68843f
C13434 VDD.n4449 GND 0.04999f
C13435 VDD.n4450 GND 0.05074f
C13436 VDD.n4451 GND 0.06295f
C13437 VDD.n4452 GND 0.0536f
C13438 VDD.n4453 GND 0.02522f
C13439 VDD.n4454 GND 0.04999f
C13440 VDD.n4455 GND 0.5126f
C13441 VDD.n4456 GND 0.02522f
C13442 VDD.n4457 GND 0.04999f
C13443 VDD.n4458 GND 0.5126f
C13444 VDD.n4459 GND 0.04999f
C13445 VDD.n4460 GND 0.05074f
C13446 VDD.n4461 GND 0.06295f
C13447 VDD.n4462 GND 0.0536f
C13448 VDD.n4463 GND 0.02522f
C13449 VDD.n4464 GND 0.04999f
C13450 VDD.n4465 GND 0.5126f
C13451 VDD.n4466 GND 0.02522f
C13452 VDD.n4467 GND 0.04999f
C13453 VDD.n4468 GND 0.5126f
C13454 VDD.n4469 GND 0.04999f
C13455 VDD.n4470 GND 0.05074f
C13456 VDD.n4471 GND 0.06295f
C13457 VDD.n4472 GND 0.0536f
C13458 VDD.n4473 GND 0.02522f
C13459 VDD.n4474 GND 0.04999f
C13460 VDD.n4475 GND 0.68843f
C13461 VDD.n4476 GND 0.02522f
C13462 VDD.n4477 GND 0.04999f
C13463 VDD.n4478 GND 0.68843f
C13464 VDD.n4479 GND 0.04999f
C13465 VDD.n4480 GND 0.05074f
C13466 VDD.n4481 GND 0.06295f
C13467 VDD.n4482 GND 0.0536f
C13468 VDD.n4483 GND 0.02522f
C13469 VDD.n4484 GND 0.04999f
C13470 VDD.n4485 GND 0.5126f
C13471 VDD.n4486 GND 0.02522f
C13472 VDD.n4487 GND 0.04999f
C13473 VDD.n4488 GND 0.5126f
C13474 VDD.n4489 GND 0.04999f
C13475 VDD.n4490 GND 0.05074f
C13476 VDD.n4491 GND 0.06295f
C13477 VDD.n4492 GND 0.0536f
C13478 VDD.n4493 GND 0.02522f
C13479 VDD.n4494 GND 0.04999f
C13480 VDD.n4495 GND 0.68843f
C13481 VDD.n4496 GND 0.68843f
C13482 VDD.n4497 GND 0.04999f
C13483 VDD.n4498 GND 0.02746f
C13484 VDD.n4499 GND 0.02967f
C13485 VDD.n4500 GND 0.02746f
C13486 VDD.n4501 GND 0.04999f
C13487 VDD.n4502 GND 0.68843f
C13488 VDD.n4503 GND 0.68843f
C13489 VDD.n4504 GND 0.04999f
C13490 VDD.n4505 GND 0.04999f
C13491 VDD.n4506 GND 0.02522f
C13492 VDD.n4507 GND 0.02522f
C13493 VDD.n4508 GND 0.02967f
C13494 VDD.n4509 GND 0.05074f
C13495 VDD.t215 GND 0.63568f
C13496 VDD.n4510 GND 0.05074f
C13497 VDD.n4511 GND 0.06295f
C13498 VDD.n4512 GND 0.02334f
C13499 VDD.n4513 GND 0.04152f
C13500 VDD.n4514 GND 0.03056f
C13501 VDD.n4515 GND 0.06295f
C13502 VDD.n4516 GND 0.0536f
C13503 VDD.n4517 GND 0.02522f
C13504 VDD.n4518 GND 0.04999f
C13505 VDD.n4519 GND 0.5126f
C13506 VDD.n4520 GND 0.02522f
C13507 VDD.n4521 GND 0.04999f
C13508 VDD.n4522 GND 0.5126f
C13509 VDD.n4523 GND 0.04999f
C13510 VDD.n4524 GND 0.05074f
C13511 VDD.n4525 GND 0.06295f
C13512 VDD.n4526 GND 0.0536f
C13513 VDD.n4527 GND 0.02522f
C13514 VDD.n4528 GND 0.04999f
C13515 VDD.n4529 GND 0.68843f
C13516 VDD.n4530 GND 0.02522f
C13517 VDD.n4531 GND 0.04999f
C13518 VDD.n4532 GND 0.68843f
C13519 VDD.n4533 GND 0.04999f
C13520 VDD.n4534 GND 0.05074f
C13521 VDD.n4535 GND 0.06295f
C13522 VDD.n4536 GND 0.0536f
C13523 VDD.n4537 GND 0.02522f
C13524 VDD.n4538 GND 0.04999f
C13525 VDD.n4539 GND 0.5126f
C13526 VDD.n4540 GND 0.02522f
C13527 VDD.n4541 GND 0.04999f
C13528 VDD.n4542 GND 0.5126f
C13529 VDD.n4543 GND 0.04999f
C13530 VDD.n4544 GND 0.05074f
C13531 VDD.n4545 GND 0.06295f
C13532 VDD.n4546 GND 0.0536f
C13533 VDD.n4547 GND 0.02522f
C13534 VDD.n4548 GND 0.04999f
C13535 VDD.n4549 GND 0.5126f
C13536 VDD.n4550 GND 0.02522f
C13537 VDD.n4551 GND 0.04999f
C13538 VDD.n4552 GND 0.5126f
C13539 VDD.n4553 GND 0.04999f
C13540 VDD.n4554 GND 0.05074f
C13541 VDD.n4555 GND 0.06295f
C13542 VDD.n4556 GND 0.0536f
C13543 VDD.n4557 GND 0.02522f
C13544 VDD.n4558 GND 0.04999f
C13545 VDD.n4559 GND 0.68843f
C13546 VDD.n4560 GND 0.68843f
C13547 VDD.n4561 GND 0.04999f
C13548 VDD.n4562 GND 0.02746f
C13549 VDD.n4563 GND 0.09132f
C13550 VDD.n4564 GND 0.01798f
C13551 VDD.n4565 GND 0.1514f
C13552 VDD.n4566 GND 0.02334f
C13553 VDD.n4567 GND 0.0536f
C13554 VDD.n4568 GND 0.05074f
C13555 VDD.n4569 GND 0.02967f
C13556 VDD.n4570 GND 0.02522f
C13557 VDD.n4571 GND 0.02522f
C13558 VDD.n4572 GND 0.04999f
C13559 VDD.n4573 GND 0.68843f
C13560 VDD.n4574 GND 0.04999f
C13561 VDD.n4575 GND 0.05074f
C13562 VDD.n4576 GND 0.06295f
C13563 VDD.n4577 GND 0.0536f
C13564 VDD.n4578 GND 0.02522f
C13565 VDD.n4579 GND 0.04999f
C13566 VDD.n4580 GND 0.5126f
C13567 VDD.n4581 GND 0.02522f
C13568 VDD.n4582 GND 0.04999f
C13569 VDD.n4583 GND 0.5126f
C13570 VDD.n4584 GND 0.04999f
C13571 VDD.n4585 GND 0.05074f
C13572 VDD.n4586 GND 0.06295f
C13573 VDD.n4587 GND 0.0536f
C13574 VDD.n4588 GND 0.02522f
C13575 VDD.n4589 GND 0.04999f
C13576 VDD.n4590 GND 0.5126f
C13577 VDD.n4591 GND 0.02522f
C13578 VDD.n4592 GND 0.04999f
C13579 VDD.n4593 GND 0.5126f
C13580 VDD.n4594 GND 0.04999f
C13581 VDD.n4595 GND 0.05074f
C13582 VDD.n4596 GND 0.06295f
C13583 VDD.n4597 GND 0.0536f
C13584 VDD.n4598 GND 0.02522f
C13585 VDD.n4599 GND 0.04999f
C13586 VDD.n4600 GND 0.68843f
C13587 VDD.n4601 GND 0.02522f
C13588 VDD.n4602 GND 0.04999f
C13589 VDD.n4603 GND 0.68843f
C13590 VDD.n4604 GND 0.04999f
C13591 VDD.n4605 GND 0.05074f
C13592 VDD.n4606 GND 0.06295f
C13593 VDD.n4607 GND 0.0536f
C13594 VDD.n4608 GND 0.02522f
C13595 VDD.n4609 GND 0.04999f
C13596 VDD.n4610 GND 0.5126f
C13597 VDD.n4611 GND 0.02522f
C13598 VDD.n4612 GND 0.04999f
C13599 VDD.n4613 GND 0.5126f
C13600 VDD.n4614 GND 0.04999f
C13601 VDD.n4615 GND 0.05074f
C13602 VDD.n4616 GND 0.06295f
C13603 VDD.n4617 GND 0.0536f
C13604 VDD.n4618 GND 0.02522f
C13605 VDD.n4619 GND 0.04999f
C13606 VDD.n4620 GND 0.68843f
C13607 VDD.n4621 GND 0.68843f
C13608 VDD.n4622 GND 0.04999f
C13609 VDD.n4623 GND 0.02746f
C13610 VDD.n4624 GND 0.02967f
C13611 VDD.n4625 GND 0.02746f
C13612 VDD.n4626 GND 0.04999f
C13613 VDD.n4627 GND 0.68843f
C13614 VDD.n4628 GND 0.68843f
C13615 VDD.n4629 GND 0.04999f
C13616 VDD.n4630 GND 0.04999f
C13617 VDD.n4631 GND 0.02522f
C13618 VDD.n4632 GND 0.02522f
C13619 VDD.n4633 GND 0.02967f
C13620 VDD.n4634 GND 0.05074f
C13621 VDD.t95 GND 0.63568f
C13622 VDD.n4635 GND 0.05074f
C13623 VDD.n4636 GND 0.06295f
C13624 VDD.n4637 GND 0.02334f
C13625 VDD.n4638 GND 0.04152f
C13626 VDD.n4639 GND 0.03056f
C13627 VDD.n4640 GND 0.06295f
C13628 VDD.n4641 GND 0.0536f
C13629 VDD.n4642 GND 0.02522f
C13630 VDD.n4643 GND 0.04999f
C13631 VDD.n4644 GND 0.5126f
C13632 VDD.n4645 GND 0.02522f
C13633 VDD.n4646 GND 0.04999f
C13634 VDD.n4647 GND 0.5126f
C13635 VDD.n4648 GND 0.04999f
C13636 VDD.n4649 GND 0.05074f
C13637 VDD.n4650 GND 0.06295f
C13638 VDD.n4651 GND 0.0536f
C13639 VDD.n4652 GND 0.02522f
C13640 VDD.n4653 GND 0.04999f
C13641 VDD.n4654 GND 0.68843f
C13642 VDD.n4655 GND 0.02522f
C13643 VDD.n4656 GND 0.04999f
C13644 VDD.n4657 GND 0.68843f
C13645 VDD.n4658 GND 0.04999f
C13646 VDD.n4659 GND 0.05074f
C13647 VDD.n4660 GND 0.06295f
C13648 VDD.n4661 GND 0.0536f
C13649 VDD.n4662 GND 0.02522f
C13650 VDD.n4663 GND 0.04999f
C13651 VDD.n4664 GND 0.5126f
C13652 VDD.n4665 GND 0.02522f
C13653 VDD.n4666 GND 0.04999f
C13654 VDD.n4667 GND 0.5126f
C13655 VDD.n4668 GND 0.04999f
C13656 VDD.n4669 GND 0.05074f
C13657 VDD.n4670 GND 0.06295f
C13658 VDD.n4671 GND 0.0536f
C13659 VDD.n4672 GND 0.02522f
C13660 VDD.n4673 GND 0.04999f
C13661 VDD.n4674 GND 0.5126f
C13662 VDD.n4675 GND 0.02522f
C13663 VDD.n4676 GND 0.04999f
C13664 VDD.n4677 GND 0.5126f
C13665 VDD.n4678 GND 0.04999f
C13666 VDD.n4679 GND 0.05074f
C13667 VDD.n4680 GND 0.06295f
C13668 VDD.n4681 GND 0.0536f
C13669 VDD.n4682 GND 0.02522f
C13670 VDD.n4683 GND 0.04999f
C13671 VDD.n4684 GND 0.68843f
C13672 VDD.n4685 GND 0.68843f
C13673 VDD.n4686 GND 0.04999f
C13674 VDD.n4687 GND 0.02746f
C13675 VDD.n4688 GND 0.09132f
C13676 VDD.n4689 GND 0.01798f
C13677 VDD.n4690 GND 0.1514f
C13678 VDD.n4691 GND 0.02334f
C13679 VDD.n4692 GND 0.0536f
C13680 VDD.n4693 GND 0.05074f
C13681 VDD.n4694 GND 0.02967f
C13682 VDD.n4695 GND 0.02522f
C13683 VDD.n4696 GND 0.02522f
C13684 VDD.n4697 GND 0.04999f
C13685 VDD.n4698 GND 0.68843f
C13686 VDD.n4699 GND 0.04999f
C13687 VDD.n4700 GND 0.05074f
C13688 VDD.n4701 GND 0.06295f
C13689 VDD.n4702 GND 0.0536f
C13690 VDD.n4703 GND 0.02522f
C13691 VDD.n4704 GND 0.04999f
C13692 VDD.n4705 GND 0.5126f
C13693 VDD.n4706 GND 0.02522f
C13694 VDD.n4707 GND 0.04999f
C13695 VDD.n4708 GND 0.5126f
C13696 VDD.n4709 GND 0.04999f
C13697 VDD.n4710 GND 0.05074f
C13698 VDD.n4711 GND 0.06295f
C13699 VDD.n4712 GND 0.0536f
C13700 VDD.n4713 GND 0.02522f
C13701 VDD.n4714 GND 0.04999f
C13702 VDD.n4715 GND 0.5126f
C13703 VDD.n4716 GND 0.02522f
C13704 VDD.n4717 GND 0.04999f
C13705 VDD.n4718 GND 0.5126f
C13706 VDD.n4719 GND 0.04999f
C13707 VDD.n4720 GND 0.05074f
C13708 VDD.n4721 GND 0.06295f
C13709 VDD.n4722 GND 0.0536f
C13710 VDD.n4723 GND 0.02522f
C13711 VDD.n4724 GND 0.04999f
C13712 VDD.n4725 GND 0.68843f
C13713 VDD.n4726 GND 0.02522f
C13714 VDD.n4727 GND 0.04999f
C13715 VDD.n4728 GND 0.68843f
C13716 VDD.n4729 GND 0.04999f
C13717 VDD.n4730 GND 0.05074f
C13718 VDD.n4731 GND 0.06295f
C13719 VDD.n4732 GND 0.0536f
C13720 VDD.n4733 GND 0.02522f
C13721 VDD.n4734 GND 0.04999f
C13722 VDD.n4735 GND 0.5126f
C13723 VDD.n4736 GND 0.02522f
C13724 VDD.n4737 GND 0.04999f
C13725 VDD.n4738 GND 0.5126f
C13726 VDD.n4739 GND 0.04999f
C13727 VDD.n4740 GND 0.05074f
C13728 VDD.n4741 GND 0.06295f
C13729 VDD.n4742 GND 0.0536f
C13730 VDD.n4743 GND 0.02522f
C13731 VDD.n4744 GND 0.04999f
C13732 VDD.n4745 GND 0.68843f
C13733 VDD.n4746 GND 0.68843f
C13734 VDD.n4747 GND 0.04999f
C13735 VDD.n4748 GND 0.02746f
C13736 VDD.n4749 GND 0.02967f
C13737 VDD.n4750 GND 0.02746f
C13738 VDD.n4751 GND 0.04999f
C13739 VDD.n4752 GND 0.68843f
C13740 VDD.n4753 GND 0.68843f
C13741 VDD.n4754 GND 0.04999f
C13742 VDD.n4755 GND 0.04999f
C13743 VDD.n4756 GND 0.02522f
C13744 VDD.n4757 GND 0.02522f
C13745 VDD.n4758 GND 0.02967f
C13746 VDD.n4759 GND 0.05074f
C13747 VDD.t562 GND 0.63568f
C13748 VDD.n4760 GND 0.05074f
C13749 VDD.n4761 GND 0.06295f
C13750 VDD.n4762 GND 0.02334f
C13751 VDD.n4763 GND 0.04152f
C13752 VDD.n4764 GND 0.03056f
C13753 VDD.n4765 GND 0.06295f
C13754 VDD.n4766 GND 0.0536f
C13755 VDD.n4767 GND 0.02522f
C13756 VDD.n4768 GND 0.04999f
C13757 VDD.n4769 GND 0.5126f
C13758 VDD.n4770 GND 0.02522f
C13759 VDD.n4771 GND 0.04999f
C13760 VDD.n4772 GND 0.5126f
C13761 VDD.n4773 GND 0.04999f
C13762 VDD.n4774 GND 0.05074f
C13763 VDD.n4775 GND 0.06295f
C13764 VDD.n4776 GND 0.0536f
C13765 VDD.n4777 GND 0.02522f
C13766 VDD.n4778 GND 0.04999f
C13767 VDD.n4779 GND 0.68843f
C13768 VDD.n4780 GND 0.02522f
C13769 VDD.n4781 GND 0.04999f
C13770 VDD.n4782 GND 0.68843f
C13771 VDD.n4783 GND 0.04999f
C13772 VDD.n4784 GND 0.05074f
C13773 VDD.n4785 GND 0.06295f
C13774 VDD.n4786 GND 0.0536f
C13775 VDD.n4787 GND 0.02522f
C13776 VDD.n4788 GND 0.04999f
C13777 VDD.n4789 GND 0.5126f
C13778 VDD.n4790 GND 0.02522f
C13779 VDD.n4791 GND 0.04999f
C13780 VDD.n4792 GND 0.5126f
C13781 VDD.n4793 GND 0.04999f
C13782 VDD.n4794 GND 0.05074f
C13783 VDD.n4795 GND 0.06295f
C13784 VDD.n4796 GND 0.0536f
C13785 VDD.n4797 GND 0.02522f
C13786 VDD.n4798 GND 0.04999f
C13787 VDD.n4799 GND 0.5126f
C13788 VDD.n4800 GND 0.02522f
C13789 VDD.n4801 GND 0.04999f
C13790 VDD.n4802 GND 0.5126f
C13791 VDD.n4803 GND 0.04999f
C13792 VDD.n4804 GND 0.05074f
C13793 VDD.n4805 GND 0.06295f
C13794 VDD.n4806 GND 0.0536f
C13795 VDD.n4807 GND 0.02522f
C13796 VDD.n4808 GND 0.04999f
C13797 VDD.n4809 GND 0.68843f
C13798 VDD.n4810 GND 0.68843f
C13799 VDD.n4811 GND 0.04999f
C13800 VDD.n4812 GND 0.02746f
C13801 VDD.n4813 GND 0.09132f
C13802 VDD.n4814 GND 0.01798f
C13803 VDD.n4815 GND 0.12268f
C13804 VDD.t575 GND 0.02334f
C13805 VDD.n4816 GND 0.02746f
C13806 VDD.n4817 GND 0.05074f
C13807 VDD.n4818 GND 0.02967f
C13808 VDD.n4819 GND 0.05074f
C13809 VDD.t496 GND 0.63568f
C13810 VDD.n4820 GND 0.04999f
C13811 VDD.n4821 GND 0.05074f
C13812 VDD.n4822 GND 0.05074f
C13813 VDD.n4823 GND 0.02967f
C13814 VDD.n4824 GND 0.02522f
C13815 VDD.n4825 GND 0.0536f
C13816 VDD.t693 GND 0.02334f
C13817 VDD.t497 GND 0.02334f
C13818 VDD.n4826 GND 0.13341f
C13819 VDD.n4827 GND 0.0263f
C13820 VDD.n4828 GND 0.05074f
C13821 VDD.n4829 GND 0.02967f
C13822 VDD.n4830 GND 0.02522f
C13823 VDD.t289 GND 0.63568f
C13824 VDD.n4831 GND 0.04999f
C13825 VDD.n4832 GND 0.05074f
C13826 VDD.n4833 GND 0.05074f
C13827 VDD.n4834 GND 0.02967f
C13828 VDD.n4835 GND 0.02522f
C13829 VDD.n4836 GND 0.0536f
C13830 VDD.n4837 GND 0.03166f
C13831 VDD.n4838 GND 0.05074f
C13832 VDD.n4839 GND 0.02967f
C13833 VDD.n4840 GND 0.02522f
C13834 VDD.t1004 GND 0.63568f
C13835 VDD.n4841 GND 0.04999f
C13836 VDD.n4842 GND 0.05074f
C13837 VDD.n4843 GND 0.05074f
C13838 VDD.n4844 GND 0.02967f
C13839 VDD.n4845 GND 0.02522f
C13840 VDD.n4846 GND 0.0536f
C13841 VDD.t1081 GND 0.02321f
C13842 VDD.t576 GND 0.02321f
C13843 VDD.n4847 GND 0.10855f
C13844 VDD.t1005 GND 0.02321f
C13845 VDD.t290 GND 0.02321f
C13846 VDD.n4848 GND 0.10855f
C13847 VDD.n4849 GND 0.04152f
C13848 VDD.n4850 GND 0.02334f
C13849 VDD.n4851 GND 0.05074f
C13850 VDD.n4852 GND 0.02967f
C13851 VDD.n4853 GND 0.02522f
C13852 VDD.t486 GND 0.63568f
C13853 VDD.n4854 GND 0.04999f
C13854 VDD.n4855 GND 0.05074f
C13855 VDD.n4856 GND 0.05074f
C13856 VDD.n4857 GND 0.02967f
C13857 VDD.n4858 GND 0.02522f
C13858 VDD.n4859 GND 0.0536f
C13859 VDD.t487 GND 0.02334f
C13860 VDD.t761 GND 0.02334f
C13861 VDD.n4860 GND 0.13341f
C13862 VDD.n4861 GND 0.0263f
C13863 VDD.n4862 GND 0.05074f
C13864 VDD.n4863 GND 0.02967f
C13865 VDD.n4864 GND 0.02522f
C13866 VDD.t259 GND 0.63568f
C13867 VDD.n4865 GND 0.04999f
C13868 VDD.n4866 GND 0.05074f
C13869 VDD.n4867 GND 0.05074f
C13870 VDD.n4868 GND 0.02967f
C13871 VDD.n4869 GND 0.02522f
C13872 VDD.n4870 GND 0.0536f
C13873 VDD.n4871 GND 0.03166f
C13874 VDD.n4872 GND 0.05074f
C13875 VDD.n4873 GND 0.02967f
C13876 VDD.n4874 GND 0.02522f
C13877 VDD.t84 GND 0.63568f
C13878 VDD.n4875 GND 0.04999f
C13879 VDD.n4876 GND 0.05074f
C13880 VDD.n4877 GND 0.05074f
C13881 VDD.n4878 GND 0.02967f
C13882 VDD.n4879 GND 0.02522f
C13883 VDD.n4880 GND 0.0536f
C13884 VDD.t947 GND 0.02321f
C13885 VDD.t260 GND 0.02321f
C13886 VDD.n4881 GND 0.10855f
C13887 VDD.t85 GND 0.02321f
C13888 VDD.t898 GND 0.02321f
C13889 VDD.n4882 GND 0.10855f
C13890 VDD.n4883 GND 0.04152f
C13891 VDD.n4884 GND 0.02334f
C13892 VDD.n4885 GND 0.05074f
C13893 VDD.n4886 GND 0.02967f
C13894 VDD.n4887 GND 0.02522f
C13895 VDD.t1052 GND 0.63568f
C13896 VDD.n4888 GND 0.05074f
C13897 VDD.n4889 GND 0.05074f
C13898 VDD.n4890 GND 0.09132f
C13899 VDD.t118 GND 0.63568f
C13900 VDD.n4891 GND 0.04999f
C13901 VDD.n4892 GND 0.05074f
C13902 VDD.n4893 GND 0.05074f
C13903 VDD.n4894 GND 0.02967f
C13904 VDD.n4895 GND 0.02522f
C13905 VDD.n4896 GND 0.0536f
C13906 VDD.t1053 GND 0.02334f
C13907 VDD.n4897 GND 0.0731f
C13908 VDD.n4898 GND 0.01798f
C13909 VDD.n4899 GND 0.02334f
C13910 VDD.n4900 GND 0.05074f
C13911 VDD.n4901 GND 0.02967f
C13912 VDD.n4902 GND 0.02522f
C13913 VDD.t380 GND 0.63568f
C13914 VDD.n4903 GND 0.04999f
C13915 VDD.n4904 GND 0.05074f
C13916 VDD.n4905 GND 0.05074f
C13917 VDD.n4906 GND 0.02967f
C13918 VDD.n4907 GND 0.02522f
C13919 VDD.n4908 GND 0.0536f
C13920 VDD.t381 GND 0.02321f
C13921 VDD.t119 GND 0.02321f
C13922 VDD.n4909 GND 0.10855f
C13923 VDD.t382 GND 0.02321f
C13924 VDD.t291 GND 0.02321f
C13925 VDD.n4910 GND 0.10855f
C13926 VDD.n4911 GND 0.04152f
C13927 VDD.n4912 GND 0.02334f
C13928 VDD.n4913 GND 0.05074f
C13929 VDD.n4914 GND 0.02967f
C13930 VDD.n4915 GND 0.02522f
C13931 VDD.t512 GND 0.63568f
C13932 VDD.n4916 GND 0.04999f
C13933 VDD.n4917 GND 0.05074f
C13934 VDD.n4918 GND 0.05074f
C13935 VDD.n4919 GND 0.02967f
C13936 VDD.n4920 GND 0.02522f
C13937 VDD.n4921 GND 0.0536f
C13938 VDD.t513 GND 0.02334f
C13939 VDD.t677 GND 0.02334f
C13940 VDD.n4922 GND 0.13341f
C13941 VDD.n4923 GND 0.0263f
C13942 VDD.n4924 GND 0.05074f
C13943 VDD.n4925 GND 0.02967f
C13944 VDD.n4926 GND 0.02522f
C13945 VDD.t181 GND 0.63568f
C13946 VDD.n4927 GND 0.04999f
C13947 VDD.n4928 GND 0.05074f
C13948 VDD.n4929 GND 0.05074f
C13949 VDD.n4930 GND 0.02967f
C13950 VDD.n4931 GND 0.02522f
C13951 VDD.n4932 GND 0.0536f
C13952 VDD.n4933 GND 0.03166f
C13953 VDD.n4934 GND 0.05074f
C13954 VDD.n4935 GND 0.02967f
C13955 VDD.n4936 GND 0.02522f
C13956 VDD.t183 GND 0.63568f
C13957 VDD.n4937 GND 0.04999f
C13958 VDD.n4938 GND 0.05074f
C13959 VDD.n4939 GND 0.05074f
C13960 VDD.n4940 GND 0.02967f
C13961 VDD.n4941 GND 0.02522f
C13962 VDD.n4942 GND 0.0536f
C13963 VDD.n4943 GND 0.05074f
C13964 VDD.n4944 GND 0.02967f
C13965 VDD.n4945 GND 0.02522f
C13966 VDD.n4946 GND 0.02522f
C13967 VDD.n4947 GND 0.04999f
C13968 VDD.n4948 GND 0.68843f
C13969 VDD.n4949 GND 0.04999f
C13970 VDD.n4950 GND 0.05074f
C13971 VDD.t184 GND 0.02321f
C13972 VDD.t182 GND 0.02321f
C13973 VDD.n4951 GND 0.10855f
C13974 VDD.t648 GND 0.02321f
C13975 VDD.t332 GND 0.02321f
C13976 VDD.n4952 GND 0.10855f
C13977 VDD.n4953 GND 0.06811f
C13978 VDD.n4954 GND 0.07249f
C13979 VDD.n4955 GND 0.0536f
C13980 VDD.n4956 GND 0.02522f
C13981 VDD.n4957 GND 0.04999f
C13982 VDD.n4958 GND 0.5126f
C13983 VDD.n4959 GND 0.02522f
C13984 VDD.n4960 GND 0.04999f
C13985 VDD.n4961 GND 0.5126f
C13986 VDD.n4962 GND 0.04999f
C13987 VDD.n4963 GND 0.05074f
C13988 VDD.n4964 GND 0.06295f
C13989 VDD.n4965 GND 0.0536f
C13990 VDD.n4966 GND 0.02522f
C13991 VDD.n4967 GND 0.04999f
C13992 VDD.n4968 GND 0.5126f
C13993 VDD.n4969 GND 0.02522f
C13994 VDD.n4970 GND 0.04999f
C13995 VDD.n4971 GND 0.5126f
C13996 VDD.n4972 GND 0.04999f
C13997 VDD.n4973 GND 0.05074f
C13998 VDD.n4974 GND 0.06295f
C13999 VDD.n4975 GND 0.0536f
C14000 VDD.n4976 GND 0.02522f
C14001 VDD.n4977 GND 0.04999f
C14002 VDD.n4978 GND 0.68843f
C14003 VDD.n4979 GND 0.02522f
C14004 VDD.n4980 GND 0.04999f
C14005 VDD.n4981 GND 0.68843f
C14006 VDD.n4982 GND 0.04999f
C14007 VDD.n4983 GND 0.05074f
C14008 VDD.n4984 GND 0.06295f
C14009 VDD.n4985 GND 0.0536f
C14010 VDD.n4986 GND 0.02522f
C14011 VDD.n4987 GND 0.04999f
C14012 VDD.n4988 GND 0.5126f
C14013 VDD.n4989 GND 0.02522f
C14014 VDD.n4990 GND 0.04999f
C14015 VDD.n4991 GND 0.5126f
C14016 VDD.n4992 GND 0.04999f
C14017 VDD.n4993 GND 0.05074f
C14018 VDD.n4994 GND 0.06295f
C14019 VDD.n4995 GND 0.0536f
C14020 VDD.n4996 GND 0.02522f
C14021 VDD.n4997 GND 0.04999f
C14022 VDD.n4998 GND 0.68843f
C14023 VDD.n4999 GND 0.68843f
C14024 VDD.n5000 GND 0.04999f
C14025 VDD.n5001 GND 0.02746f
C14026 VDD.n5002 GND 0.02967f
C14027 VDD.n5003 GND 0.02746f
C14028 VDD.n5004 GND 0.04999f
C14029 VDD.n5005 GND 0.68843f
C14030 VDD.n5006 GND 0.02522f
C14031 VDD.n5007 GND 0.04999f
C14032 VDD.n5008 GND 0.68843f
C14033 VDD.n5009 GND 0.04999f
C14034 VDD.n5010 GND 0.05074f
C14035 VDD.n5011 GND 0.06295f
C14036 VDD.n5012 GND 0.0536f
C14037 VDD.n5013 GND 0.02522f
C14038 VDD.n5014 GND 0.04999f
C14039 VDD.n5015 GND 0.5126f
C14040 VDD.n5016 GND 0.02522f
C14041 VDD.n5017 GND 0.04999f
C14042 VDD.n5018 GND 0.5126f
C14043 VDD.n5019 GND 0.04999f
C14044 VDD.n5020 GND 0.05074f
C14045 VDD.n5021 GND 0.06295f
C14046 VDD.n5022 GND 0.0536f
C14047 VDD.n5023 GND 0.02522f
C14048 VDD.n5024 GND 0.04999f
C14049 VDD.n5025 GND 0.5126f
C14050 VDD.n5026 GND 0.02522f
C14051 VDD.n5027 GND 0.04999f
C14052 VDD.n5028 GND 0.5126f
C14053 VDD.n5029 GND 0.04999f
C14054 VDD.n5030 GND 0.05074f
C14055 VDD.n5031 GND 0.06295f
C14056 VDD.n5032 GND 0.0536f
C14057 VDD.n5033 GND 0.02522f
C14058 VDD.n5034 GND 0.04999f
C14059 VDD.n5035 GND 0.68843f
C14060 VDD.n5036 GND 0.02522f
C14061 VDD.n5037 GND 0.04999f
C14062 VDD.n5038 GND 0.68843f
C14063 VDD.n5039 GND 0.04999f
C14064 VDD.n5040 GND 0.05074f
C14065 VDD.n5041 GND 0.06295f
C14066 VDD.n5042 GND 0.0536f
C14067 VDD.n5043 GND 0.02522f
C14068 VDD.n5044 GND 0.04999f
C14069 VDD.n5045 GND 0.5126f
C14070 VDD.n5046 GND 0.02522f
C14071 VDD.n5047 GND 0.04999f
C14072 VDD.n5048 GND 0.5126f
C14073 VDD.n5049 GND 0.04999f
C14074 VDD.n5050 GND 0.05074f
C14075 VDD.n5051 GND 0.06295f
C14076 VDD.n5052 GND 0.0536f
C14077 VDD.n5053 GND 0.02522f
C14078 VDD.n5054 GND 0.04999f
C14079 VDD.n5055 GND 0.5126f
C14080 VDD.n5056 GND 0.02522f
C14081 VDD.n5057 GND 0.04999f
C14082 VDD.n5058 GND 0.5126f
C14083 VDD.n5059 GND 0.04999f
C14084 VDD.n5060 GND 0.05074f
C14085 VDD.n5061 GND 0.06295f
C14086 VDD.n5062 GND 0.0536f
C14087 VDD.n5063 GND 0.02522f
C14088 VDD.n5064 GND 0.04999f
C14089 VDD.n5065 GND 0.68843f
C14090 VDD.n5066 GND 0.04999f
C14091 VDD.n5067 GND 0.68843f
C14092 VDD.t574 GND 0.74438f
C14093 VDD.n5069 GND 0.62973f
C14094 VDD.n5070 GND 0.02746f
C14095 VDD.n5071 GND 0.09132f
C14096 VDD.n5072 GND 0.01798f
C14097 VDD.n5073 GND 0.0731f
C14098 VDD.t930 GND 0.02321f
C14099 VDD.t432 GND 0.02321f
C14100 VDD.n5074 GND 0.10855f
C14101 VDD.t350 GND 0.02321f
C14102 VDD.t850 GND 0.02321f
C14103 VDD.n5075 GND 0.10855f
C14104 VDD.n5076 GND 0.04152f
C14105 VDD.n5077 GND 0.0536f
C14106 VDD.n5078 GND 0.05074f
C14107 VDD.n5079 GND 0.0536f
C14108 VDD.n5080 GND 0.04999f
C14109 VDD.n5081 GND 0.04999f
C14110 VDD.n5082 GND 0.68843f
C14111 VDD.n5083 GND 0.02522f
C14112 VDD.n5084 GND 0.02522f
C14113 VDD.n5085 GND 0.02967f
C14114 VDD.n5086 GND 0.05074f
C14115 VDD.n5087 GND 0.04999f
C14116 VDD.t431 GND 0.63568f
C14117 VDD.n5088 GND 0.05074f
C14118 VDD.n5089 GND 0.05074f
C14119 VDD.n5090 GND 0.02967f
C14120 VDD.n5091 GND 0.02522f
C14121 VDD.n5092 GND 0.03166f
C14122 VDD.n5093 GND 0.0536f
C14123 VDD.n5094 GND 0.05074f
C14124 VDD.n5095 GND 0.02967f
C14125 VDD.n5096 GND 0.02522f
C14126 VDD.n5097 GND 0.04999f
C14127 VDD.t433 GND 0.63568f
C14128 VDD.n5098 GND 0.05074f
C14129 VDD.n5099 GND 0.05074f
C14130 VDD.n5100 GND 0.02967f
C14131 VDD.n5101 GND 0.02522f
C14132 VDD.n5102 GND 0.0263f
C14133 VDD.n5103 GND 0.0536f
C14134 VDD.n5104 GND 0.05074f
C14135 VDD.n5105 GND 0.02967f
C14136 VDD.n5106 GND 0.02522f
C14137 VDD.n5107 GND 0.04999f
C14138 VDD.t330 GND 0.63568f
C14139 VDD.n5108 GND 0.05074f
C14140 VDD.n5109 GND 0.05074f
C14141 VDD.n5110 GND 0.02967f
C14142 VDD.n5111 GND 0.02522f
C14143 VDD.t434 GND 0.02334f
C14144 VDD.t707 GND 0.02334f
C14145 VDD.n5112 GND 0.13341f
C14146 VDD.n5113 GND 0.02334f
C14147 VDD.n5114 GND 0.0536f
C14148 VDD.n5115 GND 0.05074f
C14149 VDD.n5116 GND 0.02967f
C14150 VDD.n5117 GND 0.02522f
C14151 VDD.n5118 GND 0.04999f
C14152 VDD.t228 GND 0.63568f
C14153 VDD.n5119 GND 0.05074f
C14154 VDD.n5120 GND 0.05074f
C14155 VDD.n5121 GND 0.02967f
C14156 VDD.n5122 GND 0.02522f
C14157 VDD.t331 GND 0.02321f
C14158 VDD.t229 GND 0.02321f
C14159 VDD.n5123 GND 0.10855f
C14160 VDD.t851 GND 0.02321f
C14161 VDD.t286 GND 0.02321f
C14162 VDD.n5124 GND 0.10855f
C14163 VDD.n5125 GND 0.04152f
C14164 VDD.n5126 GND 0.02334f
C14165 VDD.n5127 GND 0.0536f
C14166 VDD.n5128 GND 0.05074f
C14167 VDD.n5129 GND 0.02967f
C14168 VDD.n5130 GND 0.02522f
C14169 VDD.t1076 GND 0.63568f
C14170 VDD.n5131 GND 0.05074f
C14171 VDD.n5132 GND 0.05074f
C14172 VDD.n5133 GND 0.09132f
C14173 VDD.n5134 GND 0.04999f
C14174 VDD.t226 GND 0.63568f
C14175 VDD.n5135 GND 0.05074f
C14176 VDD.n5136 GND 0.05074f
C14177 VDD.n5137 GND 0.02967f
C14178 VDD.n5138 GND 0.02522f
C14179 VDD.t1077 GND 0.02334f
C14180 VDD.n5139 GND 0.01798f
C14181 VDD.n5140 GND 0.0731f
C14182 VDD.n5141 GND 0.02334f
C14183 VDD.n5142 GND 0.0536f
C14184 VDD.n5143 GND 0.05074f
C14185 VDD.n5144 GND 0.02967f
C14186 VDD.n5145 GND 0.02522f
C14187 VDD.n5146 GND 0.04999f
C14188 VDD.t162 GND 0.63568f
C14189 VDD.n5147 GND 0.05074f
C14190 VDD.n5148 GND 0.05074f
C14191 VDD.n5149 GND 0.02967f
C14192 VDD.n5150 GND 0.02522f
C14193 VDD.t287 GND 0.02321f
C14194 VDD.t163 GND 0.02321f
C14195 VDD.n5151 GND 0.10855f
C14196 VDD.t227 GND 0.02321f
C14197 VDD.t612 GND 0.02321f
C14198 VDD.n5152 GND 0.10855f
C14199 VDD.n5153 GND 0.04152f
C14200 VDD.n5154 GND 0.03166f
C14201 VDD.n5155 GND 0.0536f
C14202 VDD.n5156 GND 0.05074f
C14203 VDD.n5157 GND 0.02967f
C14204 VDD.n5158 GND 0.02522f
C14205 VDD.n5159 GND 0.04999f
C14206 VDD.t510 GND 0.63568f
C14207 VDD.n5160 GND 0.05074f
C14208 VDD.n5161 GND 0.05074f
C14209 VDD.n5162 GND 0.02967f
C14210 VDD.n5163 GND 0.02522f
C14211 VDD.n5164 GND 0.0263f
C14212 VDD.n5165 GND 0.0536f
C14213 VDD.n5166 GND 0.05074f
C14214 VDD.n5167 GND 0.02967f
C14215 VDD.n5168 GND 0.02522f
C14216 VDD.n5169 GND 0.04999f
C14217 VDD.t1030 GND 0.63568f
C14218 VDD.n5170 GND 0.05074f
C14219 VDD.n5171 GND 0.05074f
C14220 VDD.n5172 GND 0.02967f
C14221 VDD.n5173 GND 0.02522f
C14222 VDD.t511 GND 0.02334f
C14223 VDD.t675 GND 0.02334f
C14224 VDD.n5174 GND 0.13341f
C14225 VDD.n5175 GND 0.02334f
C14226 VDD.n5176 GND 0.0536f
C14227 VDD.n5177 GND 0.05074f
C14228 VDD.n5178 GND 0.02967f
C14229 VDD.n5179 GND 0.02522f
C14230 VDD.n5180 GND 0.04999f
C14231 VDD.t390 GND 0.63568f
C14232 VDD.n5181 GND 0.05074f
C14233 VDD.n5182 GND 0.05074f
C14234 VDD.n5183 GND 0.02967f
C14235 VDD.n5184 GND 0.02522f
C14236 VDD.t1095 GND 0.02321f
C14237 VDD.t780 GND 0.02321f
C14238 VDD.n5185 GND 0.10855f
C14239 VDD.t1031 GND 0.02321f
C14240 VDD.t391 GND 0.02321f
C14241 VDD.n5186 GND 0.10855f
C14242 VDD.n5187 GND 0.04152f
C14243 VDD.n5188 GND 0.03166f
C14244 VDD.n5189 GND 0.0536f
C14245 VDD.n5190 GND 0.05074f
C14246 VDD.n5191 GND 0.02967f
C14247 VDD.n5192 GND 0.02522f
C14248 VDD.n5193 GND 0.04999f
C14249 VDD.t457 GND 0.63568f
C14250 VDD.n5194 GND 0.05074f
C14251 VDD.n5195 GND 0.05074f
C14252 VDD.n5196 GND 0.02967f
C14253 VDD.n5197 GND 0.02522f
C14254 VDD.n5198 GND 0.0263f
C14255 VDD.n5199 GND 0.0536f
C14256 VDD.n5200 GND 0.05074f
C14257 VDD.n5201 GND 0.02967f
C14258 VDD.n5202 GND 0.02522f
C14259 VDD.t919 GND 0.74438f
C14260 VDD.n5203 GND 0.05074f
C14261 VDD.n5204 GND 0.05074f
C14262 VDD.n5205 GND 0.02967f
C14263 VDD.n5207 GND 0.62973f
C14264 VDD.n5208 GND 0.02746f
C14265 VDD.t753 GND 0.02334f
C14266 VDD.t458 GND 0.02334f
C14267 VDD.n5209 GND 0.13341f
C14268 VDD.t920 GND 0.02334f
C14269 VDD.t306 GND 0.02321f
C14270 VDD.t587 GND 0.02321f
C14271 VDD.n5210 GND 0.10855f
C14272 VDD.t918 GND 0.02321f
C14273 VDD.t321 GND 0.02321f
C14274 VDD.n5211 GND 0.10855f
C14275 VDD.n5212 GND 0.04152f
C14276 VDD.n5213 GND 0.0536f
C14277 VDD.n5214 GND 0.05074f
C14278 VDD.n5215 GND 0.0536f
C14279 VDD.n5216 GND 0.04999f
C14280 VDD.n5217 GND 0.04999f
C14281 VDD.n5218 GND 0.68843f
C14282 VDD.n5219 GND 0.02522f
C14283 VDD.n5220 GND 0.02522f
C14284 VDD.n5221 GND 0.02967f
C14285 VDD.n5222 GND 0.05074f
C14286 VDD.n5223 GND 0.04999f
C14287 VDD.t320 GND 0.63568f
C14288 VDD.n5224 GND 0.05074f
C14289 VDD.n5225 GND 0.05074f
C14290 VDD.n5226 GND 0.02967f
C14291 VDD.n5227 GND 0.02522f
C14292 VDD.n5228 GND 0.03166f
C14293 VDD.n5229 GND 0.0536f
C14294 VDD.n5230 GND 0.05074f
C14295 VDD.n5231 GND 0.02967f
C14296 VDD.n5232 GND 0.02522f
C14297 VDD.n5233 GND 0.04999f
C14298 VDD.t482 GND 0.63568f
C14299 VDD.n5234 GND 0.05074f
C14300 VDD.n5235 GND 0.05074f
C14301 VDD.n5236 GND 0.02967f
C14302 VDD.n5237 GND 0.02522f
C14303 VDD.n5238 GND 0.0263f
C14304 VDD.n5239 GND 0.0536f
C14305 VDD.n5240 GND 0.05074f
C14306 VDD.n5241 GND 0.02967f
C14307 VDD.n5242 GND 0.02522f
C14308 VDD.n5243 GND 0.04999f
C14309 VDD.t378 GND 0.63568f
C14310 VDD.n5244 GND 0.05074f
C14311 VDD.n5245 GND 0.05074f
C14312 VDD.n5246 GND 0.02967f
C14313 VDD.n5247 GND 0.02522f
C14314 VDD.t483 GND 0.02334f
C14315 VDD.t757 GND 0.02334f
C14316 VDD.n5248 GND 0.13341f
C14317 VDD.n5249 GND 0.02334f
C14318 VDD.n5250 GND 0.0536f
C14319 VDD.n5251 GND 0.05074f
C14320 VDD.n5252 GND 0.02967f
C14321 VDD.n5253 GND 0.02522f
C14322 VDD.n5254 GND 0.04999f
C14323 VDD.t316 GND 0.63568f
C14324 VDD.n5255 GND 0.05074f
C14325 VDD.n5256 GND 0.05074f
C14326 VDD.n5257 GND 0.02967f
C14327 VDD.n5258 GND 0.02522f
C14328 VDD.t379 GND 0.02321f
C14329 VDD.t376 GND 0.02321f
C14330 VDD.n5259 GND 0.10855f
C14331 VDD.t543 GND 0.02321f
C14332 VDD.t317 GND 0.02321f
C14333 VDD.n5260 GND 0.10855f
C14334 VDD.n5261 GND 0.04152f
C14335 VDD.n5262 GND 0.02334f
C14336 VDD.n5263 GND 0.0536f
C14337 VDD.n5264 GND 0.05074f
C14338 VDD.n5265 GND 0.02967f
C14339 VDD.n5266 GND 0.02522f
C14340 VDD.t1058 GND 0.63568f
C14341 VDD.n5267 GND 0.05074f
C14342 VDD.n5268 GND 0.05074f
C14343 VDD.n5269 GND 0.09132f
C14344 VDD.n5270 GND 0.04999f
C14345 VDD.t314 GND 0.63568f
C14346 VDD.n5271 GND 0.05074f
C14347 VDD.n5272 GND 0.05074f
C14348 VDD.n5273 GND 0.02967f
C14349 VDD.n5274 GND 0.02522f
C14350 VDD.t1059 GND 0.02334f
C14351 VDD.n5275 GND 0.01798f
C14352 VDD.n5276 GND 0.0731f
C14353 VDD.n5277 GND 0.02334f
C14354 VDD.n5278 GND 0.0536f
C14355 VDD.n5279 GND 0.05074f
C14356 VDD.n5280 GND 0.02967f
C14357 VDD.n5281 GND 0.02522f
C14358 VDD.n5282 GND 0.04999f
C14359 VDD.t366 GND 0.63568f
C14360 VDD.n5283 GND 0.05074f
C14361 VDD.n5284 GND 0.05074f
C14362 VDD.n5285 GND 0.02967f
C14363 VDD.n5286 GND 0.02522f
C14364 VDD.t315 GND 0.02321f
C14365 VDD.t661 GND 0.02321f
C14366 VDD.n5287 GND 0.10855f
C14367 VDD.t377 GND 0.02321f
C14368 VDD.t367 GND 0.02321f
C14369 VDD.n5288 GND 0.10855f
C14370 VDD.n5289 GND 0.04152f
C14371 VDD.n5290 GND 0.03166f
C14372 VDD.n5291 GND 0.0536f
C14373 VDD.n5292 GND 0.05074f
C14374 VDD.n5293 GND 0.02967f
C14375 VDD.n5294 GND 0.02522f
C14376 VDD.n5295 GND 0.04999f
C14377 VDD.t520 GND 0.63568f
C14378 VDD.n5296 GND 0.05074f
C14379 VDD.n5297 GND 0.05074f
C14380 VDD.n5298 GND 0.02967f
C14381 VDD.n5299 GND 0.02522f
C14382 VDD.n5300 GND 0.0263f
C14383 VDD.n5301 GND 0.0536f
C14384 VDD.n5302 GND 0.05074f
C14385 VDD.n5303 GND 0.02967f
C14386 VDD.n5304 GND 0.02522f
C14387 VDD.n5305 GND 0.04999f
C14388 VDD.t1032 GND 0.63568f
C14389 VDD.n5306 GND 0.05074f
C14390 VDD.n5307 GND 0.05074f
C14391 VDD.n5308 GND 0.02967f
C14392 VDD.n5309 GND 0.02522f
C14393 VDD.t521 GND 0.02334f
C14394 VDD.t681 GND 0.02334f
C14395 VDD.n5310 GND 0.13341f
C14396 VDD.n5311 GND 0.02334f
C14397 VDD.n5312 GND 0.0536f
C14398 VDD.n5313 GND 0.05074f
C14399 VDD.n5314 GND 0.02967f
C14400 VDD.n5315 GND 0.02522f
C14401 VDD.n5316 GND 0.04999f
C14402 VDD.t835 GND 0.63568f
C14403 VDD.n5317 GND 0.05074f
C14404 VDD.n5318 GND 0.05074f
C14405 VDD.n5319 GND 0.02967f
C14406 VDD.n5320 GND 0.02522f
C14407 VDD.t1033 GND 0.02321f
C14408 VDD.t836 GND 0.02321f
C14409 VDD.n5321 GND 0.10855f
C14410 VDD.t1078 GND 0.02321f
C14411 VDD.t904 GND 0.02321f
C14412 VDD.n5322 GND 0.10855f
C14413 VDD.n5323 GND 0.04152f
C14414 VDD.n5324 GND 0.03166f
C14415 VDD.n5325 GND 0.0536f
C14416 VDD.n5326 GND 0.05074f
C14417 VDD.n5327 GND 0.02967f
C14418 VDD.n5328 GND 0.02522f
C14419 VDD.n5329 GND 0.04999f
C14420 VDD.t465 GND 0.63568f
C14421 VDD.n5330 GND 0.05074f
C14422 VDD.n5331 GND 0.05074f
C14423 VDD.n5332 GND 0.02967f
C14424 VDD.n5333 GND 0.02522f
C14425 VDD.n5334 GND 0.0263f
C14426 VDD.n5335 GND 0.0536f
C14427 VDD.n5336 GND 0.05074f
C14428 VDD.n5337 GND 0.02967f
C14429 VDD.n5338 GND 0.02522f
C14430 VDD.t840 GND 0.74438f
C14431 VDD.n5339 GND 0.05074f
C14432 VDD.n5340 GND 0.05074f
C14433 VDD.n5341 GND 0.02967f
C14434 VDD.n5343 GND 0.62973f
C14435 VDD.n5344 GND 0.02746f
C14436 VDD.t759 GND 0.02334f
C14437 VDD.t466 GND 0.02334f
C14438 VDD.n5345 GND 0.13341f
C14439 VDD.t841 GND 0.02334f
C14440 VDD.t313 GND 0.02321f
C14441 VDD.t34 GND 0.02321f
C14442 VDD.n5346 GND 0.10855f
C14443 VDD.t837 GND 0.02321f
C14444 VDD.t195 GND 0.02321f
C14445 VDD.n5347 GND 0.10855f
C14446 VDD.n5348 GND 0.04152f
C14447 VDD.n5349 GND 0.0536f
C14448 VDD.n5350 GND 0.05074f
C14449 VDD.n5351 GND 0.0536f
C14450 VDD.n5352 GND 0.04999f
C14451 VDD.n5353 GND 0.04999f
C14452 VDD.n5354 GND 0.68843f
C14453 VDD.n5355 GND 0.02522f
C14454 VDD.n5356 GND 0.02522f
C14455 VDD.n5357 GND 0.02967f
C14456 VDD.n5358 GND 0.05074f
C14457 VDD.n5359 GND 0.04999f
C14458 VDD.t33 GND 0.63568f
C14459 VDD.n5360 GND 0.05074f
C14460 VDD.n5361 GND 0.05074f
C14461 VDD.n5362 GND 0.02967f
C14462 VDD.n5363 GND 0.02522f
C14463 VDD.n5364 GND 0.03166f
C14464 VDD.n5365 GND 0.0536f
C14465 VDD.n5366 GND 0.05074f
C14466 VDD.n5367 GND 0.02967f
C14467 VDD.n5368 GND 0.02522f
C14468 VDD.n5369 GND 0.04999f
C14469 VDD.t492 GND 0.63568f
C14470 VDD.n5370 GND 0.05074f
C14471 VDD.n5371 GND 0.05074f
C14472 VDD.n5372 GND 0.02967f
C14473 VDD.n5373 GND 0.02522f
C14474 VDD.n5374 GND 0.0263f
C14475 VDD.n5375 GND 0.0536f
C14476 VDD.n5376 GND 0.05074f
C14477 VDD.n5377 GND 0.02967f
C14478 VDD.n5378 GND 0.02522f
C14479 VDD.n5379 GND 0.04999f
C14480 VDD.t139 GND 0.63568f
C14481 VDD.n5380 GND 0.05074f
C14482 VDD.n5381 GND 0.05074f
C14483 VDD.n5382 GND 0.02967f
C14484 VDD.n5383 GND 0.02522f
C14485 VDD.t493 GND 0.02334f
C14486 VDD.t663 GND 0.02334f
C14487 VDD.n5384 GND 0.13341f
C14488 VDD.n5385 GND 0.02334f
C14489 VDD.n5386 GND 0.0536f
C14490 VDD.n5387 GND 0.05074f
C14491 VDD.n5388 GND 0.02967f
C14492 VDD.n5389 GND 0.02522f
C14493 VDD.n5390 GND 0.04999f
C14494 VDD.t208 GND 0.63568f
C14495 VDD.n5391 GND 0.05074f
C14496 VDD.n5392 GND 0.05074f
C14497 VDD.n5393 GND 0.02967f
C14498 VDD.n5394 GND 0.02522f
C14499 VDD.t140 GND 0.02321f
C14500 VDD.t282 GND 0.02321f
C14501 VDD.n5395 GND 0.10855f
C14502 VDD.t551 GND 0.02321f
C14503 VDD.t209 GND 0.02321f
C14504 VDD.n5396 GND 0.10855f
C14505 VDD.n5397 GND 0.04152f
C14506 VDD.n5398 GND 0.02334f
C14507 VDD.n5399 GND 0.0536f
C14508 VDD.n5400 GND 0.05074f
C14509 VDD.n5401 GND 0.02967f
C14510 VDD.n5402 GND 0.02522f
C14511 VDD.t1084 GND 0.63568f
C14512 VDD.n5403 GND 0.05074f
C14513 VDD.n5404 GND 0.05074f
C14514 VDD.n5405 GND 0.09132f
C14515 VDD.n5406 GND 0.04999f
C14516 VDD.t280 GND 0.63568f
C14517 VDD.n5407 GND 0.05074f
C14518 VDD.n5408 GND 0.05074f
C14519 VDD.n5409 GND 0.02967f
C14520 VDD.n5410 GND 0.02522f
C14521 VDD.t1085 GND 0.02334f
C14522 VDD.n5411 GND 0.01798f
C14523 VDD.n5412 GND 0.0731f
C14524 VDD.n5413 GND 0.02334f
C14525 VDD.n5414 GND 0.0536f
C14526 VDD.n5415 GND 0.05074f
C14527 VDD.n5416 GND 0.02967f
C14528 VDD.n5417 GND 0.02522f
C14529 VDD.n5418 GND 0.04999f
C14530 VDD.t17 GND 0.63568f
C14531 VDD.n5419 GND 0.05074f
C14532 VDD.n5420 GND 0.05074f
C14533 VDD.n5421 GND 0.02967f
C14534 VDD.n5422 GND 0.02522f
C14535 VDD.t585 GND 0.02321f
C14536 VDD.t274 GND 0.02321f
C14537 VDD.n5423 GND 0.10855f
C14538 VDD.t281 GND 0.02321f
C14539 VDD.t18 GND 0.02321f
C14540 VDD.n5424 GND 0.10855f
C14541 VDD.n5425 GND 0.04152f
C14542 VDD.n5426 GND 0.03166f
C14543 VDD.n5427 GND 0.0536f
C14544 VDD.n5428 GND 0.05074f
C14545 VDD.n5429 GND 0.02967f
C14546 VDD.n5430 GND 0.02522f
C14547 VDD.n5431 GND 0.04999f
C14548 VDD.t475 GND 0.63568f
C14549 VDD.n5432 GND 0.05074f
C14550 VDD.n5433 GND 0.05074f
C14551 VDD.n5434 GND 0.02967f
C14552 VDD.n5435 GND 0.02522f
C14553 VDD.n5436 GND 0.0263f
C14554 VDD.n5437 GND 0.0536f
C14555 VDD.n5438 GND 0.05074f
C14556 VDD.n5439 GND 0.02967f
C14557 VDD.n5440 GND 0.02522f
C14558 VDD.n5441 GND 0.04999f
C14559 VDD.t1060 GND 0.63568f
C14560 VDD.n5442 GND 0.05074f
C14561 VDD.n5443 GND 0.05074f
C14562 VDD.n5444 GND 0.02967f
C14563 VDD.n5445 GND 0.02522f
C14564 VDD.t476 GND 0.02334f
C14565 VDD.t745 GND 0.02334f
C14566 VDD.n5446 GND 0.13341f
C14567 VDD.n5447 GND 0.02334f
C14568 VDD.n5448 GND 0.0536f
C14569 VDD.n5449 GND 0.05074f
C14570 VDD.n5450 GND 0.02967f
C14571 VDD.n5451 GND 0.02522f
C14572 VDD.n5452 GND 0.04999f
C14573 VDD.t425 GND 0.63568f
C14574 VDD.n5453 GND 0.05074f
C14575 VDD.n5454 GND 0.05074f
C14576 VDD.n5455 GND 0.02967f
C14577 VDD.n5456 GND 0.02522f
C14578 VDD.t1061 GND 0.02321f
C14579 VDD.t804 GND 0.02321f
C14580 VDD.n5457 GND 0.10855f
C14581 VDD.t1093 GND 0.02321f
C14582 VDD.t426 GND 0.02321f
C14583 VDD.n5458 GND 0.10855f
C14584 VDD.n5459 GND 0.04152f
C14585 VDD.n5460 GND 0.03166f
C14586 VDD.n5461 GND 0.0536f
C14587 VDD.n5462 GND 0.05074f
C14588 VDD.n5463 GND 0.02967f
C14589 VDD.n5464 GND 0.02522f
C14590 VDD.n5465 GND 0.04999f
C14591 VDD.t478 GND 0.63568f
C14592 VDD.n5466 GND 0.05074f
C14593 VDD.n5467 GND 0.05074f
C14594 VDD.n5468 GND 0.02967f
C14595 VDD.n5469 GND 0.02522f
C14596 VDD.n5470 GND 0.0263f
C14597 VDD.n5471 GND 0.0536f
C14598 VDD.n5472 GND 0.05074f
C14599 VDD.n5473 GND 0.02967f
C14600 VDD.n5474 GND 0.02522f
C14601 VDD.t23 GND 0.74438f
C14602 VDD.n5475 GND 0.05074f
C14603 VDD.n5476 GND 0.05074f
C14604 VDD.n5477 GND 0.02967f
C14605 VDD.n5479 GND 0.62973f
C14606 VDD.n5480 GND 0.02746f
C14607 VDD.t673 GND 0.02334f
C14608 VDD.t479 GND 0.02334f
C14609 VDD.n5481 GND 0.13341f
C14610 VDD.t24 GND 0.02334f
C14611 VDD.t47 GND 0.02321f
C14612 VDD.t254 GND 0.02321f
C14613 VDD.n5482 GND 0.10855f
C14614 VDD.t130 GND 0.02321f
C14615 VDD.t656 GND 0.02321f
C14616 VDD.n5483 GND 0.10855f
C14617 VDD.n5484 GND 0.04152f
C14618 VDD.n5485 GND 0.0536f
C14619 VDD.n5486 GND 0.05074f
C14620 VDD.n5487 GND 0.0536f
C14621 VDD.n5488 GND 0.04999f
C14622 VDD.n5489 GND 0.04999f
C14623 VDD.n5490 GND 0.68843f
C14624 VDD.n5491 GND 0.02522f
C14625 VDD.n5492 GND 0.02522f
C14626 VDD.n5493 GND 0.02967f
C14627 VDD.n5494 GND 0.05074f
C14628 VDD.n5495 GND 0.04999f
C14629 VDD.t253 GND 0.63568f
C14630 VDD.n5496 GND 0.05074f
C14631 VDD.n5497 GND 0.05074f
C14632 VDD.n5498 GND 0.02967f
C14633 VDD.n5499 GND 0.02522f
C14634 VDD.n5500 GND 0.03166f
C14635 VDD.n5501 GND 0.0536f
C14636 VDD.n5502 GND 0.05074f
C14637 VDD.n5503 GND 0.02967f
C14638 VDD.n5504 GND 0.02522f
C14639 VDD.n5505 GND 0.04999f
C14640 VDD.t459 GND 0.63568f
C14641 VDD.n5506 GND 0.05074f
C14642 VDD.n5507 GND 0.05074f
C14643 VDD.n5508 GND 0.02967f
C14644 VDD.n5509 GND 0.02522f
C14645 VDD.n5510 GND 0.0263f
C14646 VDD.n5511 GND 0.0536f
C14647 VDD.n5512 GND 0.05074f
C14648 VDD.n5513 GND 0.02967f
C14649 VDD.n5514 GND 0.02522f
C14650 VDD.n5515 GND 0.04999f
C14651 VDD.t237 GND 0.63568f
C14652 VDD.n5516 GND 0.05074f
C14653 VDD.n5517 GND 0.05074f
C14654 VDD.n5518 GND 0.02967f
C14655 VDD.n5519 GND 0.02522f
C14656 VDD.t460 GND 0.02334f
C14657 VDD.t735 GND 0.02334f
C14658 VDD.n5520 GND 0.13341f
C14659 VDD.n5521 GND 0.02334f
C14660 VDD.n5522 GND 0.0536f
C14661 VDD.n5523 GND 0.05074f
C14662 VDD.n5524 GND 0.02967f
C14663 VDD.n5525 GND 0.02522f
C14664 VDD.n5526 GND 0.04999f
C14665 VDD.t257 GND 0.63568f
C14666 VDD.n5527 GND 0.05074f
C14667 VDD.n5528 GND 0.05074f
C14668 VDD.n5529 GND 0.02967f
C14669 VDD.n5530 GND 0.02522f
C14670 VDD.t238 GND 0.02321f
C14671 VDD.t891 GND 0.02321f
C14672 VDD.n5531 GND 0.10855f
C14673 VDD.t960 GND 0.02321f
C14674 VDD.t258 GND 0.02321f
C14675 VDD.n5532 GND 0.10855f
C14676 VDD.n5533 GND 0.04152f
C14677 VDD.n5534 GND 0.02334f
C14678 VDD.n5535 GND 0.0536f
C14679 VDD.n5536 GND 0.05074f
C14680 VDD.n5537 GND 0.02967f
C14681 VDD.n5538 GND 0.02522f
C14682 VDD.t1096 GND 0.63568f
C14683 VDD.n5539 GND 0.05074f
C14684 VDD.n5540 GND 0.05074f
C14685 VDD.n5541 GND 0.09132f
C14686 VDD.n5542 GND 0.04999f
C14687 VDD.t135 GND 0.63568f
C14688 VDD.n5543 GND 0.05074f
C14689 VDD.n5544 GND 0.05074f
C14690 VDD.n5545 GND 0.02967f
C14691 VDD.n5546 GND 0.02522f
C14692 VDD.t1097 GND 0.02334f
C14693 VDD.n5547 GND 0.01798f
C14694 VDD.n5548 GND 0.0731f
C14695 VDD.n5549 GND 0.02334f
C14696 VDD.n5550 GND 0.0536f
C14697 VDD.n5551 GND 0.05074f
C14698 VDD.n5552 GND 0.02967f
C14699 VDD.n5553 GND 0.02522f
C14700 VDD.n5554 GND 0.04999f
C14701 VDD.t794 GND 0.63568f
C14702 VDD.n5555 GND 0.05074f
C14703 VDD.n5556 GND 0.05074f
C14704 VDD.n5557 GND 0.02967f
C14705 VDD.n5558 GND 0.02522f
C14706 VDD.t136 GND 0.02321f
C14707 VDD.t983 GND 0.02321f
C14708 VDD.n5559 GND 0.10855f
C14709 VDD.t908 GND 0.02321f
C14710 VDD.t795 GND 0.02321f
C14711 VDD.n5560 GND 0.10855f
C14712 VDD.n5561 GND 0.04152f
C14713 VDD.n5562 GND 0.03166f
C14714 VDD.n5563 GND 0.0536f
C14715 VDD.n5564 GND 0.05074f
C14716 VDD.n5565 GND 0.02967f
C14717 VDD.n5566 GND 0.02522f
C14718 VDD.n5567 GND 0.04999f
C14719 VDD.t490 GND 0.63568f
C14720 VDD.n5568 GND 0.05074f
C14721 VDD.n5569 GND 0.05074f
C14722 VDD.n5570 GND 0.02967f
C14723 VDD.n5571 GND 0.02522f
C14724 VDD.n5572 GND 0.0263f
C14725 VDD.n5573 GND 0.0536f
C14726 VDD.n5574 GND 0.05074f
C14727 VDD.n5575 GND 0.02967f
C14728 VDD.n5576 GND 0.02522f
C14729 VDD.n5577 GND 0.04999f
C14730 VDD.t1002 GND 0.63568f
C14731 VDD.n5578 GND 0.05074f
C14732 VDD.n5579 GND 0.05074f
C14733 VDD.n5580 GND 0.02967f
C14734 VDD.n5581 GND 0.02522f
C14735 VDD.t491 GND 0.02334f
C14736 VDD.t763 GND 0.02334f
C14737 VDD.n5582 GND 0.13341f
C14738 VDD.n5583 GND 0.02334f
C14739 VDD.n5584 GND 0.0536f
C14740 VDD.n5585 GND 0.05074f
C14741 VDD.n5586 GND 0.02967f
C14742 VDD.n5587 GND 0.02522f
C14743 VDD.n5588 GND 0.04999f
C14744 VDD.t871 GND 0.63568f
C14745 VDD.n5589 GND 0.05074f
C14746 VDD.n5590 GND 0.05074f
C14747 VDD.n5591 GND 0.02967f
C14748 VDD.n5592 GND 0.02522f
C14749 VDD.t1003 GND 0.02321f
C14750 VDD.t872 GND 0.02321f
C14751 VDD.n5593 GND 0.10855f
C14752 VDD.t1047 GND 0.02321f
C14753 VDD.t886 GND 0.02321f
C14754 VDD.n5594 GND 0.10855f
C14755 VDD.n5595 GND 0.04152f
C14756 VDD.n5596 GND 0.03166f
C14757 VDD.n5597 GND 0.0536f
C14758 VDD.n5598 GND 0.05074f
C14759 VDD.n5599 GND 0.02967f
C14760 VDD.n5600 GND 0.02522f
C14761 VDD.n5601 GND 0.04999f
C14762 VDD.t443 GND 0.63568f
C14763 VDD.n5602 GND 0.05074f
C14764 VDD.n5603 GND 0.05074f
C14765 VDD.n5604 GND 0.02967f
C14766 VDD.n5605 GND 0.02522f
C14767 VDD.n5606 GND 0.0263f
C14768 VDD.n5607 GND 0.0536f
C14769 VDD.n5608 GND 0.05074f
C14770 VDD.n5609 GND 0.02967f
C14771 VDD.n5610 GND 0.02522f
C14772 VDD.t621 GND 0.74438f
C14773 VDD.n5611 GND 0.05074f
C14774 VDD.n5612 GND 0.05074f
C14775 VDD.n5613 GND 0.02967f
C14776 VDD.n5615 GND 0.62973f
C14777 VDD.n5616 GND 0.02746f
C14778 VDD.t737 GND 0.02334f
C14779 VDD.t444 GND 0.02334f
C14780 VDD.n5617 GND 0.13341f
C14781 VDD.t622 GND 0.02334f
C14782 VDD.t365 GND 0.02321f
C14783 VDD.t252 GND 0.02321f
C14784 VDD.n5618 GND 0.10855f
C14785 VDD.t623 GND 0.02321f
C14786 VDD.t110 GND 0.02321f
C14787 VDD.n5619 GND 0.10855f
C14788 VDD.n5620 GND 0.04152f
C14789 VDD.n5621 GND 0.0536f
C14790 VDD.n5622 GND 0.05074f
C14791 VDD.n5623 GND 0.0536f
C14792 VDD.n5624 GND 0.04999f
C14793 VDD.n5625 GND 0.04999f
C14794 VDD.n5626 GND 0.68843f
C14795 VDD.n5627 GND 0.02522f
C14796 VDD.n5628 GND 0.02522f
C14797 VDD.n5629 GND 0.02967f
C14798 VDD.n5630 GND 0.05074f
C14799 VDD.n5631 GND 0.04999f
C14800 VDD.t109 GND 0.63568f
C14801 VDD.n5632 GND 0.05074f
C14802 VDD.n5633 GND 0.05074f
C14803 VDD.n5634 GND 0.02967f
C14804 VDD.n5635 GND 0.02522f
C14805 VDD.n5636 GND 0.03166f
C14806 VDD.n5637 GND 0.0536f
C14807 VDD.n5638 GND 0.05074f
C14808 VDD.n5639 GND 0.02967f
C14809 VDD.n5640 GND 0.02522f
C14810 VDD.n5641 GND 0.04999f
C14811 VDD.t506 GND 0.63568f
C14812 VDD.n5642 GND 0.05074f
C14813 VDD.n5643 GND 0.05074f
C14814 VDD.n5644 GND 0.02967f
C14815 VDD.n5645 GND 0.02522f
C14816 VDD.n5646 GND 0.0263f
C14817 VDD.n5647 GND 0.0536f
C14818 VDD.n5648 GND 0.05074f
C14819 VDD.n5649 GND 0.02967f
C14820 VDD.n5650 GND 0.02522f
C14821 VDD.n5651 GND 0.04999f
C14822 VDD.t552 GND 0.63568f
C14823 VDD.n5652 GND 0.05074f
C14824 VDD.n5653 GND 0.05074f
C14825 VDD.n5654 GND 0.02967f
C14826 VDD.n5655 GND 0.02522f
C14827 VDD.t507 GND 0.02334f
C14828 VDD.t679 GND 0.02334f
C14829 VDD.n5656 GND 0.13341f
C14830 VDD.n5657 GND 0.02334f
C14831 VDD.n5658 GND 0.0536f
C14832 VDD.n5659 GND 0.05074f
C14833 VDD.n5660 GND 0.02967f
C14834 VDD.n5661 GND 0.02522f
C14835 VDD.n5662 GND 0.04999f
C14836 VDD.t145 GND 0.63568f
C14837 VDD.n5663 GND 0.05074f
C14838 VDD.n5664 GND 0.05074f
C14839 VDD.n5665 GND 0.02967f
C14840 VDD.n5666 GND 0.02522f
C14841 VDD.t553 GND 0.02321f
C14842 VDD.t268 GND 0.02321f
C14843 VDD.n5667 GND 0.10855f
C14844 VDD.t554 GND 0.02321f
C14845 VDD.t146 GND 0.02321f
C14846 VDD.n5668 GND 0.10855f
C14847 VDD.n5669 GND 0.04152f
C14848 VDD.n5670 GND 0.02334f
C14849 VDD.n5671 GND 0.0536f
C14850 VDD.n5672 GND 0.05074f
C14851 VDD.n5673 GND 0.02967f
C14852 VDD.n5674 GND 0.02522f
C14853 VDD.t1054 GND 0.63568f
C14854 VDD.n5675 GND 0.05074f
C14855 VDD.n5676 GND 0.05074f
C14856 VDD.n5677 GND 0.09132f
C14857 VDD.n5678 GND 0.04999f
C14858 VDD.t147 GND 0.63568f
C14859 VDD.n5679 GND 0.05074f
C14860 VDD.n5680 GND 0.05074f
C14861 VDD.n5681 GND 0.02967f
C14862 VDD.n5682 GND 0.02522f
C14863 VDD.t1055 GND 0.02334f
C14864 VDD.n5683 GND 0.01798f
C14865 VDD.n5684 GND 0.0731f
C14866 VDD.n5685 GND 0.02334f
C14867 VDD.n5686 GND 0.0536f
C14868 VDD.n5687 GND 0.05074f
C14869 VDD.n5688 GND 0.02967f
C14870 VDD.n5689 GND 0.02522f
C14871 VDD.n5690 GND 0.04999f
C14872 VDD.t116 GND 0.63568f
C14873 VDD.n5691 GND 0.05074f
C14874 VDD.n5692 GND 0.05074f
C14875 VDD.n5693 GND 0.02967f
C14876 VDD.n5694 GND 0.02522f
C14877 VDD.t148 GND 0.02321f
C14878 VDD.t117 GND 0.02321f
C14879 VDD.n5695 GND 0.10855f
C14880 VDD.t820 GND 0.02321f
C14881 VDD.t869 GND 0.02321f
C14882 VDD.n5696 GND 0.10855f
C14883 VDD.n5697 GND 0.04152f
C14884 VDD.n5698 GND 0.03166f
C14885 VDD.n5699 GND 0.0536f
C14886 VDD.n5700 GND 0.05074f
C14887 VDD.n5701 GND 0.02967f
C14888 VDD.n5702 GND 0.02522f
C14889 VDD.n5703 GND 0.04999f
C14890 VDD.t453 GND 0.63568f
C14891 VDD.n5704 GND 0.05074f
C14892 VDD.n5705 GND 0.05074f
C14893 VDD.n5706 GND 0.02967f
C14894 VDD.n5707 GND 0.02522f
C14895 VDD.n5708 GND 0.0263f
C14896 VDD.n5709 GND 0.0536f
C14897 VDD.n5710 GND 0.05074f
C14898 VDD.n5711 GND 0.02967f
C14899 VDD.n5712 GND 0.02522f
C14900 VDD.n5713 GND 0.04999f
C14901 VDD.t1028 GND 0.63568f
C14902 VDD.n5714 GND 0.05074f
C14903 VDD.n5715 GND 0.05074f
C14904 VDD.n5716 GND 0.02967f
C14905 VDD.n5717 GND 0.02522f
C14906 VDD.t454 GND 0.02334f
C14907 VDD.t721 GND 0.02334f
C14908 VDD.n5718 GND 0.13341f
C14909 VDD.n5719 GND 0.02334f
C14910 VDD.n5720 GND 0.0536f
C14911 VDD.n5721 GND 0.05074f
C14912 VDD.n5722 GND 0.02967f
C14913 VDD.n5723 GND 0.02522f
C14914 VDD.n5724 GND 0.04999f
C14915 VDD.t368 GND 0.63568f
C14916 VDD.n5725 GND 0.05074f
C14917 VDD.n5726 GND 0.05074f
C14918 VDD.n5727 GND 0.02967f
C14919 VDD.n5728 GND 0.02522f
C14920 VDD.t1029 GND 0.02321f
C14921 VDD.t369 GND 0.02321f
C14922 VDD.n5729 GND 0.10855f
C14923 VDD.t1070 GND 0.02321f
C14924 VDD.t980 GND 0.02321f
C14925 VDD.n5730 GND 0.10855f
C14926 VDD.n5731 GND 0.04152f
C14927 VDD.n5732 GND 0.03166f
C14928 VDD.n5733 GND 0.0536f
C14929 VDD.n5734 GND 0.05074f
C14930 VDD.n5735 GND 0.02967f
C14931 VDD.n5736 GND 0.02522f
C14932 VDD.n5737 GND 0.04999f
C14933 VDD.t463 GND 0.63568f
C14934 VDD.n5738 GND 0.05074f
C14935 VDD.n5739 GND 0.05074f
C14936 VDD.n5740 GND 0.02967f
C14937 VDD.n5741 GND 0.02522f
C14938 VDD.n5742 GND 0.0263f
C14939 VDD.n5743 GND 0.0536f
C14940 VDD.n5744 GND 0.05074f
C14941 VDD.n5745 GND 0.02967f
C14942 VDD.n5746 GND 0.02522f
C14943 VDD.t916 GND 0.74438f
C14944 VDD.n5747 GND 0.05074f
C14945 VDD.n5748 GND 0.05074f
C14946 VDD.n5749 GND 0.02967f
C14947 VDD.n5751 GND 0.62973f
C14948 VDD.n5752 GND 0.02746f
C14949 VDD.t755 GND 0.02334f
C14950 VDD.t464 GND 0.02334f
C14951 VDD.n5753 GND 0.13341f
C14952 VDD.t917 GND 0.02334f
C14953 VDD.t142 GND 0.02321f
C14954 VDD.t424 GND 0.02321f
C14955 VDD.n5754 GND 0.10855f
C14956 VDD.t372 GND 0.02321f
C14957 VDD.t264 GND 0.02321f
C14958 VDD.n5755 GND 0.10855f
C14959 VDD.n5756 GND 0.04152f
C14960 VDD.n5757 GND 0.0536f
C14961 VDD.n5758 GND 0.05074f
C14962 VDD.n5759 GND 0.0536f
C14963 VDD.n5760 GND 0.04999f
C14964 VDD.n5761 GND 0.04999f
C14965 VDD.n5762 GND 0.68843f
C14966 VDD.n5763 GND 0.02522f
C14967 VDD.n5764 GND 0.02522f
C14968 VDD.n5765 GND 0.02967f
C14969 VDD.n5766 GND 0.05074f
C14970 VDD.n5767 GND 0.04999f
C14971 VDD.t263 GND 0.63568f
C14972 VDD.n5768 GND 0.05074f
C14973 VDD.n5769 GND 0.05074f
C14974 VDD.n5770 GND 0.02967f
C14975 VDD.n5771 GND 0.02522f
C14976 VDD.n5772 GND 0.03166f
C14977 VDD.n5773 GND 0.0536f
C14978 VDD.n5774 GND 0.05074f
C14979 VDD.n5775 GND 0.02967f
C14980 VDD.n5776 GND 0.02522f
C14981 VDD.n5777 GND 0.04999f
C14982 VDD.t435 GND 0.63568f
C14983 VDD.n5778 GND 0.05074f
C14984 VDD.n5779 GND 0.05074f
C14985 VDD.n5780 GND 0.02967f
C14986 VDD.n5781 GND 0.02522f
C14987 VDD.n5782 GND 0.0263f
C14988 VDD.n5783 GND 0.0536f
C14989 VDD.n5784 GND 0.05074f
C14990 VDD.n5785 GND 0.02967f
C14991 VDD.n5786 GND 0.02522f
C14992 VDD.n5787 GND 0.04999f
C14993 VDD.t827 GND 0.63568f
C14994 VDD.n5788 GND 0.05074f
C14995 VDD.n5789 GND 0.05074f
C14996 VDD.n5790 GND 0.02967f
C14997 VDD.n5791 GND 0.02522f
C14998 VDD.t436 GND 0.02334f
C14999 VDD.t705 GND 0.02334f
C15000 VDD.n5792 GND 0.13341f
C15001 VDD.n5793 GND 0.02334f
C15002 VDD.n5794 GND 0.0536f
C15003 VDD.n5795 GND 0.05074f
C15004 VDD.n5796 GND 0.02967f
C15005 VDD.n5797 GND 0.02522f
C15006 VDD.n5798 GND 0.04999f
C15007 VDD.t944 GND 0.63568f
C15008 VDD.n5799 GND 0.05074f
C15009 VDD.n5800 GND 0.05074f
C15010 VDD.n5801 GND 0.02967f
C15011 VDD.n5802 GND 0.02522f
C15012 VDD.t829 GND 0.02321f
C15013 VDD.t987 GND 0.02321f
C15014 VDD.n5803 GND 0.10855f
C15015 VDD.t828 GND 0.02321f
C15016 VDD.t945 GND 0.02321f
C15017 VDD.n5804 GND 0.10855f
C15018 VDD.n5805 GND 0.04152f
C15019 VDD.n5806 GND 0.02334f
C15020 VDD.n5807 GND 0.0536f
C15021 VDD.n5808 GND 0.05074f
C15022 VDD.n5809 GND 0.02967f
C15023 VDD.n5810 GND 0.02522f
C15024 VDD.t1079 GND 0.63568f
C15025 VDD.n5811 GND 0.05074f
C15026 VDD.n5812 GND 0.05074f
C15027 VDD.n5813 GND 0.09132f
C15028 VDD.n5814 GND 0.04999f
C15029 VDD.t632 GND 0.63568f
C15030 VDD.n5815 GND 0.05074f
C15031 VDD.n5816 GND 0.05074f
C15032 VDD.n5817 GND 0.02967f
C15033 VDD.n5818 GND 0.02522f
C15034 VDD.t1080 GND 0.02334f
C15035 VDD.n5819 GND 0.01798f
C15036 VDD.n5820 GND 0.0731f
C15037 VDD.n5821 GND 0.02334f
C15038 VDD.n5822 GND 0.0536f
C15039 VDD.n5823 GND 0.05074f
C15040 VDD.n5824 GND 0.02967f
C15041 VDD.n5825 GND 0.02522f
C15042 VDD.n5826 GND 0.04999f
C15043 VDD.t187 GND 0.63568f
C15044 VDD.n5827 GND 0.05074f
C15045 VDD.n5828 GND 0.05074f
C15046 VDD.n5829 GND 0.02967f
C15047 VDD.n5830 GND 0.02522f
C15048 VDD.t946 GND 0.02321f
C15049 VDD.t188 GND 0.02321f
C15050 VDD.n5831 GND 0.10855f
C15051 VDD.t633 GND 0.02321f
C15052 VDD.t978 GND 0.02321f
C15053 VDD.n5832 GND 0.10855f
C15054 VDD.n5833 GND 0.04152f
C15055 VDD.n5834 GND 0.03166f
C15056 VDD.n5835 GND 0.0536f
C15057 VDD.n5836 GND 0.05074f
C15058 VDD.n5837 GND 0.02967f
C15059 VDD.n5838 GND 0.02522f
C15060 VDD.n5839 GND 0.04999f
C15061 VDD.t471 GND 0.63568f
C15062 VDD.n5840 GND 0.05074f
C15063 VDD.n5841 GND 0.05074f
C15064 VDD.n5842 GND 0.02967f
C15065 VDD.n5843 GND 0.02522f
C15066 VDD.n5844 GND 0.0263f
C15067 VDD.n5845 GND 0.0536f
C15068 VDD.n5846 GND 0.05074f
C15069 VDD.n5847 GND 0.02967f
C15070 VDD.n5848 GND 0.02522f
C15071 VDD.n5849 GND 0.04999f
C15072 VDD.t1056 GND 0.63568f
C15073 VDD.n5850 GND 0.05074f
C15074 VDD.n5851 GND 0.05074f
C15075 VDD.n5852 GND 0.02967f
C15076 VDD.n5853 GND 0.02522f
C15077 VDD.t472 GND 0.02334f
C15078 VDD.t741 GND 0.02334f
C15079 VDD.n5854 GND 0.13341f
C15080 VDD.n5855 GND 0.02334f
C15081 VDD.n5856 GND 0.0536f
C15082 VDD.n5857 GND 0.05074f
C15083 VDD.n5858 GND 0.02967f
C15084 VDD.n5859 GND 0.02522f
C15085 VDD.n5860 GND 0.04999f
C15086 VDD.t341 GND 0.63568f
C15087 VDD.n5861 GND 0.05074f
C15088 VDD.n5862 GND 0.05074f
C15089 VDD.n5863 GND 0.02967f
C15090 VDD.n5864 GND 0.02522f
C15091 VDD.t1057 GND 0.02321f
C15092 VDD.t342 GND 0.02321f
C15093 VDD.n5865 GND 0.10855f
C15094 VDD.t1088 GND 0.02321f
C15095 VDD.t414 GND 0.02321f
C15096 VDD.n5866 GND 0.10855f
C15097 VDD.n5867 GND 0.04152f
C15098 VDD.n5868 GND 0.03166f
C15099 VDD.n5869 GND 0.0536f
C15100 VDD.n5870 GND 0.05074f
C15101 VDD.n5871 GND 0.02967f
C15102 VDD.n5872 GND 0.02522f
C15103 VDD.n5873 GND 0.04999f
C15104 VDD.t516 GND 0.63568f
C15105 VDD.n5874 GND 0.05074f
C15106 VDD.n5875 GND 0.05074f
C15107 VDD.n5876 GND 0.02967f
C15108 VDD.n5877 GND 0.02522f
C15109 VDD.n5878 GND 0.0263f
C15110 VDD.n5879 GND 0.0536f
C15111 VDD.n5880 GND 0.05074f
C15112 VDD.n5881 GND 0.02967f
C15113 VDD.n5882 GND 0.02522f
C15114 VDD.t881 GND 0.74438f
C15115 VDD.n5883 GND 0.05074f
C15116 VDD.n5884 GND 0.05074f
C15117 VDD.n5885 GND 0.02967f
C15118 VDD.n5887 GND 0.62973f
C15119 VDD.n5888 GND 0.02746f
C15120 VDD.t709 GND 0.02334f
C15121 VDD.t517 GND 0.02334f
C15122 VDD.n5889 GND 0.13341f
C15123 VDD.t882 GND 0.02334f
C15124 VDD.t819 GND 0.02321f
C15125 VDD.t38 GND 0.02321f
C15126 VDD.n5890 GND 0.10855f
C15127 VDD.t246 GND 0.02321f
C15128 VDD.t411 GND 0.02321f
C15129 VDD.n5891 GND 0.10855f
C15130 VDD.n5892 GND 0.04152f
C15131 VDD.n5893 GND 0.0536f
C15132 VDD.n5894 GND 0.05074f
C15133 VDD.n5895 GND 0.0536f
C15134 VDD.n5896 GND 0.04999f
C15135 VDD.n5897 GND 0.04999f
C15136 VDD.n5898 GND 0.68843f
C15137 VDD.n5899 GND 0.02522f
C15138 VDD.n5900 GND 0.02522f
C15139 VDD.n5901 GND 0.02967f
C15140 VDD.n5902 GND 0.05074f
C15141 VDD.n5903 GND 0.04999f
C15142 VDD.t37 GND 0.63568f
C15143 VDD.n5904 GND 0.05074f
C15144 VDD.n5905 GND 0.05074f
C15145 VDD.n5906 GND 0.02967f
C15146 VDD.n5907 GND 0.02522f
C15147 VDD.n5908 GND 0.03166f
C15148 VDD.n5909 GND 0.0536f
C15149 VDD.n5910 GND 0.05074f
C15150 VDD.n5911 GND 0.02967f
C15151 VDD.n5912 GND 0.02522f
C15152 VDD.n5913 GND 0.04999f
C15153 VDD.t530 GND 0.63568f
C15154 VDD.n5914 GND 0.05074f
C15155 VDD.n5915 GND 0.05074f
C15156 VDD.n5916 GND 0.02967f
C15157 VDD.n5917 GND 0.02522f
C15158 VDD.n5918 GND 0.0263f
C15159 VDD.n5919 GND 0.0536f
C15160 VDD.n5920 GND 0.05074f
C15161 VDD.n5921 GND 0.02967f
C15162 VDD.n5922 GND 0.02522f
C15163 VDD.n5923 GND 0.04999f
C15164 VDD.t56 GND 0.63568f
C15165 VDD.n5924 GND 0.05074f
C15166 VDD.n5925 GND 0.05074f
C15167 VDD.n5926 GND 0.02967f
C15168 VDD.n5927 GND 0.02522f
C15169 VDD.t727 GND 0.02334f
C15170 VDD.t531 GND 0.02334f
C15171 VDD.n5928 GND 0.13341f
C15172 VDD.n5929 GND 0.02334f
C15173 VDD.n5930 GND 0.0536f
C15174 VDD.n5931 GND 0.05074f
C15175 VDD.n5932 GND 0.02967f
C15176 VDD.n5933 GND 0.02522f
C15177 VDD.n5934 GND 0.04999f
C15178 VDD.t322 GND 0.63568f
C15179 VDD.n5935 GND 0.05074f
C15180 VDD.n5936 GND 0.05074f
C15181 VDD.n5937 GND 0.02967f
C15182 VDD.n5938 GND 0.02522f
C15183 VDD.t295 GND 0.02321f
C15184 VDD.t973 GND 0.02321f
C15185 VDD.n5939 GND 0.10855f
C15186 VDD.t57 GND 0.02321f
C15187 VDD.t323 GND 0.02321f
C15188 VDD.n5940 GND 0.10855f
C15189 VDD.n5941 GND 0.04152f
C15190 VDD.n5942 GND 0.02334f
C15191 VDD.n5943 GND 0.0536f
C15192 VDD.n5944 GND 0.05074f
C15193 VDD.n5945 GND 0.02967f
C15194 VDD.n5946 GND 0.02522f
C15195 VDD.t1024 GND 0.63568f
C15196 VDD.n5947 GND 0.05074f
C15197 VDD.n5948 GND 0.05074f
C15198 VDD.n5949 GND 0.09132f
C15199 VDD.n5950 GND 0.04999f
C15200 VDD.t324 GND 0.63568f
C15201 VDD.n5951 GND 0.05074f
C15202 VDD.n5952 GND 0.05074f
C15203 VDD.n5953 GND 0.02967f
C15204 VDD.n5954 GND 0.02522f
C15205 VDD.t1025 GND 0.02334f
C15206 VDD.n5955 GND 0.01798f
C15207 VDD.n5956 GND 0.0731f
C15208 VDD.n5957 GND 0.02334f
C15209 VDD.n5958 GND 0.0536f
C15210 VDD.n5959 GND 0.05074f
C15211 VDD.n5960 GND 0.02967f
C15212 VDD.n5961 GND 0.02522f
C15213 VDD.n5962 GND 0.04999f
C15214 VDD.t202 GND 0.63568f
C15215 VDD.n5963 GND 0.05074f
C15216 VDD.n5964 GND 0.05074f
C15217 VDD.n5965 GND 0.02967f
C15218 VDD.n5966 GND 0.02522f
C15219 VDD.t325 GND 0.02321f
C15220 VDD.t203 GND 0.02321f
C15221 VDD.n5967 GND 0.10855f
C15222 VDD.t974 GND 0.02321f
C15223 VDD.t860 GND 0.02321f
C15224 VDD.n5968 GND 0.10855f
C15225 VDD.n5969 GND 0.04152f
C15226 VDD.n5970 GND 0.03166f
C15227 VDD.n5971 GND 0.0536f
C15228 VDD.n5972 GND 0.05074f
C15229 VDD.n5973 GND 0.02967f
C15230 VDD.n5974 GND 0.02522f
C15231 VDD.n5975 GND 0.04999f
C15232 VDD.t534 GND 0.63568f
C15233 VDD.n5976 GND 0.05074f
C15234 VDD.n5977 GND 0.05074f
C15235 VDD.n5978 GND 0.02967f
C15236 VDD.n5979 GND 0.02522f
C15237 VDD.n5980 GND 0.0263f
C15238 VDD.n5981 GND 0.0536f
C15239 VDD.n5982 GND 0.05074f
C15240 VDD.n5983 GND 0.02967f
C15241 VDD.n5984 GND 0.02522f
C15242 VDD.n5985 GND 0.04999f
C15243 VDD.t1000 GND 0.63568f
C15244 VDD.n5986 GND 0.05074f
C15245 VDD.n5987 GND 0.05074f
C15246 VDD.n5988 GND 0.02967f
C15247 VDD.n5989 GND 0.02522f
C15248 VDD.t729 GND 0.02334f
C15249 VDD.t535 GND 0.02334f
C15250 VDD.n5990 GND 0.13341f
C15251 VDD.n5991 GND 0.02334f
C15252 VDD.n5992 GND 0.0536f
C15253 VDD.n5993 GND 0.05074f
C15254 VDD.n5994 GND 0.02967f
C15255 VDD.n5995 GND 0.02522f
C15256 VDD.n5996 GND 0.04999f
C15257 VDD.t185 GND 0.63568f
C15258 VDD.n5997 GND 0.05074f
C15259 VDD.n5998 GND 0.05074f
C15260 VDD.n5999 GND 0.02967f
C15261 VDD.n6000 GND 0.02522f
C15262 VDD.t1001 GND 0.02321f
C15263 VDD.t887 GND 0.02321f
C15264 VDD.n6001 GND 0.10855f
C15265 VDD.t1044 GND 0.02321f
C15266 VDD.t186 GND 0.02321f
C15267 VDD.n6002 GND 0.10855f
C15268 VDD.n6003 GND 0.04152f
C15269 VDD.n6004 GND 0.03166f
C15270 VDD.n6005 GND 0.0536f
C15271 VDD.n6006 GND 0.05074f
C15272 VDD.n6007 GND 0.02967f
C15273 VDD.n6008 GND 0.02522f
C15274 VDD.n6009 GND 0.04999f
C15275 VDD.t494 GND 0.63568f
C15276 VDD.n6010 GND 0.05074f
C15277 VDD.n6011 GND 0.05074f
C15278 VDD.n6012 GND 0.02967f
C15279 VDD.n6013 GND 0.02522f
C15280 VDD.n6014 GND 0.0263f
C15281 VDD.n6015 GND 0.0536f
C15282 VDD.n6016 GND 0.05074f
C15283 VDD.n6017 GND 0.02967f
C15284 VDD.n6018 GND 0.02522f
C15285 VDD.t888 GND 0.74438f
C15286 VDD.n6019 GND 0.05074f
C15287 VDD.n6020 GND 0.05074f
C15288 VDD.n6021 GND 0.02967f
C15289 VDD.n6023 GND 0.62973f
C15290 VDD.n6024 GND 0.02746f
C15291 VDD.t495 GND 0.02334f
C15292 VDD.t667 GND 0.02334f
C15293 VDD.n6025 GND 0.13341f
C15294 VDD.t889 GND 0.02334f
C15295 VDD.n6026 GND 0.0731f
C15296 VDD.n6027 GND 0.01798f
C15297 VDD.n6028 GND 0.09132f
C15298 VDD.n6029 GND 0.02746f
C15299 VDD.n6030 GND 0.04999f
C15300 VDD.n6031 GND 0.68843f
C15301 VDD.n6032 GND 0.02522f
C15302 VDD.n6033 GND 0.04999f
C15303 VDD.n6034 GND 0.68843f
C15304 VDD.n6035 GND 0.04999f
C15305 VDD.n6036 GND 0.05074f
C15306 VDD.n6037 GND 0.06295f
C15307 VDD.n6038 GND 0.0536f
C15308 VDD.n6039 GND 0.02522f
C15309 VDD.n6040 GND 0.04999f
C15310 VDD.n6041 GND 0.5126f
C15311 VDD.n6042 GND 0.02522f
C15312 VDD.n6043 GND 0.04999f
C15313 VDD.n6044 GND 0.5126f
C15314 VDD.n6045 GND 0.04999f
C15315 VDD.n6046 GND 0.05074f
C15316 VDD.n6047 GND 0.06295f
C15317 VDD.n6048 GND 0.0536f
C15318 VDD.n6049 GND 0.02522f
C15319 VDD.n6050 GND 0.04999f
C15320 VDD.n6051 GND 0.5126f
C15321 VDD.n6052 GND 0.02522f
C15322 VDD.n6053 GND 0.04999f
C15323 VDD.n6054 GND 0.5126f
C15324 VDD.n6055 GND 0.04999f
C15325 VDD.n6056 GND 0.05074f
C15326 VDD.n6057 GND 0.06295f
C15327 VDD.n6058 GND 0.0536f
C15328 VDD.n6059 GND 0.02522f
C15329 VDD.n6060 GND 0.04999f
C15330 VDD.n6061 GND 0.68843f
C15331 VDD.n6062 GND 0.02522f
C15332 VDD.n6063 GND 0.04999f
C15333 VDD.n6064 GND 0.68843f
C15334 VDD.n6065 GND 0.04999f
C15335 VDD.n6066 GND 0.05074f
C15336 VDD.n6067 GND 0.06295f
C15337 VDD.n6068 GND 0.0536f
C15338 VDD.n6069 GND 0.02522f
C15339 VDD.n6070 GND 0.04999f
C15340 VDD.n6071 GND 0.5126f
C15341 VDD.n6072 GND 0.02522f
C15342 VDD.n6073 GND 0.04999f
C15343 VDD.n6074 GND 0.5126f
C15344 VDD.n6075 GND 0.04999f
C15345 VDD.n6076 GND 0.05074f
C15346 VDD.n6077 GND 0.06295f
C15347 VDD.n6078 GND 0.0536f
C15348 VDD.n6079 GND 0.02522f
C15349 VDD.n6080 GND 0.04999f
C15350 VDD.n6081 GND 0.5126f
C15351 VDD.n6082 GND 0.02522f
C15352 VDD.n6083 GND 0.04999f
C15353 VDD.n6084 GND 0.5126f
C15354 VDD.n6085 GND 0.04999f
C15355 VDD.n6086 GND 0.05074f
C15356 VDD.n6087 GND 0.06295f
C15357 VDD.n6088 GND 0.0536f
C15358 VDD.n6089 GND 0.02522f
C15359 VDD.n6090 GND 0.04999f
C15360 VDD.n6091 GND 0.68843f
C15361 VDD.n6092 GND 0.68843f
C15362 VDD.n6093 GND 0.04999f
C15363 VDD.n6094 GND 0.02746f
C15364 VDD.n6095 GND 0.02967f
C15365 VDD.n6096 GND 0.02746f
C15366 VDD.n6097 GND 0.04999f
C15367 VDD.n6098 GND 0.68843f
C15368 VDD.n6099 GND 0.02522f
C15369 VDD.n6100 GND 0.04999f
C15370 VDD.n6101 GND 0.68843f
C15371 VDD.n6102 GND 0.04999f
C15372 VDD.n6103 GND 0.05074f
C15373 VDD.n6104 GND 0.06295f
C15374 VDD.n6105 GND 0.0536f
C15375 VDD.n6106 GND 0.02522f
C15376 VDD.n6107 GND 0.04999f
C15377 VDD.n6108 GND 0.5126f
C15378 VDD.n6109 GND 0.02522f
C15379 VDD.n6110 GND 0.04999f
C15380 VDD.n6111 GND 0.5126f
C15381 VDD.n6112 GND 0.04999f
C15382 VDD.n6113 GND 0.05074f
C15383 VDD.n6114 GND 0.06295f
C15384 VDD.n6115 GND 0.0536f
C15385 VDD.n6116 GND 0.02522f
C15386 VDD.n6117 GND 0.04999f
C15387 VDD.n6118 GND 0.68843f
C15388 VDD.n6119 GND 0.02522f
C15389 VDD.n6120 GND 0.04999f
C15390 VDD.n6121 GND 0.68843f
C15391 VDD.n6122 GND 0.04999f
C15392 VDD.n6123 GND 0.05074f
C15393 VDD.n6124 GND 0.06295f
C15394 VDD.n6125 GND 0.0536f
C15395 VDD.n6126 GND 0.02522f
C15396 VDD.n6127 GND 0.04999f
C15397 VDD.n6128 GND 0.5126f
C15398 VDD.n6129 GND 0.02522f
C15399 VDD.n6130 GND 0.04999f
C15400 VDD.n6131 GND 0.5126f
C15401 VDD.n6132 GND 0.04999f
C15402 VDD.n6133 GND 0.05074f
C15403 VDD.n6134 GND 0.06295f
C15404 VDD.n6135 GND 0.0536f
C15405 VDD.n6136 GND 0.02522f
C15406 VDD.n6137 GND 0.04999f
C15407 VDD.n6138 GND 0.5126f
C15408 VDD.n6139 GND 0.5126f
C15409 VDD.n6140 GND 0.04999f
C15410 VDD.n6141 GND 0.04999f
C15411 VDD.n6142 GND 0.02522f
C15412 VDD.n6143 GND 0.02522f
C15413 VDD.n6144 GND 0.02967f
C15414 VDD.n6145 GND 0.05074f
C15415 VDD.t245 GND 0.63568f
C15416 VDD.n6146 GND 0.05074f
C15417 VDD.n6147 GND 0.06295f
C15418 VDD.n6148 GND 0.10164f
C15419 VDD.n6149 GND 0.0731f
C15420 VDD.n6150 GND 0.01798f
C15421 VDD.n6151 GND 0.09132f
C15422 VDD.n6152 GND 0.02746f
C15423 VDD.n6153 GND 0.04999f
C15424 VDD.n6154 GND 0.68843f
C15425 VDD.n6155 GND 0.02522f
C15426 VDD.n6156 GND 0.04999f
C15427 VDD.n6157 GND 0.68843f
C15428 VDD.n6158 GND 0.04999f
C15429 VDD.n6159 GND 0.05074f
C15430 VDD.n6160 GND 0.06295f
C15431 VDD.n6161 GND 0.0536f
C15432 VDD.n6162 GND 0.02522f
C15433 VDD.n6163 GND 0.04999f
C15434 VDD.n6164 GND 0.5126f
C15435 VDD.n6165 GND 0.02522f
C15436 VDD.n6166 GND 0.04999f
C15437 VDD.n6167 GND 0.5126f
C15438 VDD.n6168 GND 0.04999f
C15439 VDD.n6169 GND 0.05074f
C15440 VDD.n6170 GND 0.06295f
C15441 VDD.n6171 GND 0.0536f
C15442 VDD.n6172 GND 0.02522f
C15443 VDD.n6173 GND 0.04999f
C15444 VDD.n6174 GND 0.5126f
C15445 VDD.n6175 GND 0.02522f
C15446 VDD.n6176 GND 0.04999f
C15447 VDD.n6177 GND 0.5126f
C15448 VDD.n6178 GND 0.04999f
C15449 VDD.n6179 GND 0.05074f
C15450 VDD.n6180 GND 0.06295f
C15451 VDD.n6181 GND 0.0536f
C15452 VDD.n6182 GND 0.02522f
C15453 VDD.n6183 GND 0.04999f
C15454 VDD.n6184 GND 0.68843f
C15455 VDD.n6185 GND 0.02522f
C15456 VDD.n6186 GND 0.04999f
C15457 VDD.n6187 GND 0.68843f
C15458 VDD.n6188 GND 0.04999f
C15459 VDD.n6189 GND 0.05074f
C15460 VDD.n6190 GND 0.06295f
C15461 VDD.n6191 GND 0.0536f
C15462 VDD.n6192 GND 0.02522f
C15463 VDD.n6193 GND 0.04999f
C15464 VDD.n6194 GND 0.5126f
C15465 VDD.n6195 GND 0.02522f
C15466 VDD.n6196 GND 0.04999f
C15467 VDD.n6197 GND 0.5126f
C15468 VDD.n6198 GND 0.04999f
C15469 VDD.n6199 GND 0.05074f
C15470 VDD.n6200 GND 0.06295f
C15471 VDD.n6201 GND 0.0536f
C15472 VDD.n6202 GND 0.02522f
C15473 VDD.n6203 GND 0.04999f
C15474 VDD.n6204 GND 0.5126f
C15475 VDD.n6205 GND 0.02522f
C15476 VDD.n6206 GND 0.04999f
C15477 VDD.n6207 GND 0.5126f
C15478 VDD.n6208 GND 0.04999f
C15479 VDD.n6209 GND 0.05074f
C15480 VDD.n6210 GND 0.06295f
C15481 VDD.n6211 GND 0.0536f
C15482 VDD.n6212 GND 0.02522f
C15483 VDD.n6213 GND 0.04999f
C15484 VDD.n6214 GND 0.68843f
C15485 VDD.n6215 GND 0.68843f
C15486 VDD.n6216 GND 0.04999f
C15487 VDD.n6217 GND 0.02746f
C15488 VDD.n6218 GND 0.02967f
C15489 VDD.n6219 GND 0.02746f
C15490 VDD.n6220 GND 0.04999f
C15491 VDD.n6221 GND 0.68843f
C15492 VDD.n6222 GND 0.02522f
C15493 VDD.n6223 GND 0.04999f
C15494 VDD.n6224 GND 0.68843f
C15495 VDD.n6225 GND 0.04999f
C15496 VDD.n6226 GND 0.05074f
C15497 VDD.n6227 GND 0.06295f
C15498 VDD.n6228 GND 0.0536f
C15499 VDD.n6229 GND 0.02522f
C15500 VDD.n6230 GND 0.04999f
C15501 VDD.n6231 GND 0.5126f
C15502 VDD.n6232 GND 0.02522f
C15503 VDD.n6233 GND 0.04999f
C15504 VDD.n6234 GND 0.5126f
C15505 VDD.n6235 GND 0.04999f
C15506 VDD.n6236 GND 0.05074f
C15507 VDD.n6237 GND 0.06295f
C15508 VDD.n6238 GND 0.0536f
C15509 VDD.n6239 GND 0.02522f
C15510 VDD.n6240 GND 0.04999f
C15511 VDD.n6241 GND 0.68843f
C15512 VDD.n6242 GND 0.02522f
C15513 VDD.n6243 GND 0.04999f
C15514 VDD.n6244 GND 0.68843f
C15515 VDD.n6245 GND 0.04999f
C15516 VDD.n6246 GND 0.05074f
C15517 VDD.n6247 GND 0.06295f
C15518 VDD.n6248 GND 0.0536f
C15519 VDD.n6249 GND 0.02522f
C15520 VDD.n6250 GND 0.04999f
C15521 VDD.n6251 GND 0.5126f
C15522 VDD.n6252 GND 0.02522f
C15523 VDD.n6253 GND 0.04999f
C15524 VDD.n6254 GND 0.5126f
C15525 VDD.n6255 GND 0.04999f
C15526 VDD.n6256 GND 0.05074f
C15527 VDD.n6257 GND 0.06295f
C15528 VDD.n6258 GND 0.0536f
C15529 VDD.n6259 GND 0.02522f
C15530 VDD.n6260 GND 0.04999f
C15531 VDD.n6261 GND 0.5126f
C15532 VDD.n6262 GND 0.5126f
C15533 VDD.n6263 GND 0.04999f
C15534 VDD.n6264 GND 0.04999f
C15535 VDD.n6265 GND 0.02522f
C15536 VDD.n6266 GND 0.02522f
C15537 VDD.n6267 GND 0.02967f
C15538 VDD.n6268 GND 0.05074f
C15539 VDD.t141 GND 0.63568f
C15540 VDD.n6269 GND 0.05074f
C15541 VDD.n6270 GND 0.06295f
C15542 VDD.n6271 GND 0.10164f
C15543 VDD.n6272 GND 0.0731f
C15544 VDD.n6273 GND 0.01798f
C15545 VDD.n6274 GND 0.09132f
C15546 VDD.n6275 GND 0.02746f
C15547 VDD.n6276 GND 0.04999f
C15548 VDD.n6277 GND 0.68843f
C15549 VDD.n6278 GND 0.02522f
C15550 VDD.n6279 GND 0.04999f
C15551 VDD.n6280 GND 0.68843f
C15552 VDD.n6281 GND 0.04999f
C15553 VDD.n6282 GND 0.05074f
C15554 VDD.n6283 GND 0.06295f
C15555 VDD.n6284 GND 0.0536f
C15556 VDD.n6285 GND 0.02522f
C15557 VDD.n6286 GND 0.04999f
C15558 VDD.n6287 GND 0.5126f
C15559 VDD.n6288 GND 0.02522f
C15560 VDD.n6289 GND 0.04999f
C15561 VDD.n6290 GND 0.5126f
C15562 VDD.n6291 GND 0.04999f
C15563 VDD.n6292 GND 0.05074f
C15564 VDD.n6293 GND 0.06295f
C15565 VDD.n6294 GND 0.0536f
C15566 VDD.n6295 GND 0.02522f
C15567 VDD.n6296 GND 0.04999f
C15568 VDD.n6297 GND 0.5126f
C15569 VDD.n6298 GND 0.02522f
C15570 VDD.n6299 GND 0.04999f
C15571 VDD.n6300 GND 0.5126f
C15572 VDD.n6301 GND 0.04999f
C15573 VDD.n6302 GND 0.05074f
C15574 VDD.n6303 GND 0.06295f
C15575 VDD.n6304 GND 0.0536f
C15576 VDD.n6305 GND 0.02522f
C15577 VDD.n6306 GND 0.04999f
C15578 VDD.n6307 GND 0.68843f
C15579 VDD.n6308 GND 0.02522f
C15580 VDD.n6309 GND 0.04999f
C15581 VDD.n6310 GND 0.68843f
C15582 VDD.n6311 GND 0.04999f
C15583 VDD.n6312 GND 0.05074f
C15584 VDD.n6313 GND 0.06295f
C15585 VDD.n6314 GND 0.0536f
C15586 VDD.n6315 GND 0.02522f
C15587 VDD.n6316 GND 0.04999f
C15588 VDD.n6317 GND 0.5126f
C15589 VDD.n6318 GND 0.02522f
C15590 VDD.n6319 GND 0.04999f
C15591 VDD.n6320 GND 0.5126f
C15592 VDD.n6321 GND 0.04999f
C15593 VDD.n6322 GND 0.05074f
C15594 VDD.n6323 GND 0.06295f
C15595 VDD.n6324 GND 0.0536f
C15596 VDD.n6325 GND 0.02522f
C15597 VDD.n6326 GND 0.04999f
C15598 VDD.n6327 GND 0.5126f
C15599 VDD.n6328 GND 0.02522f
C15600 VDD.n6329 GND 0.04999f
C15601 VDD.n6330 GND 0.5126f
C15602 VDD.n6331 GND 0.04999f
C15603 VDD.n6332 GND 0.05074f
C15604 VDD.n6333 GND 0.06295f
C15605 VDD.n6334 GND 0.0536f
C15606 VDD.n6335 GND 0.02522f
C15607 VDD.n6336 GND 0.04999f
C15608 VDD.n6337 GND 0.68843f
C15609 VDD.n6338 GND 0.68843f
C15610 VDD.n6339 GND 0.04999f
C15611 VDD.n6340 GND 0.02746f
C15612 VDD.n6341 GND 0.02967f
C15613 VDD.n6342 GND 0.02746f
C15614 VDD.n6343 GND 0.04999f
C15615 VDD.n6344 GND 0.68843f
C15616 VDD.n6345 GND 0.02522f
C15617 VDD.n6346 GND 0.04999f
C15618 VDD.n6347 GND 0.68843f
C15619 VDD.n6348 GND 0.04999f
C15620 VDD.n6349 GND 0.05074f
C15621 VDD.n6350 GND 0.06295f
C15622 VDD.n6351 GND 0.0536f
C15623 VDD.n6352 GND 0.02522f
C15624 VDD.n6353 GND 0.04999f
C15625 VDD.n6354 GND 0.5126f
C15626 VDD.n6355 GND 0.02522f
C15627 VDD.n6356 GND 0.04999f
C15628 VDD.n6357 GND 0.5126f
C15629 VDD.n6358 GND 0.04999f
C15630 VDD.n6359 GND 0.05074f
C15631 VDD.n6360 GND 0.06295f
C15632 VDD.n6361 GND 0.0536f
C15633 VDD.n6362 GND 0.02522f
C15634 VDD.n6363 GND 0.04999f
C15635 VDD.n6364 GND 0.68843f
C15636 VDD.n6365 GND 0.02522f
C15637 VDD.n6366 GND 0.04999f
C15638 VDD.n6367 GND 0.68843f
C15639 VDD.n6368 GND 0.04999f
C15640 VDD.n6369 GND 0.05074f
C15641 VDD.n6370 GND 0.06295f
C15642 VDD.n6371 GND 0.0536f
C15643 VDD.n6372 GND 0.02522f
C15644 VDD.n6373 GND 0.04999f
C15645 VDD.n6374 GND 0.5126f
C15646 VDD.n6375 GND 0.02522f
C15647 VDD.n6376 GND 0.04999f
C15648 VDD.n6377 GND 0.5126f
C15649 VDD.n6378 GND 0.04999f
C15650 VDD.n6379 GND 0.05074f
C15651 VDD.n6380 GND 0.06295f
C15652 VDD.n6381 GND 0.0536f
C15653 VDD.n6382 GND 0.02522f
C15654 VDD.n6383 GND 0.04999f
C15655 VDD.n6384 GND 0.5126f
C15656 VDD.n6385 GND 0.5126f
C15657 VDD.n6386 GND 0.04999f
C15658 VDD.n6387 GND 0.04999f
C15659 VDD.n6388 GND 0.02522f
C15660 VDD.n6389 GND 0.02522f
C15661 VDD.n6390 GND 0.02967f
C15662 VDD.n6391 GND 0.05074f
C15663 VDD.t364 GND 0.63568f
C15664 VDD.n6392 GND 0.05074f
C15665 VDD.n6393 GND 0.06295f
C15666 VDD.n6394 GND 0.10164f
C15667 VDD.n6395 GND 0.0731f
C15668 VDD.n6396 GND 0.01798f
C15669 VDD.n6397 GND 0.09132f
C15670 VDD.n6398 GND 0.02746f
C15671 VDD.n6399 GND 0.04999f
C15672 VDD.n6400 GND 0.68843f
C15673 VDD.n6401 GND 0.02522f
C15674 VDD.n6402 GND 0.04999f
C15675 VDD.n6403 GND 0.68843f
C15676 VDD.n6404 GND 0.04999f
C15677 VDD.n6405 GND 0.05074f
C15678 VDD.n6406 GND 0.06295f
C15679 VDD.n6407 GND 0.0536f
C15680 VDD.n6408 GND 0.02522f
C15681 VDD.n6409 GND 0.04999f
C15682 VDD.n6410 GND 0.5126f
C15683 VDD.n6411 GND 0.02522f
C15684 VDD.n6412 GND 0.04999f
C15685 VDD.n6413 GND 0.5126f
C15686 VDD.n6414 GND 0.04999f
C15687 VDD.n6415 GND 0.05074f
C15688 VDD.n6416 GND 0.06295f
C15689 VDD.n6417 GND 0.0536f
C15690 VDD.n6418 GND 0.02522f
C15691 VDD.n6419 GND 0.04999f
C15692 VDD.n6420 GND 0.5126f
C15693 VDD.n6421 GND 0.02522f
C15694 VDD.n6422 GND 0.04999f
C15695 VDD.n6423 GND 0.5126f
C15696 VDD.n6424 GND 0.04999f
C15697 VDD.n6425 GND 0.05074f
C15698 VDD.n6426 GND 0.06295f
C15699 VDD.n6427 GND 0.0536f
C15700 VDD.n6428 GND 0.02522f
C15701 VDD.n6429 GND 0.04999f
C15702 VDD.n6430 GND 0.68843f
C15703 VDD.n6431 GND 0.02522f
C15704 VDD.n6432 GND 0.04999f
C15705 VDD.n6433 GND 0.68843f
C15706 VDD.n6434 GND 0.04999f
C15707 VDD.n6435 GND 0.05074f
C15708 VDD.n6436 GND 0.06295f
C15709 VDD.n6437 GND 0.0536f
C15710 VDD.n6438 GND 0.02522f
C15711 VDD.n6439 GND 0.04999f
C15712 VDD.n6440 GND 0.5126f
C15713 VDD.n6441 GND 0.02522f
C15714 VDD.n6442 GND 0.04999f
C15715 VDD.n6443 GND 0.5126f
C15716 VDD.n6444 GND 0.04999f
C15717 VDD.n6445 GND 0.05074f
C15718 VDD.n6446 GND 0.06295f
C15719 VDD.n6447 GND 0.0536f
C15720 VDD.n6448 GND 0.02522f
C15721 VDD.n6449 GND 0.04999f
C15722 VDD.n6450 GND 0.5126f
C15723 VDD.n6451 GND 0.02522f
C15724 VDD.n6452 GND 0.04999f
C15725 VDD.n6453 GND 0.5126f
C15726 VDD.n6454 GND 0.04999f
C15727 VDD.n6455 GND 0.05074f
C15728 VDD.n6456 GND 0.06295f
C15729 VDD.n6457 GND 0.0536f
C15730 VDD.n6458 GND 0.02522f
C15731 VDD.n6459 GND 0.04999f
C15732 VDD.n6460 GND 0.68843f
C15733 VDD.n6461 GND 0.68843f
C15734 VDD.n6462 GND 0.04999f
C15735 VDD.n6463 GND 0.02746f
C15736 VDD.n6464 GND 0.02967f
C15737 VDD.n6465 GND 0.02746f
C15738 VDD.n6466 GND 0.04999f
C15739 VDD.n6467 GND 0.68843f
C15740 VDD.n6468 GND 0.02522f
C15741 VDD.n6469 GND 0.04999f
C15742 VDD.n6470 GND 0.68843f
C15743 VDD.n6471 GND 0.04999f
C15744 VDD.n6472 GND 0.05074f
C15745 VDD.n6473 GND 0.06295f
C15746 VDD.n6474 GND 0.0536f
C15747 VDD.n6475 GND 0.02522f
C15748 VDD.n6476 GND 0.04999f
C15749 VDD.n6477 GND 0.5126f
C15750 VDD.n6478 GND 0.02522f
C15751 VDD.n6479 GND 0.04999f
C15752 VDD.n6480 GND 0.5126f
C15753 VDD.n6481 GND 0.04999f
C15754 VDD.n6482 GND 0.05074f
C15755 VDD.n6483 GND 0.06295f
C15756 VDD.n6484 GND 0.0536f
C15757 VDD.n6485 GND 0.02522f
C15758 VDD.n6486 GND 0.04999f
C15759 VDD.n6487 GND 0.68843f
C15760 VDD.n6488 GND 0.02522f
C15761 VDD.n6489 GND 0.04999f
C15762 VDD.n6490 GND 0.68843f
C15763 VDD.n6491 GND 0.04999f
C15764 VDD.n6492 GND 0.05074f
C15765 VDD.n6493 GND 0.06295f
C15766 VDD.n6494 GND 0.0536f
C15767 VDD.n6495 GND 0.02522f
C15768 VDD.n6496 GND 0.04999f
C15769 VDD.n6497 GND 0.5126f
C15770 VDD.n6498 GND 0.02522f
C15771 VDD.n6499 GND 0.04999f
C15772 VDD.n6500 GND 0.5126f
C15773 VDD.n6501 GND 0.04999f
C15774 VDD.n6502 GND 0.05074f
C15775 VDD.n6503 GND 0.06295f
C15776 VDD.n6504 GND 0.0536f
C15777 VDD.n6505 GND 0.02522f
C15778 VDD.n6506 GND 0.04999f
C15779 VDD.n6507 GND 0.5126f
C15780 VDD.n6508 GND 0.5126f
C15781 VDD.n6509 GND 0.04999f
C15782 VDD.n6510 GND 0.04999f
C15783 VDD.n6511 GND 0.02522f
C15784 VDD.n6512 GND 0.02522f
C15785 VDD.n6513 GND 0.02967f
C15786 VDD.n6514 GND 0.05074f
C15787 VDD.t46 GND 0.63568f
C15788 VDD.n6515 GND 0.05074f
C15789 VDD.n6516 GND 0.06295f
C15790 VDD.n6517 GND 0.10164f
C15791 VDD.n6518 GND 0.0731f
C15792 VDD.n6519 GND 0.01798f
C15793 VDD.n6520 GND 0.09132f
C15794 VDD.n6521 GND 0.02746f
C15795 VDD.n6522 GND 0.04999f
C15796 VDD.n6523 GND 0.68843f
C15797 VDD.n6524 GND 0.02522f
C15798 VDD.n6525 GND 0.04999f
C15799 VDD.n6526 GND 0.68843f
C15800 VDD.n6527 GND 0.04999f
C15801 VDD.n6528 GND 0.05074f
C15802 VDD.n6529 GND 0.06295f
C15803 VDD.n6530 GND 0.0536f
C15804 VDD.n6531 GND 0.02522f
C15805 VDD.n6532 GND 0.04999f
C15806 VDD.n6533 GND 0.5126f
C15807 VDD.n6534 GND 0.02522f
C15808 VDD.n6535 GND 0.04999f
C15809 VDD.n6536 GND 0.5126f
C15810 VDD.n6537 GND 0.04999f
C15811 VDD.n6538 GND 0.05074f
C15812 VDD.n6539 GND 0.06295f
C15813 VDD.n6540 GND 0.0536f
C15814 VDD.n6541 GND 0.02522f
C15815 VDD.n6542 GND 0.04999f
C15816 VDD.n6543 GND 0.5126f
C15817 VDD.n6544 GND 0.02522f
C15818 VDD.n6545 GND 0.04999f
C15819 VDD.n6546 GND 0.5126f
C15820 VDD.n6547 GND 0.04999f
C15821 VDD.n6548 GND 0.05074f
C15822 VDD.n6549 GND 0.06295f
C15823 VDD.n6550 GND 0.0536f
C15824 VDD.n6551 GND 0.02522f
C15825 VDD.n6552 GND 0.04999f
C15826 VDD.n6553 GND 0.68843f
C15827 VDD.n6554 GND 0.02522f
C15828 VDD.n6555 GND 0.04999f
C15829 VDD.n6556 GND 0.68843f
C15830 VDD.n6557 GND 0.04999f
C15831 VDD.n6558 GND 0.05074f
C15832 VDD.n6559 GND 0.06295f
C15833 VDD.n6560 GND 0.0536f
C15834 VDD.n6561 GND 0.02522f
C15835 VDD.n6562 GND 0.04999f
C15836 VDD.n6563 GND 0.5126f
C15837 VDD.n6564 GND 0.02522f
C15838 VDD.n6565 GND 0.04999f
C15839 VDD.n6566 GND 0.5126f
C15840 VDD.n6567 GND 0.04999f
C15841 VDD.n6568 GND 0.05074f
C15842 VDD.n6569 GND 0.06295f
C15843 VDD.n6570 GND 0.0536f
C15844 VDD.n6571 GND 0.02522f
C15845 VDD.n6572 GND 0.04999f
C15846 VDD.n6573 GND 0.5126f
C15847 VDD.n6574 GND 0.02522f
C15848 VDD.n6575 GND 0.04999f
C15849 VDD.n6576 GND 0.5126f
C15850 VDD.n6577 GND 0.04999f
C15851 VDD.n6578 GND 0.05074f
C15852 VDD.n6579 GND 0.06295f
C15853 VDD.n6580 GND 0.0536f
C15854 VDD.n6581 GND 0.02522f
C15855 VDD.n6582 GND 0.04999f
C15856 VDD.n6583 GND 0.68843f
C15857 VDD.n6584 GND 0.68843f
C15858 VDD.n6585 GND 0.04999f
C15859 VDD.n6586 GND 0.02746f
C15860 VDD.n6587 GND 0.02967f
C15861 VDD.n6588 GND 0.02746f
C15862 VDD.n6589 GND 0.04999f
C15863 VDD.n6590 GND 0.68843f
C15864 VDD.n6591 GND 0.02522f
C15865 VDD.n6592 GND 0.04999f
C15866 VDD.n6593 GND 0.68843f
C15867 VDD.n6594 GND 0.04999f
C15868 VDD.n6595 GND 0.05074f
C15869 VDD.n6596 GND 0.06295f
C15870 VDD.n6597 GND 0.0536f
C15871 VDD.n6598 GND 0.02522f
C15872 VDD.n6599 GND 0.04999f
C15873 VDD.n6600 GND 0.5126f
C15874 VDD.n6601 GND 0.02522f
C15875 VDD.n6602 GND 0.04999f
C15876 VDD.n6603 GND 0.5126f
C15877 VDD.n6604 GND 0.04999f
C15878 VDD.n6605 GND 0.05074f
C15879 VDD.n6606 GND 0.06295f
C15880 VDD.n6607 GND 0.0536f
C15881 VDD.n6608 GND 0.02522f
C15882 VDD.n6609 GND 0.04999f
C15883 VDD.n6610 GND 0.68843f
C15884 VDD.n6611 GND 0.02522f
C15885 VDD.n6612 GND 0.04999f
C15886 VDD.n6613 GND 0.68843f
C15887 VDD.n6614 GND 0.04999f
C15888 VDD.n6615 GND 0.05074f
C15889 VDD.n6616 GND 0.06295f
C15890 VDD.n6617 GND 0.0536f
C15891 VDD.n6618 GND 0.02522f
C15892 VDD.n6619 GND 0.04999f
C15893 VDD.n6620 GND 0.5126f
C15894 VDD.n6621 GND 0.02522f
C15895 VDD.n6622 GND 0.04999f
C15896 VDD.n6623 GND 0.5126f
C15897 VDD.n6624 GND 0.04999f
C15898 VDD.n6625 GND 0.05074f
C15899 VDD.n6626 GND 0.06295f
C15900 VDD.n6627 GND 0.0536f
C15901 VDD.n6628 GND 0.02522f
C15902 VDD.n6629 GND 0.04999f
C15903 VDD.n6630 GND 0.5126f
C15904 VDD.n6631 GND 0.5126f
C15905 VDD.n6632 GND 0.04999f
C15906 VDD.n6633 GND 0.04999f
C15907 VDD.n6634 GND 0.02522f
C15908 VDD.n6635 GND 0.02522f
C15909 VDD.n6636 GND 0.02967f
C15910 VDD.n6637 GND 0.05074f
C15911 VDD.t312 GND 0.63568f
C15912 VDD.n6638 GND 0.05074f
C15913 VDD.n6639 GND 0.06295f
C15914 VDD.n6640 GND 0.10164f
C15915 VDD.n6641 GND 0.0731f
C15916 VDD.n6642 GND 0.01798f
C15917 VDD.n6643 GND 0.09132f
C15918 VDD.n6644 GND 0.02746f
C15919 VDD.n6645 GND 0.04999f
C15920 VDD.n6646 GND 0.68843f
C15921 VDD.n6647 GND 0.02522f
C15922 VDD.n6648 GND 0.04999f
C15923 VDD.n6649 GND 0.68843f
C15924 VDD.n6650 GND 0.04999f
C15925 VDD.n6651 GND 0.05074f
C15926 VDD.n6652 GND 0.06295f
C15927 VDD.n6653 GND 0.0536f
C15928 VDD.n6654 GND 0.02522f
C15929 VDD.n6655 GND 0.04999f
C15930 VDD.n6656 GND 0.5126f
C15931 VDD.n6657 GND 0.02522f
C15932 VDD.n6658 GND 0.04999f
C15933 VDD.n6659 GND 0.5126f
C15934 VDD.n6660 GND 0.04999f
C15935 VDD.n6661 GND 0.05074f
C15936 VDD.n6662 GND 0.06295f
C15937 VDD.n6663 GND 0.0536f
C15938 VDD.n6664 GND 0.02522f
C15939 VDD.n6665 GND 0.04999f
C15940 VDD.n6666 GND 0.5126f
C15941 VDD.n6667 GND 0.02522f
C15942 VDD.n6668 GND 0.04999f
C15943 VDD.n6669 GND 0.5126f
C15944 VDD.n6670 GND 0.04999f
C15945 VDD.n6671 GND 0.05074f
C15946 VDD.n6672 GND 0.06295f
C15947 VDD.n6673 GND 0.0536f
C15948 VDD.n6674 GND 0.02522f
C15949 VDD.n6675 GND 0.04999f
C15950 VDD.n6676 GND 0.68843f
C15951 VDD.n6677 GND 0.02522f
C15952 VDD.n6678 GND 0.04999f
C15953 VDD.n6679 GND 0.68843f
C15954 VDD.n6680 GND 0.04999f
C15955 VDD.n6681 GND 0.05074f
C15956 VDD.n6682 GND 0.06295f
C15957 VDD.n6683 GND 0.0536f
C15958 VDD.n6684 GND 0.02522f
C15959 VDD.n6685 GND 0.04999f
C15960 VDD.n6686 GND 0.5126f
C15961 VDD.n6687 GND 0.02522f
C15962 VDD.n6688 GND 0.04999f
C15963 VDD.n6689 GND 0.5126f
C15964 VDD.n6690 GND 0.04999f
C15965 VDD.n6691 GND 0.05074f
C15966 VDD.n6692 GND 0.06295f
C15967 VDD.n6693 GND 0.0536f
C15968 VDD.n6694 GND 0.02522f
C15969 VDD.n6695 GND 0.04999f
C15970 VDD.n6696 GND 0.5126f
C15971 VDD.n6697 GND 0.02522f
C15972 VDD.n6698 GND 0.04999f
C15973 VDD.n6699 GND 0.5126f
C15974 VDD.n6700 GND 0.04999f
C15975 VDD.n6701 GND 0.05074f
C15976 VDD.n6702 GND 0.06295f
C15977 VDD.n6703 GND 0.0536f
C15978 VDD.n6704 GND 0.02522f
C15979 VDD.n6705 GND 0.04999f
C15980 VDD.n6706 GND 0.68843f
C15981 VDD.n6707 GND 0.68843f
C15982 VDD.n6708 GND 0.04999f
C15983 VDD.n6709 GND 0.02746f
C15984 VDD.n6710 GND 0.02967f
C15985 VDD.n6711 GND 0.02746f
C15986 VDD.n6712 GND 0.04999f
C15987 VDD.n6713 GND 0.68843f
C15988 VDD.n6714 GND 0.02522f
C15989 VDD.n6715 GND 0.04999f
C15990 VDD.n6716 GND 0.68843f
C15991 VDD.n6717 GND 0.04999f
C15992 VDD.n6718 GND 0.05074f
C15993 VDD.n6719 GND 0.06295f
C15994 VDD.n6720 GND 0.0536f
C15995 VDD.n6721 GND 0.02522f
C15996 VDD.n6722 GND 0.04999f
C15997 VDD.n6723 GND 0.5126f
C15998 VDD.n6724 GND 0.02522f
C15999 VDD.n6725 GND 0.04999f
C16000 VDD.n6726 GND 0.5126f
C16001 VDD.n6727 GND 0.04999f
C16002 VDD.n6728 GND 0.05074f
C16003 VDD.n6729 GND 0.06295f
C16004 VDD.n6730 GND 0.0536f
C16005 VDD.n6731 GND 0.02522f
C16006 VDD.n6732 GND 0.04999f
C16007 VDD.n6733 GND 0.68843f
C16008 VDD.n6734 GND 0.02522f
C16009 VDD.n6735 GND 0.04999f
C16010 VDD.n6736 GND 0.68843f
C16011 VDD.n6737 GND 0.04999f
C16012 VDD.n6738 GND 0.05074f
C16013 VDD.n6739 GND 0.06295f
C16014 VDD.n6740 GND 0.0536f
C16015 VDD.n6741 GND 0.02522f
C16016 VDD.n6742 GND 0.04999f
C16017 VDD.n6743 GND 0.5126f
C16018 VDD.n6744 GND 0.02522f
C16019 VDD.n6745 GND 0.04999f
C16020 VDD.n6746 GND 0.5126f
C16021 VDD.n6747 GND 0.04999f
C16022 VDD.n6748 GND 0.05074f
C16023 VDD.n6749 GND 0.06295f
C16024 VDD.n6750 GND 0.0536f
C16025 VDD.n6751 GND 0.02522f
C16026 VDD.n6752 GND 0.04999f
C16027 VDD.n6753 GND 0.5126f
C16028 VDD.n6754 GND 0.5126f
C16029 VDD.n6755 GND 0.04999f
C16030 VDD.n6756 GND 0.04999f
C16031 VDD.n6757 GND 0.02522f
C16032 VDD.n6758 GND 0.02522f
C16033 VDD.n6759 GND 0.02967f
C16034 VDD.n6760 GND 0.05074f
C16035 VDD.t305 GND 0.63568f
C16036 VDD.n6761 GND 0.05074f
C16037 VDD.n6762 GND 0.06295f
C16038 VDD.n6763 GND 0.10164f
C16039 VDD.n6764 GND 0.0731f
C16040 VDD.n6765 GND 0.01798f
C16041 VDD.n6766 GND 0.09132f
C16042 VDD.n6767 GND 0.02746f
C16043 VDD.n6768 GND 0.04999f
C16044 VDD.n6769 GND 0.68843f
C16045 VDD.n6770 GND 0.02522f
C16046 VDD.n6771 GND 0.04999f
C16047 VDD.n6772 GND 0.68843f
C16048 VDD.n6773 GND 0.04999f
C16049 VDD.n6774 GND 0.05074f
C16050 VDD.n6775 GND 0.06295f
C16051 VDD.n6776 GND 0.0536f
C16052 VDD.n6777 GND 0.02522f
C16053 VDD.n6778 GND 0.04999f
C16054 VDD.n6779 GND 0.5126f
C16055 VDD.n6780 GND 0.02522f
C16056 VDD.n6781 GND 0.04999f
C16057 VDD.n6782 GND 0.5126f
C16058 VDD.n6783 GND 0.04999f
C16059 VDD.n6784 GND 0.05074f
C16060 VDD.n6785 GND 0.06295f
C16061 VDD.n6786 GND 0.0536f
C16062 VDD.n6787 GND 0.02522f
C16063 VDD.n6788 GND 0.04999f
C16064 VDD.n6789 GND 0.5126f
C16065 VDD.n6790 GND 0.02522f
C16066 VDD.n6791 GND 0.04999f
C16067 VDD.n6792 GND 0.5126f
C16068 VDD.n6793 GND 0.04999f
C16069 VDD.n6794 GND 0.05074f
C16070 VDD.n6795 GND 0.06295f
C16071 VDD.n6796 GND 0.0536f
C16072 VDD.n6797 GND 0.02522f
C16073 VDD.n6798 GND 0.04999f
C16074 VDD.n6799 GND 0.68843f
C16075 VDD.n6800 GND 0.02522f
C16076 VDD.n6801 GND 0.04999f
C16077 VDD.n6802 GND 0.68843f
C16078 VDD.n6803 GND 0.04999f
C16079 VDD.n6804 GND 0.05074f
C16080 VDD.n6805 GND 0.06295f
C16081 VDD.n6806 GND 0.0536f
C16082 VDD.n6807 GND 0.02522f
C16083 VDD.n6808 GND 0.04999f
C16084 VDD.n6809 GND 0.5126f
C16085 VDD.n6810 GND 0.02522f
C16086 VDD.n6811 GND 0.04999f
C16087 VDD.n6812 GND 0.5126f
C16088 VDD.n6813 GND 0.04999f
C16089 VDD.n6814 GND 0.05074f
C16090 VDD.n6815 GND 0.06295f
C16091 VDD.n6816 GND 0.0536f
C16092 VDD.n6817 GND 0.02522f
C16093 VDD.n6818 GND 0.04999f
C16094 VDD.n6819 GND 0.5126f
C16095 VDD.n6820 GND 0.02522f
C16096 VDD.n6821 GND 0.04999f
C16097 VDD.n6822 GND 0.5126f
C16098 VDD.n6823 GND 0.04999f
C16099 VDD.n6824 GND 0.05074f
C16100 VDD.n6825 GND 0.06295f
C16101 VDD.n6826 GND 0.0536f
C16102 VDD.n6827 GND 0.02522f
C16103 VDD.n6828 GND 0.04999f
C16104 VDD.n6829 GND 0.68843f
C16105 VDD.n6830 GND 0.68843f
C16106 VDD.n6831 GND 0.04999f
C16107 VDD.n6832 GND 0.02746f
C16108 VDD.n6833 GND 0.02967f
C16109 VDD.n6834 GND 0.02746f
C16110 VDD.n6835 GND 0.04999f
C16111 VDD.n6836 GND 0.68843f
C16112 VDD.n6837 GND 0.02522f
C16113 VDD.n6838 GND 0.04999f
C16114 VDD.n6839 GND 0.68843f
C16115 VDD.n6840 GND 0.04999f
C16116 VDD.n6841 GND 0.05074f
C16117 VDD.n6842 GND 0.06295f
C16118 VDD.n6843 GND 0.0536f
C16119 VDD.n6844 GND 0.02522f
C16120 VDD.n6845 GND 0.04999f
C16121 VDD.n6846 GND 0.5126f
C16122 VDD.n6847 GND 0.02522f
C16123 VDD.n6848 GND 0.04999f
C16124 VDD.n6849 GND 0.5126f
C16125 VDD.n6850 GND 0.04999f
C16126 VDD.n6851 GND 0.05074f
C16127 VDD.n6852 GND 0.06295f
C16128 VDD.n6853 GND 0.0536f
C16129 VDD.n6854 GND 0.02522f
C16130 VDD.n6855 GND 0.04999f
C16131 VDD.n6856 GND 0.68843f
C16132 VDD.n6857 GND 0.02522f
C16133 VDD.n6858 GND 0.04999f
C16134 VDD.n6859 GND 0.68843f
C16135 VDD.n6860 GND 0.04999f
C16136 VDD.n6861 GND 0.05074f
C16137 VDD.n6862 GND 0.06295f
C16138 VDD.n6863 GND 0.0536f
C16139 VDD.n6864 GND 0.02522f
C16140 VDD.n6865 GND 0.04999f
C16141 VDD.n6866 GND 0.5126f
C16142 VDD.n6867 GND 0.02522f
C16143 VDD.n6868 GND 0.04999f
C16144 VDD.n6869 GND 0.5126f
C16145 VDD.n6870 GND 0.04999f
C16146 VDD.n6871 GND 0.05074f
C16147 VDD.n6872 GND 0.06295f
C16148 VDD.n6873 GND 0.0536f
C16149 VDD.n6874 GND 0.02522f
C16150 VDD.n6875 GND 0.04999f
C16151 VDD.n6876 GND 0.5126f
C16152 VDD.n6877 GND 0.5126f
C16153 VDD.n6878 GND 0.04999f
C16154 VDD.n6879 GND 0.04999f
C16155 VDD.n6880 GND 0.02522f
C16156 VDD.n6881 GND 0.02522f
C16157 VDD.n6882 GND 0.02967f
C16158 VDD.n6883 GND 0.05074f
C16159 VDD.t349 GND 0.63568f
C16160 VDD.n6884 GND 0.05074f
C16161 VDD.n6885 GND 0.06295f
C16162 VDD.n6886 GND 0.07292f
C16163 VDD.n6887 GND 1.23109f
C16164 VDD.t951 GND 0.02321f
C16165 VDD.t1009 GND 0.02321f
C16166 VDD.n6889 GND 0.10855f
C16167 VDD.n6890 GND 0.03131f
C16168 VDD.n6891 GND 0.02746f
C16169 VDD.n6892 GND 0.02746f
C16170 VDD.n6893 GND 0.04999f
C16171 VDD.n6894 GND 0.04999f
C16172 VDD.t301 GND 0.33785f
C16173 VDD.n6895 GND 0.05074f
C16174 VDD.n6896 GND 0.05074f
C16175 VDD.t302 GND 0.02334f
C16176 VDD.n6897 GND 0.09798f
C16177 VDD.n6898 GND 0.09593f
C16178 VDD.n6900 GND 0.35737f
C16179 VDD.n6901 GND 0.02746f
C16180 VDD.n6902 GND 0.02967f
C16181 VDD.n6903 GND 0.02746f
C16182 VDD.n6904 GND 0.04999f
C16183 VDD.n6905 GND 0.33547f
C16184 VDD.n6906 GND 0.33547f
C16185 VDD.t1008 GND 0.33785f
C16186 VDD.n6907 GND 0.05074f
C16187 VDD.n6908 GND 0.05074f
C16188 VDD.t277 GND 0.02321f
C16189 VDD.t774 GND 0.02321f
C16190 VDD.n6909 GND 0.10855f
C16191 VDD.n6910 GND 0.03131f
C16192 VDD.n6911 GND 0.02746f
C16193 VDD.n6912 GND 0.05074f
C16194 VDD.n6913 GND 0.02967f
C16195 VDD.n6914 GND 0.05074f
C16196 VDD.n6915 GND 0.35737f
C16197 VDD.t276 GND 0.33785f
C16198 VDD.t773 GND 0.33785f
C16199 VDD.n6917 GND 0.05074f
C16200 VDD.n6918 GND 0.05074f
C16201 VDD.t584 GND 0.02334f
C16202 VDD.n6919 GND 0.0731f
C16203 VDD.n6920 GND 0.02746f
C16204 VDD.n6921 GND 0.05074f
C16205 VDD.n6922 GND 0.02967f
C16206 VDD.n6923 GND 0.05074f
C16207 VDD.n6924 GND 0.35737f
C16208 VDD.t583 GND 0.33785f
C16209 VDD.t399 GND 0.30977f
C16210 VDD.n6926 GND 0.05074f
C16211 VDD.n6927 GND 0.05074f
C16212 VDD.n6928 GND 0.09132f
C16213 VDD.t1040 GND 0.33785f
C16214 VDD.n6929 GND 0.05074f
C16215 VDD.n6930 GND 0.05074f
C16216 VDD.t400 GND 0.02321f
C16217 VDD.t1041 GND 0.02321f
C16218 VDD.n6931 GND 0.10855f
C16219 VDD.n6932 GND 0.02334f
C16220 VDD.n6933 GND 0.03131f
C16221 VDD.t792 GND 0.02321f
C16222 VDD.t799 GND 0.02321f
C16223 VDD.n6934 GND 0.10855f
C16224 VDD.n6935 GND 0.03131f
C16225 VDD.n6936 GND 0.02746f
C16226 VDD.n6937 GND 0.05074f
C16227 VDD.n6938 GND 0.02967f
C16228 VDD.n6939 GND 0.05074f
C16229 VDD.n6940 GND 0.35737f
C16230 VDD.t791 GND 0.33785f
C16231 VDD.t798 GND 0.33785f
C16232 VDD.n6942 GND 0.05074f
C16233 VDD.n6943 GND 0.05074f
C16234 VDD.t190 GND 0.02334f
C16235 VDD.n6944 GND 0.0731f
C16236 VDD.n6945 GND 0.02746f
C16237 VDD.n6946 GND 0.05074f
C16238 VDD.n6947 GND 0.02967f
C16239 VDD.n6948 GND 0.05074f
C16240 VDD.n6949 GND 0.35737f
C16241 VDD.t189 GND 0.33785f
C16242 VDD.t420 GND 0.30977f
C16243 VDD.n6951 GND 0.05074f
C16244 VDD.n6952 GND 0.05074f
C16245 VDD.n6953 GND 0.09132f
C16246 VDD.t1012 GND 0.33785f
C16247 VDD.n6954 GND 0.05074f
C16248 VDD.n6955 GND 0.05074f
C16249 VDD.t421 GND 0.02321f
C16250 VDD.t1013 GND 0.02321f
C16251 VDD.n6956 GND 0.10855f
C16252 VDD.n6957 GND 0.02334f
C16253 VDD.n6958 GND 0.03131f
C16254 VDD.t72 GND 0.02321f
C16255 VDD.t127 GND 0.02321f
C16256 VDD.n6959 GND 0.10855f
C16257 VDD.n6960 GND 0.03131f
C16258 VDD.n6961 GND 0.02746f
C16259 VDD.n6962 GND 0.05074f
C16260 VDD.n6963 GND 0.02967f
C16261 VDD.n6964 GND 0.05074f
C16262 VDD.n6965 GND 0.35737f
C16263 VDD.t71 GND 0.33785f
C16264 VDD.t126 GND 0.33785f
C16265 VDD.n6967 GND 0.05074f
C16266 VDD.n6968 GND 0.05074f
C16267 VDD.t932 GND 0.02334f
C16268 VDD.n6969 GND 0.0731f
C16269 VDD.n6970 GND 0.02746f
C16270 VDD.n6971 GND 0.05074f
C16271 VDD.n6972 GND 0.02967f
C16272 VDD.n6973 GND 0.05074f
C16273 VDD.n6974 GND 0.35737f
C16274 VDD.t931 GND 0.33785f
C16275 VDD.t954 GND 0.30977f
C16276 VDD.n6976 GND 0.05074f
C16277 VDD.n6977 GND 0.05074f
C16278 VDD.n6978 GND 0.09132f
C16279 VDD.t1036 GND 0.33785f
C16280 VDD.n6979 GND 0.05074f
C16281 VDD.n6980 GND 0.05074f
C16282 VDD.t955 GND 0.02321f
C16283 VDD.t1037 GND 0.02321f
C16284 VDD.n6981 GND 0.10855f
C16285 VDD.n6982 GND 0.02334f
C16286 VDD.n6983 GND 0.03131f
C16287 VDD.t969 GND 0.02321f
C16288 VDD.t940 GND 0.02321f
C16289 VDD.n6984 GND 0.10855f
C16290 VDD.n6985 GND 0.03131f
C16291 VDD.n6986 GND 0.02746f
C16292 VDD.n6987 GND 0.05074f
C16293 VDD.n6988 GND 0.02967f
C16294 VDD.n6989 GND 0.05074f
C16295 VDD.n6990 GND 0.35737f
C16296 VDD.t968 GND 0.33785f
C16297 VDD.t939 GND 0.33785f
C16298 VDD.n6992 GND 0.05074f
C16299 VDD.n6993 GND 0.05074f
C16300 VDD.n6994 GND 0.02334f
C16301 VDD.n6995 GND 0.09132f
C16302 VDD.n6997 GND 0.35737f
C16303 VDD.n6998 GND 0.02746f
C16304 VDD.n6999 GND 0.02967f
C16305 VDD.n7000 GND 0.02746f
C16306 VDD.n7001 GND 0.04999f
C16307 VDD.n7002 GND 0.24979f
C16308 VDD.n7003 GND 0.24979f
C16309 VDD.n7004 GND 0.04999f
C16310 VDD.n7005 GND 0.02746f
C16311 VDD.n7006 GND 0.09132f
C16312 VDD.n7007 GND 0.34336f
C16313 VDD.n7008 GND 0.02334f
C16314 VDD.n7009 GND 0.09132f
C16315 VDD.n7011 GND 0.35737f
C16316 VDD.n7012 GND 0.02746f
C16317 VDD.n7013 GND 0.02967f
C16318 VDD.n7014 GND 0.02746f
C16319 VDD.n7015 GND 0.04999f
C16320 VDD.n7016 GND 0.24979f
C16321 VDD.n7017 GND 0.24979f
C16322 VDD.n7018 GND 0.04999f
C16323 VDD.n7019 GND 0.02746f
C16324 VDD.n7020 GND 0.02967f
C16325 VDD.n7021 GND 0.02746f
C16326 VDD.n7022 GND 0.04999f
C16327 VDD.n7023 GND 0.33547f
C16328 VDD.n7024 GND 0.33547f
C16329 VDD.n7025 GND 0.04999f
C16330 VDD.n7026 GND 0.02746f
C16331 VDD.n7027 GND 0.09132f
C16332 VDD.n7028 GND 0.33799f
C16333 VDD.n7029 GND 0.02334f
C16334 VDD.n7030 GND 0.09132f
C16335 VDD.n7032 GND 0.35737f
C16336 VDD.n7033 GND 0.02746f
C16337 VDD.n7034 GND 0.02967f
C16338 VDD.n7035 GND 0.02746f
C16339 VDD.n7036 GND 0.04999f
C16340 VDD.n7037 GND 0.24979f
C16341 VDD.n7038 GND 0.24979f
C16342 VDD.n7039 GND 0.04999f
C16343 VDD.n7040 GND 0.02746f
C16344 VDD.n7041 GND 0.09132f
C16345 VDD.n7042 GND 0.34336f
C16346 VDD.n7043 GND 0.02334f
C16347 VDD.n7044 GND 0.09132f
C16348 VDD.n7046 GND 0.35737f
C16349 VDD.n7047 GND 0.02746f
C16350 VDD.n7048 GND 0.02967f
C16351 VDD.n7049 GND 0.02746f
C16352 VDD.n7050 GND 0.04999f
C16353 VDD.n7051 GND 0.24979f
C16354 VDD.n7052 GND 0.24979f
C16355 VDD.n7053 GND 0.04999f
C16356 VDD.n7054 GND 0.02746f
C16357 VDD.n7055 GND 0.02967f
C16358 VDD.n7056 GND 0.02746f
C16359 VDD.n7057 GND 0.04999f
C16360 VDD.n7058 GND 0.33547f
C16361 VDD.n7059 GND 0.33547f
C16362 VDD.n7060 GND 0.04999f
C16363 VDD.n7061 GND 0.02746f
C16364 VDD.n7062 GND 0.09132f
C16365 VDD.n7063 GND 0.33799f
C16366 VDD.n7064 GND 0.02334f
C16367 VDD.n7065 GND 0.09132f
C16368 VDD.n7067 GND 0.35737f
C16369 VDD.n7068 GND 0.02746f
C16370 VDD.n7069 GND 0.02967f
C16371 VDD.n7070 GND 0.02746f
C16372 VDD.n7071 GND 0.04999f
C16373 VDD.n7072 GND 0.24979f
C16374 VDD.n7073 GND 0.24979f
C16375 VDD.n7074 GND 0.04999f
C16376 VDD.n7075 GND 0.02746f
C16377 VDD.n7076 GND 0.09132f
C16378 VDD.n7077 GND 0.34336f
C16379 VDD.n7078 GND 0.02334f
C16380 VDD.n7079 GND 0.09132f
C16381 VDD.n7081 GND 0.35737f
C16382 VDD.n7082 GND 0.02746f
C16383 VDD.n7083 GND 0.02967f
C16384 VDD.n7084 GND 0.02746f
C16385 VDD.n7085 GND 0.04999f
C16386 VDD.n7086 GND 0.24979f
C16387 VDD.n7087 GND 0.24979f
C16388 VDD.n7088 GND 0.04999f
C16389 VDD.n7089 GND 0.02746f
C16390 VDD.n7090 GND 0.02967f
C16391 VDD.n7091 GND 0.02746f
C16392 VDD.n7092 GND 0.04999f
C16393 VDD.n7093 GND 0.33547f
C16394 VDD.n7094 GND 0.33547f
C16395 VDD.n7095 GND 0.04999f
C16396 VDD.n7096 GND 0.02746f
C16397 VDD.n7097 GND 0.09132f
C16398 VDD.n7098 GND 0.33799f
C16399 VDD.n7099 GND 0.02334f
C16400 VDD.n7100 GND 0.09132f
C16401 VDD.n7102 GND 0.35737f
C16402 VDD.n7103 GND 0.02746f
C16403 VDD.n7104 GND 0.02967f
C16404 VDD.n7105 GND 0.02746f
C16405 VDD.n7106 GND 0.04999f
C16406 VDD.n7107 GND 0.24979f
C16407 VDD.n7108 GND 0.24979f
C16408 VDD.n7109 GND 0.04999f
C16409 VDD.n7110 GND 0.02746f
C16410 VDD.n7111 GND 0.09132f
C16411 VDD.n7112 GND 0.34336f
C16412 VDD.n7113 GND 0.02334f
C16413 VDD.n7114 GND 0.09132f
C16414 VDD.n7116 GND 0.35737f
C16415 VDD.n7117 GND 0.02746f
C16416 VDD.n7118 GND 0.02967f
C16417 VDD.n7119 GND 0.02746f
C16418 VDD.n7120 GND 0.04999f
C16419 VDD.n7121 GND 0.24979f
C16420 VDD.n7122 GND 0.24979f
C16421 VDD.n7123 GND 0.02967f
C16422 VDD.n7124 GND 0.05074f
C16423 VDD.t950 GND 0.30977f
C16424 VDD.n7125 GND 0.05074f
C16425 VDD.n7126 GND 0.09132f
C16426 VDD.n7127 GND 0.02241f
C16427 VDD.n7128 GND 0.0768f
C16428 VDD.n7130 GND 2.13433f
C16429 VDD.n7131 GND 0.14251f
C16430 VDD.n7132 GND 0.02334f
C16431 VDD.n7133 GND 0.0536f
C16432 VDD.n7134 GND 0.05074f
C16433 VDD.n7135 GND 0.02967f
C16434 VDD.n7136 GND 0.02522f
C16435 VDD.n7137 GND 0.02522f
C16436 VDD.n7138 GND 0.04999f
C16437 VDD.n7139 GND 0.68843f
C16438 VDD.n7140 GND 0.04999f
C16439 VDD.n7141 GND 0.05074f
C16440 VDD.n7142 GND 0.06295f
C16441 VDD.n7143 GND 0.0536f
C16442 VDD.n7144 GND 0.02522f
C16443 VDD.n7145 GND 0.04999f
C16444 VDD.n7146 GND 0.5126f
C16445 VDD.n7147 GND 0.02522f
C16446 VDD.n7148 GND 0.04999f
C16447 VDD.n7149 GND 0.5126f
C16448 VDD.n7150 GND 0.04999f
C16449 VDD.n7151 GND 0.05074f
C16450 VDD.n7152 GND 0.06295f
C16451 VDD.n7153 GND 0.0536f
C16452 VDD.n7154 GND 0.02522f
C16453 VDD.n7155 GND 0.04999f
C16454 VDD.n7156 GND 0.5126f
C16455 VDD.n7157 GND 0.02522f
C16456 VDD.n7158 GND 0.04999f
C16457 VDD.n7159 GND 0.5126f
C16458 VDD.n7160 GND 0.04999f
C16459 VDD.n7161 GND 0.05074f
C16460 VDD.n7162 GND 0.06295f
C16461 VDD.n7163 GND 0.0536f
C16462 VDD.n7164 GND 0.02522f
C16463 VDD.n7165 GND 0.04999f
C16464 VDD.n7166 GND 0.68843f
C16465 VDD.n7167 GND 0.02522f
C16466 VDD.n7168 GND 0.04999f
C16467 VDD.n7169 GND 0.68843f
C16468 VDD.n7170 GND 0.04999f
C16469 VDD.n7171 GND 0.05074f
C16470 VDD.n7172 GND 0.06295f
C16471 VDD.n7173 GND 0.0536f
C16472 VDD.n7174 GND 0.02522f
C16473 VDD.n7175 GND 0.04999f
C16474 VDD.n7176 GND 0.5126f
C16475 VDD.n7177 GND 0.02522f
C16476 VDD.n7178 GND 0.04999f
C16477 VDD.n7179 GND 0.5126f
C16478 VDD.n7180 GND 0.04999f
C16479 VDD.n7181 GND 0.05074f
C16480 VDD.n7182 GND 0.06295f
C16481 VDD.n7183 GND 0.0536f
C16482 VDD.n7184 GND 0.02522f
C16483 VDD.n7185 GND 0.04999f
C16484 VDD.n7186 GND 0.68843f
C16485 VDD.n7187 GND 0.68843f
C16486 VDD.n7188 GND 0.04999f
C16487 VDD.n7189 GND 0.02746f
C16488 VDD.n7190 GND 0.02967f
C16489 VDD.n7191 GND 0.02746f
C16490 VDD.n7192 GND 0.04999f
C16491 VDD.n7193 GND 0.68843f
C16492 VDD.n7194 GND 0.68843f
C16493 VDD.n7195 GND 0.04999f
C16494 VDD.n7196 GND 0.04999f
C16495 VDD.n7197 GND 0.02522f
C16496 VDD.n7198 GND 0.02522f
C16497 VDD.n7199 GND 0.02967f
C16498 VDD.n7200 GND 0.05074f
C16499 VDD.t35 GND 0.63568f
C16500 VDD.n7201 GND 0.05074f
C16501 VDD.n7202 GND 0.06295f
C16502 VDD.n7203 GND 0.02334f
C16503 VDD.n7204 GND 0.04152f
C16504 VDD.n7205 GND 0.03056f
C16505 VDD.n7206 GND 0.06295f
C16506 VDD.n7207 GND 0.0536f
C16507 VDD.n7208 GND 0.02522f
C16508 VDD.n7209 GND 0.04999f
C16509 VDD.n7210 GND 0.5126f
C16510 VDD.n7211 GND 0.02522f
C16511 VDD.n7212 GND 0.04999f
C16512 VDD.n7213 GND 0.5126f
C16513 VDD.n7214 GND 0.04999f
C16514 VDD.n7215 GND 0.05074f
C16515 VDD.n7216 GND 0.06295f
C16516 VDD.n7217 GND 0.0536f
C16517 VDD.n7218 GND 0.02522f
C16518 VDD.n7219 GND 0.04999f
C16519 VDD.n7220 GND 0.68843f
C16520 VDD.n7221 GND 0.02522f
C16521 VDD.n7222 GND 0.04999f
C16522 VDD.n7223 GND 0.68843f
C16523 VDD.n7224 GND 0.04999f
C16524 VDD.n7225 GND 0.05074f
C16525 VDD.n7226 GND 0.06295f
C16526 VDD.n7227 GND 0.0536f
C16527 VDD.n7228 GND 0.02522f
C16528 VDD.n7229 GND 0.04999f
C16529 VDD.n7230 GND 0.5126f
C16530 VDD.n7231 GND 0.02522f
C16531 VDD.n7232 GND 0.04999f
C16532 VDD.n7233 GND 0.5126f
C16533 VDD.n7234 GND 0.04999f
C16534 VDD.n7235 GND 0.05074f
C16535 VDD.n7236 GND 0.06295f
C16536 VDD.n7237 GND 0.0536f
C16537 VDD.n7238 GND 0.02522f
C16538 VDD.n7239 GND 0.04999f
C16539 VDD.n7240 GND 0.5126f
C16540 VDD.n7241 GND 0.02522f
C16541 VDD.n7242 GND 0.04999f
C16542 VDD.n7243 GND 0.5126f
C16543 VDD.n7244 GND 0.04999f
C16544 VDD.n7245 GND 0.05074f
C16545 VDD.n7246 GND 0.06295f
C16546 VDD.n7247 GND 0.0536f
C16547 VDD.n7248 GND 0.02522f
C16548 VDD.n7249 GND 0.04999f
C16549 VDD.n7250 GND 0.68843f
C16550 VDD.n7251 GND 0.68843f
C16551 VDD.n7252 GND 0.04999f
C16552 VDD.n7253 GND 0.02746f
C16553 VDD.n7254 GND 0.09132f
C16554 VDD.n7255 GND 0.01798f
C16555 VDD.n7256 GND 0.071f
C16556 VDD.n7257 GND 0.47442f
C16557 VDD.t608 GND 0.02334f
C16558 VDD.n7258 GND 0.02746f
C16559 VDD.n7259 GND 0.05074f
C16560 VDD.n7260 GND 0.02967f
C16561 VDD.n7261 GND 0.05074f
C16562 VDD.n7262 GND 0.62973f
C16563 VDD.t607 GND 0.74438f
C16564 VDD.n7264 GND 0.04999f
C16565 VDD.t155 GND 0.63568f
C16566 VDD.n7265 GND 0.05074f
C16567 VDD.n7266 GND 0.05074f
C16568 VDD.n7267 GND 0.02967f
C16569 VDD.n7268 GND 0.02522f
C16570 VDD.t355 GND 0.02334f
C16571 VDD.t156 GND 0.02334f
C16572 VDD.n7269 GND 0.13341f
C16573 VDD.n7270 GND 0.0263f
C16574 VDD.n7271 GND 0.0536f
C16575 VDD.n7272 GND 0.05074f
C16576 VDD.n7273 GND 0.02967f
C16577 VDD.n7274 GND 0.02522f
C16578 VDD.n7275 GND 0.04999f
C16579 VDD.t337 GND 0.63568f
C16580 VDD.n7276 GND 0.05074f
C16581 VDD.n7277 GND 0.05074f
C16582 VDD.n7278 GND 0.02967f
C16583 VDD.n7279 GND 0.02522f
C16584 VDD.n7280 GND 0.03166f
C16585 VDD.n7281 GND 0.0536f
C16586 VDD.n7282 GND 0.05074f
C16587 VDD.n7283 GND 0.02967f
C16588 VDD.n7284 GND 0.02522f
C16589 VDD.n7285 GND 0.04999f
C16590 VDD.t911 GND 0.63568f
C16591 VDD.n7286 GND 0.05074f
C16592 VDD.n7287 GND 0.05074f
C16593 VDD.n7288 GND 0.02967f
C16594 VDD.n7289 GND 0.02522f
C16595 VDD.t338 GND 0.02321f
C16596 VDD.t912 GND 0.02321f
C16597 VDD.n7290 GND 0.10855f
C16598 VDD.t981 GND 0.02321f
C16599 VDD.t915 GND 0.02321f
C16600 VDD.n7291 GND 0.10855f
C16601 VDD.n7292 GND 0.04152f
C16602 VDD.n7293 GND 0.02334f
C16603 VDD.n7294 GND 0.0536f
C16604 VDD.n7295 GND 0.05074f
C16605 VDD.n7296 GND 0.02967f
C16606 VDD.n7297 GND 0.02522f
C16607 VDD.n7298 GND 0.04999f
C16608 VDD.t13 GND 0.63568f
C16609 VDD.n7299 GND 0.05074f
C16610 VDD.n7300 GND 0.05074f
C16611 VDD.n7301 GND 0.02967f
C16612 VDD.n7302 GND 0.02522f
C16613 VDD.t561 GND 0.02334f
C16614 VDD.t14 GND 0.02334f
C16615 VDD.n7303 GND 0.13341f
C16616 VDD.n7304 GND 0.0263f
C16617 VDD.n7305 GND 0.0536f
C16618 VDD.n7306 GND 0.05074f
C16619 VDD.n7307 GND 0.02967f
C16620 VDD.n7308 GND 0.02522f
C16621 VDD.n7309 GND 0.04999f
C16622 VDD.t112 GND 0.63568f
C16623 VDD.n7310 GND 0.05074f
C16624 VDD.n7311 GND 0.05074f
C16625 VDD.n7312 GND 0.02967f
C16626 VDD.n7313 GND 0.02522f
C16627 VDD.n7314 GND 0.03166f
C16628 VDD.n7315 GND 0.0536f
C16629 VDD.n7316 GND 0.05074f
C16630 VDD.n7317 GND 0.02967f
C16631 VDD.n7318 GND 0.02522f
C16632 VDD.n7319 GND 0.04999f
C16633 VDD.t948 GND 0.63568f
C16634 VDD.n7320 GND 0.05074f
C16635 VDD.n7321 GND 0.05074f
C16636 VDD.n7322 GND 0.02967f
C16637 VDD.n7323 GND 0.02522f
C16638 VDD.t288 GND 0.02321f
C16639 VDD.t949 GND 0.02321f
C16640 VDD.n7324 GND 0.10855f
C16641 VDD.t113 GND 0.02321f
C16642 VDD.t972 GND 0.02321f
C16643 VDD.n7325 GND 0.10855f
C16644 VDD.n7326 GND 0.04152f
C16645 VDD.n7327 GND 0.02334f
C16646 VDD.n7328 GND 0.0536f
C16647 VDD.n7329 GND 0.05074f
C16648 VDD.n7330 GND 0.02967f
C16649 VDD.n7331 GND 0.02522f
C16650 VDD.t913 GND 0.63568f
C16651 VDD.n7332 GND 0.05074f
C16652 VDD.n7333 GND 0.05074f
C16653 VDD.n7334 GND 0.09132f
C16654 VDD.n7335 GND 0.04999f
C16655 VDD.t222 GND 0.63568f
C16656 VDD.n7336 GND 0.05074f
C16657 VDD.n7337 GND 0.05074f
C16658 VDD.n7338 GND 0.02967f
C16659 VDD.n7339 GND 0.02522f
C16660 VDD.t914 GND 0.02334f
C16661 VDD.n7340 GND 0.0731f
C16662 VDD.n7341 GND 0.01798f
C16663 VDD.n7342 GND 0.02334f
C16664 VDD.n7343 GND 0.0536f
C16665 VDD.n7344 GND 0.05074f
C16666 VDD.n7345 GND 0.02967f
C16667 VDD.n7346 GND 0.02522f
C16668 VDD.n7347 GND 0.04999f
C16669 VDD.t48 GND 0.63568f
C16670 VDD.n7348 GND 0.05074f
C16671 VDD.n7349 GND 0.05074f
C16672 VDD.n7350 GND 0.02967f
C16673 VDD.n7351 GND 0.02522f
C16674 VDD.t971 GND 0.02321f
C16675 VDD.t50 GND 0.02321f
C16676 VDD.n7352 GND 0.10855f
C16677 VDD.t223 GND 0.02321f
C16678 VDD.t49 GND 0.02321f
C16679 VDD.n7353 GND 0.10855f
C16680 VDD.n7354 GND 0.04152f
C16681 VDD.n7355 GND 0.02334f
C16682 VDD.n7356 GND 0.0536f
C16683 VDD.n7357 GND 0.05074f
C16684 VDD.n7358 GND 0.02967f
C16685 VDD.n7359 GND 0.02522f
C16686 VDD.n7360 GND 0.04999f
C16687 VDD.t639 GND 0.63568f
C16688 VDD.n7361 GND 0.05074f
C16689 VDD.n7362 GND 0.05074f
C16690 VDD.n7363 GND 0.02967f
C16691 VDD.n7364 GND 0.02522f
C16692 VDD.t970 GND 0.02334f
C16693 VDD.t640 GND 0.02334f
C16694 VDD.n7365 GND 0.13341f
C16695 VDD.n7366 GND 0.0263f
C16696 VDD.n7367 GND 0.0536f
C16697 VDD.n7368 GND 0.05074f
C16698 VDD.n7369 GND 0.02967f
C16699 VDD.n7370 GND 0.02522f
C16700 VDD.n7371 GND 0.04999f
C16701 VDD.t652 GND 0.63568f
C16702 VDD.n7372 GND 0.05074f
C16703 VDD.n7373 GND 0.05074f
C16704 VDD.n7374 GND 0.02967f
C16705 VDD.n7375 GND 0.02522f
C16706 VDD.n7376 GND 0.03166f
C16707 VDD.n7377 GND 0.0536f
C16708 VDD.n7378 GND 0.05074f
C16709 VDD.n7379 GND 0.02967f
C16710 VDD.n7380 GND 0.02522f
C16711 VDD.n7381 GND 0.04999f
C16712 VDD.t544 GND 0.63568f
C16713 VDD.n7382 GND 0.05074f
C16714 VDD.n7383 GND 0.05074f
C16715 VDD.n7384 GND 0.02967f
C16716 VDD.n7385 GND 0.02522f
C16717 VDD.t653 GND 0.02321f
C16718 VDD.t874 GND 0.02321f
C16719 VDD.n7386 GND 0.10855f
C16720 VDD.t803 GND 0.02321f
C16721 VDD.t545 GND 0.02321f
C16722 VDD.n7387 GND 0.10855f
C16723 VDD.n7388 GND 0.04152f
C16724 VDD.n7389 GND 0.02334f
C16725 VDD.n7390 GND 0.0536f
C16726 VDD.n7391 GND 0.05074f
C16727 VDD.n7392 GND 0.02967f
C16728 VDD.n7393 GND 0.02522f
C16729 VDD.n7394 GND 0.02522f
C16730 VDD.n7395 GND 0.04999f
C16731 VDD.n7396 GND 0.68843f
C16732 VDD.n7397 GND 0.04999f
C16733 VDD.n7398 GND 0.05074f
C16734 VDD.n7399 GND 0.06295f
C16735 VDD.n7400 GND 0.0536f
C16736 VDD.n7401 GND 0.02522f
C16737 VDD.n7402 GND 0.04999f
C16738 VDD.n7403 GND 0.5126f
C16739 VDD.n7404 GND 0.02522f
C16740 VDD.n7405 GND 0.04999f
C16741 VDD.n7406 GND 0.5126f
C16742 VDD.n7407 GND 0.04999f
C16743 VDD.n7408 GND 0.05074f
C16744 VDD.n7409 GND 0.06295f
C16745 VDD.n7410 GND 0.0536f
C16746 VDD.n7411 GND 0.02522f
C16747 VDD.n7412 GND 0.04999f
C16748 VDD.n7413 GND 0.5126f
C16749 VDD.n7414 GND 0.02522f
C16750 VDD.n7415 GND 0.04999f
C16751 VDD.n7416 GND 0.5126f
C16752 VDD.n7417 GND 0.04999f
C16753 VDD.n7418 GND 0.05074f
C16754 VDD.n7419 GND 0.06295f
C16755 VDD.n7420 GND 0.0536f
C16756 VDD.n7421 GND 0.02522f
C16757 VDD.n7422 GND 0.04999f
C16758 VDD.n7423 GND 0.68843f
C16759 VDD.n7424 GND 0.02522f
C16760 VDD.n7425 GND 0.04999f
C16761 VDD.n7426 GND 0.68843f
C16762 VDD.n7427 GND 0.04999f
C16763 VDD.n7428 GND 0.05074f
C16764 VDD.n7429 GND 0.06295f
C16765 VDD.n7430 GND 0.0536f
C16766 VDD.n7431 GND 0.02522f
C16767 VDD.n7432 GND 0.04999f
C16768 VDD.n7433 GND 0.5126f
C16769 VDD.n7434 GND 0.02522f
C16770 VDD.n7435 GND 0.04999f
C16771 VDD.n7436 GND 0.5126f
C16772 VDD.n7437 GND 0.04999f
C16773 VDD.n7438 GND 0.05074f
C16774 VDD.n7439 GND 0.06295f
C16775 VDD.n7440 GND 0.0536f
C16776 VDD.n7441 GND 0.02522f
C16777 VDD.n7442 GND 0.04999f
C16778 VDD.n7443 GND 0.68843f
C16779 VDD.n7444 GND 0.68843f
C16780 VDD.n7445 GND 0.04999f
C16781 VDD.n7446 GND 0.02746f
C16782 VDD.n7447 GND 0.02967f
C16783 VDD.n7448 GND 0.02746f
C16784 VDD.n7449 GND 0.04999f
C16785 VDD.n7450 GND 0.68843f
C16786 VDD.n7451 GND 0.02522f
C16787 VDD.n7452 GND 0.04999f
C16788 VDD.n7453 GND 0.68843f
C16789 VDD.n7454 GND 0.04999f
C16790 VDD.n7455 GND 0.05074f
C16791 VDD.n7456 GND 0.06295f
C16792 VDD.n7457 GND 0.0536f
C16793 VDD.n7458 GND 0.02522f
C16794 VDD.n7459 GND 0.04999f
C16795 VDD.n7460 GND 0.5126f
C16796 VDD.n7461 GND 0.02522f
C16797 VDD.n7462 GND 0.04999f
C16798 VDD.n7463 GND 0.5126f
C16799 VDD.n7464 GND 0.04999f
C16800 VDD.n7465 GND 0.05074f
C16801 VDD.n7466 GND 0.06295f
C16802 VDD.n7467 GND 0.0536f
C16803 VDD.n7468 GND 0.02522f
C16804 VDD.n7469 GND 0.04999f
C16805 VDD.n7470 GND 0.5126f
C16806 VDD.n7471 GND 0.02522f
C16807 VDD.n7472 GND 0.04999f
C16808 VDD.n7473 GND 0.5126f
C16809 VDD.n7474 GND 0.04999f
C16810 VDD.n7475 GND 0.05074f
C16811 VDD.n7476 GND 0.06295f
C16812 VDD.n7477 GND 0.0536f
C16813 VDD.n7478 GND 0.02522f
C16814 VDD.n7479 GND 0.04999f
C16815 VDD.n7480 GND 0.68843f
C16816 VDD.n7481 GND 0.02522f
C16817 VDD.n7482 GND 0.04999f
C16818 VDD.n7483 GND 0.68843f
C16819 VDD.n7484 GND 0.04999f
C16820 VDD.n7485 GND 0.05074f
C16821 VDD.n7486 GND 0.06295f
C16822 VDD.n7487 GND 0.0536f
C16823 VDD.n7488 GND 0.02522f
C16824 VDD.n7489 GND 0.04999f
C16825 VDD.n7490 GND 0.5126f
C16826 VDD.n7491 GND 0.02522f
C16827 VDD.n7492 GND 0.04999f
C16828 VDD.n7493 GND 0.5126f
C16829 VDD.n7494 GND 0.04999f
C16830 VDD.n7495 GND 0.05074f
C16831 VDD.n7496 GND 0.06295f
C16832 VDD.n7497 GND 0.0536f
C16833 VDD.n7498 GND 0.02522f
C16834 VDD.n7499 GND 0.04999f
C16835 VDD.n7500 GND 0.5126f
C16836 VDD.n7501 GND 0.02522f
C16837 VDD.n7502 GND 0.04999f
C16838 VDD.n7503 GND 0.5126f
C16839 VDD.n7504 GND 0.04999f
C16840 VDD.n7505 GND 0.05074f
C16841 VDD.n7506 GND 0.06295f
C16842 VDD.n7507 GND 0.0536f
C16843 VDD.n7508 GND 0.02522f
C16844 VDD.n7509 GND 0.04999f
C16845 VDD.n7510 GND 0.68843f
C16846 VDD.n7511 GND 0.68843f
C16847 VDD.n7512 GND 0.04999f
C16848 VDD.n7513 GND 0.02746f
C16849 VDD.n7514 GND 0.09132f
C16850 VDD.n7515 GND 0.01798f
C16851 VDD.n7516 GND 0.09868f
C16852 VDD.n7517 GND 0.89643f
C16853 VDD.n7518 GND 0.3275f
C16854 VDD.n7519 GND 0.09868f
C16855 VDD.t251 GND 0.02334f
C16856 VDD.t242 GND 0.02334f
C16857 VDD.n7520 GND 0.13341f
C16858 VDD.n7521 GND 0.01798f
C16859 VDD.n7522 GND 0.09132f
C16860 VDD.n7523 GND 0.02746f
C16861 VDD.n7524 GND 0.04999f
C16862 VDD.n7525 GND 0.68843f
C16863 VDD.n7526 GND 0.02522f
C16864 VDD.n7527 GND 0.04999f
C16865 VDD.n7528 GND 0.68843f
C16866 VDD.n7529 GND 0.04999f
C16867 VDD.n7530 GND 0.05074f
C16868 VDD.n7531 GND 0.06295f
C16869 VDD.n7532 GND 0.0536f
C16870 VDD.n7533 GND 0.02522f
C16871 VDD.n7534 GND 0.04999f
C16872 VDD.n7535 GND 0.5126f
C16873 VDD.n7536 GND 0.02522f
C16874 VDD.n7537 GND 0.04999f
C16875 VDD.n7538 GND 0.5126f
C16876 VDD.n7539 GND 0.04999f
C16877 VDD.n7540 GND 0.05074f
C16878 VDD.n7541 GND 0.06295f
C16879 VDD.n7542 GND 0.0536f
C16880 VDD.n7543 GND 0.02522f
C16881 VDD.n7544 GND 0.04999f
C16882 VDD.n7545 GND 0.5126f
C16883 VDD.n7546 GND 0.02522f
C16884 VDD.n7547 GND 0.04999f
C16885 VDD.n7548 GND 0.5126f
C16886 VDD.n7549 GND 0.04999f
C16887 VDD.n7550 GND 0.05074f
C16888 VDD.n7551 GND 0.06295f
C16889 VDD.n7552 GND 0.0536f
C16890 VDD.n7553 GND 0.02522f
C16891 VDD.n7554 GND 0.04999f
C16892 VDD.n7555 GND 0.68843f
C16893 VDD.n7556 GND 0.68843f
C16894 VDD.n7557 GND 0.02522f
C16895 VDD.n7558 GND 0.02522f
C16896 VDD.n7559 GND 0.02967f
C16897 VDD.n7560 GND 0.05074f
C16898 VDD.n7561 GND 0.04999f
C16899 VDD.t224 GND 0.63568f
C16900 VDD.n7562 GND 0.05074f
C16901 VDD.n7563 GND 0.05074f
C16902 VDD.n7564 GND 0.02967f
C16903 VDD.n7565 GND 0.02522f
C16904 VDD.n7566 GND 0.0536f
C16905 VDD.n7567 GND 0.05074f
C16906 VDD.n7568 GND 0.02967f
C16907 VDD.n7569 GND 0.02522f
C16908 VDD.n7570 GND 0.04999f
C16909 VDD.t578 GND 0.63568f
C16910 VDD.n7571 GND 0.05074f
C16911 VDD.n7572 GND 0.05074f
C16912 VDD.n7573 GND 0.02967f
C16913 VDD.n7574 GND 0.02522f
C16914 VDD.t823 GND 0.02321f
C16915 VDD.t579 GND 0.02321f
C16916 VDD.n7575 GND 0.10855f
C16917 VDD.t225 GND 0.02321f
C16918 VDD.t637 GND 0.02321f
C16919 VDD.n7576 GND 0.10855f
C16920 VDD.n7577 GND 0.04152f
C16921 VDD.n7578 GND 0.02334f
C16922 VDD.n7579 GND 0.0536f
C16923 VDD.n7580 GND 0.05074f
C16924 VDD.n7581 GND 0.02967f
C16925 VDD.n7582 GND 0.02522f
C16926 VDD.t832 GND 0.63568f
C16927 VDD.n7583 GND 0.05074f
C16928 VDD.n7584 GND 0.05074f
C16929 VDD.n7585 GND 0.09132f
C16930 VDD.n7586 GND 0.04999f
C16931 VDD.t580 GND 0.63568f
C16932 VDD.n7587 GND 0.05074f
C16933 VDD.n7588 GND 0.05074f
C16934 VDD.n7589 GND 0.02967f
C16935 VDD.n7590 GND 0.02522f
C16936 VDD.t833 GND 0.02334f
C16937 VDD.n7591 GND 0.0731f
C16938 VDD.n7592 GND 0.01798f
C16939 VDD.n7593 GND 0.02334f
C16940 VDD.n7594 GND 0.0536f
C16941 VDD.n7595 GND 0.05074f
C16942 VDD.n7596 GND 0.02967f
C16943 VDD.n7597 GND 0.02522f
C16944 VDD.n7598 GND 0.04999f
C16945 VDD.t405 GND 0.63568f
C16946 VDD.n7599 GND 0.05074f
C16947 VDD.n7600 GND 0.05074f
C16948 VDD.n7601 GND 0.02967f
C16949 VDD.n7602 GND 0.02522f
C16950 VDD.t636 GND 0.02321f
C16951 VDD.t406 GND 0.02321f
C16952 VDD.n7603 GND 0.10855f
C16953 VDD.t581 GND 0.02321f
C16954 VDD.t407 GND 0.02321f
C16955 VDD.n7604 GND 0.10855f
C16956 VDD.n7605 GND 0.04152f
C16957 VDD.n7606 GND 0.02334f
C16958 VDD.n7607 GND 0.0536f
C16959 VDD.n7608 GND 0.05074f
C16960 VDD.n7609 GND 0.02967f
C16961 VDD.n7610 GND 0.02522f
C16962 VDD.n7611 GND 0.04999f
C16963 VDD.t73 GND 0.63568f
C16964 VDD.n7612 GND 0.05074f
C16965 VDD.n7613 GND 0.05074f
C16966 VDD.n7614 GND 0.02967f
C16967 VDD.n7615 GND 0.02522f
C16968 VDD.t74 GND 0.02334f
C16969 VDD.t210 GND 0.02334f
C16970 VDD.n7616 GND 0.13341f
C16971 VDD.n7617 GND 0.0263f
C16972 VDD.n7618 GND 0.0536f
C16973 VDD.n7619 GND 0.05074f
C16974 VDD.n7620 GND 0.02967f
C16975 VDD.n7621 GND 0.02522f
C16976 VDD.n7622 GND 0.04999f
C16977 VDD.t403 GND 0.63568f
C16978 VDD.n7623 GND 0.05074f
C16979 VDD.n7624 GND 0.05074f
C16980 VDD.n7625 GND 0.02967f
C16981 VDD.n7626 GND 0.02522f
C16982 VDD.n7627 GND 0.03166f
C16983 VDD.n7628 GND 0.0536f
C16984 VDD.n7629 GND 0.05074f
C16985 VDD.n7630 GND 0.02967f
C16986 VDD.n7631 GND 0.02522f
C16987 VDD.n7632 GND 0.04999f
C16988 VDD.t856 GND 0.63568f
C16989 VDD.n7633 GND 0.05074f
C16990 VDD.n7634 GND 0.05074f
C16991 VDD.n7635 GND 0.02967f
C16992 VDD.n7636 GND 0.02522f
C16993 VDD.t845 GND 0.02321f
C16994 VDD.t857 GND 0.02321f
C16995 VDD.n7637 GND 0.10855f
C16996 VDD.t404 GND 0.02321f
C16997 VDD.t901 GND 0.02321f
C16998 VDD.n7638 GND 0.10855f
C16999 VDD.n7639 GND 0.04152f
C17000 VDD.n7640 GND 0.02334f
C17001 VDD.n7641 GND 0.0536f
C17002 VDD.n7642 GND 0.05074f
C17003 VDD.n7643 GND 0.02967f
C17004 VDD.n7644 GND 0.02522f
C17005 VDD.n7645 GND 0.02522f
C17006 VDD.n7646 GND 0.04999f
C17007 VDD.n7647 GND 0.68843f
C17008 VDD.n7648 GND 0.04999f
C17009 VDD.n7649 GND 0.05074f
C17010 VDD.n7650 GND 0.06295f
C17011 VDD.n7651 GND 0.0536f
C17012 VDD.n7652 GND 0.02522f
C17013 VDD.n7653 GND 0.04999f
C17014 VDD.n7654 GND 0.5126f
C17015 VDD.n7655 GND 0.02522f
C17016 VDD.n7656 GND 0.04999f
C17017 VDD.n7657 GND 0.5126f
C17018 VDD.n7658 GND 0.04999f
C17019 VDD.n7659 GND 0.05074f
C17020 VDD.n7660 GND 0.06295f
C17021 VDD.n7661 GND 0.0536f
C17022 VDD.n7662 GND 0.02522f
C17023 VDD.n7663 GND 0.04999f
C17024 VDD.n7664 GND 0.5126f
C17025 VDD.n7665 GND 0.02522f
C17026 VDD.n7666 GND 0.04999f
C17027 VDD.n7667 GND 0.5126f
C17028 VDD.n7668 GND 0.04999f
C17029 VDD.n7669 GND 0.05074f
C17030 VDD.n7670 GND 0.06295f
C17031 VDD.n7671 GND 0.0536f
C17032 VDD.n7672 GND 0.02522f
C17033 VDD.n7673 GND 0.04999f
C17034 VDD.n7674 GND 0.68843f
C17035 VDD.n7675 GND 0.02522f
C17036 VDD.n7676 GND 0.04999f
C17037 VDD.n7677 GND 0.68843f
C17038 VDD.n7678 GND 0.04999f
C17039 VDD.n7679 GND 0.05074f
C17040 VDD.n7680 GND 0.06295f
C17041 VDD.n7681 GND 0.0536f
C17042 VDD.n7682 GND 0.02522f
C17043 VDD.n7683 GND 0.04999f
C17044 VDD.n7684 GND 0.5126f
C17045 VDD.n7685 GND 0.02522f
C17046 VDD.n7686 GND 0.04999f
C17047 VDD.n7687 GND 0.5126f
C17048 VDD.n7688 GND 0.04999f
C17049 VDD.n7689 GND 0.05074f
C17050 VDD.n7690 GND 0.06295f
C17051 VDD.n7691 GND 0.0536f
C17052 VDD.n7692 GND 0.02522f
C17053 VDD.n7693 GND 0.04999f
C17054 VDD.n7694 GND 0.68843f
C17055 VDD.n7695 GND 0.68843f
C17056 VDD.n7696 GND 0.04999f
C17057 VDD.n7697 GND 0.02746f
C17058 VDD.n7698 GND 0.02967f
C17059 VDD.n7699 GND 0.02746f
C17060 VDD.n7700 GND 0.04999f
C17061 VDD.n7701 GND 0.68843f
C17062 VDD.n7702 GND 0.02522f
C17063 VDD.n7703 GND 0.04999f
C17064 VDD.n7704 GND 0.68843f
C17065 VDD.n7705 GND 0.04999f
C17066 VDD.n7706 GND 0.05074f
C17067 VDD.n7707 GND 0.06295f
C17068 VDD.n7708 GND 0.0536f
C17069 VDD.n7709 GND 0.02522f
C17070 VDD.n7710 GND 0.04999f
C17071 VDD.n7711 GND 0.5126f
C17072 VDD.n7712 GND 0.02522f
C17073 VDD.n7713 GND 0.04999f
C17074 VDD.n7714 GND 0.5126f
C17075 VDD.n7715 GND 0.04999f
C17076 VDD.n7716 GND 0.05074f
C17077 VDD.n7717 GND 0.06295f
C17078 VDD.n7718 GND 0.0536f
C17079 VDD.n7719 GND 0.02522f
C17080 VDD.n7720 GND 0.04999f
C17081 VDD.n7721 GND 0.5126f
C17082 VDD.n7722 GND 0.5126f
C17083 VDD.n7723 GND 0.04999f
C17084 VDD.n7724 GND 0.04999f
C17085 VDD.n7725 GND 0.02522f
C17086 VDD.n7726 GND 0.02522f
C17087 VDD.n7727 GND 0.02967f
C17088 VDD.n7728 GND 0.05074f
C17089 VDD.t239 GND 0.63568f
C17090 VDD.n7729 GND 0.05074f
C17091 VDD.n7730 GND 0.06295f
C17092 VDD.n7731 GND 0.0263f
C17093 VDD.n7732 GND 0.13341f
C17094 Nand_Gate_4.A.t10 GND 0.27993f
C17095 Nand_Gate_4.A.n0 GND 0.08177f
C17096 Nand_Gate_4.A.n1 GND 0.03548f
C17097 Nand_Gate_4.A.n2 GND 0.15601f
C17098 Nand_Gate_4.A.t4 GND 0.1302f
C17099 Nand_Gate_4.A.n3 GND 0.04085f
C17100 Nand_Gate_4.A.t2 GND 0.03651f
C17101 Nand_Gate_4.A.n4 GND 0.159f
C17102 Nand_Gate_4.A.n5 GND 0.03942f
C17103 Nand_Gate_4.A.t5 GND 0.27994f
C17104 Nand_Gate_4.A.n6 GND 0.27511f
C17105 Nand_Gate_4.A.n7 GND 0.03007f
C17106 Nand_Gate_4.A.t11 GND 0.14554f
C17107 Nand_Gate_4.A.n8 GND 0.04192f
C17108 Nand_Gate_4.A.n9 GND 0.01797f
C17109 Nand_Gate_4.A.n10 GND 0.03367f
C17110 Nand_Gate_4.A.n11 GND 0.04236f
C17111 Nand_Gate_4.A.t9 GND 0.27994f
C17112 Nand_Gate_4.A.n12 GND 0.27511f
C17113 Nand_Gate_4.A.n13 GND 0.03007f
C17114 Nand_Gate_4.A.t7 GND 0.14554f
C17115 Nand_Gate_4.A.n14 GND 0.04192f
C17116 Nand_Gate_4.A.n15 GND 0.01797f
C17117 Nand_Gate_4.A.n16 GND 0.03367f
C17118 Nand_Gate_4.A.n18 GND 0.12656f
C17119 Nand_Gate_4.A.n19 GND 0.03459f
C17120 Nand_Gate_4.A.n20 GND 0.09204f
C17121 Nand_Gate_4.A.t8 GND 0.14555f
C17122 Nand_Gate_4.A.n21 GND 0.14257f
C17123 Nand_Gate_4.A.n22 GND 0.03007f
C17124 Nand_Gate_4.A.t6 GND 0.27993f
C17125 Nand_Gate_4.A.n23 GND 0.08177f
C17126 Nand_Gate_4.A.n24 GND 0.02035f
C17127 Nand_Gate_4.A.n25 GND 0.0296f
C17128 Nand_Gate_4.A.n26 GND 0.14551f
C17129 Nand_Gate_4.A.n27 GND 0.25531f
C17130 Nand_Gate_4.A.n28 GND 0.15873f
C17131 Nand_Gate_4.A.n29 GND 0.34318f
C17132 Nand_Gate_4.A.n31 GND 0.04546f
C17133 Nand_Gate_4.A.n32 GND 0.02608f
C17134 Nand_Gate_4.A.t1 GND 0.03876f
C17135 Nand_Gate_4.A.t0 GND 0.03797f
C17136 Nand_Gate_4.A.n33 GND 0.21593f
C17137 Nand_Gate_4.A.n34 GND 0.07184f
C17138 Nand_Gate_4.A.t3 GND 0.03797f
C17139 Nand_Gate_4.A.n35 GND 0.05849f
C17140 Nand_Gate_4.A.n36 GND 0.10356f
C17141 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 GND 0.07037f
C17142 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 GND 0.16004f
C17143 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 GND 0.07725f
C17144 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 GND 0.2799f
C17145 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 GND 0.27418f
C17146 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 GND 0.05783f
C17147 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 GND 0.53832f
C17148 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 GND 0.15726f
C17149 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 GND 0.03913f
C17150 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 GND 0.05692f
C17151 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 GND 0.14585f
C17152 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 GND 0.14585f
C17153 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 GND 0.07581f
C17154 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 GND 0.07318f
C17155 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 GND 0.07454f
C17156 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 GND 0.07302f
C17157 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 GND 0.41525f
C17158 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 GND 0.23391f
C17159 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 GND 0.22303f
C17160 CLK.t64 GND 0.34775f
C17161 CLK.n0 GND 0.36055f
C17162 CLK.n1 GND 0.03901f
C17163 CLK.n2 GND 0.05208f
C17164 CLK.t95 GND 0.16006f
C17165 CLK.n3 GND 0.13494f
C17166 CLK.n4 GND 0.04584f
C17167 CLK.t86 GND 0.34774f
C17168 CLK.t33 GND 0.1808f
C17169 CLK.n5 GND 0.19066f
C17170 CLK.t82 GND 0.34774f
C17171 CLK.n6 GND 0.30782f
C17172 CLK.n7 GND 0.30867f
C17173 CLK.n8 GND 0.19316f
C17174 CLK.t42 GND 0.16007f
C17175 CLK.n9 GND 0.01795f
C17176 CLK.n10 GND 0.04351f
C17177 CLK.n11 GND 0.46223f
C17178 CLK.t46 GND 0.34775f
C17179 CLK.n12 GND 0.36055f
C17180 CLK.n13 GND 0.03901f
C17181 CLK.n14 GND 0.05208f
C17182 CLK.t27 GND 0.16006f
C17183 CLK.n15 GND 0.13494f
C17184 CLK.n16 GND 0.04584f
C17185 CLK.t79 GND 0.34774f
C17186 CLK.t57 GND 0.1808f
C17187 CLK.n17 GND 0.19066f
C17188 CLK.t7 GND 0.34774f
C17189 CLK.n18 GND 0.30782f
C17190 CLK.n19 GND 0.30867f
C17191 CLK.n20 GND 0.19316f
C17192 CLK.t113 GND 0.16007f
C17193 CLK.n21 GND 0.01795f
C17194 CLK.n22 GND 0.04351f
C17195 CLK.n23 GND 0.161f
C17196 CLK.t9 GND 0.34775f
C17197 CLK.n24 GND 0.36055f
C17198 CLK.n25 GND 0.03901f
C17199 CLK.n26 GND 0.05208f
C17200 CLK.t117 GND 0.16006f
C17201 CLK.n27 GND 0.13494f
C17202 CLK.n28 GND 0.04584f
C17203 CLK.t36 GND 0.34774f
C17204 CLK.t88 GND 0.1808f
C17205 CLK.n29 GND 0.19066f
C17206 CLK.t73 GND 0.34774f
C17207 CLK.n30 GND 0.30782f
C17208 CLK.n31 GND 0.30867f
C17209 CLK.n32 GND 0.19316f
C17210 CLK.t70 GND 0.16007f
C17211 CLK.n33 GND 0.01795f
C17212 CLK.n34 GND 0.04351f
C17213 CLK.n35 GND 0.74111f
C17214 CLK.t71 GND 0.34775f
C17215 CLK.n36 GND 0.36055f
C17216 CLK.n37 GND 0.03901f
C17217 CLK.n38 GND 0.05208f
C17218 CLK.t54 GND 0.16006f
C17219 CLK.n39 GND 0.13494f
C17220 CLK.n40 GND 0.04584f
C17221 CLK.t112 GND 0.34774f
C17222 CLK.t28 GND 0.1808f
C17223 CLK.n41 GND 0.19066f
C17224 CLK.t101 GND 0.34774f
C17225 CLK.n42 GND 0.30782f
C17226 CLK.n43 GND 0.30867f
C17227 CLK.n44 GND 0.19316f
C17228 CLK.t19 GND 0.16007f
C17229 CLK.n45 GND 0.01795f
C17230 CLK.n46 GND 0.04351f
C17231 CLK.n48 GND 2.31789f
C17232 CLK.t99 GND 0.34775f
C17233 CLK.n49 GND 0.36055f
C17234 CLK.n50 GND 0.03901f
C17235 CLK.n51 GND 0.05208f
C17236 CLK.t84 GND 0.16006f
C17237 CLK.n52 GND 0.13494f
C17238 CLK.n53 GND 0.04584f
C17239 CLK.t14 GND 0.34774f
C17240 CLK.t55 GND 0.1808f
C17241 CLK.n54 GND 0.19066f
C17242 CLK.t4 GND 0.34774f
C17243 CLK.n55 GND 0.30782f
C17244 CLK.n56 GND 0.30867f
C17245 CLK.n57 GND 0.19316f
C17246 CLK.t38 GND 0.16007f
C17247 CLK.n58 GND 0.01795f
C17248 CLK.n59 GND 0.04351f
C17249 CLK.n61 GND 2.02899f
C17250 CLK.t41 GND 0.34775f
C17251 CLK.n62 GND 0.36055f
C17252 CLK.n63 GND 0.03901f
C17253 CLK.n64 GND 0.05208f
C17254 CLK.t114 GND 0.16006f
C17255 CLK.n65 GND 0.13494f
C17256 CLK.n66 GND 0.04584f
C17257 CLK.t76 GND 0.34774f
C17258 CLK.t11 GND 0.1808f
C17259 CLK.n67 GND 0.19066f
C17260 CLK.t66 GND 0.34774f
C17261 CLK.n68 GND 0.30782f
C17262 CLK.n69 GND 0.30867f
C17263 CLK.n70 GND 0.19316f
C17264 CLK.t63 GND 0.16007f
C17265 CLK.n71 GND 0.01795f
C17266 CLK.n72 GND 0.04351f
C17267 CLK.n74 GND 2.02899f
C17268 CLK.t65 GND 0.34775f
C17269 CLK.n75 GND 0.36055f
C17270 CLK.n76 GND 0.03901f
C17271 CLK.n77 GND 0.05208f
C17272 CLK.t51 GND 0.16006f
C17273 CLK.n78 GND 0.13494f
C17274 CLK.n79 GND 0.04584f
C17275 CLK.t109 GND 0.34774f
C17276 CLK.t25 GND 0.1808f
C17277 CLK.n80 GND 0.19066f
C17278 CLK.t92 GND 0.34774f
C17279 CLK.n81 GND 0.30782f
C17280 CLK.n82 GND 0.30867f
C17281 CLK.n83 GND 0.19316f
C17282 CLK.t16 GND 0.16007f
C17283 CLK.n84 GND 0.01795f
C17284 CLK.n85 GND 0.04351f
C17285 CLK.n87 GND 2.02899f
C17286 CLK.t91 GND 0.34775f
C17287 CLK.n88 GND 0.36055f
C17288 CLK.n89 GND 0.03901f
C17289 CLK.n90 GND 0.05208f
C17290 CLK.t80 GND 0.16006f
C17291 CLK.n91 GND 0.13494f
C17292 CLK.n92 GND 0.04584f
C17293 CLK.t12 GND 0.34774f
C17294 CLK.t52 GND 0.1808f
C17295 CLK.n93 GND 0.19066f
C17296 CLK.t32 GND 0.34774f
C17297 CLK.n94 GND 0.30782f
C17298 CLK.n95 GND 0.30867f
C17299 CLK.n96 GND 0.19316f
C17300 CLK.t30 GND 0.16007f
C17301 CLK.n97 GND 0.01795f
C17302 CLK.n98 GND 0.04351f
C17303 CLK.n100 GND 2.02899f
C17304 CLK.t20 GND 0.34775f
C17305 CLK.n101 GND 0.36055f
C17306 CLK.n102 GND 0.03901f
C17307 CLK.n103 GND 0.05208f
C17308 CLK.t13 GND 0.16006f
C17309 CLK.n104 GND 0.13494f
C17310 CLK.n105 GND 0.04584f
C17311 CLK.t50 GND 0.34774f
C17312 CLK.t31 GND 0.1808f
C17313 CLK.n106 GND 0.19066f
C17314 CLK.t104 GND 0.34774f
C17315 CLK.n107 GND 0.30782f
C17316 CLK.n108 GND 0.30867f
C17317 CLK.n109 GND 0.19316f
C17318 CLK.t83 GND 0.16007f
C17319 CLK.n110 GND 0.01795f
C17320 CLK.n111 GND 0.04351f
C17321 CLK.n113 GND 1.6993f
C17322 CLK.n114 GND 1.33849f
C17323 CLK.n115 GND 3.26289f
C17324 CLK.t77 GND 0.1808f
C17325 CLK.t3 GND 0.34774f
C17326 CLK.n116 GND 0.10158f
C17327 CLK.n117 GND 0.04344f
C17328 CLK.n118 GND 0.08021f
C17329 CLK.n119 GND 1.49061f
C17330 CLK.t105 GND 0.1808f
C17331 CLK.t21 GND 0.34774f
C17332 CLK.n120 GND 0.10158f
C17333 CLK.n121 GND 0.04344f
C17334 CLK.n122 GND 0.08021f
C17335 CLK.n123 GND 0.04177f
C17336 CLK.n124 GND 2.2385f
C17337 CLK.t18 GND 0.1808f
C17338 CLK.n125 GND 0.19316f
C17339 CLK.t49 GND 0.34774f
C17340 CLK.n126 GND 0.78151f
C17341 CLK.n127 GND 1.66232f
C17342 CLK.t44 GND 0.1808f
C17343 CLK.n128 GND 0.19316f
C17344 CLK.t81 GND 0.34774f
C17345 CLK.n129 GND 0.1094f
C17346 CLK.n130 GND 2.33217f
C17347 CLK.t87 GND 0.1808f
C17348 CLK.n131 GND 0.19316f
C17349 CLK.t48 GND 0.34774f
C17350 CLK.n132 GND 0.1094f
C17351 CLK.n133 GND 1.80643f
C17352 CLK.t34 GND 0.1808f
C17353 CLK.n134 GND 0.19316f
C17354 CLK.t43 GND 0.34774f
C17355 CLK.n135 GND 1.30135f
C17356 CLK.n136 GND 4.44918f
C17357 CLK.n137 GND 4.34264f
C17358 CLK.t74 GND 0.1808f
C17359 CLK.t115 GND 0.34774f
C17360 CLK.n138 GND 0.10158f
C17361 CLK.n139 GND 0.04344f
C17362 CLK.n140 GND 0.08021f
C17363 CLK.n141 GND 0.04177f
C17364 CLK.n142 GND 2.54051f
C17365 CLK.t110 GND 0.1808f
C17366 CLK.t61 GND 0.34774f
C17367 CLK.n143 GND 0.10158f
C17368 CLK.n144 GND 0.04344f
C17369 CLK.n145 GND 0.08021f
C17370 CLK.n146 GND 0.04177f
C17371 CLK.n147 GND 1.63439f
C17372 CLK.n148 GND 3.26269f
C17373 CLK.n149 GND 1.09574f
C17374 CLK.n150 GND 0.6418f
C17375 CLK.t68 GND 0.34775f
C17376 CLK.n151 GND 0.36055f
C17377 CLK.n152 GND 0.03901f
C17378 CLK.n153 GND 0.05208f
C17379 CLK.t102 GND 0.16006f
C17380 CLK.n154 GND 0.13494f
C17381 CLK.n155 GND 0.04584f
C17382 CLK.t90 GND 0.34774f
C17383 CLK.t17 GND 0.1808f
C17384 CLK.n156 GND 0.19066f
C17385 CLK.t106 GND 0.34774f
C17386 CLK.n157 GND 0.30782f
C17387 CLK.n158 GND 0.30867f
C17388 CLK.n159 GND 0.19316f
C17389 CLK.t45 GND 0.16007f
C17390 CLK.n160 GND 0.01795f
C17391 CLK.n161 GND 0.04351f
C17392 CLK.n162 GND 0.74111f
C17393 CLK.t96 GND 0.34775f
C17394 CLK.n163 GND 0.36055f
C17395 CLK.n164 GND 0.03901f
C17396 CLK.n165 GND 0.05208f
C17397 CLK.t5 GND 0.16006f
C17398 CLK.n166 GND 0.13494f
C17399 CLK.n167 GND 0.04584f
C17400 CLK.t0 GND 0.34774f
C17401 CLK.t78 GND 0.1808f
C17402 CLK.n168 GND 0.19066f
C17403 CLK.t10 GND 0.34774f
C17404 CLK.n169 GND 0.30782f
C17405 CLK.n170 GND 0.30867f
C17406 CLK.n171 GND 0.19316f
C17407 CLK.t69 GND 0.16007f
C17408 CLK.n172 GND 0.01795f
C17409 CLK.n173 GND 0.04351f
C17410 CLK.n175 GND 2.31789f
C17411 CLK.t35 GND 0.34775f
C17412 CLK.n176 GND 0.36055f
C17413 CLK.n177 GND 0.03901f
C17414 CLK.n178 GND 0.05208f
C17415 CLK.t22 GND 0.16006f
C17416 CLK.n179 GND 0.13494f
C17417 CLK.n180 GND 0.04584f
C17418 CLK.t56 GND 0.34774f
C17419 CLK.t111 GND 0.1808f
C17420 CLK.n181 GND 0.19066f
C17421 CLK.t24 GND 0.34774f
C17422 CLK.n182 GND 0.30782f
C17423 CLK.n183 GND 0.30867f
C17424 CLK.n184 GND 0.19316f
C17425 CLK.t97 GND 0.16007f
C17426 CLK.n185 GND 0.01795f
C17427 CLK.n186 GND 0.04351f
C17428 CLK.n188 GND 2.02899f
C17429 CLK.t60 GND 0.34775f
C17430 CLK.n189 GND 0.36055f
C17431 CLK.n190 GND 0.03901f
C17432 CLK.n191 GND 0.05208f
C17433 CLK.t93 GND 0.16006f
C17434 CLK.n192 GND 0.13494f
C17435 CLK.n193 GND 0.04584f
C17436 CLK.t85 GND 0.34774f
C17437 CLK.t47 GND 0.1808f
C17438 CLK.n194 GND 0.19066f
C17439 CLK.t103 GND 0.34774f
C17440 CLK.n195 GND 0.30782f
C17441 CLK.n196 GND 0.30867f
C17442 CLK.n197 GND 0.19316f
C17443 CLK.t37 GND 0.16007f
C17444 CLK.n198 GND 0.01795f
C17445 CLK.n199 GND 0.04351f
C17446 CLK.n201 GND 2.02899f
C17447 CLK.t89 GND 0.34775f
C17448 CLK.n202 GND 0.36055f
C17449 CLK.n203 GND 0.03901f
C17450 CLK.n204 GND 0.05208f
C17451 CLK.t2 GND 0.16006f
C17452 CLK.n205 GND 0.13494f
C17453 CLK.n206 GND 0.04584f
C17454 CLK.t116 GND 0.34774f
C17455 CLK.t75 GND 0.1808f
C17456 CLK.n207 GND 0.19066f
C17457 CLK.t6 GND 0.34774f
C17458 CLK.n208 GND 0.30782f
C17459 CLK.n209 GND 0.30867f
C17460 CLK.n210 GND 0.19316f
C17461 CLK.t62 GND 0.16007f
C17462 CLK.n211 GND 0.01795f
C17463 CLK.n212 GND 0.04351f
C17464 CLK.n214 GND 2.02899f
C17465 CLK.t29 GND 0.34775f
C17466 CLK.n215 GND 0.36055f
C17467 CLK.n216 GND 0.03901f
C17468 CLK.n217 GND 0.05208f
C17469 CLK.t59 GND 0.16006f
C17470 CLK.n218 GND 0.13494f
C17471 CLK.n219 GND 0.04584f
C17472 CLK.t53 GND 0.34774f
C17473 CLK.t108 GND 0.1808f
C17474 CLK.n220 GND 0.19066f
C17475 CLK.t67 GND 0.34774f
C17476 CLK.n221 GND 0.30782f
C17477 CLK.n222 GND 0.30867f
C17478 CLK.n223 GND 0.19316f
C17479 CLK.t15 GND 0.16007f
C17480 CLK.n224 GND 0.01795f
C17481 CLK.n225 GND 0.04351f
C17482 CLK.n227 GND 2.02899f
C17483 CLK.t98 GND 0.34775f
C17484 CLK.n228 GND 0.36055f
C17485 CLK.n229 GND 0.03901f
C17486 CLK.n230 GND 0.05208f
C17487 CLK.t8 GND 0.16006f
C17488 CLK.n231 GND 0.13494f
C17489 CLK.n232 GND 0.04584f
C17490 CLK.t1 GND 0.34774f
C17491 CLK.t26 GND 0.1808f
C17492 CLK.n233 GND 0.19066f
C17493 CLK.t94 GND 0.34774f
C17494 CLK.n234 GND 0.30782f
C17495 CLK.n235 GND 0.30867f
C17496 CLK.n236 GND 0.19316f
C17497 CLK.t72 GND 0.16007f
C17498 CLK.n237 GND 0.01795f
C17499 CLK.n238 GND 0.04351f
C17500 CLK.n240 GND 2.02899f
C17501 CLK.t40 GND 0.34775f
C17502 CLK.n241 GND 0.36055f
C17503 CLK.n242 GND 0.03901f
C17504 CLK.n243 GND 0.05208f
C17505 CLK.t23 GND 0.16006f
C17506 CLK.n244 GND 0.13494f
C17507 CLK.n245 GND 0.04584f
C17508 CLK.t58 GND 0.34774f
C17509 CLK.t39 GND 0.1808f
C17510 CLK.n246 GND 0.19066f
C17511 CLK.t107 GND 0.34774f
C17512 CLK.n247 GND 0.30782f
C17513 CLK.n248 GND 0.30867f
C17514 CLK.n249 GND 0.19316f
C17515 CLK.t100 GND 0.16007f
C17516 CLK.n250 GND 0.01795f
C17517 CLK.n251 GND 0.04351f
C17518 CLK.n253 GND 1.01773f
C17519 CLK.n254 GND 0.30418f
C17520 EN.t16 GND 0.26648f
C17521 EN.n0 GND 0.07676f
C17522 EN.n1 GND 0.02044f
C17523 EN.n2 GND 0.03186f
C17524 EN.t54 GND 0.51254f
C17525 EN.n3 GND 0.14973f
C17526 EN.n4 GND 0.06496f
C17527 EN.n5 GND 0.28564f
C17528 EN.t98 GND 0.23837f
C17529 EN.n6 GND 0.13678f
C17530 EN.n7 GND 0.42412f
C17531 EN.t74 GND 0.51256f
C17532 EN.n8 GND 0.51617f
C17533 EN.n9 GND 0.05506f
C17534 EN.t38 GND 0.26648f
C17535 EN.n10 GND 0.07676f
C17536 EN.n11 GND 0.02044f
C17537 EN.n12 GND 0.03186f
C17538 EN.n14 GND 0.82537f
C17539 EN.n15 GND 0.31786f
C17540 EN.n16 GND 0.05506f
C17541 EN.n17 GND 2.30076f
C17542 EN.t86 GND 0.51256f
C17543 EN.n18 GND 0.51617f
C17544 EN.n19 GND 0.05506f
C17545 EN.t106 GND 0.26648f
C17546 EN.n20 GND 0.07676f
C17547 EN.n21 GND 0.02044f
C17548 EN.n22 GND 0.03186f
C17549 EN.n23 GND 0.31786f
C17550 EN.t8 GND 0.51256f
C17551 EN.n24 GND 0.51617f
C17552 EN.n25 GND 0.05506f
C17553 EN.t29 GND 0.26648f
C17554 EN.n26 GND 0.07676f
C17555 EN.n27 GND 0.02044f
C17556 EN.n28 GND 0.03186f
C17557 EN.n30 GND 0.70792f
C17558 EN.t65 GND 0.51254f
C17559 EN.n31 GND 0.14973f
C17560 EN.n32 GND 0.06496f
C17561 EN.n33 GND 0.28564f
C17562 EN.t81 GND 0.23837f
C17563 EN.n34 GND 0.13678f
C17564 EN.n35 GND 0.31369f
C17565 EN.n36 GND 0.38752f
C17566 EN.t7 GND 0.51256f
C17567 EN.n37 GND 0.51617f
C17568 EN.n38 GND 0.05506f
C17569 EN.t26 GND 0.26648f
C17570 EN.n39 GND 0.07676f
C17571 EN.n40 GND 0.02044f
C17572 EN.n41 GND 0.03186f
C17573 EN.n42 GND 0.31786f
C17574 EN.t64 GND 0.51256f
C17575 EN.n43 GND 0.51617f
C17576 EN.n44 GND 0.05506f
C17577 EN.t49 GND 0.26648f
C17578 EN.n45 GND 0.07676f
C17579 EN.n46 GND 0.02044f
C17580 EN.n47 GND 0.03186f
C17581 EN.n49 GND 0.70792f
C17582 EN.t84 GND 0.51254f
C17583 EN.n50 GND 0.14973f
C17584 EN.n51 GND 0.06496f
C17585 EN.n52 GND 0.28564f
C17586 EN.t40 GND 0.23837f
C17587 EN.n53 GND 0.13678f
C17588 EN.n54 GND 0.31369f
C17589 EN.n55 GND 0.38752f
C17590 EN.n56 GND 2.22935f
C17591 EN.n57 GND 5.05735f
C17592 EN.t41 GND 0.51256f
C17593 EN.n58 GND 0.53143f
C17594 EN.n59 GND 0.05749f
C17595 EN.n60 GND 0.07676f
C17596 EN.t56 GND 0.2394f
C17597 EN.n61 GND 0.48121f
C17598 EN.n62 GND 0.13678f
C17599 EN.t61 GND 0.26649f
C17600 EN.n63 GND 0.24859f
C17601 EN.n64 GND 0.05506f
C17602 EN.t87 GND 0.51254f
C17603 EN.n65 GND 0.14973f
C17604 EN.n66 GND 0.04971f
C17605 EN.n67 GND 0.08397f
C17606 EN.n68 GND 0.31786f
C17607 EN.t6 GND 0.26649f
C17608 EN.n69 GND 0.24859f
C17609 EN.n70 GND 0.05506f
C17610 EN.t43 GND 0.51254f
C17611 EN.n71 GND 0.14973f
C17612 EN.n72 GND 0.04971f
C17613 EN.n73 GND 0.08397f
C17614 EN.n75 GND 0.80717f
C17615 EN.n76 GND 2.62416f
C17616 EN.n77 GND 2.4169f
C17617 EN.n78 GND 4.44397f
C17618 EN.n79 GND 7.08467f
C17619 EN.n80 GND 1.66156f
C17620 EN.n81 GND 2.30076f
C17621 EN.t27 GND 0.51256f
C17622 EN.n82 GND 0.51617f
C17623 EN.n83 GND 0.05506f
C17624 EN.t45 GND 0.26648f
C17625 EN.n84 GND 0.07676f
C17626 EN.n85 GND 0.02044f
C17627 EN.n86 GND 0.03186f
C17628 EN.n87 GND 0.31786f
C17629 EN.t83 GND 0.51256f
C17630 EN.n88 GND 0.51617f
C17631 EN.n89 GND 0.05506f
C17632 EN.t66 GND 0.26648f
C17633 EN.n90 GND 0.07676f
C17634 EN.n91 GND 0.02044f
C17635 EN.n92 GND 0.03186f
C17636 EN.n94 GND 0.70792f
C17637 EN.t102 GND 0.51254f
C17638 EN.n95 GND 0.14973f
C17639 EN.n96 GND 0.06496f
C17640 EN.n97 GND 0.28564f
C17641 EN.t60 GND 0.23837f
C17642 EN.n98 GND 0.13678f
C17643 EN.n99 GND 0.31369f
C17644 EN.n100 GND 0.38752f
C17645 EN.t11 GND 0.26648f
C17646 EN.n101 GND 0.07676f
C17647 EN.n102 GND 0.02044f
C17648 EN.n103 GND 0.03186f
C17649 EN.t70 GND 0.51254f
C17650 EN.n104 GND 0.14973f
C17651 EN.n105 GND 0.06496f
C17652 EN.n106 GND 0.28564f
C17653 EN.t35 GND 0.23837f
C17654 EN.n107 GND 0.13678f
C17655 EN.n108 GND 0.42412f
C17656 EN.t22 GND 0.51256f
C17657 EN.n109 GND 0.51617f
C17658 EN.n110 GND 0.05506f
C17659 EN.t18 GND 0.26648f
C17660 EN.n111 GND 0.07676f
C17661 EN.n112 GND 0.02044f
C17662 EN.n113 GND 0.03186f
C17663 EN.n115 GND 0.82537f
C17664 EN.n116 GND 0.31786f
C17665 EN.n117 GND 0.05506f
C17666 EN.n118 GND 0.51617f
C17667 EN.t19 GND 0.46087f
C17668 EN.n119 GND 2.30076f
C17669 EN.t4 GND 0.51256f
C17670 EN.n120 GND 0.51617f
C17671 EN.n121 GND 0.05506f
C17672 EN.t25 GND 0.26648f
C17673 EN.n122 GND 0.07676f
C17674 EN.n123 GND 0.02044f
C17675 EN.n124 GND 0.03186f
C17676 EN.n125 GND 0.31786f
C17677 EN.t0 GND 0.51256f
C17678 EN.n126 GND 0.51617f
C17679 EN.n127 GND 0.05506f
C17680 EN.t89 GND 0.26648f
C17681 EN.n128 GND 0.07676f
C17682 EN.n129 GND 0.02044f
C17683 EN.n130 GND 0.03186f
C17684 EN.n132 GND 0.70792f
C17685 EN.t32 GND 0.51254f
C17686 EN.n133 GND 0.14973f
C17687 EN.n134 GND 0.06496f
C17688 EN.n135 GND 0.28564f
C17689 EN.t77 GND 0.23837f
C17690 EN.n136 GND 0.13678f
C17691 EN.n137 GND 0.31369f
C17692 EN.n138 GND 0.38752f
C17693 EN.t12 GND 0.26649f
C17694 EN.n139 GND 0.24859f
C17695 EN.n140 GND 0.05506f
C17696 EN.t95 GND 0.51254f
C17697 EN.n141 GND 0.14973f
C17698 EN.n142 GND 0.04971f
C17699 EN.n143 GND 0.08397f
C17700 EN.n144 GND 0.31786f
C17701 EN.t10 GND 0.26649f
C17702 EN.n145 GND 0.24859f
C17703 EN.n146 GND 0.05506f
C17704 EN.t62 GND 0.51254f
C17705 EN.n147 GND 0.14973f
C17706 EN.n148 GND 0.04971f
C17707 EN.n149 GND 0.08397f
C17708 EN.n151 GND 0.70792f
C17709 EN.t20 GND 0.51256f
C17710 EN.n152 GND 0.53143f
C17711 EN.n153 GND 0.05749f
C17712 EN.n154 GND 0.07676f
C17713 EN.t42 GND 0.2394f
C17714 EN.n155 GND 0.48121f
C17715 EN.n156 GND 0.13678f
C17716 EN.n157 GND 0.24703f
C17717 EN.t93 GND 0.26648f
C17718 EN.n158 GND 0.07676f
C17719 EN.n159 GND 0.02044f
C17720 EN.n160 GND 0.03186f
C17721 EN.t3 GND 0.51254f
C17722 EN.n161 GND 0.14973f
C17723 EN.n162 GND 0.06496f
C17724 EN.n163 GND 0.28564f
C17725 EN.t37 GND 0.23837f
C17726 EN.n164 GND 0.13678f
C17727 EN.n165 GND 0.42412f
C17728 EN.t107 GND 0.51256f
C17729 EN.n166 GND 0.51617f
C17730 EN.n167 GND 0.05506f
C17731 EN.t101 GND 0.26648f
C17732 EN.n168 GND 0.07676f
C17733 EN.n169 GND 0.02044f
C17734 EN.n170 GND 0.03186f
C17735 EN.n172 GND 0.82537f
C17736 EN.n173 GND 0.31786f
C17737 EN.n174 GND 0.05506f
C17738 EN.n175 GND 0.51617f
C17739 EN.t73 GND 0.46087f
C17740 EN.t94 GND 0.26648f
C17741 EN.n176 GND 0.07676f
C17742 EN.n177 GND 0.02044f
C17743 EN.n178 GND 0.03186f
C17744 EN.t59 GND 0.51254f
C17745 EN.n179 GND 0.14973f
C17746 EN.n180 GND 0.06496f
C17747 EN.n181 GND 0.28564f
C17748 EN.t13 GND 0.23837f
C17749 EN.n182 GND 0.13678f
C17750 EN.n183 GND 0.42412f
C17751 EN.t57 GND 0.51256f
C17752 EN.n184 GND 0.51617f
C17753 EN.n185 GND 0.05506f
C17754 EN.t50 GND 0.26648f
C17755 EN.n186 GND 0.07676f
C17756 EN.n187 GND 0.02044f
C17757 EN.n188 GND 0.03186f
C17758 EN.n190 GND 0.82537f
C17759 EN.n191 GND 0.31786f
C17760 EN.n192 GND 0.05506f
C17761 EN.n193 GND 0.51617f
C17762 EN.t1 GND 0.83255f
C17763 EN.n194 GND 3.33243f
C17764 EN.n195 GND 4.67738f
C17765 EN.n196 GND 5.78002f
C17766 EN.t85 GND 0.51256f
C17767 EN.n197 GND 0.51617f
C17768 EN.n198 GND 0.05506f
C17769 EN.t104 GND 0.26648f
C17770 EN.n199 GND 0.07676f
C17771 EN.n200 GND 0.02044f
C17772 EN.n201 GND 0.03186f
C17773 EN.n202 GND 0.31786f
C17774 EN.t58 GND 0.51256f
C17775 EN.n203 GND 0.51617f
C17776 EN.n204 GND 0.05506f
C17777 EN.t71 GND 0.26648f
C17778 EN.n205 GND 0.07676f
C17779 EN.n206 GND 0.02044f
C17780 EN.n207 GND 0.03186f
C17781 EN.n209 GND 0.70792f
C17782 EN.t2 GND 0.51254f
C17783 EN.n210 GND 0.14973f
C17784 EN.n211 GND 0.06496f
C17785 EN.n212 GND 0.28564f
C17786 EN.t21 GND 0.23837f
C17787 EN.n213 GND 0.13678f
C17788 EN.n214 GND 0.31369f
C17789 EN.n215 GND 0.38752f
C17790 EN.t15 GND 0.26648f
C17791 EN.n216 GND 0.07676f
C17792 EN.n217 GND 0.02044f
C17793 EN.n218 GND 0.03186f
C17794 EN.t33 GND 0.51254f
C17795 EN.n219 GND 0.14973f
C17796 EN.n220 GND 0.06496f
C17797 EN.n221 GND 0.28564f
C17798 EN.t88 GND 0.23837f
C17799 EN.n222 GND 0.13678f
C17800 EN.n223 GND 0.42412f
C17801 EN.t28 GND 0.51256f
C17802 EN.n224 GND 0.51617f
C17803 EN.n225 GND 0.05506f
C17804 EN.t23 GND 0.26648f
C17805 EN.n226 GND 0.07676f
C17806 EN.n227 GND 0.02044f
C17807 EN.n228 GND 0.03186f
C17808 EN.n230 GND 0.82537f
C17809 EN.n231 GND 0.31786f
C17810 EN.n232 GND 0.05506f
C17811 EN.n233 GND 0.51617f
C17812 EN.t91 GND 0.46087f
C17813 EN.n234 GND 4.67738f
C17814 EN.n235 GND 5.05946f
C17815 EN.n236 GND 2.41971f
C17816 EN.n237 GND 2.30076f
C17817 EN.n238 GND 5.05946f
C17818 EN.t72 GND 0.26648f
C17819 EN.n239 GND 0.07676f
C17820 EN.n240 GND 0.02044f
C17821 EN.n241 GND 0.03186f
C17822 EN.t52 GND 0.51254f
C17823 EN.n242 GND 0.14973f
C17824 EN.n243 GND 0.06496f
C17825 EN.n244 GND 0.28564f
C17826 EN.t9 GND 0.23837f
C17827 EN.n245 GND 0.13678f
C17828 EN.n246 GND 0.42412f
C17829 EN.t82 GND 0.51256f
C17830 EN.n247 GND 0.51617f
C17831 EN.n248 GND 0.05506f
C17832 EN.t47 GND 0.26648f
C17833 EN.n249 GND 0.07676f
C17834 EN.n250 GND 0.02044f
C17835 EN.n251 GND 0.03186f
C17836 EN.n253 GND 0.82537f
C17837 EN.n254 GND 0.31786f
C17838 EN.n255 GND 0.05506f
C17839 EN.n256 GND 0.51617f
C17840 EN.t48 GND 0.46087f
C17841 EN.n257 GND 4.67738f
C17842 EN.n258 GND 2.30076f
C17843 EN.t63 GND 0.51256f
C17844 EN.n259 GND 0.51617f
C17845 EN.n260 GND 0.05506f
C17846 EN.t80 GND 0.26648f
C17847 EN.n261 GND 0.07676f
C17848 EN.n262 GND 0.02044f
C17849 EN.n263 GND 0.03186f
C17850 EN.n264 GND 0.31786f
C17851 EN.t31 GND 0.51256f
C17852 EN.n265 GND 0.51617f
C17853 EN.n266 GND 0.05506f
C17854 EN.t46 GND 0.26648f
C17855 EN.n267 GND 0.07676f
C17856 EN.n268 GND 0.02044f
C17857 EN.n269 GND 0.03186f
C17858 EN.n271 GND 0.70792f
C17859 EN.t51 GND 0.51254f
C17860 EN.n272 GND 0.14973f
C17861 EN.n273 GND 0.06496f
C17862 EN.n274 GND 0.28564f
C17863 EN.t96 GND 0.23837f
C17864 EN.n275 GND 0.13678f
C17865 EN.n276 GND 0.31369f
C17866 EN.n277 GND 0.38752f
C17867 EN.n278 GND 5.05946f
C17868 EN.t90 GND 0.26648f
C17869 EN.n279 GND 0.07676f
C17870 EN.n280 GND 0.02044f
C17871 EN.n281 GND 0.03186f
C17872 EN.t103 GND 0.51254f
C17873 EN.n282 GND 0.14973f
C17874 EN.n283 GND 0.06496f
C17875 EN.n284 GND 0.28564f
C17876 EN.t36 GND 0.23837f
C17877 EN.n285 GND 0.13678f
C17878 EN.n286 GND 0.42412f
C17879 EN.t99 GND 0.51256f
C17880 EN.n287 GND 0.51617f
C17881 EN.n288 GND 0.05506f
C17882 EN.t97 GND 0.26648f
C17883 EN.n289 GND 0.07676f
C17884 EN.n290 GND 0.02044f
C17885 EN.n291 GND 0.03186f
C17886 EN.n293 GND 0.82537f
C17887 EN.n294 GND 0.31786f
C17888 EN.n295 GND 0.05506f
C17889 EN.n296 GND 0.51617f
C17890 EN.t69 GND 0.46087f
C17891 EN.n297 GND 4.67738f
C17892 EN.n298 GND 2.30076f
C17893 EN.n299 GND 2.30076f
C17894 EN.n300 GND 4.67738f
C17895 EN.n301 GND 5.05946f
C17896 EN.n302 GND 2.30076f
C17897 EN.t68 GND 0.51256f
C17898 EN.n303 GND 0.51617f
C17899 EN.n304 GND 0.05506f
C17900 EN.t55 GND 0.26648f
C17901 EN.n305 GND 0.07676f
C17902 EN.n306 GND 0.02044f
C17903 EN.n307 GND 0.03186f
C17904 EN.n308 GND 0.31786f
C17905 EN.t100 GND 0.51256f
C17906 EN.n309 GND 0.51617f
C17907 EN.n310 GND 0.05506f
C17908 EN.t17 GND 0.26648f
C17909 EN.n311 GND 0.07676f
C17910 EN.n312 GND 0.02044f
C17911 EN.n313 GND 0.03186f
C17912 EN.n315 GND 0.70792f
C17913 EN.t24 GND 0.51254f
C17914 EN.n316 GND 0.14973f
C17915 EN.n317 GND 0.06496f
C17916 EN.n318 GND 0.28564f
C17917 EN.t76 GND 0.23837f
C17918 EN.n319 GND 0.13678f
C17919 EN.n320 GND 0.31369f
C17920 EN.n321 GND 0.38752f
C17921 EN.t67 GND 0.26648f
C17922 EN.n322 GND 0.07676f
C17923 EN.n323 GND 0.02044f
C17924 EN.n324 GND 0.03186f
C17925 EN.t5 GND 0.51254f
C17926 EN.n325 GND 0.14973f
C17927 EN.n326 GND 0.06496f
C17928 EN.n327 GND 0.28564f
C17929 EN.t39 GND 0.23837f
C17930 EN.n328 GND 0.13678f
C17931 EN.n329 GND 0.42412f
C17932 EN.t78 GND 0.51256f
C17933 EN.n330 GND 0.51617f
C17934 EN.n331 GND 0.05506f
C17935 EN.t92 GND 0.26648f
C17936 EN.n332 GND 0.07676f
C17937 EN.n333 GND 0.02044f
C17938 EN.n334 GND 0.03186f
C17939 EN.n336 GND 0.82537f
C17940 EN.n337 GND 0.31786f
C17941 EN.n338 GND 0.05506f
C17942 EN.n339 GND 0.51617f
C17943 EN.t44 GND 0.46087f
C17944 EN.n340 GND 4.67738f
C17945 EN.n341 GND 5.05946f
C17946 EN.n342 GND 2.30076f
C17947 EN.n343 GND 2.41971f
C17948 EN.n344 GND 5.05946f
C17949 EN.t75 GND 0.26648f
C17950 EN.n345 GND 0.07676f
C17951 EN.n346 GND 0.02044f
C17952 EN.n347 GND 0.03186f
C17953 EN.t34 GND 0.51254f
C17954 EN.n348 GND 0.14973f
C17955 EN.n349 GND 0.06496f
C17956 EN.n350 GND 0.28564f
C17957 EN.t79 GND 0.23837f
C17958 EN.n351 GND 0.13678f
C17959 EN.n352 GND 0.42412f
C17960 EN.t30 GND 0.51256f
C17961 EN.n353 GND 0.51617f
C17962 EN.n354 GND 0.05506f
C17963 EN.t14 GND 0.26648f
C17964 EN.n355 GND 0.07676f
C17965 EN.n356 GND 0.02044f
C17966 EN.n357 GND 0.03186f
C17967 EN.n359 GND 0.82537f
C17968 EN.n360 GND 0.31786f
C17969 EN.n361 GND 0.05506f
C17970 EN.n362 GND 0.51617f
C17971 EN.t53 GND 0.46087f
C17972 EN.n363 GND 4.67738f
C17973 EN.n364 GND 2.41971f
C17974 EN.n365 GND 1.27874f
C17975 EN.t105 GND 0.46087f
C17976 EN.n366 GND 0.51617f
C17977 CDAC8_0.switch_7.Z.t1 GND 0.03153f
C17978 CDAC8_0.switch_7.Z.t2 GND 0.03153f
C17979 CDAC8_0.switch_7.Z.n0 GND 0.1139f
C17980 CDAC8_0.switch_7.Z.n1 GND 0.26217f
C17981 CDAC8_0.switch_7.Z.t0 GND 0.0331f
C17982 CDAC8_0.switch_7.Z.n2 GND 2.15463f
C17983 CDAC8_0.switch_7.Z.n3 GND 0.71546f
C17984 CDAC8_0.switch_7.Z.t71 GND 5.56982f
C17985 CDAC8_0.switch_7.Z.n4 GND 1.29151f
C17986 CDAC8_0.switch_7.Z.n5 GND 0.84008f
C17987 CDAC8_0.switch_7.Z.t14 GND 5.56982f
C17988 CDAC8_0.switch_7.Z.n6 GND 1.29151f
C17989 CDAC8_0.switch_7.Z.t62 GND 5.56982f
C17990 CDAC8_0.switch_7.Z.n7 GND 1.29151f
C17991 CDAC8_0.switch_7.Z.n8 GND 0.71546f
C17992 CDAC8_0.switch_7.Z.n9 GND 1.0316f
C17993 CDAC8_0.switch_7.Z.t68 GND 5.56982f
C17994 CDAC8_0.switch_7.Z.n10 GND 1.29151f
C17995 CDAC8_0.switch_7.Z.t121 GND 5.56982f
C17996 CDAC8_0.switch_7.Z.n11 GND 1.29151f
C17997 CDAC8_0.switch_7.Z.t51 GND 5.56982f
C17998 CDAC8_0.switch_7.Z.n12 GND 1.29151f
C17999 CDAC8_0.switch_7.Z.n13 GND 1.0316f
C18000 CDAC8_0.switch_7.Z.t103 GND 5.56982f
C18001 CDAC8_0.switch_7.Z.n14 GND 1.29151f
C18002 CDAC8_0.switch_7.Z.n15 GND 1.0316f
C18003 CDAC8_0.switch_7.Z.t106 GND 5.56982f
C18004 CDAC8_0.switch_7.Z.n16 GND 1.43374f
C18005 CDAC8_0.switch_7.Z.t81 GND 5.56982f
C18006 CDAC8_0.switch_7.Z.n17 GND 1.63966f
C18007 CDAC8_0.switch_7.Z.n18 GND 1.0316f
C18008 CDAC8_0.switch_7.Z.t57 GND 5.56982f
C18009 CDAC8_0.switch_7.Z.n19 GND 1.29151f
C18010 CDAC8_0.switch_7.Z.n20 GND 0.84008f
C18011 CDAC8_0.switch_7.Z.t17 GND 5.56982f
C18012 CDAC8_0.switch_7.Z.n21 GND 1.29151f
C18013 CDAC8_0.switch_7.Z.n22 GND 0.84008f
C18014 CDAC8_0.switch_7.Z.t12 GND 5.56982f
C18015 CDAC8_0.switch_7.Z.n23 GND 1.29151f
C18016 CDAC8_0.switch_7.Z.n24 GND 0.84008f
C18017 CDAC8_0.switch_7.Z.t125 GND 5.56982f
C18018 CDAC8_0.switch_7.Z.n25 GND 1.29151f
C18019 CDAC8_0.switch_7.Z.n26 GND 0.84008f
C18020 CDAC8_0.switch_7.Z.t117 GND 5.6506f
C18021 CDAC8_0.switch_7.Z.t98 GND 5.6506f
C18022 CDAC8_0.switch_7.Z.t58 GND 5.56982f
C18023 CDAC8_0.switch_7.Z.n27 GND 1.29151f
C18024 CDAC8_0.switch_7.Z.n28 GND 1.0316f
C18025 CDAC8_0.switch_7.Z.t39 GND 5.56982f
C18026 CDAC8_0.switch_7.Z.n29 GND 1.29151f
C18027 CDAC8_0.switch_7.Z.n30 GND 1.0316f
C18028 CDAC8_0.switch_7.Z.t113 GND 5.56982f
C18029 CDAC8_0.switch_7.Z.n31 GND 1.29151f
C18030 CDAC8_0.switch_7.Z.n32 GND 1.0316f
C18031 CDAC8_0.switch_7.Z.t120 GND 5.56982f
C18032 CDAC8_0.switch_7.Z.n33 GND 1.29151f
C18033 CDAC8_0.switch_7.Z.n34 GND 1.0316f
C18034 CDAC8_0.switch_7.Z.t92 GND 5.56982f
C18035 CDAC8_0.switch_7.Z.n35 GND 1.29151f
C18036 CDAC8_0.switch_7.Z.n36 GND 2.08272f
C18037 CDAC8_0.switch_7.Z.t36 GND 5.6506f
C18038 CDAC8_0.switch_7.Z.n37 GND 0.60909f
C18039 CDAC8_0.switch_7.Z.t100 GND 5.56982f
C18040 CDAC8_0.switch_7.Z.n38 GND 1.29151f
C18041 CDAC8_0.switch_7.Z.n39 GND 0.60909f
C18042 CDAC8_0.switch_7.Z.t48 GND 5.56982f
C18043 CDAC8_0.switch_7.Z.n40 GND 1.29151f
C18044 CDAC8_0.switch_7.Z.n41 GND 0.60909f
C18045 CDAC8_0.switch_7.Z.t54 GND 5.56982f
C18046 CDAC8_0.switch_7.Z.n42 GND 1.29151f
C18047 CDAC8_0.switch_7.Z.n43 GND 0.60909f
C18048 CDAC8_0.switch_7.Z.t29 GND 5.56982f
C18049 CDAC8_0.switch_7.Z.n44 GND 1.29151f
C18050 CDAC8_0.switch_7.Z.n45 GND 1.66021f
C18051 CDAC8_0.switch_7.Z.n46 GND 0.84008f
C18052 CDAC8_0.switch_7.Z.t129 GND 5.6506f
C18053 CDAC8_0.switch_7.Z.n47 GND 2.08272f
C18054 CDAC8_0.switch_7.Z.n48 GND 0.84008f
C18055 CDAC8_0.switch_7.Z.n49 GND 1.66021f
C18056 CDAC8_0.switch_7.Z.t111 GND 5.56982f
C18057 CDAC8_0.switch_7.Z.n50 GND 1.29151f
C18058 CDAC8_0.switch_7.Z.n51 GND 0.60909f
C18059 CDAC8_0.switch_7.Z.n52 GND 0.84008f
C18060 CDAC8_0.switch_7.Z.n53 GND 1.0316f
C18061 CDAC8_0.switch_7.Z.t23 GND 5.56982f
C18062 CDAC8_0.switch_7.Z.n54 GND 1.29151f
C18063 CDAC8_0.switch_7.Z.n55 GND 1.0316f
C18064 CDAC8_0.switch_7.Z.n56 GND 0.84008f
C18065 CDAC8_0.switch_7.Z.n57 GND 0.60909f
C18066 CDAC8_0.switch_7.Z.t5 GND 5.56982f
C18067 CDAC8_0.switch_7.Z.n58 GND 1.29151f
C18068 CDAC8_0.switch_7.Z.n59 GND 0.60909f
C18069 CDAC8_0.switch_7.Z.n60 GND 0.84008f
C18070 CDAC8_0.switch_7.Z.n61 GND 1.0316f
C18071 CDAC8_0.switch_7.Z.t66 GND 5.56982f
C18072 CDAC8_0.switch_7.Z.n62 GND 1.29151f
C18073 CDAC8_0.switch_7.Z.t85 GND 5.56982f
C18074 CDAC8_0.switch_7.Z.n63 GND 1.29151f
C18075 CDAC8_0.switch_7.Z.n64 GND 1.0316f
C18076 CDAC8_0.switch_7.Z.n65 GND 0.84008f
C18077 CDAC8_0.switch_7.Z.n66 GND 0.60909f
C18078 CDAC8_0.switch_7.Z.t74 GND 5.56982f
C18079 CDAC8_0.switch_7.Z.n67 GND 1.29151f
C18080 CDAC8_0.switch_7.Z.n68 GND 0.60909f
C18081 CDAC8_0.switch_7.Z.n69 GND 0.84008f
C18082 CDAC8_0.switch_7.Z.n70 GND 0.84008f
C18083 CDAC8_0.switch_7.Z.n71 GND 0.60909f
C18084 CDAC8_0.switch_7.Z.t114 GND 5.56982f
C18085 CDAC8_0.switch_7.Z.n72 GND 1.29151f
C18086 CDAC8_0.switch_7.Z.n73 GND 0.60909f
C18087 CDAC8_0.switch_7.Z.n74 GND 0.87801f
C18088 CDAC8_0.switch_7.Z.n75 GND 1.0316f
C18089 CDAC8_0.switch_7.Z.t97 GND 5.56982f
C18090 CDAC8_0.switch_7.Z.n76 GND 1.29151f
C18091 CDAC8_0.switch_7.Z.n77 GND 0.60909f
C18092 CDAC8_0.switch_7.Z.t91 GND 5.56982f
C18093 CDAC8_0.switch_7.Z.n78 GND 1.29151f
C18094 CDAC8_0.switch_7.Z.t42 GND 5.56982f
C18095 CDAC8_0.switch_7.Z.n79 GND 1.29151f
C18096 CDAC8_0.switch_7.Z.n80 GND 0.84008f
C18097 CDAC8_0.switch_7.Z.t35 GND 5.56982f
C18098 CDAC8_0.switch_7.Z.n81 GND 1.29151f
C18099 CDAC8_0.switch_7.Z.t46 GND 5.56982f
C18100 CDAC8_0.switch_7.Z.n82 GND 1.29151f
C18101 CDAC8_0.switch_7.Z.n83 GND 0.84008f
C18102 CDAC8_0.switch_7.Z.t55 GND 5.56982f
C18103 CDAC8_0.switch_7.Z.n84 GND 1.29151f
C18104 CDAC8_0.switch_7.Z.n85 GND 0.84008f
C18105 CDAC8_0.switch_7.Z.t122 GND 5.56982f
C18106 CDAC8_0.switch_7.Z.n86 GND 1.29151f
C18107 CDAC8_0.switch_7.Z.n87 GND 0.84008f
C18108 CDAC8_0.switch_7.Z.t104 GND 5.56982f
C18109 CDAC8_0.switch_7.Z.n88 GND 1.29151f
C18110 CDAC8_0.switch_7.Z.n89 GND 0.84008f
C18111 CDAC8_0.switch_7.Z.t9 GND 5.79883f
C18112 CDAC8_0.switch_7.Z.n90 GND 0.71546f
C18113 CDAC8_0.switch_7.Z.t15 GND 5.56982f
C18114 CDAC8_0.switch_7.Z.n91 GND 1.29151f
C18115 CDAC8_0.switch_7.Z.n92 GND 0.84008f
C18116 CDAC8_0.switch_7.Z.t59 GND 5.56982f
C18117 CDAC8_0.switch_7.Z.n93 GND 1.29151f
C18118 CDAC8_0.switch_7.Z.t72 GND 5.56982f
C18119 CDAC8_0.switch_7.Z.n94 GND 1.29151f
C18120 CDAC8_0.switch_7.Z.n95 GND 0.84008f
C18121 CDAC8_0.switch_7.Z.t31 GND 5.56982f
C18122 CDAC8_0.switch_7.Z.n96 GND 1.29151f
C18123 CDAC8_0.switch_7.Z.n97 GND 0.84008f
C18124 CDAC8_0.switch_7.Z.t24 GND 5.56982f
C18125 CDAC8_0.switch_7.Z.n98 GND 1.29151f
C18126 CDAC8_0.switch_7.Z.n99 GND 0.84008f
C18127 CDAC8_0.switch_7.Z.t79 GND 5.56982f
C18128 CDAC8_0.switch_7.Z.n100 GND 1.29151f
C18129 CDAC8_0.switch_7.Z.n101 GND 0.84008f
C18130 CDAC8_0.switch_7.Z.t40 GND 5.79883f
C18131 CDAC8_0.switch_7.Z.t19 GND 5.79883f
C18132 CDAC8_0.switch_7.Z.n102 GND 2.24889f
C18133 CDAC8_0.switch_7.Z.t47 GND 5.56982f
C18134 CDAC8_0.switch_7.Z.n103 GND 1.29151f
C18135 CDAC8_0.switch_7.Z.t126 GND 5.56982f
C18136 CDAC8_0.switch_7.Z.n104 GND 1.29151f
C18137 CDAC8_0.switch_7.Z.n105 GND 1.0316f
C18138 CDAC8_0.switch_7.Z.t130 GND 5.56982f
C18139 CDAC8_0.switch_7.Z.n106 GND 1.29151f
C18140 CDAC8_0.switch_7.Z.n107 GND 1.0316f
C18141 CDAC8_0.switch_7.Z.t73 GND 5.56982f
C18142 CDAC8_0.switch_7.Z.n108 GND 1.29151f
C18143 CDAC8_0.switch_7.Z.n109 GND 1.0316f
C18144 CDAC8_0.switch_7.Z.t56 GND 5.56982f
C18145 CDAC8_0.switch_7.Z.n110 GND 1.29151f
C18146 CDAC8_0.switch_7.Z.n111 GND 1.0316f
C18147 CDAC8_0.switch_7.Z.t60 GND 5.56982f
C18148 CDAC8_0.switch_7.Z.n112 GND 1.29151f
C18149 CDAC8_0.switch_7.Z.n113 GND 1.0316f
C18150 CDAC8_0.switch_7.Z.t41 GND 5.56982f
C18151 CDAC8_0.switch_7.Z.n114 GND 1.29151f
C18152 CDAC8_0.switch_7.Z.n115 GND 1.0316f
C18153 CDAC8_0.switch_7.Z.t7 GND 5.56982f
C18154 CDAC8_0.switch_7.Z.n116 GND 1.29151f
C18155 CDAC8_0.switch_7.Z.t110 GND 5.56982f
C18156 CDAC8_0.switch_7.Z.n117 GND 1.29151f
C18157 CDAC8_0.switch_7.Z.n118 GND 1.0316f
C18158 CDAC8_0.switch_7.Z.t27 GND 5.56982f
C18159 CDAC8_0.switch_7.Z.n119 GND 1.29151f
C18160 CDAC8_0.switch_7.Z.t116 GND 5.56982f
C18161 CDAC8_0.switch_7.Z.n120 GND 1.29151f
C18162 CDAC8_0.switch_7.Z.n121 GND 1.0316f
C18163 CDAC8_0.switch_7.Z.n122 GND 0.71546f
C18164 CDAC8_0.switch_7.Z.t115 GND 5.56982f
C18165 CDAC8_0.switch_7.Z.n123 GND 1.29151f
C18166 CDAC8_0.switch_7.Z.n124 GND 0.84008f
C18167 CDAC8_0.switch_7.Z.t32 GND 5.56982f
C18168 CDAC8_0.switch_7.Z.n125 GND 1.29151f
C18169 CDAC8_0.switch_7.Z.n126 GND 0.84008f
C18170 CDAC8_0.switch_7.Z.t45 GND 5.56982f
C18171 CDAC8_0.switch_7.Z.n127 GND 1.29151f
C18172 CDAC8_0.switch_7.Z.n128 GND 0.84008f
C18173 CDAC8_0.switch_7.Z.t112 GND 5.56982f
C18174 CDAC8_0.switch_7.Z.n129 GND 1.29151f
C18175 CDAC8_0.switch_7.Z.n130 GND 0.84008f
C18176 CDAC8_0.switch_7.Z.t25 GND 5.56982f
C18177 CDAC8_0.switch_7.Z.n131 GND 1.29151f
C18178 CDAC8_0.switch_7.Z.n132 GND 0.84008f
C18179 CDAC8_0.switch_7.Z.t90 GND 5.6506f
C18180 CDAC8_0.switch_7.Z.t8 GND 5.6506f
C18181 CDAC8_0.switch_7.Z.t88 GND 5.56982f
C18182 CDAC8_0.switch_7.Z.n133 GND 1.29151f
C18183 CDAC8_0.switch_7.Z.n134 GND 1.0316f
C18184 CDAC8_0.switch_7.Z.t96 GND 5.56982f
C18185 CDAC8_0.switch_7.Z.n135 GND 1.29151f
C18186 CDAC8_0.switch_7.Z.n136 GND 1.0316f
C18187 CDAC8_0.switch_7.Z.t75 GND 5.56982f
C18188 CDAC8_0.switch_7.Z.n137 GND 1.29151f
C18189 CDAC8_0.switch_7.Z.n138 GND 1.0316f
C18190 CDAC8_0.switch_7.Z.t26 GND 5.56982f
C18191 CDAC8_0.switch_7.Z.n139 GND 1.29151f
C18192 CDAC8_0.switch_7.Z.n140 GND 1.0316f
C18193 CDAC8_0.switch_7.Z.t33 GND 5.56982f
C18194 CDAC8_0.switch_7.Z.n141 GND 1.29151f
C18195 CDAC8_0.switch_7.Z.n142 GND 1.0316f
C18196 CDAC8_0.switch_7.Z.t4 GND 5.56982f
C18197 CDAC8_0.switch_7.Z.n143 GND 1.29151f
C18198 CDAC8_0.switch_7.Z.n144 GND 2.08272f
C18199 CDAC8_0.switch_7.Z.t70 GND 5.6506f
C18200 CDAC8_0.switch_7.Z.n145 GND 0.60909f
C18201 CDAC8_0.switch_7.Z.t34 GND 5.56982f
C18202 CDAC8_0.switch_7.Z.n146 GND 1.29151f
C18203 CDAC8_0.switch_7.Z.n147 GND 0.60909f
C18204 CDAC8_0.switch_7.Z.t13 GND 5.56982f
C18205 CDAC8_0.switch_7.Z.n148 GND 1.29151f
C18206 CDAC8_0.switch_7.Z.n149 GND 0.60909f
C18207 CDAC8_0.switch_7.Z.t87 GND 5.56982f
C18208 CDAC8_0.switch_7.Z.n150 GND 1.29151f
C18209 CDAC8_0.switch_7.Z.n151 GND 0.60909f
C18210 CDAC8_0.switch_7.Z.t93 GND 5.56982f
C18211 CDAC8_0.switch_7.Z.n152 GND 1.29151f
C18212 CDAC8_0.switch_7.Z.n153 GND 0.60909f
C18213 CDAC8_0.switch_7.Z.t67 GND 5.56982f
C18214 CDAC8_0.switch_7.Z.n154 GND 1.29151f
C18215 CDAC8_0.switch_7.Z.n155 GND 1.66021f
C18216 CDAC8_0.switch_7.Z.n156 GND 0.84008f
C18217 CDAC8_0.switch_7.Z.t30 GND 5.6506f
C18218 CDAC8_0.switch_7.Z.n157 GND 1.66021f
C18219 CDAC8_0.switch_7.Z.n158 GND 0.84008f
C18220 CDAC8_0.switch_7.Z.n159 GND 2.08272f
C18221 CDAC8_0.switch_7.Z.t86 GND 5.56982f
C18222 CDAC8_0.switch_7.Z.n160 GND 1.29151f
C18223 CDAC8_0.switch_7.Z.n161 GND 1.0316f
C18224 CDAC8_0.switch_7.Z.n162 GND 0.84008f
C18225 CDAC8_0.switch_7.Z.n163 GND 0.60909f
C18226 CDAC8_0.switch_7.Z.t50 GND 5.56982f
C18227 CDAC8_0.switch_7.Z.n164 GND 1.29151f
C18228 CDAC8_0.switch_7.Z.n165 GND 0.60909f
C18229 CDAC8_0.switch_7.Z.n166 GND 0.84008f
C18230 CDAC8_0.switch_7.Z.n167 GND 1.0316f
C18231 CDAC8_0.switch_7.Z.t107 GND 5.56982f
C18232 CDAC8_0.switch_7.Z.n168 GND 1.29151f
C18233 CDAC8_0.switch_7.Z.n169 GND 1.0316f
C18234 CDAC8_0.switch_7.Z.n170 GND 0.84008f
C18235 CDAC8_0.switch_7.Z.n171 GND 0.60909f
C18236 CDAC8_0.switch_7.Z.t95 GND 5.56982f
C18237 CDAC8_0.switch_7.Z.n172 GND 1.29151f
C18238 CDAC8_0.switch_7.Z.n173 GND 0.60909f
C18239 CDAC8_0.switch_7.Z.n174 GND 0.84008f
C18240 CDAC8_0.switch_7.Z.n175 GND 1.0316f
C18241 CDAC8_0.switch_7.Z.t49 GND 5.56982f
C18242 CDAC8_0.switch_7.Z.n176 GND 1.29151f
C18243 CDAC8_0.switch_7.Z.t44 GND 5.56982f
C18244 CDAC8_0.switch_7.Z.n177 GND 1.29151f
C18245 CDAC8_0.switch_7.Z.n178 GND 1.0316f
C18246 CDAC8_0.switch_7.Z.n179 GND 0.84008f
C18247 CDAC8_0.switch_7.Z.n180 GND 0.60909f
C18248 CDAC8_0.switch_7.Z.t108 GND 5.56982f
C18249 CDAC8_0.switch_7.Z.n181 GND 1.29151f
C18250 CDAC8_0.switch_7.Z.n182 GND 0.60909f
C18251 CDAC8_0.switch_7.Z.n183 GND 0.84008f
C18252 CDAC8_0.switch_7.Z.n184 GND 0.84008f
C18253 CDAC8_0.switch_7.Z.n185 GND 0.60909f
C18254 CDAC8_0.switch_7.Z.t53 GND 5.56982f
C18255 CDAC8_0.switch_7.Z.n186 GND 1.29151f
C18256 CDAC8_0.switch_7.Z.n187 GND 0.60909f
C18257 CDAC8_0.switch_7.Z.n188 GND 0.84008f
C18258 CDAC8_0.switch_7.Z.t69 GND 5.56982f
C18259 CDAC8_0.switch_7.Z.n189 GND 1.17522f
C18260 CDAC8_0.switch_7.Z.t65 GND 5.56982f
C18261 CDAC8_0.switch_7.Z.n190 GND 1.29151f
C18262 CDAC8_0.switch_7.Z.n191 GND 1.0316f
C18263 CDAC8_0.switch_7.Z.n192 GND 0.84008f
C18264 CDAC8_0.switch_7.Z.n193 GND 0.60909f
C18265 CDAC8_0.switch_7.Z.t131 GND 5.56982f
C18266 CDAC8_0.switch_7.Z.n194 GND 1.29151f
C18267 CDAC8_0.switch_7.Z.n195 GND 0.60909f
C18268 CDAC8_0.switch_7.Z.n196 GND 0.84008f
C18269 CDAC8_0.switch_7.Z.n197 GND 0.84008f
C18270 CDAC8_0.switch_7.Z.n198 GND 0.60909f
C18271 CDAC8_0.switch_7.Z.t102 GND 5.56982f
C18272 CDAC8_0.switch_7.Z.n199 GND 1.29151f
C18273 CDAC8_0.switch_7.Z.n200 GND 0.60909f
C18274 CDAC8_0.switch_7.Z.t124 GND 5.56982f
C18275 CDAC8_0.switch_7.Z.n201 GND 1.29151f
C18276 CDAC8_0.switch_7.Z.n202 GND 0.60909f
C18277 CDAC8_0.switch_7.Z.t119 GND 5.56982f
C18278 CDAC8_0.switch_7.Z.n203 GND 1.29151f
C18279 CDAC8_0.switch_7.Z.n204 GND 0.60909f
C18280 CDAC8_0.switch_7.Z.t11 GND 5.56982f
C18281 CDAC8_0.switch_7.Z.n205 GND 1.29151f
C18282 CDAC8_0.switch_7.Z.n206 GND 0.60909f
C18283 CDAC8_0.switch_7.Z.t63 GND 5.56982f
C18284 CDAC8_0.switch_7.Z.n207 GND 1.29151f
C18285 CDAC8_0.switch_7.Z.n208 GND 0.60909f
C18286 CDAC8_0.switch_7.Z.t61 GND 5.56982f
C18287 CDAC8_0.switch_7.Z.n209 GND 1.29151f
C18288 CDAC8_0.switch_7.Z.t80 GND 5.79883f
C18289 CDAC8_0.switch_7.Z.n210 GND 1.82639f
C18290 CDAC8_0.switch_7.Z.n211 GND 0.84008f
C18291 CDAC8_0.switch_7.Z.t101 GND 5.79883f
C18292 CDAC8_0.switch_7.Z.n212 GND 2.24889f
C18293 CDAC8_0.switch_7.Z.n213 GND 0.84008f
C18294 CDAC8_0.switch_7.Z.n214 GND 1.82639f
C18295 CDAC8_0.switch_7.Z.t18 GND 5.56982f
C18296 CDAC8_0.switch_7.Z.n215 GND 1.29151f
C18297 CDAC8_0.switch_7.Z.n216 GND 0.60909f
C18298 CDAC8_0.switch_7.Z.n217 GND 0.84008f
C18299 CDAC8_0.switch_7.Z.n218 GND 1.0316f
C18300 CDAC8_0.switch_7.Z.t83 GND 5.56982f
C18301 CDAC8_0.switch_7.Z.n219 GND 1.29151f
C18302 CDAC8_0.switch_7.Z.n220 GND 1.0316f
C18303 CDAC8_0.switch_7.Z.n221 GND 0.84008f
C18304 CDAC8_0.switch_7.Z.n222 GND 0.60909f
C18305 CDAC8_0.switch_7.Z.t94 GND 5.56982f
C18306 CDAC8_0.switch_7.Z.n223 GND 1.29151f
C18307 CDAC8_0.switch_7.Z.n224 GND 0.60909f
C18308 CDAC8_0.switch_7.Z.n225 GND 0.84008f
C18309 CDAC8_0.switch_7.Z.n226 GND 1.0316f
C18310 CDAC8_0.switch_7.Z.t10 GND 5.56982f
C18311 CDAC8_0.switch_7.Z.n227 GND 1.29151f
C18312 CDAC8_0.switch_7.Z.n228 GND 1.0316f
C18313 CDAC8_0.switch_7.Z.n229 GND 0.84008f
C18314 CDAC8_0.switch_7.Z.n230 GND 0.60909f
C18315 CDAC8_0.switch_7.Z.t78 GND 5.56982f
C18316 CDAC8_0.switch_7.Z.n231 GND 1.29151f
C18317 CDAC8_0.switch_7.Z.n232 GND 0.60909f
C18318 CDAC8_0.switch_7.Z.n233 GND 0.84008f
C18319 CDAC8_0.switch_7.Z.n234 GND 1.0316f
C18320 CDAC8_0.switch_7.Z.t123 GND 5.56982f
C18321 CDAC8_0.switch_7.Z.n235 GND 1.17522f
C18322 CDAC8_0.switch_7.Z.n236 GND 3.78828f
C18323 CDAC8_0.switch_7.Z.n237 GND 3.78828f
C18324 CDAC8_0.switch_7.Z.t128 GND 5.56982f
C18325 CDAC8_0.switch_7.Z.n238 GND 1.17522f
C18326 CDAC8_0.switch_7.Z.n239 GND 1.0316f
C18327 CDAC8_0.switch_7.Z.t21 GND 5.56982f
C18328 CDAC8_0.switch_7.Z.n240 GND 1.29151f
C18329 CDAC8_0.switch_7.Z.n241 GND 1.0316f
C18330 CDAC8_0.switch_7.Z.t16 GND 5.56982f
C18331 CDAC8_0.switch_7.Z.n242 GND 1.29151f
C18332 CDAC8_0.switch_7.Z.n243 GND 1.0316f
C18333 CDAC8_0.switch_7.Z.t38 GND 5.56982f
C18334 CDAC8_0.switch_7.Z.n244 GND 1.29151f
C18335 CDAC8_0.switch_7.Z.n245 GND 1.0316f
C18336 CDAC8_0.switch_7.Z.t89 GND 5.56982f
C18337 CDAC8_0.switch_7.Z.n246 GND 1.29151f
C18338 CDAC8_0.switch_7.Z.n247 GND 1.0316f
C18339 CDAC8_0.switch_7.Z.t84 GND 5.56982f
C18340 CDAC8_0.switch_7.Z.n248 GND 1.29151f
C18341 CDAC8_0.switch_7.Z.t105 GND 5.79883f
C18342 CDAC8_0.switch_7.Z.n249 GND 2.24889f
C18343 CDAC8_0.switch_7.Z.n250 GND 0.60909f
C18344 CDAC8_0.switch_7.Z.t82 GND 5.56982f
C18345 CDAC8_0.switch_7.Z.n251 GND 1.29151f
C18346 CDAC8_0.switch_7.Z.n252 GND 0.60909f
C18347 CDAC8_0.switch_7.Z.t77 GND 5.56982f
C18348 CDAC8_0.switch_7.Z.n253 GND 1.29151f
C18349 CDAC8_0.switch_7.Z.n254 GND 0.60909f
C18350 CDAC8_0.switch_7.Z.t99 GND 5.56982f
C18351 CDAC8_0.switch_7.Z.n255 GND 1.29151f
C18352 CDAC8_0.switch_7.Z.n256 GND 0.60909f
C18353 CDAC8_0.switch_7.Z.t28 GND 5.56982f
C18354 CDAC8_0.switch_7.Z.n257 GND 1.29151f
C18355 CDAC8_0.switch_7.Z.n258 GND 0.60909f
C18356 CDAC8_0.switch_7.Z.t22 GND 5.56982f
C18357 CDAC8_0.switch_7.Z.n259 GND 1.29151f
C18358 CDAC8_0.switch_7.Z.t43 GND 5.79883f
C18359 CDAC8_0.switch_7.Z.n260 GND 1.82639f
C18360 CDAC8_0.switch_7.Z.n261 GND 0.84008f
C18361 CDAC8_0.switch_7.Z.t127 GND 5.79883f
C18362 CDAC8_0.switch_7.Z.n262 GND 1.82639f
C18363 CDAC8_0.switch_7.Z.n263 GND 0.84008f
C18364 CDAC8_0.switch_7.Z.n264 GND 2.24889f
C18365 CDAC8_0.switch_7.Z.t118 GND 5.56982f
C18366 CDAC8_0.switch_7.Z.n265 GND 1.29151f
C18367 CDAC8_0.switch_7.Z.n266 GND 1.0316f
C18368 CDAC8_0.switch_7.Z.n267 GND 0.84008f
C18369 CDAC8_0.switch_7.Z.n268 GND 0.60909f
C18370 CDAC8_0.switch_7.Z.t109 GND 5.56982f
C18371 CDAC8_0.switch_7.Z.n269 GND 1.29151f
C18372 CDAC8_0.switch_7.Z.n270 GND 0.60909f
C18373 CDAC8_0.switch_7.Z.n271 GND 0.84008f
C18374 CDAC8_0.switch_7.Z.n272 GND 1.0316f
C18375 CDAC8_0.switch_7.Z.t64 GND 5.56982f
C18376 CDAC8_0.switch_7.Z.n273 GND 1.29151f
C18377 CDAC8_0.switch_7.Z.n274 GND 1.0316f
C18378 CDAC8_0.switch_7.Z.n275 GND 0.84008f
C18379 CDAC8_0.switch_7.Z.n276 GND 0.60909f
C18380 CDAC8_0.switch_7.Z.t37 GND 5.56982f
C18381 CDAC8_0.switch_7.Z.n277 GND 1.29151f
C18382 CDAC8_0.switch_7.Z.n278 GND 0.60909f
C18383 CDAC8_0.switch_7.Z.n279 GND 0.84008f
C18384 CDAC8_0.switch_7.Z.n280 GND 1.0316f
C18385 CDAC8_0.switch_7.Z.t52 GND 5.56982f
C18386 CDAC8_0.switch_7.Z.n281 GND 1.29151f
C18387 CDAC8_0.switch_7.Z.n282 GND 1.0316f
C18388 CDAC8_0.switch_7.Z.n283 GND 0.84008f
C18389 CDAC8_0.switch_7.Z.n284 GND 0.60909f
C18390 CDAC8_0.switch_7.Z.t20 GND 5.56982f
C18391 CDAC8_0.switch_7.Z.n285 GND 1.29151f
C18392 CDAC8_0.switch_7.Z.n286 GND 0.60909f
C18393 CDAC8_0.switch_7.Z.n287 GND 0.84008f
C18394 CDAC8_0.switch_7.Z.n288 GND 0.84008f
C18395 CDAC8_0.switch_7.Z.n289 GND 0.60909f
C18396 CDAC8_0.switch_7.Z.t6 GND 5.56982f
C18397 CDAC8_0.switch_7.Z.n290 GND 1.29151f
C18398 CDAC8_0.switch_7.Z.n291 GND 0.60909f
C18399 CDAC8_0.switch_7.Z.n292 GND 0.84008f
C18400 CDAC8_0.switch_7.Z.n293 GND 1.0316f
C18401 CDAC8_0.switch_7.Z.t76 GND 5.56982f
C18402 CDAC8_0.switch_7.Z.n294 GND 1.17522f
C18403 CDAC8_0.switch_7.Z.n295 GND 2.11533f
C18404 CDAC8_0.switch_7.Z.n296 GND 3.3587f
C18405 CDAC8_0.switch_7.Z.n297 GND 0.13264f
C18406 CDAC8_0.switch_7.Z.t3 GND 0.03308f
.ends

