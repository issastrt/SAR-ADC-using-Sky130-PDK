magic
tech sky130A
magscale 1 2
timestamp 1756538730
<< error_p >>
rect -158 -2000 -100 2000
rect 100 -2000 158 2000
<< pwell >>
rect -328 2235 328 2258
rect -328 2147 -307 2235
rect -306 2147 328 2235
rect -328 -2258 328 2147
<< mvnmos >>
rect -100 -2000 100 2000
<< mvndiff >>
rect -158 1988 -100 2000
rect -158 -1988 -146 1988
rect -112 -1988 -100 1988
rect -158 -2000 -100 -1988
rect 100 1988 158 2000
rect 100 -1988 112 1988
rect 146 -1988 158 1988
rect 100 -2000 158 -1988
<< mvndiffc >>
rect -146 -1988 -112 1988
rect 112 -1988 146 1988
<< poly >>
rect -100 2072 100 2088
rect -100 2038 -84 2072
rect 84 2038 100 2072
rect -100 2000 100 2038
rect -100 -2038 100 -2000
rect -100 -2072 -84 -2038
rect 84 -2072 100 -2038
rect -100 -2088 100 -2072
<< polycont >>
rect -84 2038 84 2072
rect -84 -2072 84 -2038
<< locali >>
rect -100 2038 -84 2072
rect 84 2038 100 2072
rect -146 1988 -112 2004
rect -146 -2004 -112 -1988
rect 112 1988 146 2004
rect 112 -2004 146 -1988
rect -100 -2072 -84 -2038
rect 84 -2072 100 -2038
<< viali >>
rect -84 2038 84 2072
rect -146 -1988 -112 1988
rect 112 -1988 146 1988
rect -84 -2072 84 -2038
<< metal1 >>
rect -96 2072 96 2078
rect -96 2038 -84 2072
rect 84 2038 96 2072
rect -96 2032 96 2038
rect -152 1988 -106 2000
rect -152 -1988 -146 1988
rect -112 -1988 -106 1988
rect -152 -2000 -106 -1988
rect 106 1988 152 2000
rect 106 -1988 112 1988
rect 146 -1988 152 1988
rect 106 -2000 152 -1988
rect -96 -2038 96 -2032
rect -96 -2072 -84 -2038
rect 84 -2072 96 -2038
rect -96 -2078 96 -2072
<< properties >>
string FIXED_BBOX -262 -2192 262 2192
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_g5v0d10v5_53M7DK parameters
<< end >>
