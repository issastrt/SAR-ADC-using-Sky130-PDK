** sch_path: /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_22-00-39/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.418235294000 8.5u 0.418235294000 8.500001u 0.420000000000 17u 0.420000000000 17.000001u 0.421764705875 25.5u
+ 0.421764705875 25.500001u 0.423529411750 34u 0.423529411750 34.000001u 0.425294117625 42.5u 0.425294117625 42.500001u 0.427058823500 51u
+ 0.427058823500 51.000001u 0.428823529375 59.5u 0.428823529375 59.500001u 0.430588235250 68u 0.430588235250 68.000001u 0.432352941125 76.5u
+ 0.432352941125 76.500001u 0.434117647000 85u 0.434117647000 85.000001u 0.435882352875 93.5u 0.435882352875 93.500001u 0.437647058750 102u
+ 0.437647058750 102.000001u 0.439411764625 110.5u 0.439411764625 110.500001u 0.441176470500 119u 0.441176470500 119.000001u 0.442941176375 127.5u
+ 0.442941176375 127.500001u 0.444705882250 136u 0.444705882250 136.000001u 0.446470588125 144.5u 0.446470588125 144.500001u 0.448235294000 153u
+ 0.448235294000 153.000001u 0.450000000000 161.5u 0.450000000000 161.500001u 0.451764705875 170u 0.451764705875 170.000001u 0.453529411750 178.5u
+ 0.453529411750 178.500001u 0.455294117625 187u 0.455294117625 187.000001u 0.457058823500 195.5u 0.457058823500 195.500001u 0.458823529375 204u
+ 0.458823529375 204.000001u 0.460588235250 212.5u 0.460588235250 212.500001u 0.462352941125 221u 0.462352941125 221.000001u 0.464117647000 229.5u
+ 0.464117647000 229.500001u 0.465882352875 238u 0.465882352875 238.000001u 0.467647058750 246.5u 0.467647058750 246.500001u 0.469411764625 255u
+ 0.469411764625 255.000001u 0.471176470500 263.5u 0.471176470500 263.500001u 0.472941176375 272u 0.472941176375 272.000001u 0.474705882250 280.5u
+ 0.474705882250 280.500001u 0.476470588125 289u 0.476470588125 289.000001u 0.478235294000 297.5u 0.478235294000 297.500001u 0.480000000000 306u
+ 0.480000000000 306.000001u 0.481764705875 314.5u 0.481764705875 314.500001u 0.483529411750 323u 0.483529411750 323.000001u 0.485294117625 331.5u
+ 0.485294117625 331.500001u 0.487058823500 340u 0.487058823500 340.000001u 0.488823529375 348.5u 0.488823529375 348.500001u 0.490588235250 357u
+ 0.490588235250 357.000001u 0.492352941125 365.5u 0.492352941125 365.500001u 0.494117647000 374u 0.494117647000 374.000001u 0.495882352875 382.5u
+ 0.495882352875 382.500001u 0.497647058750 391u 0.497647058750 391.000001u 0.499411764625 399.5u 0.499411764625 399.500001u 0.501176470500 408u
+ 0.501176470500 408.000001u 0.502941176375 416.5u 0.502941176375 416.500001u 0.504705882250 425u 0.504705882250 425.000001u 0.506470588125 433.5u
+ 0.506470588125 433.500001u 0.508235294000 442u 0.508235294000 442.000001u 0.510000000000 450.5u 0.510000000000 450.500001u 0.511764705875 459u
+ 0.511764705875 459.000001u 0.513529411750 467.5u 0.513529411750 467.500001u 0.515294117625 476u 0.515294117625 476.000001u 0.517058823500 484.5u
+ 0.517058823500 484.500001u 0.518823529375 493u 0.518823529375 493.000001u 0.520588235250 501.5u 0.520588235250 501.500001u 0.522352941125 510u
+ 0.522352941125 510.000001u 0.524117647000 518.5u 0.524117647000 518.500001u 0.525882352875 527u 0.525882352875 527.000001u 0.527647058750 535.5u
+ 0.527647058750 535.500001u 0.529411764625 544u 0.529411764625 544.000001u 0.531176470500 552.5u 0.531176470500 552.500001u 0.532941176375 561u
+ 0.532941176375 561.000001u 0.534705882250 569.5u 0.534705882250 569.500001u 0.536470588125 578u 0.536470588125 578.000001u 0.538235294000 586.5u
+ 0.538235294000 586.500001u 0.540000000000 595u 0.540000000000 595.000001u 0.541764705875 603.5u 0.541764705875 603.500001u 0.543529411750 612u
+ 0.543529411750 612.000001u 0.545294117625 620.5u 0.545294117625 620.500001u 0.547058823500 629u 0.547058823500 629.000001u 0.548823529375 637.5u
+ 0.548823529375 637.500001u 0.550588235250 646u 0.550588235250 646.000001u 0.552352941125 654.5u 0.552352941125 654.500001u 0.554117647000 663u
+ 0.554117647000 663.000001u 0.555882352875 671.5u 0.555882352875 671.500001u 0.557647058750 680u 0.557647058750)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/madra/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 680u uic
  wrdata /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_22-00-39/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
