** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_02-12-45/parameters/SNDR/run_4/sndr_enob_fom.sch
**.subckt sndr_enob_fom
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VVin Vin GND SIN(0.9 0.85 229.7794 0 0 45)
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
R1 net1 GND 0.01 m=1
**** begin user architecture code

.control
tran 0.5u 272u uic
set wr_singlescale
wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_02-12-45/parameters/SNDR/run_4/sndr_enob_fom_4.data -I(VVDD) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0) V(Vin)
quit
.endc



* CACE gensim simulation file sndr_enob_fom_4
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice sf

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
