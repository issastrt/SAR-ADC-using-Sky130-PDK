magic
tech sky130A
magscale 1 2
timestamp 1757231656
<< metal1 >>
rect 7136 46724 7200 46730
rect 7136 46721 7142 46724
rect 6634 46675 7142 46721
rect 7136 46672 7142 46675
rect 7194 46721 7200 46724
rect 11080 46724 11144 46730
rect 11080 46721 11086 46724
rect 7194 46675 11086 46721
rect 7194 46672 7200 46675
rect 7136 46666 7200 46672
rect 11080 46672 11086 46675
rect 11138 46721 11144 46724
rect 15024 46724 15088 46730
rect 15024 46721 15030 46724
rect 11138 46675 15030 46721
rect 11138 46672 11144 46675
rect 11080 46666 11144 46672
rect 15024 46672 15030 46675
rect 15082 46721 15088 46724
rect 18968 46724 19032 46730
rect 18968 46721 18974 46724
rect 15082 46675 18974 46721
rect 15082 46672 15088 46675
rect 15024 46666 15088 46672
rect 18968 46672 18974 46675
rect 19026 46721 19032 46724
rect 22912 46724 22976 46730
rect 22912 46721 22918 46724
rect 19026 46675 22918 46721
rect 19026 46672 19032 46675
rect 18968 46666 19032 46672
rect 22912 46672 22918 46675
rect 22970 46721 22976 46724
rect 26856 46724 26920 46730
rect 26856 46721 26862 46724
rect 22970 46675 26862 46721
rect 22970 46672 22976 46675
rect 22912 46666 22976 46672
rect 26856 46672 26862 46675
rect 26914 46721 26920 46724
rect 30800 46724 30864 46730
rect 30800 46721 30806 46724
rect 26914 46675 30806 46721
rect 26914 46672 26920 46675
rect 26856 46666 26920 46672
rect 30800 46672 30806 46675
rect 30858 46721 30864 46724
rect 34744 46724 34808 46730
rect 34744 46721 34750 46724
rect 30858 46675 34750 46721
rect 30858 46672 30864 46675
rect 30800 46666 30864 46672
rect 34744 46672 34750 46675
rect 34802 46721 34808 46724
rect 34802 46675 36214 46721
rect 34802 46672 34808 46675
rect 34744 46666 34808 46672
rect 7597 45865 8257 45911
rect 11541 45865 12201 45911
rect 15485 45865 16145 45911
rect 19429 45865 20089 45911
rect 23373 45865 24033 45911
rect 27317 45865 27977 45911
rect 31261 45865 31921 45911
rect 35205 45865 35865 45911
rect 7281 45590 7345 45596
rect 7281 45538 7287 45590
rect 7339 45538 7345 45590
rect 7281 45532 7345 45538
rect 11225 45590 11289 45596
rect 11225 45538 11231 45590
rect 11283 45538 11289 45590
rect 11225 45532 11289 45538
rect 15169 45590 15233 45596
rect 15169 45538 15175 45590
rect 15227 45538 15233 45590
rect 15169 45532 15233 45538
rect 19113 45590 19177 45596
rect 19113 45538 19119 45590
rect 19171 45538 19177 45590
rect 19113 45532 19177 45538
rect 23057 45590 23121 45596
rect 23057 45538 23063 45590
rect 23115 45538 23121 45590
rect 23057 45532 23121 45538
rect 27001 45590 27065 45596
rect 27001 45538 27007 45590
rect 27059 45538 27065 45590
rect 27001 45532 27065 45538
rect 30945 45590 31009 45596
rect 30945 45538 30951 45590
rect 31003 45538 31009 45590
rect 30945 45532 31009 45538
rect 34889 45590 34953 45596
rect 34889 45538 34895 45590
rect 34947 45538 34953 45590
rect 34889 45532 34953 45538
rect 362 44942 426 44948
rect 362 44890 368 44942
rect 420 44939 426 44942
rect 2794 44942 2858 44948
rect 2794 44939 2800 44942
rect 420 44893 2800 44939
rect 420 44890 426 44893
rect 362 44884 426 44890
rect 2794 44890 2800 44893
rect 2852 44939 2858 44942
rect 5226 44942 5290 44948
rect 5226 44939 5232 44942
rect 2852 44893 5232 44939
rect 2852 44890 2858 44893
rect 2794 44884 2858 44890
rect 5226 44890 5232 44893
rect 5284 44939 5290 44942
rect 7426 44942 7490 44948
rect 7426 44939 7432 44942
rect 5284 44893 7432 44939
rect 5284 44890 5290 44893
rect 5226 44884 5290 44890
rect 7426 44890 7432 44893
rect 7484 44939 7490 44942
rect 7658 44942 7722 44948
rect 7658 44939 7664 44942
rect 7484 44893 7664 44939
rect 7484 44890 7490 44893
rect 7426 44884 7490 44890
rect 7658 44890 7664 44893
rect 7716 44939 7722 44942
rect 10090 44942 10154 44948
rect 10090 44939 10096 44942
rect 7716 44893 10096 44939
rect 7716 44890 7722 44893
rect 7658 44884 7722 44890
rect 10090 44890 10096 44893
rect 10148 44939 10154 44942
rect 11370 44942 11434 44948
rect 11370 44939 11376 44942
rect 10148 44893 11376 44939
rect 10148 44890 10154 44893
rect 10090 44884 10154 44890
rect 11370 44890 11376 44893
rect 11428 44939 11434 44942
rect 12522 44942 12586 44948
rect 12522 44939 12528 44942
rect 11428 44893 12528 44939
rect 11428 44890 11434 44893
rect 11370 44884 11434 44890
rect 12522 44890 12528 44893
rect 12580 44939 12586 44942
rect 14954 44942 15018 44948
rect 14954 44939 14960 44942
rect 12580 44893 14960 44939
rect 12580 44890 12586 44893
rect 12522 44884 12586 44890
rect 14954 44890 14960 44893
rect 15012 44939 15018 44942
rect 15314 44942 15378 44948
rect 15314 44939 15320 44942
rect 15012 44893 15320 44939
rect 15012 44890 15018 44893
rect 14954 44884 15018 44890
rect 15314 44890 15320 44893
rect 15372 44939 15378 44942
rect 17386 44942 17450 44948
rect 17386 44939 17392 44942
rect 15372 44893 17392 44939
rect 15372 44890 15378 44893
rect 15314 44884 15378 44890
rect 17386 44890 17392 44893
rect 17444 44939 17450 44942
rect 19258 44942 19322 44948
rect 19258 44939 19264 44942
rect 17444 44893 19264 44939
rect 17444 44890 17450 44893
rect 17386 44884 17450 44890
rect 19258 44890 19264 44893
rect 19316 44939 19322 44942
rect 19818 44942 19882 44948
rect 19818 44939 19824 44942
rect 19316 44893 19824 44939
rect 19316 44890 19322 44893
rect 19258 44884 19322 44890
rect 19818 44890 19824 44893
rect 19876 44939 19882 44942
rect 22250 44942 22314 44948
rect 22250 44939 22256 44942
rect 19876 44893 22256 44939
rect 19876 44890 19882 44893
rect 19818 44884 19882 44890
rect 22250 44890 22256 44893
rect 22308 44939 22314 44942
rect 23202 44942 23266 44948
rect 23202 44939 23208 44942
rect 22308 44893 23208 44939
rect 22308 44890 22314 44893
rect 22250 44884 22314 44890
rect 23202 44890 23208 44893
rect 23260 44939 23266 44942
rect 24682 44942 24746 44948
rect 24682 44939 24688 44942
rect 23260 44893 24688 44939
rect 23260 44890 23266 44893
rect 23202 44884 23266 44890
rect 24682 44890 24688 44893
rect 24740 44939 24746 44942
rect 27146 44942 27210 44948
rect 27146 44939 27152 44942
rect 24740 44893 27152 44939
rect 24740 44890 24746 44893
rect 24682 44884 24746 44890
rect 27146 44890 27152 44893
rect 27204 44939 27210 44942
rect 29546 44942 29610 44948
rect 29546 44939 29552 44942
rect 27204 44893 29552 44939
rect 27204 44890 27210 44893
rect 27146 44884 27210 44890
rect 29546 44890 29552 44893
rect 29604 44939 29610 44942
rect 31090 44942 31154 44948
rect 31090 44939 31096 44942
rect 29604 44893 31096 44939
rect 29604 44890 29610 44893
rect 29546 44884 29610 44890
rect 31090 44890 31096 44893
rect 31148 44939 31154 44942
rect 31978 44942 32042 44948
rect 31978 44939 31984 44942
rect 31148 44893 31984 44939
rect 31148 44890 31154 44893
rect 31090 44884 31154 44890
rect 31978 44890 31984 44893
rect 32036 44939 32042 44942
rect 34410 44942 34474 44948
rect 34410 44939 34416 44942
rect 32036 44893 34416 44939
rect 32036 44890 32042 44893
rect 31978 44884 32042 44890
rect 34410 44890 34416 44893
rect 34468 44939 34474 44942
rect 35034 44942 35098 44948
rect 35034 44939 35040 44942
rect 34468 44893 35040 44939
rect 34468 44890 34474 44893
rect 34410 44884 34474 44890
rect 35034 44890 35040 44893
rect 35092 44939 35098 44942
rect 36842 44942 36906 44948
rect 36842 44939 36848 44942
rect 35092 44893 36848 44939
rect 35092 44890 35098 44893
rect 35034 44884 35098 44890
rect 36842 44890 36848 44893
rect 36900 44939 36906 44942
rect 39274 44942 39338 44948
rect 39274 44939 39280 44942
rect 36900 44893 39280 44939
rect 36900 44890 36906 44893
rect 36842 44884 36906 44890
rect 39274 44890 39280 44893
rect 39332 44939 39338 44942
rect 41706 44942 41770 44948
rect 41706 44939 41712 44942
rect 39332 44893 41712 44939
rect 39332 44890 39338 44893
rect 39274 44884 39338 44890
rect 41706 44890 41712 44893
rect 41764 44890 41770 44942
rect 41706 44884 41770 44890
<< via1 >>
rect 7142 46672 7194 46724
rect 11086 46672 11138 46724
rect 15030 46672 15082 46724
rect 18974 46672 19026 46724
rect 22918 46672 22970 46724
rect 26862 46672 26914 46724
rect 30806 46672 30858 46724
rect 34750 46672 34802 46724
rect 7287 45538 7339 45590
rect 11231 45538 11283 45590
rect 15175 45538 15227 45590
rect 19119 45538 19171 45590
rect 23063 45538 23115 45590
rect 27007 45538 27059 45590
rect 30951 45538 31003 45590
rect 34895 45538 34947 45590
rect 368 44890 420 44942
rect 2800 44890 2852 44942
rect 5232 44890 5284 44942
rect 7432 44890 7484 44942
rect 7664 44890 7716 44942
rect 10096 44890 10148 44942
rect 11376 44890 11428 44942
rect 12528 44890 12580 44942
rect 14960 44890 15012 44942
rect 15320 44890 15372 44942
rect 17392 44890 17444 44942
rect 19264 44890 19316 44942
rect 19824 44890 19876 44942
rect 22256 44890 22308 44942
rect 23208 44890 23260 44942
rect 24688 44890 24740 44942
rect 27152 44890 27204 44942
rect 29552 44890 29604 44942
rect 31096 44890 31148 44942
rect 31984 44890 32036 44942
rect 34416 44890 34468 44942
rect 35040 44890 35092 44942
rect 36848 44890 36900 44942
rect 39280 44890 39332 44942
rect 41712 44890 41764 44942
<< metal2 >>
rect 7131 46726 7205 46735
rect 7131 46670 7140 46726
rect 7196 46670 7205 46726
rect 7131 46661 7205 46670
rect 11075 46726 11149 46735
rect 11075 46670 11084 46726
rect 11140 46670 11149 46726
rect 11075 46661 11149 46670
rect 15019 46726 15093 46735
rect 15019 46670 15028 46726
rect 15084 46670 15093 46726
rect 15019 46661 15093 46670
rect 18963 46726 19037 46735
rect 18963 46670 18972 46726
rect 19028 46670 19037 46726
rect 18963 46661 19037 46670
rect 22907 46726 22981 46735
rect 22907 46670 22916 46726
rect 22972 46670 22981 46726
rect 22907 46661 22981 46670
rect 26851 46726 26925 46735
rect 26851 46670 26860 46726
rect 26916 46670 26925 46726
rect 26851 46661 26925 46670
rect 30795 46726 30869 46735
rect 30795 46670 30804 46726
rect 30860 46670 30869 46726
rect 30795 46661 30869 46670
rect 34739 46726 34813 46735
rect 34739 46670 34748 46726
rect 34804 46670 34813 46726
rect 34739 46661 34813 46670
rect 7276 45592 7350 45601
rect 7276 45536 7285 45592
rect 7341 45536 7350 45592
rect 7276 45527 7350 45536
rect 11220 45592 11294 45601
rect 11220 45536 11229 45592
rect 11285 45536 11294 45592
rect 11220 45527 11294 45536
rect 15164 45592 15238 45601
rect 15164 45536 15173 45592
rect 15229 45536 15238 45592
rect 15164 45527 15238 45536
rect 19108 45592 19182 45601
rect 19108 45536 19117 45592
rect 19173 45536 19182 45592
rect 19108 45527 19182 45536
rect 23052 45592 23126 45601
rect 23052 45536 23061 45592
rect 23117 45536 23126 45592
rect 23052 45527 23126 45536
rect 26996 45592 27070 45601
rect 26996 45536 27005 45592
rect 27061 45536 27070 45592
rect 26996 45527 27070 45536
rect 30940 45592 31014 45601
rect 30940 45536 30949 45592
rect 31005 45536 31014 45592
rect 30940 45527 31014 45536
rect 34884 45592 34958 45601
rect 34884 45536 34893 45592
rect 34949 45536 34958 45592
rect 34884 45527 34958 45536
rect 357 44944 431 44953
rect 357 44888 366 44944
rect 422 44888 431 44944
rect 357 44879 431 44888
rect 2789 44944 2863 44953
rect 2789 44888 2798 44944
rect 2854 44888 2863 44944
rect 2789 44879 2863 44888
rect 5221 44944 5295 44953
rect 5221 44888 5230 44944
rect 5286 44888 5295 44944
rect 5221 44879 5295 44888
rect 7421 44944 7495 44953
rect 7421 44888 7430 44944
rect 7486 44888 7495 44944
rect 7421 44879 7495 44888
rect 7653 44944 7727 44953
rect 7653 44888 7662 44944
rect 7718 44888 7727 44944
rect 7653 44879 7727 44888
rect 10085 44944 10159 44953
rect 10085 44888 10094 44944
rect 10150 44888 10159 44944
rect 10085 44879 10159 44888
rect 11365 44944 11439 44953
rect 11365 44888 11374 44944
rect 11430 44888 11439 44944
rect 11365 44879 11439 44888
rect 12517 44944 12591 44953
rect 12517 44888 12526 44944
rect 12582 44888 12591 44944
rect 12517 44879 12591 44888
rect 14949 44944 15023 44953
rect 14949 44888 14958 44944
rect 15014 44888 15023 44944
rect 14949 44879 15023 44888
rect 15309 44944 15383 44953
rect 15309 44888 15318 44944
rect 15374 44888 15383 44944
rect 15309 44879 15383 44888
rect 17381 44944 17455 44953
rect 17381 44888 17390 44944
rect 17446 44888 17455 44944
rect 17381 44879 17455 44888
rect 19253 44944 19327 44953
rect 19253 44888 19262 44944
rect 19318 44888 19327 44944
rect 19253 44879 19327 44888
rect 19813 44944 19887 44953
rect 19813 44888 19822 44944
rect 19878 44888 19887 44944
rect 19813 44879 19887 44888
rect 22245 44944 22319 44953
rect 22245 44888 22254 44944
rect 22310 44888 22319 44944
rect 22245 44879 22319 44888
rect 23197 44944 23271 44953
rect 23197 44888 23206 44944
rect 23262 44888 23271 44944
rect 23197 44879 23271 44888
rect 24677 44944 24751 44953
rect 24677 44888 24686 44944
rect 24742 44888 24751 44944
rect 24677 44879 24751 44888
rect 27141 44944 27215 44953
rect 27141 44888 27150 44944
rect 27206 44888 27215 44944
rect 27141 44879 27215 44888
rect 29541 44944 29615 44953
rect 29541 44888 29550 44944
rect 29606 44888 29615 44944
rect 29541 44879 29615 44888
rect 31085 44944 31159 44953
rect 31085 44888 31094 44944
rect 31150 44888 31159 44944
rect 31085 44879 31159 44888
rect 31973 44944 32047 44953
rect 31973 44888 31982 44944
rect 32038 44888 32047 44944
rect 31973 44879 32047 44888
rect 34405 44944 34479 44953
rect 34405 44888 34414 44944
rect 34470 44888 34479 44944
rect 34405 44879 34479 44888
rect 35029 44944 35103 44953
rect 35029 44888 35038 44944
rect 35094 44888 35103 44944
rect 35029 44879 35103 44888
rect 36837 44944 36911 44953
rect 36837 44888 36846 44944
rect 36902 44888 36911 44944
rect 36837 44879 36911 44888
rect 39269 44944 39343 44953
rect 39269 44888 39278 44944
rect 39334 44888 39343 44944
rect 39269 44879 39343 44888
rect 41701 44944 41775 44953
rect 41701 44888 41710 44944
rect 41766 44888 41775 44944
rect 41701 44879 41775 44888
<< via2 >>
rect 7140 46724 7196 46726
rect 7140 46672 7142 46724
rect 7142 46672 7194 46724
rect 7194 46672 7196 46724
rect 7140 46670 7196 46672
rect 11084 46724 11140 46726
rect 11084 46672 11086 46724
rect 11086 46672 11138 46724
rect 11138 46672 11140 46724
rect 11084 46670 11140 46672
rect 15028 46724 15084 46726
rect 15028 46672 15030 46724
rect 15030 46672 15082 46724
rect 15082 46672 15084 46724
rect 15028 46670 15084 46672
rect 18972 46724 19028 46726
rect 18972 46672 18974 46724
rect 18974 46672 19026 46724
rect 19026 46672 19028 46724
rect 18972 46670 19028 46672
rect 22916 46724 22972 46726
rect 22916 46672 22918 46724
rect 22918 46672 22970 46724
rect 22970 46672 22972 46724
rect 22916 46670 22972 46672
rect 26860 46724 26916 46726
rect 26860 46672 26862 46724
rect 26862 46672 26914 46724
rect 26914 46672 26916 46724
rect 26860 46670 26916 46672
rect 30804 46724 30860 46726
rect 30804 46672 30806 46724
rect 30806 46672 30858 46724
rect 30858 46672 30860 46724
rect 30804 46670 30860 46672
rect 34748 46724 34804 46726
rect 34748 46672 34750 46724
rect 34750 46672 34802 46724
rect 34802 46672 34804 46724
rect 34748 46670 34804 46672
rect 7285 45590 7341 45592
rect 7285 45538 7287 45590
rect 7287 45538 7339 45590
rect 7339 45538 7341 45590
rect 7285 45536 7341 45538
rect 11229 45590 11285 45592
rect 11229 45538 11231 45590
rect 11231 45538 11283 45590
rect 11283 45538 11285 45590
rect 11229 45536 11285 45538
rect 15173 45590 15229 45592
rect 15173 45538 15175 45590
rect 15175 45538 15227 45590
rect 15227 45538 15229 45590
rect 15173 45536 15229 45538
rect 19117 45590 19173 45592
rect 19117 45538 19119 45590
rect 19119 45538 19171 45590
rect 19171 45538 19173 45590
rect 19117 45536 19173 45538
rect 23061 45590 23117 45592
rect 23061 45538 23063 45590
rect 23063 45538 23115 45590
rect 23115 45538 23117 45590
rect 23061 45536 23117 45538
rect 27005 45590 27061 45592
rect 27005 45538 27007 45590
rect 27007 45538 27059 45590
rect 27059 45538 27061 45590
rect 27005 45536 27061 45538
rect 30949 45590 31005 45592
rect 30949 45538 30951 45590
rect 30951 45538 31003 45590
rect 31003 45538 31005 45590
rect 30949 45536 31005 45538
rect 34893 45590 34949 45592
rect 34893 45538 34895 45590
rect 34895 45538 34947 45590
rect 34947 45538 34949 45590
rect 34893 45536 34949 45538
rect 366 44942 422 44944
rect 366 44890 368 44942
rect 368 44890 420 44942
rect 420 44890 422 44942
rect 366 44888 422 44890
rect 2798 44942 2854 44944
rect 2798 44890 2800 44942
rect 2800 44890 2852 44942
rect 2852 44890 2854 44942
rect 2798 44888 2854 44890
rect 5230 44942 5286 44944
rect 5230 44890 5232 44942
rect 5232 44890 5284 44942
rect 5284 44890 5286 44942
rect 5230 44888 5286 44890
rect 7430 44942 7486 44944
rect 7430 44890 7432 44942
rect 7432 44890 7484 44942
rect 7484 44890 7486 44942
rect 7430 44888 7486 44890
rect 7662 44942 7718 44944
rect 7662 44890 7664 44942
rect 7664 44890 7716 44942
rect 7716 44890 7718 44942
rect 7662 44888 7718 44890
rect 10094 44942 10150 44944
rect 10094 44890 10096 44942
rect 10096 44890 10148 44942
rect 10148 44890 10150 44942
rect 10094 44888 10150 44890
rect 11374 44942 11430 44944
rect 11374 44890 11376 44942
rect 11376 44890 11428 44942
rect 11428 44890 11430 44942
rect 11374 44888 11430 44890
rect 12526 44942 12582 44944
rect 12526 44890 12528 44942
rect 12528 44890 12580 44942
rect 12580 44890 12582 44942
rect 12526 44888 12582 44890
rect 14958 44942 15014 44944
rect 14958 44890 14960 44942
rect 14960 44890 15012 44942
rect 15012 44890 15014 44942
rect 14958 44888 15014 44890
rect 15318 44942 15374 44944
rect 15318 44890 15320 44942
rect 15320 44890 15372 44942
rect 15372 44890 15374 44942
rect 15318 44888 15374 44890
rect 17390 44942 17446 44944
rect 17390 44890 17392 44942
rect 17392 44890 17444 44942
rect 17444 44890 17446 44942
rect 17390 44888 17446 44890
rect 19262 44942 19318 44944
rect 19262 44890 19264 44942
rect 19264 44890 19316 44942
rect 19316 44890 19318 44942
rect 19262 44888 19318 44890
rect 19822 44942 19878 44944
rect 19822 44890 19824 44942
rect 19824 44890 19876 44942
rect 19876 44890 19878 44942
rect 19822 44888 19878 44890
rect 22254 44942 22310 44944
rect 22254 44890 22256 44942
rect 22256 44890 22308 44942
rect 22308 44890 22310 44942
rect 22254 44888 22310 44890
rect 23206 44942 23262 44944
rect 23206 44890 23208 44942
rect 23208 44890 23260 44942
rect 23260 44890 23262 44942
rect 23206 44888 23262 44890
rect 24686 44942 24742 44944
rect 24686 44890 24688 44942
rect 24688 44890 24740 44942
rect 24740 44890 24742 44942
rect 24686 44888 24742 44890
rect 27150 44942 27206 44944
rect 27150 44890 27152 44942
rect 27152 44890 27204 44942
rect 27204 44890 27206 44942
rect 27150 44888 27206 44890
rect 29550 44942 29606 44944
rect 29550 44890 29552 44942
rect 29552 44890 29604 44942
rect 29604 44890 29606 44942
rect 29550 44888 29606 44890
rect 31094 44942 31150 44944
rect 31094 44890 31096 44942
rect 31096 44890 31148 44942
rect 31148 44890 31150 44942
rect 31094 44888 31150 44890
rect 31982 44942 32038 44944
rect 31982 44890 31984 44942
rect 31984 44890 32036 44942
rect 32036 44890 32038 44942
rect 31982 44888 32038 44890
rect 34414 44942 34470 44944
rect 34414 44890 34416 44942
rect 34416 44890 34468 44942
rect 34468 44890 34470 44942
rect 34414 44888 34470 44890
rect 35038 44942 35094 44944
rect 35038 44890 35040 44942
rect 35040 44890 35092 44942
rect 35092 44890 35094 44942
rect 35038 44888 35094 44890
rect 36846 44942 36902 44944
rect 36846 44890 36848 44942
rect 36848 44890 36900 44942
rect 36900 44890 36902 44942
rect 36846 44888 36902 44890
rect 39278 44942 39334 44944
rect 39278 44890 39280 44942
rect 39280 44890 39332 44942
rect 39332 44890 39334 44942
rect 39278 44888 39334 44890
rect 41710 44942 41766 44944
rect 41710 44890 41712 44942
rect 41712 44890 41764 44942
rect 41764 44890 41766 44942
rect 41710 44888 41766 44890
<< metal3 >>
rect 7135 46726 7201 46731
rect 7135 46670 7140 46726
rect 7196 46670 7201 46726
rect 7135 46665 7201 46670
rect 11079 46726 11145 46731
rect 11079 46670 11084 46726
rect 11140 46670 11145 46726
rect 11079 46665 11145 46670
rect 15023 46726 15089 46731
rect 15023 46670 15028 46726
rect 15084 46670 15089 46726
rect 15023 46665 15089 46670
rect 18967 46726 19033 46731
rect 18967 46670 18972 46726
rect 19028 46670 19033 46726
rect 18967 46665 19033 46670
rect 22911 46726 22977 46731
rect 22911 46670 22916 46726
rect 22972 46670 22977 46726
rect 22911 46665 22977 46670
rect 26855 46726 26921 46731
rect 26855 46670 26860 46726
rect 26916 46670 26921 46726
rect 26855 46665 26921 46670
rect 30799 46726 30865 46731
rect 30799 46670 30804 46726
rect 30860 46670 30865 46726
rect 30799 46665 30865 46670
rect 34743 46726 34809 46731
rect 34743 46670 34748 46726
rect 34804 46670 34809 46726
rect 34743 46665 34809 46670
rect 7138 46094 7198 46665
rect 11082 46094 11142 46665
rect 15026 46094 15086 46665
rect 18970 46094 19030 46665
rect 22914 46094 22974 46665
rect 26858 46094 26918 46665
rect 30802 46094 30862 46665
rect 34746 46094 34806 46665
rect 7280 45592 7346 45597
rect 7280 45536 7285 45592
rect 7341 45536 7346 45592
rect 7280 45531 7346 45536
rect 361 44944 427 44949
rect 361 44888 366 44944
rect 422 44888 427 44944
rect 361 44883 427 44888
rect 2793 44944 2859 44949
rect 2793 44888 2798 44944
rect 2854 44888 2859 44944
rect 2793 44883 2859 44888
rect 5225 44944 5291 44949
rect 5225 44888 5230 44944
rect 5286 44888 5291 44944
rect 5225 44883 5291 44888
rect 364 43314 424 44883
rect 2796 43314 2856 44883
rect 5228 43314 5288 44883
rect 7283 44826 7343 45531
rect 7428 44949 7488 45737
rect 11224 45592 11290 45597
rect 11224 45536 11229 45592
rect 11285 45536 11290 45592
rect 11224 45531 11290 45536
rect 7425 44944 7491 44949
rect 7425 44888 7430 44944
rect 7486 44888 7491 44944
rect 7425 44883 7491 44888
rect 7657 44944 7723 44949
rect 7657 44888 7662 44944
rect 7718 44888 7723 44944
rect 7657 44883 7723 44888
rect 10089 44944 10155 44949
rect 10089 44888 10094 44944
rect 10150 44888 10155 44944
rect 10089 44883 10155 44888
rect 7275 44820 7351 44826
rect 7275 44756 7281 44820
rect 7345 44756 7351 44820
rect 7275 44750 7351 44756
rect 7660 43314 7720 44883
rect 10092 43314 10152 44883
rect 11227 44698 11287 45531
rect 11372 44949 11432 45737
rect 15168 45592 15234 45597
rect 15168 45536 15173 45592
rect 15229 45536 15234 45592
rect 15168 45531 15234 45536
rect 11369 44944 11435 44949
rect 11369 44888 11374 44944
rect 11430 44888 11435 44944
rect 11369 44883 11435 44888
rect 12521 44944 12587 44949
rect 12521 44888 12526 44944
rect 12582 44888 12587 44944
rect 12521 44883 12587 44888
rect 14953 44944 15019 44949
rect 14953 44888 14958 44944
rect 15014 44888 15019 44944
rect 14953 44883 15019 44888
rect 11219 44692 11295 44698
rect 11219 44628 11225 44692
rect 11289 44628 11295 44692
rect 11219 44622 11295 44628
rect 12524 43314 12584 44883
rect 14956 43314 15016 44883
rect 15171 44570 15231 45531
rect 15316 44949 15376 45737
rect 19112 45592 19178 45597
rect 19112 45536 19117 45592
rect 19173 45536 19178 45592
rect 19112 45531 19178 45536
rect 15313 44944 15379 44949
rect 15313 44888 15318 44944
rect 15374 44888 15379 44944
rect 15313 44883 15379 44888
rect 17385 44944 17451 44949
rect 17385 44888 17390 44944
rect 17446 44888 17451 44944
rect 17385 44883 17451 44888
rect 15163 44564 15239 44570
rect 15163 44500 15169 44564
rect 15233 44500 15239 44564
rect 15163 44494 15239 44500
rect 17388 43314 17448 44883
rect 19115 44442 19175 45531
rect 19260 44949 19320 45737
rect 23056 45592 23122 45597
rect 23056 45536 23061 45592
rect 23117 45536 23122 45592
rect 23056 45531 23122 45536
rect 19257 44944 19323 44949
rect 19257 44888 19262 44944
rect 19318 44888 19323 44944
rect 19257 44883 19323 44888
rect 19817 44944 19883 44949
rect 19817 44888 19822 44944
rect 19878 44888 19883 44944
rect 19817 44883 19883 44888
rect 22249 44944 22315 44949
rect 22249 44888 22254 44944
rect 22310 44888 22315 44944
rect 22249 44883 22315 44888
rect 19107 44436 19183 44442
rect 19107 44372 19113 44436
rect 19177 44372 19183 44436
rect 19107 44366 19183 44372
rect 19820 43314 19880 44883
rect 22252 43314 22312 44883
rect 23059 44314 23119 45531
rect 23204 44949 23264 45737
rect 27000 45592 27066 45597
rect 27000 45536 27005 45592
rect 27061 45536 27066 45592
rect 27000 45531 27066 45536
rect 23201 44944 23267 44949
rect 23201 44888 23206 44944
rect 23262 44888 23267 44944
rect 23201 44883 23267 44888
rect 24681 44944 24747 44949
rect 24681 44888 24686 44944
rect 24742 44888 24747 44944
rect 24681 44883 24747 44888
rect 23051 44308 23127 44314
rect 23051 44244 23057 44308
rect 23121 44244 23127 44308
rect 23051 44238 23127 44244
rect 24684 43314 24744 44883
rect 27003 44186 27063 45531
rect 27148 44949 27208 45737
rect 30944 45592 31010 45597
rect 30944 45536 30949 45592
rect 31005 45536 31010 45592
rect 30944 45531 31010 45536
rect 27145 44944 27211 44949
rect 27145 44888 27150 44944
rect 27206 44888 27211 44944
rect 27145 44883 27211 44888
rect 29545 44944 29611 44949
rect 29545 44888 29550 44944
rect 29606 44888 29611 44944
rect 29545 44883 29611 44888
rect 26995 44180 27071 44186
rect 26995 44116 27001 44180
rect 27065 44116 27071 44180
rect 26995 44110 27071 44116
rect 27148 43321 27208 44883
rect 355 43308 432 43314
rect 355 43244 361 43308
rect 426 43244 432 43308
rect 355 43238 432 43244
rect 2787 43308 2864 43314
rect 2787 43244 2793 43308
rect 2858 43244 2864 43308
rect 2787 43238 2864 43244
rect 5219 43308 5296 43314
rect 5219 43244 5225 43308
rect 5290 43244 5296 43308
rect 5219 43238 5296 43244
rect 7651 43308 7728 43314
rect 7651 43244 7657 43308
rect 7722 43244 7728 43308
rect 7651 43238 7728 43244
rect 10083 43308 10160 43314
rect 10083 43244 10089 43308
rect 10154 43244 10160 43308
rect 10083 43238 10160 43244
rect 12515 43308 12592 43314
rect 12515 43244 12521 43308
rect 12586 43244 12592 43308
rect 12515 43238 12592 43244
rect 14947 43308 15024 43314
rect 14947 43244 14953 43308
rect 15018 43244 15024 43308
rect 14947 43238 15024 43244
rect 17379 43308 17456 43314
rect 17379 43244 17385 43308
rect 17450 43244 17456 43308
rect 17379 43238 17456 43244
rect 19811 43308 19888 43314
rect 19811 43244 19817 43308
rect 19882 43244 19888 43308
rect 19811 43238 19888 43244
rect 22243 43308 22320 43314
rect 22243 43244 22249 43308
rect 22314 43244 22320 43308
rect 22243 43238 22320 43244
rect 24675 43308 24752 43314
rect 24675 43244 24681 43308
rect 24746 43244 24752 43308
rect 24675 43238 24752 43244
rect 27107 43308 27208 43321
rect 29548 43314 29608 44883
rect 30947 44058 31007 45531
rect 31092 44949 31152 45737
rect 34888 45592 34954 45597
rect 34888 45536 34893 45592
rect 34949 45536 34954 45592
rect 34888 45531 34954 45536
rect 31089 44944 31155 44949
rect 31089 44888 31094 44944
rect 31150 44888 31155 44944
rect 31089 44883 31155 44888
rect 31977 44944 32043 44949
rect 31977 44888 31982 44944
rect 32038 44888 32043 44944
rect 31977 44883 32043 44888
rect 34409 44944 34475 44949
rect 34409 44888 34414 44944
rect 34470 44888 34475 44944
rect 34409 44883 34475 44888
rect 30939 44052 31015 44058
rect 30939 43988 30945 44052
rect 31009 43988 31015 44052
rect 30939 43982 31015 43988
rect 31980 43314 32040 44883
rect 34412 43314 34472 44883
rect 34891 43930 34951 45531
rect 35036 44949 35096 45737
rect 35033 44944 35099 44949
rect 35033 44888 35038 44944
rect 35094 44888 35099 44944
rect 35033 44883 35099 44888
rect 36841 44944 36907 44949
rect 36841 44888 36846 44944
rect 36902 44888 36907 44944
rect 36841 44883 36907 44888
rect 39273 44944 39339 44949
rect 39273 44888 39278 44944
rect 39334 44888 39339 44944
rect 39273 44883 39339 44888
rect 41705 44944 41771 44949
rect 41705 44888 41710 44944
rect 41766 44888 41771 44944
rect 41705 44883 41771 44888
rect 34883 43924 34959 43930
rect 34883 43860 34889 43924
rect 34953 43860 34959 43924
rect 34883 43854 34959 43860
rect 36844 43314 36904 44883
rect 39276 43314 39336 44883
rect 41708 43314 41768 44883
rect 27107 43244 27113 43308
rect 27178 43244 27208 43308
rect 27107 43238 27208 43244
rect 29539 43308 29616 43314
rect 29539 43244 29545 43308
rect 29610 43244 29616 43308
rect 29539 43238 29616 43244
rect 31971 43308 32048 43314
rect 31971 43244 31977 43308
rect 32042 43244 32048 43308
rect 31971 43238 32048 43244
rect 34403 43308 34480 43314
rect 34403 43244 34409 43308
rect 34474 43244 34480 43308
rect 34403 43238 34480 43244
rect 36835 43308 36912 43314
rect 36835 43244 36841 43308
rect 36906 43244 36912 43308
rect 36835 43238 36912 43244
rect 39267 43308 39344 43314
rect 39267 43244 39273 43308
rect 39338 43244 39344 43308
rect 39267 43238 39344 43244
rect 41699 43308 41776 43314
rect 41699 43244 41705 43308
rect 41770 43244 41776 43308
rect 41699 43238 41776 43244
rect 364 42998 424 43238
rect 2796 42998 2856 43238
rect 5228 42998 5288 43238
rect 7660 42998 7720 43238
rect 10092 42998 10152 43238
rect 12524 42998 12584 43238
rect 14956 42998 15016 43238
rect 17388 42998 17448 43238
rect 19820 42998 19880 43238
rect 22252 42998 22312 43238
rect 24684 42998 24744 43238
rect 27116 42998 27176 43238
rect 29548 42998 29608 43238
rect 31980 42998 32040 43238
rect 34412 42998 34472 43238
rect 36844 42998 36904 43238
rect 39276 42998 39336 43238
rect 41708 42998 41768 43238
rect 1708 42673 1784 42679
rect 1708 42670 1714 42673
rect 1468 42610 1714 42670
rect 1708 42608 1714 42610
rect 1778 42608 1784 42673
rect 4140 42673 4216 42679
rect 4140 42670 4146 42673
rect 3900 42610 4146 42670
rect 1708 42602 1784 42608
rect 4140 42608 4146 42610
rect 4210 42608 4216 42673
rect 6572 42673 6648 42679
rect 6572 42670 6578 42673
rect 6332 42610 6578 42670
rect 4140 42602 4216 42608
rect 6572 42608 6578 42610
rect 6642 42608 6648 42673
rect 9004 42673 9080 42679
rect 9004 42670 9010 42673
rect 8764 42610 9010 42670
rect 6572 42602 6648 42608
rect 9004 42608 9010 42610
rect 9074 42608 9080 42673
rect 11436 42673 11512 42679
rect 11436 42670 11442 42673
rect 11196 42610 11442 42670
rect 9004 42602 9080 42608
rect 11436 42608 11442 42610
rect 11506 42608 11512 42673
rect 13868 42673 13944 42679
rect 13868 42670 13874 42673
rect 13628 42610 13874 42670
rect 11436 42602 11512 42608
rect 13868 42608 13874 42610
rect 13938 42608 13944 42673
rect 16300 42673 16376 42679
rect 16300 42670 16306 42673
rect 16060 42610 16306 42670
rect 13868 42602 13944 42608
rect 16300 42608 16306 42610
rect 16370 42608 16376 42673
rect 18732 42673 18808 42679
rect 18732 42670 18738 42673
rect 18492 42610 18738 42670
rect 16300 42602 16376 42608
rect 18732 42608 18738 42610
rect 18802 42608 18808 42673
rect 21164 42673 21240 42679
rect 21164 42670 21170 42673
rect 20924 42610 21170 42670
rect 18732 42602 18808 42608
rect 21164 42608 21170 42610
rect 21234 42608 21240 42673
rect 23596 42673 23672 42679
rect 23596 42670 23602 42673
rect 23356 42610 23602 42670
rect 21164 42602 21240 42608
rect 23596 42608 23602 42610
rect 23666 42608 23672 42673
rect 26028 42673 26104 42679
rect 26028 42670 26034 42673
rect 25788 42610 26034 42670
rect 23596 42602 23672 42608
rect 26028 42608 26034 42610
rect 26098 42608 26104 42673
rect 28460 42673 28536 42679
rect 28460 42670 28466 42673
rect 28220 42610 28466 42670
rect 26028 42602 26104 42608
rect 28460 42608 28466 42610
rect 28530 42608 28536 42673
rect 30892 42673 30968 42679
rect 30892 42670 30898 42673
rect 30652 42610 30898 42670
rect 28460 42602 28536 42608
rect 30892 42608 30898 42610
rect 30962 42608 30968 42673
rect 33324 42673 33400 42679
rect 33324 42670 33330 42673
rect 33084 42610 33330 42670
rect 30892 42602 30968 42608
rect 33324 42608 33330 42610
rect 33394 42608 33400 42673
rect 35756 42673 35832 42679
rect 35756 42670 35762 42673
rect 35516 42610 35762 42670
rect 33324 42602 33400 42608
rect 35756 42608 35762 42610
rect 35826 42608 35832 42673
rect 38188 42673 38264 42679
rect 38188 42670 38194 42673
rect 37948 42610 38194 42670
rect 35756 42602 35832 42608
rect 38188 42608 38194 42610
rect 38258 42608 38264 42673
rect 40620 42673 40696 42679
rect 40620 42670 40626 42673
rect 40380 42610 40626 42670
rect 38188 42602 38264 42608
rect 40620 42608 40626 42610
rect 40690 42608 40696 42673
rect 43052 42673 43128 42679
rect 43052 42670 43058 42673
rect 42812 42610 43058 42670
rect 40620 42602 40696 42608
rect 43052 42608 43058 42610
rect 43122 42608 43128 42673
rect 43052 42602 43128 42608
rect -280 41956 -204 41962
rect -280 41891 -274 41956
rect -210 41954 -204 41956
rect 2152 41956 2228 41962
rect -210 41894 36 41954
rect -210 41891 -204 41894
rect -280 41885 -204 41891
rect 2152 41891 2158 41956
rect 2222 41954 2228 41956
rect 4584 41956 4660 41962
rect 2222 41894 2468 41954
rect 2222 41891 2228 41894
rect 2152 41885 2228 41891
rect 4584 41891 4590 41956
rect 4654 41954 4660 41956
rect 7016 41956 7092 41962
rect 4654 41894 4900 41954
rect 4654 41891 4660 41894
rect 4584 41885 4660 41891
rect 7016 41891 7022 41956
rect 7086 41954 7092 41956
rect 9448 41956 9524 41962
rect 7086 41894 7332 41954
rect 7086 41891 7092 41894
rect 7016 41885 7092 41891
rect 9448 41891 9454 41956
rect 9518 41954 9524 41956
rect 11880 41956 11956 41962
rect 9518 41894 9764 41954
rect 9518 41891 9524 41894
rect 9448 41885 9524 41891
rect 11880 41891 11886 41956
rect 11950 41954 11956 41956
rect 14312 41956 14388 41962
rect 11950 41894 12196 41954
rect 11950 41891 11956 41894
rect 11880 41885 11956 41891
rect 14312 41891 14318 41956
rect 14382 41954 14388 41956
rect 16744 41956 16820 41962
rect 14382 41894 14628 41954
rect 14382 41891 14388 41894
rect 14312 41885 14388 41891
rect 16744 41891 16750 41956
rect 16814 41954 16820 41956
rect 19176 41956 19252 41962
rect 16814 41894 17060 41954
rect 16814 41891 16820 41894
rect 16744 41885 16820 41891
rect 19176 41891 19182 41956
rect 19246 41954 19252 41956
rect 21608 41956 21684 41962
rect 19246 41894 19492 41954
rect 19246 41891 19252 41894
rect 19176 41885 19252 41891
rect 21608 41891 21614 41956
rect 21678 41954 21684 41956
rect 24040 41956 24116 41962
rect 21678 41894 21924 41954
rect 21678 41891 21684 41894
rect 21608 41885 21684 41891
rect 24040 41891 24046 41956
rect 24110 41954 24116 41956
rect 26472 41956 26548 41962
rect 24110 41894 24356 41954
rect 24110 41891 24116 41894
rect 24040 41885 24116 41891
rect 26472 41891 26478 41956
rect 26542 41954 26548 41956
rect 28904 41956 28980 41962
rect 26542 41894 26788 41954
rect 26542 41891 26548 41894
rect 26472 41885 26548 41891
rect 28904 41891 28910 41956
rect 28974 41954 28980 41956
rect 31336 41956 31412 41962
rect 28974 41894 29220 41954
rect 28974 41891 28980 41894
rect 28904 41885 28980 41891
rect 31336 41891 31342 41956
rect 31406 41954 31412 41956
rect 33768 41956 33844 41962
rect 31406 41894 31652 41954
rect 31406 41891 31412 41894
rect 31336 41885 31412 41891
rect 33768 41891 33774 41956
rect 33838 41954 33844 41956
rect 36200 41956 36276 41962
rect 33838 41894 34084 41954
rect 33838 41891 33844 41894
rect 33768 41885 33844 41891
rect 36200 41891 36206 41956
rect 36270 41954 36276 41956
rect 38632 41956 38708 41962
rect 36270 41894 36516 41954
rect 36270 41891 36276 41894
rect 36200 41885 36276 41891
rect 38632 41891 38638 41956
rect 38702 41954 38708 41956
rect 41064 41956 41140 41962
rect 38702 41894 38948 41954
rect 38702 41891 38708 41894
rect 38632 41885 38708 41891
rect 41064 41891 41070 41956
rect 41134 41954 41140 41956
rect 41134 41894 41380 41954
rect 41134 41891 41140 41894
rect 41064 41885 41140 41891
rect 1080 41326 1140 41566
rect 3512 41326 3572 41566
rect 5944 41326 6004 41566
rect 8376 41326 8436 41566
rect 10808 41326 10868 41566
rect 13240 41326 13300 41566
rect 15672 41326 15732 41566
rect 18104 41326 18164 41566
rect 20536 41326 20596 41566
rect 22968 41326 23028 41566
rect 25400 41326 25460 41566
rect 27832 41326 27892 41566
rect 30264 41326 30324 41566
rect 32696 41326 32756 41566
rect 35128 41326 35188 41566
rect 37560 41326 37620 41566
rect 39992 41326 40052 41566
rect 42424 41326 42484 41566
rect 1072 41320 1149 41326
rect 1072 41256 1078 41320
rect 1143 41256 1149 41320
rect 1072 41250 1149 41256
rect 3504 41320 3581 41326
rect 3504 41256 3510 41320
rect 3575 41256 3581 41320
rect 3504 41250 3581 41256
rect 5936 41320 6013 41326
rect 5936 41256 5942 41320
rect 6007 41256 6013 41320
rect 5936 41250 6013 41256
rect 8368 41320 8445 41326
rect 8368 41256 8374 41320
rect 8439 41256 8445 41320
rect 8368 41250 8445 41256
rect 10800 41320 10877 41326
rect 10800 41256 10806 41320
rect 10871 41256 10877 41320
rect 10800 41250 10877 41256
rect 13232 41320 13309 41326
rect 13232 41256 13238 41320
rect 13303 41256 13309 41320
rect 13232 41250 13309 41256
rect 15664 41320 15741 41326
rect 15664 41256 15670 41320
rect 15735 41256 15741 41320
rect 15664 41250 15741 41256
rect 18096 41320 18173 41326
rect 18096 41256 18102 41320
rect 18167 41256 18173 41320
rect 18096 41250 18173 41256
rect 20528 41320 20605 41326
rect 20528 41256 20534 41320
rect 20599 41256 20605 41320
rect 20528 41250 20605 41256
rect 22960 41320 23037 41326
rect 22960 41256 22966 41320
rect 23031 41256 23037 41320
rect 22960 41250 23037 41256
rect 25392 41320 25469 41326
rect 25392 41256 25398 41320
rect 25463 41256 25469 41320
rect 25392 41250 25469 41256
rect 27824 41320 27901 41326
rect 27824 41256 27830 41320
rect 27895 41256 27901 41320
rect 27824 41250 27901 41256
rect 30256 41320 30333 41326
rect 30256 41256 30262 41320
rect 30327 41256 30333 41320
rect 30256 41250 30333 41256
rect 32688 41320 32765 41326
rect 32688 41256 32694 41320
rect 32759 41256 32765 41320
rect 32688 41250 32765 41256
rect 35120 41320 35197 41326
rect 35120 41256 35126 41320
rect 35191 41256 35197 41320
rect 35120 41250 35197 41256
rect 37552 41320 37629 41326
rect 37552 41256 37558 41320
rect 37623 41256 37629 41320
rect 37552 41250 37629 41256
rect 39984 41320 40061 41326
rect 39984 41256 39990 41320
rect 40055 41256 40061 41320
rect 39984 41250 40061 41256
rect 42416 41320 42493 41326
rect 42416 41256 42422 41320
rect 42487 41256 42493 41320
rect 42416 41250 42493 41256
rect -632 41005 -556 41011
rect -632 40941 -626 41005
rect -562 41003 -556 41005
rect -562 40943 40380 41003
rect -562 40941 -556 40943
rect -632 40935 -556 40941
rect 355 40876 432 40882
rect 355 40812 361 40876
rect 426 40812 432 40876
rect 355 40806 432 40812
rect 364 40566 424 40806
rect 2796 40566 2856 40943
rect 5228 40566 5288 40602
rect 7660 40566 7720 40943
rect 10092 40566 10152 40602
rect 12524 40566 12584 40943
rect 14956 40566 15016 40602
rect 17388 40566 17448 40943
rect 19820 40566 19880 40602
rect 22252 40566 22312 40943
rect 24684 40566 24744 40602
rect 27116 40566 27176 40943
rect 29548 40566 29608 40602
rect 31980 40566 32040 40943
rect 34412 40566 34472 40602
rect 36844 40566 36904 40943
rect 41699 40876 41776 40882
rect 41699 40812 41705 40876
rect 41770 40812 41776 40876
rect 41699 40806 41776 40812
rect 39276 40566 39336 40602
rect 41708 40566 41768 40806
rect 1708 40241 1784 40247
rect 1708 40238 1714 40241
rect 1468 40178 1714 40238
rect 1708 40176 1714 40178
rect 1778 40176 1784 40241
rect 43052 40241 43128 40247
rect 43052 40238 43058 40241
rect 42812 40178 43058 40238
rect 1708 40170 1784 40176
rect 43052 40176 43058 40178
rect 43122 40176 43128 40241
rect 43052 40170 43128 40176
rect -280 39524 -204 39530
rect -280 39459 -274 39524
rect -210 39522 -204 39524
rect 41064 39524 41140 39530
rect -210 39462 36 39522
rect -210 39459 -204 39462
rect -280 39453 -204 39459
rect 41064 39459 41070 39524
rect 41134 39522 41140 39524
rect 41134 39462 41380 39522
rect 41134 39459 41140 39462
rect 41064 39453 41140 39459
rect 1080 38894 1140 39134
rect 3512 39098 3572 39134
rect 1072 38888 1149 38894
rect 1072 38824 1078 38888
rect 1143 38824 1149 38888
rect 1072 38818 1149 38824
rect 2788 38759 2864 38765
rect 2788 38757 2794 38759
rect 2468 38697 2794 38757
rect 2788 38695 2794 38697
rect 2858 38757 2864 38759
rect 5944 38757 6004 39134
rect 8376 39098 8436 39134
rect 7652 38759 7728 38765
rect 7652 38757 7658 38759
rect 2858 38697 7658 38757
rect 2858 38695 2864 38697
rect 2788 38689 2864 38695
rect 7652 38695 7658 38697
rect 7722 38757 7728 38759
rect 10808 38757 10868 39134
rect 13240 39098 13300 39134
rect 12516 38759 12592 38765
rect 12516 38757 12522 38759
rect 7722 38697 12522 38757
rect 7722 38695 7728 38697
rect 7652 38689 7728 38695
rect 12516 38695 12522 38697
rect 12586 38757 12592 38759
rect 15672 38757 15732 39134
rect 18104 39098 18164 39134
rect 17380 38759 17456 38765
rect 17380 38757 17386 38759
rect 12586 38697 17386 38757
rect 12586 38695 12592 38697
rect 12516 38689 12592 38695
rect 17380 38695 17386 38697
rect 17450 38757 17456 38759
rect 20536 38757 20596 39134
rect 22968 39098 23028 39134
rect 22244 38759 22320 38765
rect 22244 38757 22250 38759
rect 17450 38697 22250 38757
rect 17450 38695 17456 38697
rect 17380 38689 17456 38695
rect 22244 38695 22250 38697
rect 22314 38757 22320 38759
rect 25400 38757 25460 39134
rect 27832 39098 27892 39134
rect 27108 38759 27184 38765
rect 27108 38757 27114 38759
rect 22314 38697 27114 38757
rect 22314 38695 22320 38697
rect 22244 38689 22320 38695
rect 27108 38695 27114 38697
rect 27178 38757 27184 38759
rect 30264 38757 30324 39134
rect 32696 39098 32756 39134
rect 31972 38759 32048 38765
rect 31972 38757 31978 38759
rect 27178 38697 31978 38757
rect 27178 38695 27184 38697
rect 27108 38689 27184 38695
rect 31972 38695 31978 38697
rect 32042 38757 32048 38759
rect 35128 38757 35188 39134
rect 37560 39098 37620 39134
rect 36836 38759 36912 38765
rect 36836 38757 36842 38759
rect 32042 38697 36842 38757
rect 32042 38695 32048 38697
rect 31972 38689 32048 38695
rect 36836 38695 36842 38697
rect 36906 38757 36912 38759
rect 39992 38757 40052 39134
rect 42424 38894 42484 39134
rect 42416 38888 42493 38894
rect 42416 38824 42422 38888
rect 42487 38824 42493 38888
rect 42416 38818 42493 38824
rect 43404 38759 43480 38765
rect 43404 38757 43410 38759
rect 36906 38697 43410 38757
rect 36906 38695 36912 38697
rect 36836 38689 36912 38695
rect 43404 38695 43410 38697
rect 43474 38695 43480 38759
rect 43404 38689 43480 38695
rect 2468 38511 40380 38571
rect 355 38444 432 38450
rect 355 38380 361 38444
rect 426 38380 432 38444
rect 355 38374 432 38380
rect 2788 38444 2864 38450
rect 2788 38380 2794 38444
rect 2858 38380 2864 38444
rect 2788 38374 2864 38380
rect 7652 38444 7728 38450
rect 7652 38380 7658 38444
rect 7722 38380 7728 38444
rect 7652 38374 7728 38380
rect 12516 38444 12592 38450
rect 12516 38380 12522 38444
rect 12586 38380 12592 38444
rect 12516 38374 12592 38380
rect 17380 38444 17456 38450
rect 17380 38380 17386 38444
rect 17450 38380 17456 38444
rect 17380 38374 17456 38380
rect 22244 38444 22320 38450
rect 22244 38380 22250 38444
rect 22314 38380 22320 38444
rect 22244 38374 22320 38380
rect 27108 38444 27184 38450
rect 27108 38380 27114 38444
rect 27178 38380 27184 38444
rect 27108 38374 27184 38380
rect 31972 38444 32048 38450
rect 31972 38380 31978 38444
rect 32042 38380 32048 38444
rect 31972 38374 32048 38380
rect 36836 38444 36912 38450
rect 36836 38380 36842 38444
rect 36906 38380 36912 38444
rect 36836 38374 36912 38380
rect 41699 38444 41776 38450
rect 41699 38380 41705 38444
rect 41770 38380 41776 38444
rect 41699 38374 41776 38380
rect 364 38134 424 38374
rect 2796 38134 2856 38374
rect 5228 38134 5288 38170
rect 7660 38134 7720 38374
rect 10092 38134 10152 38170
rect 12524 38134 12584 38374
rect 14956 38134 15016 38170
rect 17388 38134 17448 38374
rect 19820 38134 19880 38170
rect 22252 38134 22312 38374
rect 24684 38134 24744 38170
rect 27116 38134 27176 38374
rect 29548 38134 29608 38170
rect 31980 38134 32040 38374
rect 34412 38134 34472 38170
rect 36844 38134 36904 38374
rect 39276 38134 39336 38170
rect 41708 38134 41768 38374
rect 1708 37809 1784 37815
rect 1708 37806 1714 37809
rect 1468 37746 1714 37806
rect 1708 37744 1714 37746
rect 1778 37744 1784 37809
rect 43052 37809 43128 37815
rect 43052 37806 43058 37809
rect 42812 37746 43058 37806
rect 1708 37738 1784 37744
rect 43052 37744 43058 37746
rect 43122 37744 43128 37809
rect 43052 37738 43128 37744
rect -280 37092 -204 37098
rect -280 37027 -274 37092
rect -210 37090 -204 37092
rect 41064 37092 41140 37098
rect -210 37030 36 37090
rect -210 37027 -204 37030
rect -280 37021 -204 37027
rect 41064 37027 41070 37092
rect 41134 37090 41140 37092
rect 41134 37030 41380 37090
rect 41134 37027 41140 37030
rect 41064 37021 41140 37027
rect 1080 36462 1140 36702
rect 3512 36666 3572 36702
rect 1072 36456 1149 36462
rect 1072 36392 1078 36456
rect 1143 36392 1149 36456
rect 1072 36386 1149 36392
rect 5944 36325 6004 36702
rect 8376 36666 8436 36702
rect 10808 36325 10868 36702
rect 13240 36666 13300 36702
rect 15672 36325 15732 36702
rect 18104 36666 18164 36702
rect 20536 36325 20596 36702
rect 22968 36666 23028 36702
rect 25400 36325 25460 36702
rect 27832 36666 27892 36702
rect 30264 36325 30324 36702
rect 32696 36666 32756 36702
rect 35128 36325 35188 36702
rect 37560 36666 37620 36702
rect 39992 36325 40052 36702
rect 42424 36462 42484 36702
rect 42416 36456 42493 36462
rect 42416 36392 42422 36456
rect 42487 36392 42493 36456
rect 42416 36386 42493 36392
rect 43528 36327 43604 36333
rect 43528 36325 43534 36327
rect 2468 36265 43534 36325
rect 43528 36263 43534 36265
rect 43598 36263 43604 36327
rect 43528 36257 43604 36263
rect -632 36141 -556 36147
rect -632 36077 -626 36141
rect -562 36139 -556 36141
rect -562 36079 40380 36139
rect -562 36077 -556 36079
rect -632 36071 -556 36077
rect 355 36012 432 36018
rect 355 35948 361 36012
rect 426 35948 432 36012
rect 355 35942 432 35948
rect 364 35702 424 35942
rect 2796 35702 2856 36079
rect 5228 35702 5288 35738
rect 7660 35702 7720 36079
rect 10092 35702 10152 35738
rect 12524 35702 12584 36079
rect 14956 35702 15016 35738
rect 17388 35702 17448 36079
rect 19820 35702 19880 35738
rect 22252 35702 22312 36079
rect 24684 35702 24744 35738
rect 27116 35702 27176 36079
rect 29548 35702 29608 35738
rect 31980 35702 32040 36079
rect 34412 35702 34472 35738
rect 36844 35702 36904 36079
rect 41699 36012 41776 36018
rect 41699 35948 41705 36012
rect 41770 35948 41776 36012
rect 41699 35942 41776 35948
rect 39276 35702 39336 35738
rect 41708 35702 41768 35942
rect 1708 35377 1784 35383
rect 1708 35374 1714 35377
rect 1468 35314 1714 35374
rect 1708 35312 1714 35314
rect 1778 35312 1784 35377
rect 43052 35377 43128 35383
rect 43052 35374 43058 35377
rect 42812 35314 43058 35374
rect 1708 35306 1784 35312
rect 43052 35312 43058 35314
rect 43122 35312 43128 35377
rect 43052 35306 43128 35312
rect -280 34660 -204 34666
rect -280 34595 -274 34660
rect -210 34658 -204 34660
rect 41064 34660 41140 34666
rect -210 34598 36 34658
rect -210 34595 -204 34598
rect -280 34589 -204 34595
rect 41064 34595 41070 34660
rect 41134 34658 41140 34660
rect 41134 34598 41380 34658
rect 41134 34595 41140 34598
rect 41064 34589 41140 34595
rect 1080 34030 1140 34270
rect 3512 34234 3572 34270
rect 1072 34024 1149 34030
rect 1072 33960 1078 34024
rect 1143 33960 1149 34024
rect 1072 33954 1149 33960
rect 2788 33895 2864 33901
rect 2788 33893 2794 33895
rect 2468 33833 2794 33893
rect 2788 33831 2794 33833
rect 2858 33893 2864 33895
rect 5944 33893 6004 34270
rect 8376 34234 8436 34270
rect 7652 33895 7728 33901
rect 7652 33893 7658 33895
rect 2858 33833 7658 33893
rect 2858 33831 2864 33833
rect 2788 33825 2864 33831
rect 7652 33831 7658 33833
rect 7722 33893 7728 33895
rect 10808 33893 10868 34270
rect 13240 34234 13300 34270
rect 12516 33895 12592 33901
rect 12516 33893 12522 33895
rect 7722 33833 12522 33893
rect 7722 33831 7728 33833
rect 7652 33825 7728 33831
rect 12516 33831 12522 33833
rect 12586 33893 12592 33895
rect 15672 33893 15732 34270
rect 18104 34234 18164 34270
rect 17380 33895 17456 33901
rect 17380 33893 17386 33895
rect 12586 33833 17386 33893
rect 12586 33831 12592 33833
rect 12516 33825 12592 33831
rect 17380 33831 17386 33833
rect 17450 33893 17456 33895
rect 20536 33893 20596 34270
rect 22968 34234 23028 34270
rect 22244 33895 22320 33901
rect 22244 33893 22250 33895
rect 17450 33833 22250 33893
rect 17450 33831 17456 33833
rect 17380 33825 17456 33831
rect 22244 33831 22250 33833
rect 22314 33893 22320 33895
rect 25400 33893 25460 34270
rect 27832 34234 27892 34270
rect 27108 33895 27184 33901
rect 27108 33893 27114 33895
rect 22314 33833 27114 33893
rect 22314 33831 22320 33833
rect 22244 33825 22320 33831
rect 27108 33831 27114 33833
rect 27178 33893 27184 33895
rect 30264 33893 30324 34270
rect 32696 34234 32756 34270
rect 31972 33895 32048 33901
rect 31972 33893 31978 33895
rect 27178 33833 31978 33893
rect 27178 33831 27184 33833
rect 27108 33825 27184 33831
rect 31972 33831 31978 33833
rect 32042 33893 32048 33895
rect 35128 33893 35188 34270
rect 37560 34234 37620 34270
rect 36836 33895 36912 33901
rect 36836 33893 36842 33895
rect 32042 33833 36842 33893
rect 32042 33831 32048 33833
rect 31972 33825 32048 33831
rect 36836 33831 36842 33833
rect 36906 33893 36912 33895
rect 39992 33893 40052 34270
rect 42424 34030 42484 34270
rect 42416 34024 42493 34030
rect 42416 33960 42422 34024
rect 42487 33960 42493 34024
rect 42416 33954 42493 33960
rect 43404 33895 43480 33901
rect 43404 33893 43410 33895
rect 36906 33833 43410 33893
rect 36906 33831 36912 33833
rect 36836 33825 36912 33831
rect 43404 33831 43410 33833
rect 43474 33831 43480 33895
rect 43404 33825 43480 33831
rect 2468 33647 40380 33707
rect 355 33580 432 33586
rect 355 33516 361 33580
rect 426 33516 432 33580
rect 355 33510 432 33516
rect 2788 33580 2864 33586
rect 2788 33516 2794 33580
rect 2858 33516 2864 33580
rect 2788 33510 2864 33516
rect 7652 33580 7728 33586
rect 7652 33516 7658 33580
rect 7722 33516 7728 33580
rect 7652 33510 7728 33516
rect 12516 33580 12592 33586
rect 12516 33516 12522 33580
rect 12586 33516 12592 33580
rect 12516 33510 12592 33516
rect 17380 33580 17456 33586
rect 17380 33516 17386 33580
rect 17450 33516 17456 33580
rect 17380 33510 17456 33516
rect 22244 33580 22320 33586
rect 22244 33516 22250 33580
rect 22314 33516 22320 33580
rect 22244 33510 22320 33516
rect 27108 33580 27184 33586
rect 27108 33516 27114 33580
rect 27178 33516 27184 33580
rect 27108 33510 27184 33516
rect 31972 33580 32048 33586
rect 31972 33516 31978 33580
rect 32042 33516 32048 33580
rect 31972 33510 32048 33516
rect 36836 33580 36912 33586
rect 36836 33516 36842 33580
rect 36906 33516 36912 33580
rect 36836 33510 36912 33516
rect 41699 33580 41776 33586
rect 41699 33516 41705 33580
rect 41770 33516 41776 33580
rect 41699 33510 41776 33516
rect 364 33270 424 33510
rect 2796 33270 2856 33510
rect 5228 33270 5288 33306
rect 7660 33270 7720 33510
rect 10092 33270 10152 33306
rect 12524 33270 12584 33510
rect 14956 33270 15016 33306
rect 17388 33270 17448 33510
rect 19820 33270 19880 33306
rect 22252 33270 22312 33510
rect 24684 33270 24744 33306
rect 27116 33270 27176 33510
rect 29548 33270 29608 33306
rect 31980 33270 32040 33510
rect 34412 33270 34472 33306
rect 36844 33270 36904 33510
rect 39276 33270 39336 33306
rect 41708 33270 41768 33510
rect 1708 32945 1784 32951
rect 1708 32942 1714 32945
rect 1468 32882 1714 32942
rect 1708 32880 1714 32882
rect 1778 32880 1784 32945
rect 43052 32945 43128 32951
rect 43052 32942 43058 32945
rect 42812 32882 43058 32942
rect 1708 32874 1784 32880
rect 43052 32880 43058 32882
rect 43122 32880 43128 32945
rect 43052 32874 43128 32880
rect -280 32228 -204 32234
rect -280 32163 -274 32228
rect -210 32226 -204 32228
rect 41064 32228 41140 32234
rect -210 32166 36 32226
rect -210 32163 -204 32166
rect -280 32157 -204 32163
rect 41064 32163 41070 32228
rect 41134 32226 41140 32228
rect 41134 32166 41380 32226
rect 41134 32163 41140 32166
rect 41064 32157 41140 32163
rect 1080 31598 1140 31838
rect 3512 31802 3572 31838
rect 1072 31592 1149 31598
rect 1072 31528 1078 31592
rect 1143 31528 1149 31592
rect 1072 31522 1149 31528
rect 5944 31461 6004 31838
rect 8376 31802 8436 31838
rect 10808 31461 10868 31838
rect 13240 31802 13300 31838
rect 15672 31461 15732 31838
rect 18104 31802 18164 31838
rect 20536 31461 20596 31838
rect 22968 31802 23028 31838
rect 25400 31461 25460 31838
rect 27832 31802 27892 31838
rect 30264 31461 30324 31838
rect 32696 31802 32756 31838
rect 35128 31461 35188 31838
rect 37560 31802 37620 31838
rect 39992 31461 40052 31838
rect 42424 31598 42484 31838
rect 42416 31592 42493 31598
rect 42416 31528 42422 31592
rect 42487 31528 42493 31592
rect 42416 31522 42493 31528
rect 43528 31463 43604 31469
rect 43528 31461 43534 31463
rect 2468 31401 43534 31461
rect 43528 31399 43534 31401
rect 43598 31399 43604 31463
rect 43528 31393 43604 31399
rect -632 31277 -556 31283
rect -632 31213 -626 31277
rect -562 31275 -556 31277
rect -562 31215 40380 31275
rect -562 31213 -556 31215
rect -632 31207 -556 31213
rect 355 31148 432 31154
rect 355 31084 361 31148
rect 426 31084 432 31148
rect 355 31078 432 31084
rect 364 30838 424 31078
rect 2796 30838 2856 31215
rect 5228 30838 5288 30874
rect 7660 30838 7720 31215
rect 10092 30838 10152 30874
rect 12524 30838 12584 31215
rect 14956 30838 15016 30874
rect 17388 30838 17448 31215
rect 19820 30838 19880 30874
rect 22252 30838 22312 31215
rect 24684 30838 24744 30874
rect 27116 30838 27176 31215
rect 29548 30838 29608 30874
rect 31980 30838 32040 31215
rect 34412 30838 34472 30874
rect 36844 30838 36904 31215
rect 41699 31148 41776 31154
rect 41699 31084 41705 31148
rect 41770 31084 41776 31148
rect 41699 31078 41776 31084
rect 39276 30838 39336 30874
rect 41708 30838 41768 31078
rect 1708 30513 1784 30519
rect 1708 30510 1714 30513
rect 1468 30450 1714 30510
rect 1708 30448 1714 30450
rect 1778 30448 1784 30513
rect 43052 30513 43128 30519
rect 43052 30510 43058 30513
rect 42812 30450 43058 30510
rect 1708 30442 1784 30448
rect 43052 30448 43058 30450
rect 43122 30448 43128 30513
rect 43052 30442 43128 30448
rect -280 29796 -204 29802
rect -280 29731 -274 29796
rect -210 29794 -204 29796
rect 41064 29796 41140 29802
rect -210 29734 36 29794
rect -210 29731 -204 29734
rect -280 29725 -204 29731
rect 41064 29731 41070 29796
rect 41134 29794 41140 29796
rect 41134 29734 41380 29794
rect 41134 29731 41140 29734
rect 41064 29725 41140 29731
rect 1080 29166 1140 29406
rect 3512 29370 3572 29406
rect 1072 29160 1149 29166
rect 1072 29096 1078 29160
rect 1143 29096 1149 29160
rect 1072 29090 1149 29096
rect 2788 29031 2864 29037
rect 2788 29029 2794 29031
rect 2468 28969 2794 29029
rect 2788 28967 2794 28969
rect 2858 29029 2864 29031
rect 5944 29029 6004 29406
rect 8376 29370 8436 29406
rect 7652 29031 7728 29037
rect 7652 29029 7658 29031
rect 2858 28969 7658 29029
rect 2858 28967 2864 28969
rect 2788 28961 2864 28967
rect 7652 28967 7658 28969
rect 7722 29029 7728 29031
rect 10808 29029 10868 29406
rect 13240 29370 13300 29406
rect 12516 29031 12592 29037
rect 12516 29029 12522 29031
rect 7722 28969 12522 29029
rect 7722 28967 7728 28969
rect 7652 28961 7728 28967
rect 12516 28967 12522 28969
rect 12586 29029 12592 29031
rect 15672 29029 15732 29406
rect 18104 29370 18164 29406
rect 17380 29031 17456 29037
rect 17380 29029 17386 29031
rect 12586 28969 17386 29029
rect 12586 28967 12592 28969
rect 12516 28961 12592 28967
rect 17380 28967 17386 28969
rect 17450 29029 17456 29031
rect 20536 29029 20596 29406
rect 22968 29370 23028 29406
rect 22244 29031 22320 29037
rect 22244 29029 22250 29031
rect 17450 28969 22250 29029
rect 17450 28967 17456 28969
rect 17380 28961 17456 28967
rect 22244 28967 22250 28969
rect 22314 29029 22320 29031
rect 25400 29029 25460 29406
rect 27832 29370 27892 29406
rect 27108 29031 27184 29037
rect 27108 29029 27114 29031
rect 22314 28969 27114 29029
rect 22314 28967 22320 28969
rect 22244 28961 22320 28967
rect 27108 28967 27114 28969
rect 27178 29029 27184 29031
rect 30264 29029 30324 29406
rect 32696 29370 32756 29406
rect 31972 29031 32048 29037
rect 31972 29029 31978 29031
rect 27178 28969 31978 29029
rect 27178 28967 27184 28969
rect 27108 28961 27184 28967
rect 31972 28967 31978 28969
rect 32042 29029 32048 29031
rect 35128 29029 35188 29406
rect 37560 29370 37620 29406
rect 36836 29031 36912 29037
rect 36836 29029 36842 29031
rect 32042 28969 36842 29029
rect 32042 28967 32048 28969
rect 31972 28961 32048 28967
rect 36836 28967 36842 28969
rect 36906 29029 36912 29031
rect 39992 29029 40052 29406
rect 42424 29166 42484 29406
rect 42416 29160 42493 29166
rect 42416 29096 42422 29160
rect 42487 29096 42493 29160
rect 42416 29090 42493 29096
rect 43404 29031 43480 29037
rect 43404 29029 43410 29031
rect 36906 28969 43410 29029
rect 36906 28967 36912 28969
rect 36836 28961 36912 28967
rect 43404 28967 43410 28969
rect 43474 28967 43480 29031
rect 43404 28961 43480 28967
rect 43652 28845 43728 28851
rect 43652 28843 43658 28845
rect 2468 28783 43658 28843
rect 355 28716 432 28722
rect 355 28652 361 28716
rect 426 28652 432 28716
rect 355 28646 432 28652
rect 2788 28716 2864 28722
rect 2788 28652 2794 28716
rect 2858 28652 2864 28716
rect 2788 28646 2864 28652
rect 7652 28716 7728 28722
rect 7652 28652 7658 28716
rect 7722 28652 7728 28716
rect 7652 28646 7728 28652
rect 364 28406 424 28646
rect 2796 28406 2856 28646
rect 5228 28406 5288 28442
rect 7660 28406 7720 28646
rect 10092 28406 10152 28783
rect 12516 28716 12592 28722
rect 12516 28652 12522 28716
rect 12586 28652 12592 28716
rect 12516 28646 12592 28652
rect 17380 28716 17456 28722
rect 17380 28652 17386 28716
rect 17450 28652 17456 28716
rect 17380 28646 17456 28652
rect 12524 28406 12584 28646
rect 14956 28406 15016 28442
rect 17388 28406 17448 28646
rect 19820 28406 19880 28783
rect 22244 28716 22320 28722
rect 22244 28652 22250 28716
rect 22314 28652 22320 28716
rect 22244 28646 22320 28652
rect 27108 28716 27184 28722
rect 27108 28652 27114 28716
rect 27178 28652 27184 28716
rect 27108 28646 27184 28652
rect 22252 28406 22312 28646
rect 24684 28406 24744 28442
rect 27116 28406 27176 28646
rect 29548 28406 29608 28783
rect 31972 28716 32048 28722
rect 31972 28652 31978 28716
rect 32042 28652 32048 28716
rect 31972 28646 32048 28652
rect 36836 28716 36912 28722
rect 36836 28652 36842 28716
rect 36906 28652 36912 28716
rect 36836 28646 36912 28652
rect 31980 28406 32040 28646
rect 34412 28406 34472 28442
rect 36844 28406 36904 28646
rect 39276 28406 39336 28783
rect 43652 28781 43658 28783
rect 43722 28781 43728 28845
rect 43652 28775 43728 28781
rect 41699 28716 41776 28722
rect 41699 28652 41705 28716
rect 41770 28652 41776 28716
rect 41699 28646 41776 28652
rect 41708 28406 41768 28646
rect 1708 28081 1784 28087
rect 1708 28078 1714 28081
rect 1468 28018 1714 28078
rect 1708 28016 1714 28018
rect 1778 28016 1784 28081
rect 43052 28081 43128 28087
rect 43052 28078 43058 28081
rect 42812 28018 43058 28078
rect 1708 28010 1784 28016
rect 43052 28016 43058 28018
rect 43122 28016 43128 28081
rect 43052 28010 43128 28016
rect -280 27364 -204 27370
rect -280 27299 -274 27364
rect -210 27362 -204 27364
rect 41064 27364 41140 27370
rect -210 27302 36 27362
rect -210 27299 -204 27302
rect -280 27293 -204 27299
rect 41064 27299 41070 27364
rect 41134 27362 41140 27364
rect 41134 27302 41380 27362
rect 41134 27299 41140 27302
rect 41064 27293 41140 27299
rect 1080 26734 1140 26974
rect 3512 26938 3572 26974
rect 1072 26728 1149 26734
rect 1072 26664 1078 26728
rect 1143 26664 1149 26728
rect 1072 26658 1149 26664
rect -756 26599 -680 26605
rect -756 26535 -750 26599
rect -686 26597 -680 26599
rect 5944 26597 6004 26974
rect 8376 26938 8436 26974
rect 13240 26938 13300 26974
rect 15672 26597 15732 26974
rect 18104 26938 18164 26974
rect 22968 26938 23028 26974
rect 25400 26597 25460 26974
rect 27832 26938 27892 26974
rect 32696 26938 32756 26974
rect 35128 26597 35188 26974
rect 37560 26938 37620 26974
rect 42424 26734 42484 26974
rect 42416 26728 42493 26734
rect 42416 26664 42422 26728
rect 42487 26664 42493 26728
rect 42416 26658 42493 26664
rect -686 26537 40380 26597
rect -686 26535 -680 26537
rect -756 26529 -680 26535
rect -632 26413 -556 26419
rect -632 26349 -626 26413
rect -562 26411 -556 26413
rect -562 26351 40380 26411
rect -562 26349 -556 26351
rect -632 26343 -556 26349
rect 355 26284 432 26290
rect 355 26220 361 26284
rect 426 26220 432 26284
rect 355 26214 432 26220
rect 364 25974 424 26214
rect 2796 25974 2856 26351
rect 5228 25974 5288 26010
rect 7660 25974 7720 26351
rect 10092 25974 10152 26010
rect 12524 25974 12584 26351
rect 14956 25974 15016 26010
rect 17388 25974 17448 26351
rect 19820 25974 19880 26010
rect 22252 25974 22312 26351
rect 24684 25974 24744 26010
rect 27116 25974 27176 26351
rect 29548 25974 29608 26010
rect 31980 25974 32040 26351
rect 34412 25974 34472 26010
rect 36844 25974 36904 26351
rect 41699 26284 41776 26290
rect 41699 26220 41705 26284
rect 41770 26220 41776 26284
rect 41699 26214 41776 26220
rect 39276 25974 39336 26010
rect 41708 25974 41768 26214
rect 1708 25649 1784 25655
rect 1708 25646 1714 25649
rect 1468 25586 1714 25646
rect 1708 25584 1714 25586
rect 1778 25584 1784 25649
rect 43052 25649 43128 25655
rect 43052 25646 43058 25649
rect 42812 25586 43058 25646
rect 1708 25578 1784 25584
rect 43052 25584 43058 25586
rect 43122 25584 43128 25649
rect 43052 25578 43128 25584
rect -280 24932 -204 24938
rect -280 24867 -274 24932
rect -210 24930 -204 24932
rect 41064 24932 41140 24938
rect -210 24870 36 24930
rect -210 24867 -204 24870
rect -280 24861 -204 24867
rect 41064 24867 41070 24932
rect 41134 24930 41140 24932
rect 41134 24870 41380 24930
rect 41134 24867 41140 24870
rect 41064 24861 41140 24867
rect 1080 24302 1140 24542
rect 3512 24506 3572 24542
rect 1072 24296 1149 24302
rect 1072 24232 1078 24296
rect 1143 24232 1149 24296
rect 1072 24226 1149 24232
rect 2788 24167 2864 24173
rect 2788 24165 2794 24167
rect 2468 24105 2794 24165
rect 2788 24103 2794 24105
rect 2858 24165 2864 24167
rect 5944 24165 6004 24542
rect 8376 24506 8436 24542
rect 7652 24167 7728 24173
rect 7652 24165 7658 24167
rect 2858 24105 7658 24165
rect 2858 24103 2864 24105
rect 2788 24097 2864 24103
rect 7652 24103 7658 24105
rect 7722 24165 7728 24167
rect 10808 24165 10868 24542
rect 13240 24506 13300 24542
rect 12516 24167 12592 24173
rect 12516 24165 12522 24167
rect 7722 24105 12522 24165
rect 7722 24103 7728 24105
rect 7652 24097 7728 24103
rect 12516 24103 12522 24105
rect 12586 24165 12592 24167
rect 15672 24165 15732 24542
rect 18104 24506 18164 24542
rect 17380 24167 17456 24173
rect 17380 24165 17386 24167
rect 12586 24105 17386 24165
rect 12586 24103 12592 24105
rect 12516 24097 12592 24103
rect 17380 24103 17386 24105
rect 17450 24165 17456 24167
rect 20536 24165 20596 24542
rect 22968 24506 23028 24542
rect 22244 24167 22320 24173
rect 22244 24165 22250 24167
rect 17450 24105 22250 24165
rect 17450 24103 17456 24105
rect 17380 24097 17456 24103
rect 22244 24103 22250 24105
rect 22314 24165 22320 24167
rect 25400 24165 25460 24542
rect 27832 24506 27892 24542
rect 27108 24167 27184 24173
rect 27108 24165 27114 24167
rect 22314 24105 27114 24165
rect 22314 24103 22320 24105
rect 22244 24097 22320 24103
rect 27108 24103 27114 24105
rect 27178 24165 27184 24167
rect 30264 24165 30324 24542
rect 32696 24506 32756 24542
rect 31972 24167 32048 24173
rect 31972 24165 31978 24167
rect 27178 24105 31978 24165
rect 27178 24103 27184 24105
rect 27108 24097 27184 24103
rect 31972 24103 31978 24105
rect 32042 24165 32048 24167
rect 35128 24165 35188 24542
rect 37560 24506 37620 24542
rect 36836 24167 36912 24173
rect 36836 24165 36842 24167
rect 32042 24105 36842 24165
rect 32042 24103 32048 24105
rect 31972 24097 32048 24103
rect 36836 24103 36842 24105
rect 36906 24165 36912 24167
rect 39992 24165 40052 24542
rect 42424 24302 42484 24542
rect 42416 24296 42493 24302
rect 42416 24232 42422 24296
rect 42487 24232 42493 24296
rect 42416 24226 42493 24232
rect 43404 24167 43480 24173
rect 43404 24165 43410 24167
rect 36906 24105 43410 24165
rect 36906 24103 36912 24105
rect 36836 24097 36912 24103
rect 43404 24103 43410 24105
rect 43474 24103 43480 24167
rect 43404 24097 43480 24103
rect -756 23981 -680 23987
rect -756 23917 -750 23981
rect -686 23979 -680 23981
rect -686 23919 40380 23979
rect -686 23917 -680 23919
rect -756 23911 -680 23917
rect 355 23852 432 23858
rect 355 23788 361 23852
rect 426 23788 432 23852
rect 355 23782 432 23788
rect 2788 23852 2864 23858
rect 2788 23788 2794 23852
rect 2858 23788 2864 23852
rect 2788 23782 2864 23788
rect 364 23542 424 23782
rect 2796 23542 2856 23782
rect 5228 23542 5288 23919
rect 7652 23852 7728 23858
rect 7652 23788 7658 23852
rect 7722 23788 7728 23852
rect 7652 23782 7728 23788
rect 12516 23852 12592 23858
rect 12516 23788 12522 23852
rect 12586 23788 12592 23852
rect 12516 23782 12592 23788
rect 7660 23542 7720 23782
rect 10092 23542 10152 23578
rect 12524 23542 12584 23782
rect 14956 23542 15016 23919
rect 17380 23852 17456 23858
rect 17380 23788 17386 23852
rect 17450 23788 17456 23852
rect 17380 23782 17456 23788
rect 22244 23852 22320 23858
rect 22244 23788 22250 23852
rect 22314 23788 22320 23852
rect 22244 23782 22320 23788
rect 17388 23542 17448 23782
rect 22252 23542 22312 23782
rect 24684 23542 24744 23919
rect 27108 23852 27184 23858
rect 27108 23788 27114 23852
rect 27178 23788 27184 23852
rect 27108 23782 27184 23788
rect 31972 23852 32048 23858
rect 31972 23788 31978 23852
rect 32042 23788 32048 23852
rect 31972 23782 32048 23788
rect 27116 23542 27176 23782
rect 29548 23542 29608 23578
rect 31980 23542 32040 23782
rect 34412 23542 34472 23919
rect 36836 23852 36912 23858
rect 36836 23788 36842 23852
rect 36906 23788 36912 23852
rect 36836 23782 36912 23788
rect 41699 23852 41776 23858
rect 41699 23788 41705 23852
rect 41770 23788 41776 23852
rect 41699 23782 41776 23788
rect 36844 23542 36904 23782
rect 39276 23542 39336 23578
rect 41708 23542 41768 23782
rect 1708 23217 1784 23223
rect 1708 23214 1714 23217
rect 1468 23154 1714 23214
rect 1708 23152 1714 23154
rect 1778 23152 1784 23217
rect 43052 23217 43128 23223
rect 43052 23214 43058 23217
rect 42812 23154 43058 23214
rect 1708 23146 1784 23152
rect 43052 23152 43058 23154
rect 43122 23152 43128 23217
rect 43052 23146 43128 23152
rect -280 22500 -204 22506
rect -280 22435 -274 22500
rect -210 22498 -204 22500
rect 41064 22500 41140 22506
rect -210 22438 36 22498
rect -210 22435 -204 22438
rect -280 22429 -204 22435
rect 41064 22435 41070 22500
rect 41134 22498 41140 22500
rect 41134 22438 41380 22498
rect 41134 22435 41140 22438
rect 41064 22429 41140 22435
rect 1080 21870 1140 22110
rect 10808 21870 10868 22074
rect 1072 21864 1149 21870
rect 1072 21800 1078 21864
rect 1143 21800 1149 21864
rect 1072 21794 1149 21800
rect 10800 21864 10876 21870
rect 10800 21799 10806 21864
rect 10870 21799 10876 21864
rect 10800 21793 10876 21799
rect 12516 21735 12592 21741
rect 12516 21733 12522 21735
rect 2468 21673 12522 21733
rect 12516 21671 12522 21673
rect 12586 21733 12592 21735
rect 30264 21733 30324 22074
rect 39992 21870 40052 22074
rect 42424 21870 42484 22110
rect 39984 21864 40060 21870
rect 39984 21799 39990 21864
rect 40054 21799 40060 21864
rect 39984 21793 40060 21799
rect 42416 21864 42493 21870
rect 42416 21800 42422 21864
rect 42487 21800 42493 21864
rect 42416 21794 42493 21800
rect 43776 21735 43852 21741
rect 43776 21733 43782 21735
rect 12586 21673 43782 21733
rect 12586 21671 12592 21673
rect 12516 21665 12592 21671
rect 43776 21671 43782 21673
rect 43846 21671 43852 21735
rect 43776 21665 43852 21671
rect -1004 21549 -928 21555
rect -1004 21485 -998 21549
rect -934 21547 -928 21549
rect 22244 21549 22320 21555
rect 22244 21547 22250 21549
rect -934 21487 22250 21547
rect -934 21485 -928 21487
rect -1004 21479 -928 21485
rect 22244 21485 22250 21487
rect 22314 21485 22320 21549
rect 22244 21479 22320 21485
rect -880 21363 -804 21369
rect -880 21299 -874 21363
rect -810 21361 -804 21363
rect 10800 21364 10876 21370
rect 10800 21361 10806 21364
rect -810 21301 10806 21361
rect -810 21299 -804 21301
rect -880 21293 -804 21299
rect 355 21234 432 21240
rect 355 21170 361 21234
rect 426 21170 432 21234
rect 355 21164 432 21170
rect 364 20924 424 21164
rect 2796 20960 2856 21301
rect 10800 21299 10806 21301
rect 10870 21361 10876 21364
rect 39984 21364 40060 21370
rect 39984 21361 39990 21364
rect 10870 21301 39990 21361
rect 10870 21299 10876 21301
rect 10800 21293 10876 21299
rect 12516 21234 12592 21240
rect 12516 21170 12522 21234
rect 12586 21170 12592 21234
rect 12516 21164 12592 21170
rect 22244 21234 22320 21240
rect 22244 21170 22250 21234
rect 22314 21170 22320 21234
rect 22244 21164 22320 21170
rect 12524 20924 12584 21164
rect 22252 20924 22312 21164
rect 31980 20960 32040 21301
rect 39984 21299 39990 21301
rect 40054 21361 40060 21364
rect 40054 21301 40380 21361
rect 40054 21299 40060 21301
rect 39984 21293 40060 21299
rect 41699 21234 41776 21240
rect 41699 21170 41705 21234
rect 41770 21170 41776 21234
rect 41699 21164 41776 21170
rect 41708 20924 41768 21164
rect 1708 20599 1784 20605
rect 1708 20596 1714 20599
rect 1468 20536 1714 20596
rect 1708 20534 1714 20536
rect 1778 20534 1784 20599
rect 43052 20599 43128 20605
rect 43052 20596 43058 20599
rect 42812 20536 43058 20596
rect 1708 20528 1784 20534
rect 43052 20534 43058 20536
rect 43122 20534 43128 20599
rect 43052 20528 43128 20534
rect -280 19882 -204 19888
rect -280 19817 -274 19882
rect -210 19880 -204 19882
rect 41064 19882 41140 19888
rect -210 19820 36 19880
rect -210 19817 -204 19820
rect -280 19811 -204 19817
rect 41064 19817 41070 19882
rect 41134 19880 41140 19882
rect 41134 19820 41380 19880
rect 41134 19817 41140 19820
rect 41064 19811 41140 19817
rect 1080 19252 1140 19492
rect 3512 19456 3572 19492
rect 5944 19252 6004 19492
rect 1072 19246 1149 19252
rect 1072 19182 1078 19246
rect 1143 19182 1149 19246
rect 1072 19176 1149 19182
rect 5936 19246 6012 19252
rect 5936 19181 5942 19246
rect 6006 19181 6012 19246
rect 5936 19175 6012 19181
rect -756 19117 -680 19123
rect -756 19053 -750 19117
rect -686 19115 -680 19117
rect 8376 19115 8436 19492
rect 10808 19252 10868 19492
rect 13240 19456 13300 19492
rect 15672 19252 15732 19492
rect 10800 19246 10876 19252
rect 10800 19181 10806 19246
rect 10870 19181 10876 19246
rect 10800 19175 10876 19181
rect 15664 19246 15740 19252
rect 15664 19181 15670 19246
rect 15734 19181 15740 19246
rect 15664 19175 15740 19181
rect 18104 19115 18164 19492
rect 20536 19252 20596 19492
rect 22968 19456 23028 19492
rect 25400 19252 25460 19492
rect 20528 19246 20604 19252
rect 20528 19181 20534 19246
rect 20598 19181 20604 19246
rect 20528 19175 20604 19181
rect 25392 19246 25468 19252
rect 25392 19181 25398 19246
rect 25462 19181 25468 19246
rect 25392 19175 25468 19181
rect 27832 19115 27892 19492
rect 30264 19252 30324 19492
rect 32696 19456 32756 19492
rect 35128 19252 35188 19492
rect 30256 19246 30332 19252
rect 30256 19181 30262 19246
rect 30326 19181 30332 19246
rect 30256 19175 30332 19181
rect 35120 19246 35196 19252
rect 35120 19181 35126 19246
rect 35190 19181 35196 19246
rect 35120 19175 35196 19181
rect 37560 19115 37620 19492
rect 39992 19252 40052 19492
rect 42424 19252 42484 19492
rect 39984 19246 40060 19252
rect 39984 19181 39990 19246
rect 40054 19181 40060 19246
rect 39984 19175 40060 19181
rect 42416 19246 42493 19252
rect 42416 19182 42422 19246
rect 42487 19182 42493 19246
rect 42416 19176 42493 19182
rect -686 19055 40380 19115
rect -686 19053 -680 19055
rect -756 19047 -680 19053
rect 5936 18932 6012 18938
rect 5936 18929 5942 18932
rect 2468 18869 5942 18929
rect 355 18802 432 18808
rect 355 18738 361 18802
rect 426 18738 432 18802
rect 355 18732 432 18738
rect 364 18492 424 18732
rect 2796 18492 2856 18869
rect 5936 18867 5942 18869
rect 6006 18929 6012 18932
rect 10800 18932 10876 18938
rect 10800 18929 10806 18932
rect 6006 18869 10806 18929
rect 6006 18867 6012 18869
rect 5936 18861 6012 18867
rect 5228 18492 5288 18528
rect 7660 18492 7720 18869
rect 10800 18867 10806 18869
rect 10870 18929 10876 18932
rect 15664 18932 15740 18938
rect 15664 18929 15670 18932
rect 10870 18869 15670 18929
rect 10870 18867 10876 18869
rect 10800 18861 10876 18867
rect 10092 18492 10152 18528
rect 12524 18492 12584 18869
rect 15664 18867 15670 18869
rect 15734 18929 15740 18932
rect 20528 18932 20604 18938
rect 20528 18929 20534 18932
rect 15734 18869 20534 18929
rect 15734 18867 15740 18869
rect 15664 18861 15740 18867
rect 14956 18492 15016 18528
rect 17388 18492 17448 18869
rect 20528 18867 20534 18869
rect 20598 18929 20604 18932
rect 25392 18932 25468 18938
rect 25392 18929 25398 18932
rect 20598 18869 25398 18929
rect 20598 18867 20604 18869
rect 20528 18861 20604 18867
rect 19820 18492 19880 18528
rect 22252 18492 22312 18869
rect 25392 18867 25398 18869
rect 25462 18929 25468 18932
rect 30256 18932 30332 18938
rect 30256 18929 30262 18932
rect 25462 18869 30262 18929
rect 25462 18867 25468 18869
rect 25392 18861 25468 18867
rect 24684 18492 24744 18528
rect 27116 18492 27176 18869
rect 30256 18867 30262 18869
rect 30326 18929 30332 18932
rect 35120 18932 35196 18938
rect 35120 18929 35126 18932
rect 30326 18869 35126 18929
rect 30326 18867 30332 18869
rect 30256 18861 30332 18867
rect 29548 18492 29608 18528
rect 31980 18492 32040 18869
rect 35120 18867 35126 18869
rect 35190 18929 35196 18932
rect 39984 18932 40060 18938
rect 39984 18929 39990 18932
rect 35190 18869 39990 18929
rect 35190 18867 35196 18869
rect 35120 18861 35196 18867
rect 34412 18492 34472 18528
rect 36844 18492 36904 18869
rect 39984 18867 39990 18869
rect 40054 18929 40060 18932
rect 43404 18931 43480 18937
rect 43404 18929 43410 18931
rect 40054 18869 43410 18929
rect 40054 18867 40060 18869
rect 39984 18861 40060 18867
rect 43404 18867 43410 18869
rect 43474 18867 43480 18931
rect 43404 18861 43480 18867
rect 41699 18802 41776 18808
rect 41699 18738 41705 18802
rect 41770 18738 41776 18802
rect 41699 18732 41776 18738
rect 39276 18492 39336 18528
rect 41708 18492 41768 18732
rect 1708 18167 1784 18173
rect 1708 18164 1714 18167
rect 1468 18104 1714 18164
rect 1708 18102 1714 18104
rect 1778 18102 1784 18167
rect 43052 18167 43128 18173
rect 43052 18164 43058 18167
rect 42812 18104 43058 18164
rect 1708 18096 1784 18102
rect 43052 18102 43058 18104
rect 43122 18102 43128 18167
rect 43052 18096 43128 18102
rect -280 17450 -204 17456
rect -280 17385 -274 17450
rect -210 17448 -204 17450
rect 41064 17450 41140 17456
rect -210 17388 36 17448
rect -210 17385 -204 17388
rect -280 17379 -204 17385
rect 41064 17385 41070 17450
rect 41134 17448 41140 17450
rect 41134 17388 41380 17448
rect 41134 17385 41140 17388
rect 41064 17379 41140 17385
rect 1080 16820 1140 17060
rect 3512 17024 3572 17060
rect 1072 16814 1149 16820
rect 1072 16750 1078 16814
rect 1143 16750 1149 16814
rect 1072 16744 1149 16750
rect -632 16685 -556 16691
rect -632 16621 -626 16685
rect -562 16683 -556 16685
rect 5944 16683 6004 17060
rect 8376 17024 8436 17060
rect 10808 16683 10868 17060
rect 13240 17024 13300 17060
rect 15672 16683 15732 17060
rect 18104 17024 18164 17060
rect 20536 16683 20596 17060
rect 22968 17024 23028 17060
rect 25400 16683 25460 17060
rect 27832 17024 27892 17060
rect 30264 16683 30324 17060
rect 32696 17024 32756 17060
rect 35128 16683 35188 17060
rect 37560 17024 37620 17060
rect 39992 16683 40052 17060
rect 42424 16820 42484 17060
rect 42416 16814 42493 16820
rect 42416 16750 42422 16814
rect 42487 16750 42493 16814
rect 42416 16744 42493 16750
rect -562 16623 40380 16683
rect -562 16621 -556 16623
rect -632 16615 -556 16621
rect -756 16499 -680 16505
rect -756 16435 -750 16499
rect -686 16497 -680 16499
rect -686 16437 40380 16497
rect -686 16435 -680 16437
rect -756 16429 -680 16435
rect 355 16370 432 16376
rect 355 16306 361 16370
rect 426 16306 432 16370
rect 355 16300 432 16306
rect 364 16060 424 16300
rect 5228 16060 5288 16096
rect 7660 16060 7720 16437
rect 10092 16060 10152 16096
rect 14956 16060 15016 16096
rect 17388 16060 17448 16437
rect 19820 16060 19880 16096
rect 24684 16060 24744 16096
rect 27116 16060 27176 16437
rect 29548 16060 29608 16096
rect 34412 16060 34472 16096
rect 36844 16060 36904 16437
rect 41699 16370 41776 16376
rect 41699 16306 41705 16370
rect 41770 16306 41776 16370
rect 41699 16300 41776 16306
rect 39276 16060 39336 16096
rect 41708 16060 41768 16300
rect 1708 15735 1784 15741
rect 1708 15732 1714 15735
rect 1468 15672 1714 15732
rect 1708 15670 1714 15672
rect 1778 15670 1784 15735
rect 43052 15735 43128 15741
rect 43052 15732 43058 15735
rect 42812 15672 43058 15732
rect 1708 15664 1784 15670
rect 43052 15670 43058 15672
rect 43122 15670 43128 15735
rect 43052 15664 43128 15670
rect -280 15018 -204 15024
rect -280 14953 -274 15018
rect -210 15016 -204 15018
rect 41064 15018 41140 15024
rect -210 14956 36 15016
rect -210 14953 -204 14956
rect -280 14947 -204 14953
rect 41064 14953 41070 15018
rect 41134 15016 41140 15018
rect 41134 14956 41380 15016
rect 41134 14953 41140 14956
rect 41064 14947 41140 14953
rect 1080 14388 1140 14628
rect 1072 14382 1149 14388
rect 1072 14318 1078 14382
rect 1143 14318 1149 14382
rect 1072 14312 1149 14318
rect 3512 14251 3572 14628
rect 5944 14388 6004 14628
rect 8376 14592 8436 14628
rect 10808 14388 10868 14628
rect 5936 14382 6012 14388
rect 5936 14317 5942 14382
rect 6006 14317 6012 14382
rect 5936 14311 6012 14317
rect 10800 14382 10876 14388
rect 10800 14317 10806 14382
rect 10870 14317 10876 14382
rect 10800 14311 10876 14317
rect 13240 14251 13300 14628
rect 15672 14388 15732 14628
rect 18104 14592 18164 14628
rect 20536 14388 20596 14628
rect 15664 14382 15740 14388
rect 15664 14317 15670 14382
rect 15734 14317 15740 14382
rect 15664 14311 15740 14317
rect 20528 14382 20604 14388
rect 20528 14317 20534 14382
rect 20598 14317 20604 14382
rect 20528 14311 20604 14317
rect 22968 14251 23028 14628
rect 25400 14388 25460 14628
rect 27832 14592 27892 14628
rect 30264 14388 30324 14628
rect 25392 14382 25468 14388
rect 25392 14317 25398 14382
rect 25462 14317 25468 14382
rect 25392 14311 25468 14317
rect 30256 14382 30332 14388
rect 30256 14317 30262 14382
rect 30326 14317 30332 14382
rect 30256 14311 30332 14317
rect 32696 14251 32756 14628
rect 35128 14388 35188 14628
rect 37560 14592 37620 14628
rect 39992 14388 40052 14628
rect 42424 14388 42484 14628
rect 35120 14382 35196 14388
rect 35120 14317 35126 14382
rect 35190 14317 35196 14382
rect 35120 14311 35196 14317
rect 39984 14382 40060 14388
rect 39984 14317 39990 14382
rect 40054 14317 40060 14382
rect 39984 14311 40060 14317
rect 42416 14382 42493 14388
rect 42416 14318 42422 14382
rect 42487 14318 42493 14382
rect 42416 14312 42493 14318
rect 43652 14253 43728 14259
rect 43652 14251 43658 14253
rect 2468 14191 43658 14251
rect 43652 14189 43658 14191
rect 43722 14189 43728 14253
rect 43652 14183 43728 14189
rect 5936 14068 6012 14074
rect 5936 14065 5942 14068
rect 2468 14005 5942 14065
rect 355 13938 432 13944
rect 355 13874 361 13938
rect 426 13874 432 13938
rect 355 13868 432 13874
rect 364 13628 424 13868
rect 2796 13628 2856 14005
rect 5936 14003 5942 14005
rect 6006 14065 6012 14068
rect 10800 14068 10876 14074
rect 10800 14065 10806 14068
rect 6006 14005 10806 14065
rect 6006 14003 6012 14005
rect 5936 13997 6012 14003
rect 5228 13628 5288 13664
rect 7660 13628 7720 14005
rect 10800 14003 10806 14005
rect 10870 14065 10876 14068
rect 15664 14068 15740 14074
rect 15664 14065 15670 14068
rect 10870 14005 15670 14065
rect 10870 14003 10876 14005
rect 10800 13997 10876 14003
rect 10092 13628 10152 13664
rect 12524 13628 12584 14005
rect 15664 14003 15670 14005
rect 15734 14065 15740 14068
rect 20528 14068 20604 14074
rect 20528 14065 20534 14068
rect 15734 14005 20534 14065
rect 15734 14003 15740 14005
rect 15664 13997 15740 14003
rect 14956 13628 15016 13664
rect 17388 13628 17448 14005
rect 20528 14003 20534 14005
rect 20598 14065 20604 14068
rect 25392 14068 25468 14074
rect 25392 14065 25398 14068
rect 20598 14005 25398 14065
rect 20598 14003 20604 14005
rect 20528 13997 20604 14003
rect 19820 13628 19880 13664
rect 22252 13628 22312 14005
rect 25392 14003 25398 14005
rect 25462 14065 25468 14068
rect 30256 14068 30332 14074
rect 30256 14065 30262 14068
rect 25462 14005 30262 14065
rect 25462 14003 25468 14005
rect 25392 13997 25468 14003
rect 24684 13628 24744 13664
rect 27116 13628 27176 14005
rect 30256 14003 30262 14005
rect 30326 14065 30332 14068
rect 35120 14068 35196 14074
rect 35120 14065 35126 14068
rect 30326 14005 35126 14065
rect 30326 14003 30332 14005
rect 30256 13997 30332 14003
rect 29548 13628 29608 13664
rect 31980 13628 32040 14005
rect 35120 14003 35126 14005
rect 35190 14065 35196 14068
rect 39984 14068 40060 14074
rect 39984 14065 39990 14068
rect 35190 14005 39990 14065
rect 35190 14003 35196 14005
rect 35120 13997 35196 14003
rect 34412 13628 34472 13664
rect 36844 13628 36904 14005
rect 39984 14003 39990 14005
rect 40054 14065 40060 14068
rect 43404 14067 43480 14073
rect 43404 14065 43410 14067
rect 40054 14005 43410 14065
rect 40054 14003 40060 14005
rect 39984 13997 40060 14003
rect 43404 14003 43410 14005
rect 43474 14003 43480 14067
rect 43404 13997 43480 14003
rect 41699 13938 41776 13944
rect 41699 13874 41705 13938
rect 41770 13874 41776 13938
rect 41699 13868 41776 13874
rect 39276 13628 39336 13664
rect 41708 13628 41768 13868
rect 1708 13303 1784 13309
rect 1708 13300 1714 13303
rect 1468 13240 1714 13300
rect 1708 13238 1714 13240
rect 1778 13238 1784 13303
rect 43052 13303 43128 13309
rect 43052 13300 43058 13303
rect 42812 13240 43058 13300
rect 1708 13232 1784 13238
rect 43052 13238 43058 13240
rect 43122 13238 43128 13303
rect 43052 13232 43128 13238
rect -280 12586 -204 12592
rect -280 12521 -274 12586
rect -210 12584 -204 12586
rect 41064 12586 41140 12592
rect -210 12524 36 12584
rect -210 12521 -204 12524
rect -280 12515 -204 12521
rect 41064 12521 41070 12586
rect 41134 12584 41140 12586
rect 41134 12524 41380 12584
rect 41134 12521 41140 12524
rect 41064 12515 41140 12521
rect 1080 11956 1140 12196
rect 3512 12160 3572 12196
rect 1072 11950 1149 11956
rect 1072 11886 1078 11950
rect 1143 11886 1149 11950
rect 1072 11880 1149 11886
rect -632 11821 -556 11827
rect -632 11757 -626 11821
rect -562 11819 -556 11821
rect 5944 11819 6004 12196
rect 8376 12160 8436 12196
rect 10808 11819 10868 12196
rect 13240 12160 13300 12196
rect 15672 11819 15732 12196
rect 18104 12160 18164 12196
rect 20536 11819 20596 12196
rect 22968 12160 23028 12196
rect 25400 11819 25460 12196
rect 27832 12160 27892 12196
rect 30264 11819 30324 12196
rect 32696 12160 32756 12196
rect 35128 11819 35188 12196
rect 37560 12160 37620 12196
rect 39992 11819 40052 12196
rect 42424 11956 42484 12196
rect 42416 11950 42493 11956
rect 42416 11886 42422 11950
rect 42487 11886 42493 11950
rect 42416 11880 42493 11886
rect -562 11759 40380 11819
rect -562 11757 -556 11759
rect -632 11751 -556 11757
rect 43528 11635 43604 11641
rect 43528 11633 43534 11635
rect 2468 11573 43534 11633
rect 355 11506 432 11512
rect 355 11442 361 11506
rect 426 11442 432 11506
rect 355 11436 432 11442
rect 364 11196 424 11436
rect 2796 11196 2856 11573
rect 5228 11196 5288 11232
rect 7660 11196 7720 11573
rect 10092 11196 10152 11232
rect 12524 11196 12584 11573
rect 14956 11196 15016 11232
rect 17388 11196 17448 11573
rect 19820 11196 19880 11232
rect 22252 11196 22312 11573
rect 24684 11196 24744 11232
rect 27116 11196 27176 11573
rect 29548 11196 29608 11232
rect 31980 11196 32040 11573
rect 34412 11196 34472 11232
rect 36844 11196 36904 11573
rect 43528 11571 43534 11573
rect 43598 11571 43604 11635
rect 43528 11565 43604 11571
rect 41699 11506 41776 11512
rect 41699 11442 41705 11506
rect 41770 11442 41776 11506
rect 41699 11436 41776 11442
rect 39276 11196 39336 11232
rect 41708 11196 41768 11436
rect 1708 10871 1784 10877
rect 1708 10868 1714 10871
rect 1468 10808 1714 10868
rect 1708 10806 1714 10808
rect 1778 10806 1784 10871
rect 43052 10871 43128 10877
rect 43052 10868 43058 10871
rect 42812 10808 43058 10868
rect 1708 10800 1784 10806
rect 43052 10806 43058 10808
rect 43122 10806 43128 10871
rect 43052 10800 43128 10806
rect -280 10154 -204 10160
rect -280 10089 -274 10154
rect -210 10152 -204 10154
rect 41064 10154 41140 10160
rect -210 10092 36 10152
rect -210 10089 -204 10092
rect -280 10083 -204 10089
rect 41064 10089 41070 10154
rect 41134 10152 41140 10154
rect 41134 10092 41380 10152
rect 41134 10089 41140 10092
rect 41064 10083 41140 10089
rect 1080 9524 1140 9764
rect 3512 9728 3572 9764
rect 5944 9524 6004 9764
rect 8376 9728 8436 9764
rect 10808 9524 10868 9764
rect 13240 9728 13300 9764
rect 15672 9524 15732 9764
rect 18104 9728 18164 9764
rect 20536 9524 20596 9764
rect 22968 9728 23028 9764
rect 25400 9524 25460 9764
rect 27832 9728 27892 9764
rect 30264 9524 30324 9764
rect 32696 9728 32756 9764
rect 35128 9524 35188 9764
rect 37560 9728 37620 9764
rect 39992 9524 40052 9764
rect 42424 9524 42484 9764
rect 1072 9518 1149 9524
rect 1072 9454 1078 9518
rect 1143 9454 1149 9518
rect 1072 9448 1149 9454
rect 5936 9518 6012 9524
rect 5936 9453 5942 9518
rect 6006 9453 6012 9518
rect 5936 9447 6012 9453
rect 10800 9518 10876 9524
rect 10800 9453 10806 9518
rect 10870 9453 10876 9518
rect 10800 9447 10876 9453
rect 15664 9518 15740 9524
rect 15664 9453 15670 9518
rect 15734 9453 15740 9518
rect 15664 9447 15740 9453
rect 20528 9518 20604 9524
rect 20528 9453 20534 9518
rect 20598 9453 20604 9518
rect 20528 9447 20604 9453
rect 25392 9518 25468 9524
rect 25392 9453 25398 9518
rect 25462 9453 25468 9518
rect 25392 9447 25468 9453
rect 30256 9518 30332 9524
rect 30256 9453 30262 9518
rect 30326 9453 30332 9518
rect 30256 9447 30332 9453
rect 35120 9518 35196 9524
rect 35120 9453 35126 9518
rect 35190 9453 35196 9518
rect 35120 9447 35196 9453
rect 39984 9518 40060 9524
rect 39984 9453 39990 9518
rect 40054 9453 40060 9518
rect 39984 9447 40060 9453
rect 42416 9518 42493 9524
rect 42416 9454 42422 9518
rect 42487 9454 42493 9518
rect 42416 9448 42493 9454
rect 2468 9327 40380 9387
rect 5936 9204 6012 9210
rect 5936 9201 5942 9204
rect 2468 9141 5942 9201
rect 355 9074 432 9080
rect 355 9010 361 9074
rect 426 9010 432 9074
rect 355 9004 432 9010
rect 364 8764 424 9004
rect 2796 8764 2856 9141
rect 5936 9139 5942 9141
rect 6006 9201 6012 9204
rect 10800 9204 10876 9210
rect 10800 9201 10806 9204
rect 6006 9141 10806 9201
rect 6006 9139 6012 9141
rect 5936 9133 6012 9139
rect 5228 8764 5288 8800
rect 7660 8764 7720 9141
rect 10800 9139 10806 9141
rect 10870 9201 10876 9204
rect 15664 9204 15740 9210
rect 15664 9201 15670 9204
rect 10870 9141 15670 9201
rect 10870 9139 10876 9141
rect 10800 9133 10876 9139
rect 10092 8764 10152 8800
rect 12524 8764 12584 9141
rect 15664 9139 15670 9141
rect 15734 9201 15740 9204
rect 20528 9204 20604 9210
rect 20528 9201 20534 9204
rect 15734 9141 20534 9201
rect 15734 9139 15740 9141
rect 15664 9133 15740 9139
rect 14956 8764 15016 8800
rect 17388 8764 17448 9141
rect 20528 9139 20534 9141
rect 20598 9201 20604 9204
rect 25392 9204 25468 9210
rect 25392 9201 25398 9204
rect 20598 9141 25398 9201
rect 20598 9139 20604 9141
rect 20528 9133 20604 9139
rect 19820 8764 19880 8800
rect 22252 8764 22312 9141
rect 25392 9139 25398 9141
rect 25462 9201 25468 9204
rect 30256 9204 30332 9210
rect 30256 9201 30262 9204
rect 25462 9141 30262 9201
rect 25462 9139 25468 9141
rect 25392 9133 25468 9139
rect 24684 8764 24744 8800
rect 27116 8764 27176 9141
rect 30256 9139 30262 9141
rect 30326 9201 30332 9204
rect 35120 9204 35196 9210
rect 35120 9201 35126 9204
rect 30326 9141 35126 9201
rect 30326 9139 30332 9141
rect 30256 9133 30332 9139
rect 29548 8764 29608 8800
rect 31980 8764 32040 9141
rect 35120 9139 35126 9141
rect 35190 9201 35196 9204
rect 39984 9204 40060 9210
rect 39984 9201 39990 9204
rect 35190 9141 39990 9201
rect 35190 9139 35196 9141
rect 35120 9133 35196 9139
rect 34412 8764 34472 8800
rect 36844 8764 36904 9141
rect 39984 9139 39990 9141
rect 40054 9201 40060 9204
rect 43404 9203 43480 9209
rect 43404 9201 43410 9203
rect 40054 9141 43410 9201
rect 40054 9139 40060 9141
rect 39984 9133 40060 9139
rect 43404 9139 43410 9141
rect 43474 9139 43480 9203
rect 43404 9133 43480 9139
rect 41699 9074 41776 9080
rect 41699 9010 41705 9074
rect 41770 9010 41776 9074
rect 41699 9004 41776 9010
rect 39276 8764 39336 8800
rect 41708 8764 41768 9004
rect 1708 8439 1784 8445
rect 1708 8436 1714 8439
rect 1468 8376 1714 8436
rect 1708 8374 1714 8376
rect 1778 8374 1784 8439
rect 43052 8439 43128 8445
rect 43052 8436 43058 8439
rect 42812 8376 43058 8436
rect 1708 8368 1784 8374
rect 43052 8374 43058 8376
rect 43122 8374 43128 8439
rect 43052 8368 43128 8374
rect -280 7722 -204 7728
rect -280 7657 -274 7722
rect -210 7720 -204 7722
rect 41064 7722 41140 7728
rect -210 7660 36 7720
rect -210 7657 -204 7660
rect -280 7651 -204 7657
rect 41064 7657 41070 7722
rect 41134 7720 41140 7722
rect 41134 7660 41380 7720
rect 41134 7657 41140 7660
rect 41064 7651 41140 7657
rect 1080 7092 1140 7332
rect 3512 7296 3572 7332
rect 1072 7086 1149 7092
rect 1072 7022 1078 7086
rect 1143 7022 1149 7086
rect 1072 7016 1149 7022
rect -632 6957 -556 6963
rect -632 6893 -626 6957
rect -562 6955 -556 6957
rect 5944 6955 6004 7332
rect 8376 7296 8436 7332
rect 10808 6955 10868 7332
rect 13240 7296 13300 7332
rect 15672 6955 15732 7332
rect 18104 7296 18164 7332
rect 20536 6955 20596 7332
rect 22968 7296 23028 7332
rect 25400 6955 25460 7332
rect 27832 7296 27892 7332
rect 30264 6955 30324 7332
rect 32696 7296 32756 7332
rect 35128 6955 35188 7332
rect 37560 7296 37620 7332
rect 39992 6955 40052 7332
rect 42424 7092 42484 7332
rect 42416 7086 42493 7092
rect 42416 7022 42422 7086
rect 42487 7022 42493 7086
rect 42416 7016 42493 7022
rect -562 6895 40380 6955
rect -562 6893 -556 6895
rect -632 6887 -556 6893
rect 43528 6771 43604 6777
rect 43528 6769 43534 6771
rect 2468 6709 43534 6769
rect 355 6642 432 6648
rect 355 6578 361 6642
rect 426 6578 432 6642
rect 355 6572 432 6578
rect 364 6332 424 6572
rect 2796 6332 2856 6709
rect 5228 6332 5288 6368
rect 7660 6332 7720 6709
rect 10092 6332 10152 6368
rect 12524 6332 12584 6709
rect 14956 6332 15016 6368
rect 17388 6332 17448 6709
rect 19820 6332 19880 6368
rect 22252 6332 22312 6709
rect 24684 6332 24744 6368
rect 27116 6332 27176 6709
rect 29548 6332 29608 6368
rect 31980 6332 32040 6709
rect 34412 6332 34472 6368
rect 36844 6332 36904 6709
rect 43528 6707 43534 6709
rect 43598 6707 43604 6771
rect 43528 6701 43604 6707
rect 41699 6642 41776 6648
rect 41699 6578 41705 6642
rect 41770 6578 41776 6642
rect 41699 6572 41776 6578
rect 39276 6332 39336 6368
rect 41708 6332 41768 6572
rect 1708 6007 1784 6013
rect 1708 6004 1714 6007
rect 1468 5944 1714 6004
rect 1708 5942 1714 5944
rect 1778 5942 1784 6007
rect 43052 6007 43128 6013
rect 43052 6004 43058 6007
rect 42812 5944 43058 6004
rect 1708 5936 1784 5942
rect 43052 5942 43058 5944
rect 43122 5942 43128 6007
rect 43052 5936 43128 5942
rect -280 5290 -204 5296
rect -280 5225 -274 5290
rect -210 5288 -204 5290
rect 41064 5290 41140 5296
rect -210 5228 36 5288
rect -210 5225 -204 5228
rect -280 5219 -204 5225
rect 41064 5225 41070 5290
rect 41134 5288 41140 5290
rect 41134 5228 41380 5288
rect 41134 5225 41140 5228
rect 41064 5219 41140 5225
rect 1080 4660 1140 4900
rect 3512 4864 3572 4900
rect 5944 4660 6004 4900
rect 8376 4864 8436 4900
rect 10808 4660 10868 4900
rect 13240 4864 13300 4900
rect 15672 4660 15732 4900
rect 18104 4864 18164 4900
rect 20536 4660 20596 4900
rect 22968 4864 23028 4900
rect 25400 4660 25460 4900
rect 27832 4864 27892 4900
rect 30264 4660 30324 4900
rect 32696 4864 32756 4900
rect 35128 4660 35188 4900
rect 37560 4864 37620 4900
rect 39992 4660 40052 4900
rect 42424 4660 42484 4900
rect 1072 4654 1149 4660
rect 1072 4590 1078 4654
rect 1143 4590 1149 4654
rect 1072 4584 1149 4590
rect 5936 4654 6012 4660
rect 5936 4589 5942 4654
rect 6006 4589 6012 4654
rect 5936 4583 6012 4589
rect 10800 4654 10876 4660
rect 10800 4589 10806 4654
rect 10870 4589 10876 4654
rect 10800 4583 10876 4589
rect 15664 4654 15740 4660
rect 15664 4589 15670 4654
rect 15734 4589 15740 4654
rect 15664 4583 15740 4589
rect 20528 4654 20604 4660
rect 20528 4589 20534 4654
rect 20598 4589 20604 4654
rect 20528 4583 20604 4589
rect 25392 4654 25468 4660
rect 25392 4589 25398 4654
rect 25462 4589 25468 4654
rect 25392 4583 25468 4589
rect 30256 4654 30332 4660
rect 30256 4589 30262 4654
rect 30326 4589 30332 4654
rect 30256 4583 30332 4589
rect 35120 4654 35196 4660
rect 35120 4589 35126 4654
rect 35190 4589 35196 4654
rect 35120 4583 35196 4589
rect 39984 4654 40060 4660
rect 39984 4589 39990 4654
rect 40054 4589 40060 4654
rect 39984 4583 40060 4589
rect 42416 4654 42493 4660
rect 42416 4590 42422 4654
rect 42487 4590 42493 4654
rect 42416 4584 42493 4590
rect 2468 4463 40380 4523
rect 5936 4340 6012 4346
rect 5936 4337 5942 4340
rect 2468 4277 5942 4337
rect 355 4210 432 4216
rect 355 4146 361 4210
rect 426 4146 432 4210
rect 355 4140 432 4146
rect 364 3900 424 4140
rect 2796 3900 2856 4277
rect 5936 4275 5942 4277
rect 6006 4337 6012 4340
rect 10800 4340 10876 4346
rect 10800 4337 10806 4340
rect 6006 4277 10806 4337
rect 6006 4275 6012 4277
rect 5936 4269 6012 4275
rect 5228 3900 5288 3936
rect 7660 3900 7720 4277
rect 10800 4275 10806 4277
rect 10870 4337 10876 4340
rect 15664 4340 15740 4346
rect 15664 4337 15670 4340
rect 10870 4277 15670 4337
rect 10870 4275 10876 4277
rect 10800 4269 10876 4275
rect 10092 3900 10152 3936
rect 12524 3900 12584 4277
rect 15664 4275 15670 4277
rect 15734 4337 15740 4340
rect 20528 4340 20604 4346
rect 20528 4337 20534 4340
rect 15734 4277 20534 4337
rect 15734 4275 15740 4277
rect 15664 4269 15740 4275
rect 14956 3900 15016 3936
rect 17388 3900 17448 4277
rect 20528 4275 20534 4277
rect 20598 4337 20604 4340
rect 25392 4340 25468 4346
rect 25392 4337 25398 4340
rect 20598 4277 25398 4337
rect 20598 4275 20604 4277
rect 20528 4269 20604 4275
rect 19820 3900 19880 3936
rect 22252 3900 22312 4277
rect 25392 4275 25398 4277
rect 25462 4337 25468 4340
rect 30256 4340 30332 4346
rect 30256 4337 30262 4340
rect 25462 4277 30262 4337
rect 25462 4275 25468 4277
rect 25392 4269 25468 4275
rect 24684 3900 24744 3936
rect 27116 3900 27176 4277
rect 30256 4275 30262 4277
rect 30326 4337 30332 4340
rect 35120 4340 35196 4346
rect 35120 4337 35126 4340
rect 30326 4277 35126 4337
rect 30326 4275 30332 4277
rect 30256 4269 30332 4275
rect 29548 3900 29608 3936
rect 31980 3900 32040 4277
rect 35120 4275 35126 4277
rect 35190 4337 35196 4340
rect 39984 4340 40060 4346
rect 39984 4337 39990 4340
rect 35190 4277 39990 4337
rect 35190 4275 35196 4277
rect 35120 4269 35196 4275
rect 34412 3900 34472 3936
rect 36844 3900 36904 4277
rect 39984 4275 39990 4277
rect 40054 4337 40060 4340
rect 43404 4340 43480 4346
rect 43404 4337 43410 4340
rect 40054 4277 43410 4337
rect 40054 4275 40060 4277
rect 39984 4269 40060 4275
rect 43404 4275 43410 4277
rect 43474 4275 43480 4340
rect 43404 4269 43480 4275
rect 41699 4210 41776 4216
rect 41699 4146 41705 4210
rect 41770 4146 41776 4210
rect 41699 4140 41776 4146
rect 39276 3900 39336 3936
rect 41708 3900 41768 4140
rect 1708 3575 1784 3581
rect 1708 3572 1714 3575
rect 1468 3512 1714 3572
rect 1708 3510 1714 3512
rect 1778 3510 1784 3575
rect 43052 3575 43128 3581
rect 43052 3572 43058 3575
rect 42812 3512 43058 3572
rect 1708 3504 1784 3510
rect 43052 3510 43058 3512
rect 43122 3510 43128 3575
rect 43052 3504 43128 3510
rect -280 2858 -204 2864
rect -280 2793 -274 2858
rect -210 2856 -204 2858
rect 41064 2858 41140 2864
rect -210 2796 36 2856
rect -210 2793 -204 2796
rect -280 2787 -204 2793
rect 41064 2793 41070 2858
rect 41134 2856 41140 2858
rect 41134 2796 41380 2856
rect 41134 2793 41140 2796
rect 41064 2787 41140 2793
rect 1080 2228 1140 2468
rect 3512 2432 3572 2468
rect 1072 2222 1149 2228
rect 1072 2158 1078 2222
rect 1143 2158 1149 2222
rect 1072 2152 1149 2158
rect -632 2093 -556 2099
rect -632 2029 -626 2093
rect -562 2091 -556 2093
rect 5944 2091 6004 2468
rect 8376 2432 8436 2468
rect 10808 2091 10868 2468
rect 13240 2432 13300 2468
rect 15672 2091 15732 2468
rect 18104 2432 18164 2468
rect 20536 2091 20596 2468
rect 22968 2432 23028 2468
rect 25400 2091 25460 2468
rect 27832 2432 27892 2468
rect 30264 2091 30324 2468
rect 32696 2432 32756 2468
rect 35128 2091 35188 2468
rect 37560 2432 37620 2468
rect 39992 2091 40052 2468
rect 42424 2228 42484 2468
rect 42416 2222 42493 2228
rect 42416 2158 42422 2222
rect 42487 2158 42493 2222
rect 42416 2152 42493 2158
rect -562 2031 40380 2091
rect -562 2029 -556 2031
rect -632 2023 -556 2029
rect 355 1778 432 1784
rect 355 1714 361 1778
rect 426 1714 432 1778
rect 355 1708 432 1714
rect 2787 1778 2864 1784
rect 2787 1714 2793 1778
rect 2858 1714 2864 1778
rect 2787 1708 2864 1714
rect 5219 1778 5296 1784
rect 5219 1714 5225 1778
rect 5290 1714 5296 1778
rect 5219 1708 5296 1714
rect 7651 1778 7728 1784
rect 7651 1714 7657 1778
rect 7722 1714 7728 1778
rect 7651 1708 7728 1714
rect 10083 1778 10160 1784
rect 10083 1714 10089 1778
rect 10154 1714 10160 1778
rect 10083 1708 10160 1714
rect 12515 1778 12592 1784
rect 12515 1714 12521 1778
rect 12586 1714 12592 1778
rect 12515 1708 12592 1714
rect 14947 1778 15024 1784
rect 14947 1714 14953 1778
rect 15018 1714 15024 1778
rect 14947 1708 15024 1714
rect 17379 1778 17456 1784
rect 17379 1714 17385 1778
rect 17450 1714 17456 1778
rect 17379 1708 17456 1714
rect 19811 1778 19888 1784
rect 19811 1714 19817 1778
rect 19882 1714 19888 1778
rect 19811 1708 19888 1714
rect 22243 1778 22320 1784
rect 22243 1714 22249 1778
rect 22314 1714 22320 1778
rect 22243 1708 22320 1714
rect 24675 1778 24752 1784
rect 24675 1714 24681 1778
rect 24746 1714 24752 1778
rect 24675 1708 24752 1714
rect 27107 1778 27184 1784
rect 27107 1714 27113 1778
rect 27178 1714 27184 1778
rect 27107 1708 27184 1714
rect 29539 1778 29616 1784
rect 29539 1714 29545 1778
rect 29610 1714 29616 1778
rect 29539 1708 29616 1714
rect 31971 1778 32048 1784
rect 31971 1714 31977 1778
rect 32042 1714 32048 1778
rect 31971 1708 32048 1714
rect 34403 1778 34480 1784
rect 34403 1714 34409 1778
rect 34474 1714 34480 1778
rect 34403 1708 34480 1714
rect 36835 1778 36912 1784
rect 36835 1714 36841 1778
rect 36906 1714 36912 1778
rect 36835 1708 36912 1714
rect 39267 1778 39344 1784
rect 39267 1714 39273 1778
rect 39338 1714 39344 1778
rect 39267 1708 39344 1714
rect 41699 1778 41776 1784
rect 41699 1714 41705 1778
rect 41770 1714 41776 1778
rect 41699 1708 41776 1714
rect 364 1468 424 1708
rect 2796 1468 2856 1708
rect 5228 1468 5288 1708
rect 7660 1468 7720 1708
rect 10092 1468 10152 1708
rect 12524 1468 12584 1708
rect 14956 1468 15016 1708
rect 17388 1468 17448 1708
rect 19820 1468 19880 1708
rect 22252 1468 22312 1708
rect 24684 1468 24744 1708
rect 27116 1468 27176 1708
rect 29548 1468 29608 1708
rect 31980 1468 32040 1708
rect 34412 1468 34472 1708
rect 36844 1468 36904 1708
rect 39276 1468 39336 1708
rect 41708 1468 41768 1708
rect 1708 1143 1784 1149
rect 1708 1140 1714 1143
rect 1468 1080 1714 1140
rect 1708 1078 1714 1080
rect 1778 1078 1784 1143
rect 4140 1143 4216 1149
rect 4140 1140 4146 1143
rect 3900 1080 4146 1140
rect 1708 1072 1784 1078
rect 4140 1078 4146 1080
rect 4210 1078 4216 1143
rect 6572 1143 6648 1149
rect 6572 1140 6578 1143
rect 6332 1080 6578 1140
rect 4140 1072 4216 1078
rect 6572 1078 6578 1080
rect 6642 1078 6648 1143
rect 9004 1143 9080 1149
rect 9004 1140 9010 1143
rect 8764 1080 9010 1140
rect 6572 1072 6648 1078
rect 9004 1078 9010 1080
rect 9074 1078 9080 1143
rect 11436 1143 11512 1149
rect 11436 1140 11442 1143
rect 11196 1080 11442 1140
rect 9004 1072 9080 1078
rect 11436 1078 11442 1080
rect 11506 1078 11512 1143
rect 13868 1143 13944 1149
rect 13868 1140 13874 1143
rect 13628 1080 13874 1140
rect 11436 1072 11512 1078
rect 13868 1078 13874 1080
rect 13938 1078 13944 1143
rect 16300 1143 16376 1149
rect 16300 1140 16306 1143
rect 16060 1080 16306 1140
rect 13868 1072 13944 1078
rect 16300 1078 16306 1080
rect 16370 1078 16376 1143
rect 18732 1143 18808 1149
rect 18732 1140 18738 1143
rect 18492 1080 18738 1140
rect 16300 1072 16376 1078
rect 18732 1078 18738 1080
rect 18802 1078 18808 1143
rect 21164 1143 21240 1149
rect 21164 1140 21170 1143
rect 20924 1080 21170 1140
rect 18732 1072 18808 1078
rect 21164 1078 21170 1080
rect 21234 1078 21240 1143
rect 23596 1143 23672 1149
rect 23596 1140 23602 1143
rect 23356 1080 23602 1140
rect 21164 1072 21240 1078
rect 23596 1078 23602 1080
rect 23666 1078 23672 1143
rect 26028 1143 26104 1149
rect 26028 1140 26034 1143
rect 25788 1080 26034 1140
rect 23596 1072 23672 1078
rect 26028 1078 26034 1080
rect 26098 1078 26104 1143
rect 28460 1143 28536 1149
rect 28460 1140 28466 1143
rect 28220 1080 28466 1140
rect 26028 1072 26104 1078
rect 28460 1078 28466 1080
rect 28530 1078 28536 1143
rect 30892 1143 30968 1149
rect 30892 1140 30898 1143
rect 30652 1080 30898 1140
rect 28460 1072 28536 1078
rect 30892 1078 30898 1080
rect 30962 1078 30968 1143
rect 33324 1143 33400 1149
rect 33324 1140 33330 1143
rect 33084 1080 33330 1140
rect 30892 1072 30968 1078
rect 33324 1078 33330 1080
rect 33394 1078 33400 1143
rect 35756 1143 35832 1149
rect 35756 1140 35762 1143
rect 35516 1080 35762 1140
rect 33324 1072 33400 1078
rect 35756 1078 35762 1080
rect 35826 1078 35832 1143
rect 38188 1143 38264 1149
rect 38188 1140 38194 1143
rect 37948 1080 38194 1140
rect 35756 1072 35832 1078
rect 38188 1078 38194 1080
rect 38258 1078 38264 1143
rect 40620 1143 40696 1149
rect 40620 1140 40626 1143
rect 40380 1080 40626 1140
rect 38188 1072 38264 1078
rect 40620 1078 40626 1080
rect 40690 1078 40696 1143
rect 43052 1143 43128 1149
rect 43052 1140 43058 1143
rect 42812 1080 43058 1140
rect 40620 1072 40696 1078
rect 43052 1078 43058 1080
rect 43122 1078 43128 1143
rect 43052 1072 43128 1078
rect -280 426 -204 432
rect -280 361 -274 426
rect -210 424 -204 426
rect 2152 426 2228 432
rect -210 364 36 424
rect -210 361 -204 364
rect -280 355 -204 361
rect 2152 361 2158 426
rect 2222 424 2228 426
rect 4584 426 4660 432
rect 2222 364 2468 424
rect 2222 361 2228 364
rect 2152 355 2228 361
rect 4584 361 4590 426
rect 4654 424 4660 426
rect 7016 426 7092 432
rect 4654 364 4900 424
rect 4654 361 4660 364
rect 4584 355 4660 361
rect 7016 361 7022 426
rect 7086 424 7092 426
rect 9448 426 9524 432
rect 7086 364 7332 424
rect 7086 361 7092 364
rect 7016 355 7092 361
rect 9448 361 9454 426
rect 9518 424 9524 426
rect 11880 426 11956 432
rect 9518 364 9764 424
rect 9518 361 9524 364
rect 9448 355 9524 361
rect 11880 361 11886 426
rect 11950 424 11956 426
rect 14312 426 14388 432
rect 11950 364 12196 424
rect 11950 361 11956 364
rect 11880 355 11956 361
rect 14312 361 14318 426
rect 14382 424 14388 426
rect 16744 426 16820 432
rect 14382 364 14628 424
rect 14382 361 14388 364
rect 14312 355 14388 361
rect 16744 361 16750 426
rect 16814 424 16820 426
rect 19176 426 19252 432
rect 16814 364 17060 424
rect 16814 361 16820 364
rect 16744 355 16820 361
rect 19176 361 19182 426
rect 19246 424 19252 426
rect 21608 426 21684 432
rect 19246 364 19492 424
rect 19246 361 19252 364
rect 19176 355 19252 361
rect 21608 361 21614 426
rect 21678 424 21684 426
rect 24040 426 24116 432
rect 21678 364 21924 424
rect 21678 361 21684 364
rect 21608 355 21684 361
rect 24040 361 24046 426
rect 24110 424 24116 426
rect 26472 426 26548 432
rect 24110 364 24356 424
rect 24110 361 24116 364
rect 24040 355 24116 361
rect 26472 361 26478 426
rect 26542 424 26548 426
rect 28904 426 28980 432
rect 26542 364 26788 424
rect 26542 361 26548 364
rect 26472 355 26548 361
rect 28904 361 28910 426
rect 28974 424 28980 426
rect 31336 426 31412 432
rect 28974 364 29220 424
rect 28974 361 28980 364
rect 28904 355 28980 361
rect 31336 361 31342 426
rect 31406 424 31412 426
rect 33768 426 33844 432
rect 31406 364 31652 424
rect 31406 361 31412 364
rect 31336 355 31412 361
rect 33768 361 33774 426
rect 33838 424 33844 426
rect 36200 426 36276 432
rect 33838 364 34084 424
rect 33838 361 33844 364
rect 33768 355 33844 361
rect 36200 361 36206 426
rect 36270 424 36276 426
rect 38632 426 38708 432
rect 36270 364 36516 424
rect 36270 361 36276 364
rect 36200 355 36276 361
rect 38632 361 38638 426
rect 38702 424 38708 426
rect 41064 426 41140 432
rect 38702 364 38948 424
rect 38702 361 38708 364
rect 38632 355 38708 361
rect 41064 361 41070 426
rect 41134 424 41140 426
rect 41134 364 41380 424
rect 41134 361 41140 364
rect 41064 355 41140 361
rect 1080 -204 1140 36
rect 3512 -204 3572 36
rect 5944 -204 6004 36
rect 8376 -204 8436 36
rect 10808 -204 10868 36
rect 13240 -204 13300 36
rect 15672 -204 15732 36
rect 18104 -204 18164 36
rect 20536 -204 20596 36
rect 22968 -204 23028 36
rect 25400 -204 25460 36
rect 27832 -204 27892 36
rect 30264 -204 30324 36
rect 32696 -204 32756 36
rect 35128 -204 35188 36
rect 37560 -204 37620 36
rect 39992 -204 40052 36
rect 42424 -204 42484 36
rect 1072 -210 1149 -204
rect 1072 -274 1078 -210
rect 1143 -274 1149 -210
rect 1072 -280 1149 -274
rect 3504 -210 3581 -204
rect 3504 -274 3510 -210
rect 3575 -274 3581 -210
rect 3504 -280 3581 -274
rect 5936 -210 6013 -204
rect 5936 -274 5942 -210
rect 6007 -274 6013 -210
rect 5936 -280 6013 -274
rect 8368 -210 8445 -204
rect 8368 -274 8374 -210
rect 8439 -274 8445 -210
rect 8368 -280 8445 -274
rect 10800 -210 10877 -204
rect 10800 -274 10806 -210
rect 10871 -274 10877 -210
rect 10800 -280 10877 -274
rect 13232 -210 13309 -204
rect 13232 -274 13238 -210
rect 13303 -274 13309 -210
rect 13232 -280 13309 -274
rect 15664 -210 15741 -204
rect 15664 -274 15670 -210
rect 15735 -274 15741 -210
rect 15664 -280 15741 -274
rect 18096 -210 18173 -204
rect 18096 -274 18102 -210
rect 18167 -274 18173 -210
rect 18096 -280 18173 -274
rect 20528 -210 20605 -204
rect 20528 -274 20534 -210
rect 20599 -274 20605 -210
rect 20528 -280 20605 -274
rect 22960 -210 23037 -204
rect 22960 -274 22966 -210
rect 23031 -274 23037 -210
rect 22960 -280 23037 -274
rect 25392 -210 25469 -204
rect 25392 -274 25398 -210
rect 25463 -274 25469 -210
rect 25392 -280 25469 -274
rect 27824 -210 27901 -204
rect 27824 -274 27830 -210
rect 27895 -274 27901 -210
rect 27824 -280 27901 -274
rect 30256 -210 30333 -204
rect 30256 -274 30262 -210
rect 30327 -274 30333 -210
rect 30256 -280 30333 -274
rect 32688 -210 32765 -204
rect 32688 -274 32694 -210
rect 32759 -274 32765 -210
rect 32688 -280 32765 -274
rect 35120 -210 35197 -204
rect 35120 -274 35126 -210
rect 35191 -274 35197 -210
rect 35120 -280 35197 -274
rect 37552 -210 37629 -204
rect 37552 -274 37558 -210
rect 37623 -274 37629 -210
rect 37552 -280 37629 -274
rect 39984 -210 40061 -204
rect 39984 -274 39990 -210
rect 40055 -274 40061 -210
rect 39984 -280 40061 -274
rect 42416 -210 42493 -204
rect 42416 -274 42422 -210
rect 42487 -274 42493 -210
rect 42416 -280 42493 -274
<< via3 >>
rect 7281 44756 7345 44820
rect 11225 44628 11289 44692
rect 15169 44500 15233 44564
rect 19113 44372 19177 44436
rect 23057 44244 23121 44308
rect 27001 44116 27065 44180
rect 361 43244 426 43308
rect 2793 43244 2858 43308
rect 5225 43244 5290 43308
rect 7657 43244 7722 43308
rect 10089 43244 10154 43308
rect 12521 43244 12586 43308
rect 14953 43244 15018 43308
rect 17385 43244 17450 43308
rect 19817 43244 19882 43308
rect 22249 43244 22314 43308
rect 24681 43244 24746 43308
rect 30945 43988 31009 44052
rect 34889 43860 34953 43924
rect 27113 43244 27178 43308
rect 29545 43244 29610 43308
rect 31977 43244 32042 43308
rect 34409 43244 34474 43308
rect 36841 43244 36906 43308
rect 39273 43244 39338 43308
rect 41705 43244 41770 43308
rect 1714 42608 1778 42673
rect 4146 42608 4210 42673
rect 6578 42608 6642 42673
rect 9010 42608 9074 42673
rect 11442 42608 11506 42673
rect 13874 42608 13938 42673
rect 16306 42608 16370 42673
rect 18738 42608 18802 42673
rect 21170 42608 21234 42673
rect 23602 42608 23666 42673
rect 26034 42608 26098 42673
rect 28466 42608 28530 42673
rect 30898 42608 30962 42673
rect 33330 42608 33394 42673
rect 35762 42608 35826 42673
rect 38194 42608 38258 42673
rect 40626 42608 40690 42673
rect 43058 42608 43122 42673
rect -274 41891 -210 41956
rect 2158 41891 2222 41956
rect 4590 41891 4654 41956
rect 7022 41891 7086 41956
rect 9454 41891 9518 41956
rect 11886 41891 11950 41956
rect 14318 41891 14382 41956
rect 16750 41891 16814 41956
rect 19182 41891 19246 41956
rect 21614 41891 21678 41956
rect 24046 41891 24110 41956
rect 26478 41891 26542 41956
rect 28910 41891 28974 41956
rect 31342 41891 31406 41956
rect 33774 41891 33838 41956
rect 36206 41891 36270 41956
rect 38638 41891 38702 41956
rect 41070 41891 41134 41956
rect 1078 41256 1143 41320
rect 3510 41256 3575 41320
rect 5942 41256 6007 41320
rect 8374 41256 8439 41320
rect 10806 41256 10871 41320
rect 13238 41256 13303 41320
rect 15670 41256 15735 41320
rect 18102 41256 18167 41320
rect 20534 41256 20599 41320
rect 22966 41256 23031 41320
rect 25398 41256 25463 41320
rect 27830 41256 27895 41320
rect 30262 41256 30327 41320
rect 32694 41256 32759 41320
rect 35126 41256 35191 41320
rect 37558 41256 37623 41320
rect 39990 41256 40055 41320
rect 42422 41256 42487 41320
rect -626 40941 -562 41005
rect 361 40812 426 40876
rect 41705 40812 41770 40876
rect 1714 40176 1778 40241
rect 43058 40176 43122 40241
rect -274 39459 -210 39524
rect 41070 39459 41134 39524
rect 1078 38824 1143 38888
rect 2794 38695 2858 38759
rect 7658 38695 7722 38759
rect 12522 38695 12586 38759
rect 17386 38695 17450 38759
rect 22250 38695 22314 38759
rect 27114 38695 27178 38759
rect 31978 38695 32042 38759
rect 36842 38695 36906 38759
rect 42422 38824 42487 38888
rect 43410 38695 43474 38759
rect 361 38380 426 38444
rect 2794 38380 2858 38444
rect 7658 38380 7722 38444
rect 12522 38380 12586 38444
rect 17386 38380 17450 38444
rect 22250 38380 22314 38444
rect 27114 38380 27178 38444
rect 31978 38380 32042 38444
rect 36842 38380 36906 38444
rect 41705 38380 41770 38444
rect 1714 37744 1778 37809
rect 43058 37744 43122 37809
rect -274 37027 -210 37092
rect 41070 37027 41134 37092
rect 1078 36392 1143 36456
rect 42422 36392 42487 36456
rect 43534 36263 43598 36327
rect -626 36077 -562 36141
rect 361 35948 426 36012
rect 41705 35948 41770 36012
rect 1714 35312 1778 35377
rect 43058 35312 43122 35377
rect -274 34595 -210 34660
rect 41070 34595 41134 34660
rect 1078 33960 1143 34024
rect 2794 33831 2858 33895
rect 7658 33831 7722 33895
rect 12522 33831 12586 33895
rect 17386 33831 17450 33895
rect 22250 33831 22314 33895
rect 27114 33831 27178 33895
rect 31978 33831 32042 33895
rect 36842 33831 36906 33895
rect 42422 33960 42487 34024
rect 43410 33831 43474 33895
rect 361 33516 426 33580
rect 2794 33516 2858 33580
rect 7658 33516 7722 33580
rect 12522 33516 12586 33580
rect 17386 33516 17450 33580
rect 22250 33516 22314 33580
rect 27114 33516 27178 33580
rect 31978 33516 32042 33580
rect 36842 33516 36906 33580
rect 41705 33516 41770 33580
rect 1714 32880 1778 32945
rect 43058 32880 43122 32945
rect -274 32163 -210 32228
rect 41070 32163 41134 32228
rect 1078 31528 1143 31592
rect 42422 31528 42487 31592
rect 43534 31399 43598 31463
rect -626 31213 -562 31277
rect 361 31084 426 31148
rect 41705 31084 41770 31148
rect 1714 30448 1778 30513
rect 43058 30448 43122 30513
rect -274 29731 -210 29796
rect 41070 29731 41134 29796
rect 1078 29096 1143 29160
rect 2794 28967 2858 29031
rect 7658 28967 7722 29031
rect 12522 28967 12586 29031
rect 17386 28967 17450 29031
rect 22250 28967 22314 29031
rect 27114 28967 27178 29031
rect 31978 28967 32042 29031
rect 36842 28967 36906 29031
rect 42422 29096 42487 29160
rect 43410 28967 43474 29031
rect 361 28652 426 28716
rect 2794 28652 2858 28716
rect 7658 28652 7722 28716
rect 12522 28652 12586 28716
rect 17386 28652 17450 28716
rect 22250 28652 22314 28716
rect 27114 28652 27178 28716
rect 31978 28652 32042 28716
rect 36842 28652 36906 28716
rect 43658 28781 43722 28845
rect 41705 28652 41770 28716
rect 1714 28016 1778 28081
rect 43058 28016 43122 28081
rect -274 27299 -210 27364
rect 41070 27299 41134 27364
rect 1078 26664 1143 26728
rect -750 26535 -686 26599
rect 42422 26664 42487 26728
rect -626 26349 -562 26413
rect 361 26220 426 26284
rect 41705 26220 41770 26284
rect 1714 25584 1778 25649
rect 43058 25584 43122 25649
rect -274 24867 -210 24932
rect 41070 24867 41134 24932
rect 1078 24232 1143 24296
rect 2794 24103 2858 24167
rect 7658 24103 7722 24167
rect 12522 24103 12586 24167
rect 17386 24103 17450 24167
rect 22250 24103 22314 24167
rect 27114 24103 27178 24167
rect 31978 24103 32042 24167
rect 36842 24103 36906 24167
rect 42422 24232 42487 24296
rect 43410 24103 43474 24167
rect -750 23917 -686 23981
rect 361 23788 426 23852
rect 2794 23788 2858 23852
rect 7658 23788 7722 23852
rect 12522 23788 12586 23852
rect 17386 23788 17450 23852
rect 22250 23788 22314 23852
rect 27114 23788 27178 23852
rect 31978 23788 32042 23852
rect 36842 23788 36906 23852
rect 41705 23788 41770 23852
rect 1714 23152 1778 23217
rect 43058 23152 43122 23217
rect -274 22435 -210 22500
rect 41070 22435 41134 22500
rect 1078 21800 1143 21864
rect 10806 21799 10870 21864
rect 12522 21671 12586 21735
rect 39990 21799 40054 21864
rect 42422 21800 42487 21864
rect 43782 21671 43846 21735
rect -998 21485 -934 21549
rect 22250 21485 22314 21549
rect -874 21299 -810 21363
rect 361 21170 426 21234
rect 10806 21299 10870 21364
rect 12522 21170 12586 21234
rect 22250 21170 22314 21234
rect 39990 21299 40054 21364
rect 41705 21170 41770 21234
rect 1714 20534 1778 20599
rect 43058 20534 43122 20599
rect -274 19817 -210 19882
rect 41070 19817 41134 19882
rect 1078 19182 1143 19246
rect 5942 19181 6006 19246
rect -750 19053 -686 19117
rect 10806 19181 10870 19246
rect 15670 19181 15734 19246
rect 20534 19181 20598 19246
rect 25398 19181 25462 19246
rect 30262 19181 30326 19246
rect 35126 19181 35190 19246
rect 39990 19181 40054 19246
rect 42422 19182 42487 19246
rect 361 18738 426 18802
rect 5942 18867 6006 18932
rect 10806 18867 10870 18932
rect 15670 18867 15734 18932
rect 20534 18867 20598 18932
rect 25398 18867 25462 18932
rect 30262 18867 30326 18932
rect 35126 18867 35190 18932
rect 39990 18867 40054 18932
rect 43410 18867 43474 18931
rect 41705 18738 41770 18802
rect 1714 18102 1778 18167
rect 43058 18102 43122 18167
rect -274 17385 -210 17450
rect 41070 17385 41134 17450
rect 1078 16750 1143 16814
rect -626 16621 -562 16685
rect 42422 16750 42487 16814
rect -750 16435 -686 16499
rect 361 16306 426 16370
rect 41705 16306 41770 16370
rect 1714 15670 1778 15735
rect 43058 15670 43122 15735
rect -274 14953 -210 15018
rect 41070 14953 41134 15018
rect 1078 14318 1143 14382
rect 5942 14317 6006 14382
rect 10806 14317 10870 14382
rect 15670 14317 15734 14382
rect 20534 14317 20598 14382
rect 25398 14317 25462 14382
rect 30262 14317 30326 14382
rect 35126 14317 35190 14382
rect 39990 14317 40054 14382
rect 42422 14318 42487 14382
rect 43658 14189 43722 14253
rect 361 13874 426 13938
rect 5942 14003 6006 14068
rect 10806 14003 10870 14068
rect 15670 14003 15734 14068
rect 20534 14003 20598 14068
rect 25398 14003 25462 14068
rect 30262 14003 30326 14068
rect 35126 14003 35190 14068
rect 39990 14003 40054 14068
rect 43410 14003 43474 14067
rect 41705 13874 41770 13938
rect 1714 13238 1778 13303
rect 43058 13238 43122 13303
rect -274 12521 -210 12586
rect 41070 12521 41134 12586
rect 1078 11886 1143 11950
rect -626 11757 -562 11821
rect 42422 11886 42487 11950
rect 361 11442 426 11506
rect 43534 11571 43598 11635
rect 41705 11442 41770 11506
rect 1714 10806 1778 10871
rect 43058 10806 43122 10871
rect -274 10089 -210 10154
rect 41070 10089 41134 10154
rect 1078 9454 1143 9518
rect 5942 9453 6006 9518
rect 10806 9453 10870 9518
rect 15670 9453 15734 9518
rect 20534 9453 20598 9518
rect 25398 9453 25462 9518
rect 30262 9453 30326 9518
rect 35126 9453 35190 9518
rect 39990 9453 40054 9518
rect 42422 9454 42487 9518
rect 361 9010 426 9074
rect 5942 9139 6006 9204
rect 10806 9139 10870 9204
rect 15670 9139 15734 9204
rect 20534 9139 20598 9204
rect 25398 9139 25462 9204
rect 30262 9139 30326 9204
rect 35126 9139 35190 9204
rect 39990 9139 40054 9204
rect 43410 9139 43474 9203
rect 41705 9010 41770 9074
rect 1714 8374 1778 8439
rect 43058 8374 43122 8439
rect -274 7657 -210 7722
rect 41070 7657 41134 7722
rect 1078 7022 1143 7086
rect -626 6893 -562 6957
rect 42422 7022 42487 7086
rect 361 6578 426 6642
rect 43534 6707 43598 6771
rect 41705 6578 41770 6642
rect 1714 5942 1778 6007
rect 43058 5942 43122 6007
rect -274 5225 -210 5290
rect 41070 5225 41134 5290
rect 1078 4590 1143 4654
rect 5942 4589 6006 4654
rect 10806 4589 10870 4654
rect 15670 4589 15734 4654
rect 20534 4589 20598 4654
rect 25398 4589 25462 4654
rect 30262 4589 30326 4654
rect 35126 4589 35190 4654
rect 39990 4589 40054 4654
rect 42422 4590 42487 4654
rect 361 4146 426 4210
rect 5942 4275 6006 4340
rect 10806 4275 10870 4340
rect 15670 4275 15734 4340
rect 20534 4275 20598 4340
rect 25398 4275 25462 4340
rect 30262 4275 30326 4340
rect 35126 4275 35190 4340
rect 39990 4275 40054 4340
rect 43410 4275 43474 4340
rect 41705 4146 41770 4210
rect 1714 3510 1778 3575
rect 43058 3510 43122 3575
rect -274 2793 -210 2858
rect 41070 2793 41134 2858
rect 1078 2158 1143 2222
rect -626 2029 -562 2093
rect 42422 2158 42487 2222
rect 361 1714 426 1778
rect 2793 1714 2858 1778
rect 5225 1714 5290 1778
rect 7657 1714 7722 1778
rect 10089 1714 10154 1778
rect 12521 1714 12586 1778
rect 14953 1714 15018 1778
rect 17385 1714 17450 1778
rect 19817 1714 19882 1778
rect 22249 1714 22314 1778
rect 24681 1714 24746 1778
rect 27113 1714 27178 1778
rect 29545 1714 29610 1778
rect 31977 1714 32042 1778
rect 34409 1714 34474 1778
rect 36841 1714 36906 1778
rect 39273 1714 39338 1778
rect 41705 1714 41770 1778
rect 1714 1078 1778 1143
rect 4146 1078 4210 1143
rect 6578 1078 6642 1143
rect 9010 1078 9074 1143
rect 11442 1078 11506 1143
rect 13874 1078 13938 1143
rect 16306 1078 16370 1143
rect 18738 1078 18802 1143
rect 21170 1078 21234 1143
rect 23602 1078 23666 1143
rect 26034 1078 26098 1143
rect 28466 1078 28530 1143
rect 30898 1078 30962 1143
rect 33330 1078 33394 1143
rect 35762 1078 35826 1143
rect 38194 1078 38258 1143
rect 40626 1078 40690 1143
rect 43058 1078 43122 1143
rect -274 361 -210 426
rect 2158 361 2222 426
rect 4590 361 4654 426
rect 7022 361 7086 426
rect 9454 361 9518 426
rect 11886 361 11950 426
rect 14318 361 14382 426
rect 16750 361 16814 426
rect 19182 361 19246 426
rect 21614 361 21678 426
rect 24046 361 24110 426
rect 26478 361 26542 426
rect 28910 361 28974 426
rect 31342 361 31406 426
rect 33774 361 33838 426
rect 36206 361 36270 426
rect 38638 361 38702 426
rect 41070 361 41134 426
rect 1078 -274 1143 -210
rect 3510 -274 3575 -210
rect 5942 -274 6007 -210
rect 8374 -274 8439 -210
rect 10806 -274 10871 -210
rect 13238 -274 13303 -210
rect 15670 -274 15735 -210
rect 18102 -274 18167 -210
rect 20534 -274 20599 -210
rect 22966 -274 23031 -210
rect 25398 -274 25463 -210
rect 27830 -274 27895 -210
rect 30262 -274 30327 -210
rect 32694 -274 32759 -210
rect 35126 -274 35191 -210
rect 37558 -274 37623 -210
rect 39990 -274 40055 -210
rect 42422 -274 42487 -210
<< metal4 >>
rect 7280 44820 7346 44821
rect 7280 44818 7281 44820
rect -996 44758 7281 44818
rect -996 21550 -936 44758
rect 7280 44756 7281 44758
rect 7345 44756 7346 44820
rect 7280 44755 7346 44756
rect 11224 44692 11290 44693
rect 11224 44628 11225 44692
rect 11289 44690 11290 44692
rect 11289 44630 43844 44690
rect 11289 44628 11290 44630
rect 11224 44627 11290 44628
rect 15168 44564 15234 44565
rect 15168 44562 15169 44564
rect -872 44502 15169 44562
rect -999 21549 -933 21550
rect -999 21485 -998 21549
rect -934 21485 -933 21549
rect -999 21484 -933 21485
rect -872 21364 -812 44502
rect 15168 44500 15169 44502
rect 15233 44500 15234 44564
rect 15168 44499 15234 44500
rect 19112 44436 19178 44437
rect 19112 44372 19113 44436
rect 19177 44434 19178 44436
rect 19177 44374 43720 44434
rect 19177 44372 19178 44374
rect 19112 44371 19178 44372
rect 23056 44308 23122 44309
rect 23056 44306 23057 44308
rect -748 44246 23057 44306
rect -748 26600 -688 44246
rect 23056 44244 23057 44246
rect 23121 44244 23122 44308
rect 23056 44243 23122 44244
rect 27000 44180 27066 44181
rect 27000 44116 27001 44180
rect 27065 44178 27066 44180
rect 27065 44118 43596 44178
rect 27065 44116 27066 44118
rect 27000 44115 27066 44116
rect 30944 44052 31010 44053
rect 30944 44050 30945 44052
rect -624 43990 30945 44050
rect -624 41006 -564 43990
rect 30944 43988 30945 43990
rect 31009 43988 31010 44052
rect 30944 43987 31010 43988
rect 34888 43924 34954 43925
rect 34888 43860 34889 43924
rect 34953 43922 34954 43924
rect 34953 43862 43472 43922
rect 34953 43860 34954 43862
rect 34888 43859 34954 43860
rect 360 43308 427 43309
rect 360 43244 361 43308
rect 426 43306 427 43308
rect 722 43306 782 43430
rect 426 43246 782 43306
rect 426 43244 427 43246
rect 360 43243 427 43244
rect 722 42931 782 43246
rect 2792 43308 2859 43309
rect 2792 43244 2793 43308
rect 2858 43306 2859 43308
rect 5224 43308 5291 43309
rect 2858 43246 3214 43306
rect 2858 43244 2859 43246
rect 2792 43243 2859 43244
rect 3154 42931 3214 43246
rect 5224 43244 5225 43308
rect 5290 43306 5291 43308
rect 7656 43308 7723 43309
rect 5290 43246 5646 43306
rect 5290 43244 5291 43246
rect 5224 43243 5291 43244
rect 5586 42931 5646 43246
rect 7656 43244 7657 43308
rect 7722 43306 7723 43308
rect 10088 43308 10155 43309
rect 7722 43246 8078 43306
rect 7722 43244 7723 43246
rect 7656 43243 7723 43244
rect 8018 42931 8078 43246
rect 10088 43244 10089 43308
rect 10154 43306 10155 43308
rect 12520 43308 12587 43309
rect 10154 43246 10510 43306
rect 10154 43244 10155 43246
rect 10088 43243 10155 43244
rect 10450 42931 10510 43246
rect 12520 43244 12521 43308
rect 12586 43306 12587 43308
rect 14952 43308 15019 43309
rect 12586 43246 12942 43306
rect 12586 43244 12587 43246
rect 12520 43243 12587 43244
rect 12882 42931 12942 43246
rect 14952 43244 14953 43308
rect 15018 43306 15019 43308
rect 17384 43308 17451 43309
rect 15018 43246 15374 43306
rect 15018 43244 15019 43246
rect 14952 43243 15019 43244
rect 15314 42931 15374 43246
rect 17384 43244 17385 43308
rect 17450 43306 17451 43308
rect 19816 43308 19883 43309
rect 17450 43246 17806 43306
rect 17450 43244 17451 43246
rect 17384 43243 17451 43244
rect 17746 42931 17806 43246
rect 19816 43244 19817 43308
rect 19882 43306 19883 43308
rect 22248 43308 22315 43309
rect 19882 43246 20238 43306
rect 19882 43244 19883 43246
rect 19816 43243 19883 43244
rect 20178 42931 20238 43246
rect 22248 43244 22249 43308
rect 22314 43306 22315 43308
rect 24680 43308 24747 43309
rect 22314 43246 22670 43306
rect 22314 43244 22315 43246
rect 22248 43243 22315 43244
rect 22610 42931 22670 43246
rect 24680 43244 24681 43308
rect 24746 43306 24747 43308
rect 27112 43308 27179 43309
rect 24746 43246 25102 43306
rect 24746 43244 24747 43246
rect 24680 43243 24747 43244
rect 25042 42931 25102 43246
rect 27112 43244 27113 43308
rect 27178 43306 27179 43308
rect 29544 43308 29611 43309
rect 27178 43246 27534 43306
rect 27178 43244 27179 43246
rect 27112 43243 27179 43244
rect 27474 42931 27534 43246
rect 29544 43244 29545 43308
rect 29610 43306 29611 43308
rect 31976 43308 32043 43309
rect 29610 43246 29966 43306
rect 29610 43244 29611 43246
rect 29544 43243 29611 43244
rect 29906 42931 29966 43246
rect 31976 43244 31977 43308
rect 32042 43306 32043 43308
rect 34408 43308 34475 43309
rect 32042 43246 32398 43306
rect 32042 43244 32043 43246
rect 31976 43243 32043 43244
rect 32338 42931 32398 43246
rect 34408 43244 34409 43308
rect 34474 43306 34475 43308
rect 36840 43308 36907 43309
rect 34474 43246 34830 43306
rect 34474 43244 34475 43246
rect 34408 43243 34475 43244
rect 34770 42931 34830 43246
rect 36840 43244 36841 43308
rect 36906 43306 36907 43308
rect 39272 43308 39339 43309
rect 36906 43246 37262 43306
rect 36906 43244 36907 43246
rect 36840 43243 36907 43244
rect 37202 42931 37262 43246
rect 39272 43244 39273 43308
rect 39338 43306 39339 43308
rect 41704 43308 41771 43309
rect 39338 43246 39694 43306
rect 39338 43244 39339 43246
rect 39272 43243 39339 43244
rect 39634 42931 39694 43246
rect 41704 43244 41705 43308
rect 41770 43306 41771 43308
rect 42066 43306 42126 43404
rect 41770 43246 42126 43306
rect 41770 43244 41771 43246
rect 41704 43243 41771 43244
rect 42066 42931 42126 43246
rect 1713 42673 1779 42674
rect 1713 42608 1714 42673
rect 1778 42608 1779 42673
rect 1713 42607 1779 42608
rect 4145 42673 4211 42674
rect 4145 42608 4146 42673
rect 4210 42608 4211 42673
rect 4145 42607 4211 42608
rect 6577 42673 6643 42674
rect 6577 42608 6578 42673
rect 6642 42608 6643 42673
rect 6577 42607 6643 42608
rect 9009 42673 9075 42674
rect 9009 42608 9010 42673
rect 9074 42608 9075 42673
rect 9009 42607 9075 42608
rect 11441 42673 11507 42674
rect 11441 42608 11442 42673
rect 11506 42608 11507 42673
rect 11441 42607 11507 42608
rect 13873 42673 13939 42674
rect 13873 42608 13874 42673
rect 13938 42608 13939 42673
rect 13873 42607 13939 42608
rect 16305 42673 16371 42674
rect 16305 42608 16306 42673
rect 16370 42608 16371 42673
rect 16305 42607 16371 42608
rect 18737 42673 18803 42674
rect 18737 42608 18738 42673
rect 18802 42608 18803 42673
rect 18737 42607 18803 42608
rect 21169 42673 21235 42674
rect 21169 42608 21170 42673
rect 21234 42608 21235 42673
rect 21169 42607 21235 42608
rect 23601 42673 23667 42674
rect 23601 42608 23602 42673
rect 23666 42608 23667 42673
rect 23601 42607 23667 42608
rect 26033 42673 26099 42674
rect 26033 42608 26034 42673
rect 26098 42608 26099 42673
rect 26033 42607 26099 42608
rect 28465 42673 28531 42674
rect 28465 42608 28466 42673
rect 28530 42608 28531 42673
rect 28465 42607 28531 42608
rect 30897 42673 30963 42674
rect 30897 42608 30898 42673
rect 30962 42608 30963 42673
rect 30897 42607 30963 42608
rect 33329 42673 33395 42674
rect 33329 42608 33330 42673
rect 33394 42608 33395 42673
rect 33329 42607 33395 42608
rect 35761 42673 35827 42674
rect 35761 42608 35762 42673
rect 35826 42608 35827 42673
rect 35761 42607 35827 42608
rect 38193 42673 38259 42674
rect 38193 42608 38194 42673
rect 38258 42608 38259 42673
rect 38193 42607 38259 42608
rect 40625 42673 40691 42674
rect 40625 42608 40626 42673
rect 40690 42608 40691 42673
rect 40625 42607 40691 42608
rect 43057 42673 43123 42674
rect 43057 42608 43058 42673
rect 43122 42608 43123 42673
rect 43057 42607 43123 42608
rect 1716 42312 1776 42607
rect 4148 42312 4208 42607
rect 6580 42312 6640 42607
rect 9012 42312 9072 42607
rect 11444 42312 11504 42607
rect 13876 42312 13936 42607
rect 16308 42312 16368 42607
rect 18740 42312 18800 42607
rect 21172 42312 21232 42607
rect 23604 42312 23664 42607
rect 26036 42312 26096 42607
rect 28468 42312 28528 42607
rect 30900 42312 30960 42607
rect 33332 42312 33392 42607
rect 35764 42312 35824 42607
rect 38196 42312 38256 42607
rect 40628 42312 40688 42607
rect 43060 42312 43120 42607
rect -272 42252 103 42312
rect 1401 42252 2535 42312
rect 3833 42252 4967 42312
rect 6265 42252 7399 42312
rect 8697 42252 9831 42312
rect 11129 42252 12263 42312
rect 13561 42252 14695 42312
rect 15993 42252 17127 42312
rect 18425 42252 19559 42312
rect 20857 42252 21991 42312
rect 23289 42252 24423 42312
rect 25721 42252 26855 42312
rect 28153 42252 29287 42312
rect 30585 42252 31719 42312
rect 33017 42252 34151 42312
rect 35449 42252 36583 42312
rect 37881 42252 39015 42312
rect 40313 42252 41447 42312
rect 42745 42252 43120 42312
rect -272 41957 -212 42252
rect 2160 41957 2220 42252
rect 4592 41957 4652 42252
rect 7024 41957 7084 42252
rect 9456 41957 9516 42252
rect 11888 41957 11948 42252
rect 14320 41957 14380 42252
rect 16752 41957 16812 42252
rect 19184 41957 19244 42252
rect 21616 41957 21676 42252
rect 24048 41957 24108 42252
rect 26480 41957 26540 42252
rect 28912 41957 28972 42252
rect 31344 41957 31404 42252
rect 33776 41957 33836 42252
rect 36208 41957 36268 42252
rect 38640 41957 38700 42252
rect 41072 41957 41132 42252
rect -275 41956 -209 41957
rect -275 41891 -274 41956
rect -210 41891 -209 41956
rect -275 41890 -209 41891
rect 2157 41956 2223 41957
rect 2157 41891 2158 41956
rect 2222 41891 2223 41956
rect 2157 41890 2223 41891
rect 4589 41956 4655 41957
rect 4589 41891 4590 41956
rect 4654 41891 4655 41956
rect 4589 41890 4655 41891
rect 7021 41956 7087 41957
rect 7021 41891 7022 41956
rect 7086 41891 7087 41956
rect 7021 41890 7087 41891
rect 9453 41956 9519 41957
rect 9453 41891 9454 41956
rect 9518 41891 9519 41956
rect 9453 41890 9519 41891
rect 11885 41956 11951 41957
rect 11885 41891 11886 41956
rect 11950 41891 11951 41956
rect 11885 41890 11951 41891
rect 14317 41956 14383 41957
rect 14317 41891 14318 41956
rect 14382 41891 14383 41956
rect 14317 41890 14383 41891
rect 16749 41956 16815 41957
rect 16749 41891 16750 41956
rect 16814 41891 16815 41956
rect 16749 41890 16815 41891
rect 19181 41956 19247 41957
rect 19181 41891 19182 41956
rect 19246 41891 19247 41956
rect 19181 41890 19247 41891
rect 21613 41956 21679 41957
rect 21613 41891 21614 41956
rect 21678 41891 21679 41956
rect 21613 41890 21679 41891
rect 24045 41956 24111 41957
rect 24045 41891 24046 41956
rect 24110 41891 24111 41956
rect 24045 41890 24111 41891
rect 26477 41956 26543 41957
rect 26477 41891 26478 41956
rect 26542 41891 26543 41956
rect 26477 41890 26543 41891
rect 28909 41956 28975 41957
rect 28909 41891 28910 41956
rect 28974 41891 28975 41956
rect 28909 41890 28975 41891
rect 31341 41956 31407 41957
rect 31341 41891 31342 41956
rect 31406 41891 31407 41956
rect 31341 41890 31407 41891
rect 33773 41956 33839 41957
rect 33773 41891 33774 41956
rect 33838 41891 33839 41956
rect 33773 41890 33839 41891
rect 36205 41956 36271 41957
rect 36205 41891 36206 41956
rect 36270 41891 36271 41956
rect 36205 41890 36271 41891
rect 38637 41956 38703 41957
rect 38637 41891 38638 41956
rect 38702 41891 38703 41956
rect 38637 41890 38703 41891
rect 41069 41956 41135 41957
rect 41069 41891 41070 41956
rect 41134 41891 41135 41956
rect 41069 41890 41135 41891
rect 722 41318 782 41633
rect 1077 41320 1144 41321
rect 1077 41318 1078 41320
rect 722 41258 1078 41318
rect -627 41005 -561 41006
rect -627 40941 -626 41005
rect -562 40941 -561 41005
rect -627 40940 -561 40941
rect -624 36142 -564 40940
rect 360 40876 427 40877
rect 360 40812 361 40876
rect 426 40874 427 40876
rect 722 40874 782 41258
rect 1077 41256 1078 41258
rect 1143 41256 1144 41320
rect 3154 41318 3214 41633
rect 3509 41320 3576 41321
rect 3509 41318 3510 41320
rect 3154 41258 3510 41318
rect 1077 41255 1144 41256
rect 3509 41256 3510 41258
rect 3575 41256 3576 41320
rect 5586 41318 5646 41633
rect 5941 41320 6008 41321
rect 5941 41318 5942 41320
rect 5586 41258 5942 41318
rect 3509 41255 3576 41256
rect 5941 41256 5942 41258
rect 6007 41256 6008 41320
rect 8018 41318 8078 41633
rect 8373 41320 8440 41321
rect 8373 41318 8374 41320
rect 8018 41258 8374 41318
rect 5941 41255 6008 41256
rect 8373 41256 8374 41258
rect 8439 41256 8440 41320
rect 10450 41318 10510 41633
rect 10805 41320 10872 41321
rect 10805 41318 10806 41320
rect 10450 41258 10806 41318
rect 8373 41255 8440 41256
rect 10805 41256 10806 41258
rect 10871 41256 10872 41320
rect 12882 41318 12942 41633
rect 13237 41320 13304 41321
rect 13237 41318 13238 41320
rect 12882 41258 13238 41318
rect 10805 41255 10872 41256
rect 13237 41256 13238 41258
rect 13303 41256 13304 41320
rect 15314 41318 15374 41633
rect 15669 41320 15736 41321
rect 15669 41318 15670 41320
rect 15314 41258 15670 41318
rect 13237 41255 13304 41256
rect 15669 41256 15670 41258
rect 15735 41256 15736 41320
rect 17746 41318 17806 41633
rect 18101 41320 18168 41321
rect 18101 41318 18102 41320
rect 17746 41258 18102 41318
rect 15669 41255 15736 41256
rect 18101 41256 18102 41258
rect 18167 41256 18168 41320
rect 20178 41318 20238 41633
rect 20533 41320 20600 41321
rect 20533 41318 20534 41320
rect 20178 41258 20534 41318
rect 18101 41255 18168 41256
rect 20533 41256 20534 41258
rect 20599 41256 20600 41320
rect 22610 41318 22670 41633
rect 22965 41320 23032 41321
rect 22965 41318 22966 41320
rect 22610 41258 22966 41318
rect 20533 41255 20600 41256
rect 22965 41256 22966 41258
rect 23031 41256 23032 41320
rect 25042 41318 25102 41633
rect 25397 41320 25464 41321
rect 25397 41318 25398 41320
rect 25042 41258 25398 41318
rect 22965 41255 23032 41256
rect 25397 41256 25398 41258
rect 25463 41256 25464 41320
rect 27474 41318 27534 41633
rect 27829 41320 27896 41321
rect 27829 41318 27830 41320
rect 27474 41258 27830 41318
rect 25397 41255 25464 41256
rect 27829 41256 27830 41258
rect 27895 41256 27896 41320
rect 29906 41318 29966 41633
rect 30261 41320 30328 41321
rect 30261 41318 30262 41320
rect 29906 41258 30262 41318
rect 27829 41255 27896 41256
rect 30261 41256 30262 41258
rect 30327 41256 30328 41320
rect 32338 41318 32398 41633
rect 32693 41320 32760 41321
rect 32693 41318 32694 41320
rect 32338 41258 32694 41318
rect 30261 41255 30328 41256
rect 32693 41256 32694 41258
rect 32759 41256 32760 41320
rect 34770 41318 34830 41633
rect 35125 41320 35192 41321
rect 35125 41318 35126 41320
rect 34770 41258 35126 41318
rect 32693 41255 32760 41256
rect 35125 41256 35126 41258
rect 35191 41256 35192 41320
rect 37202 41318 37262 41633
rect 37557 41320 37624 41321
rect 37557 41318 37558 41320
rect 37202 41258 37558 41318
rect 35125 41255 35192 41256
rect 37557 41256 37558 41258
rect 37623 41256 37624 41320
rect 39634 41318 39694 41633
rect 39989 41320 40056 41321
rect 39989 41318 39990 41320
rect 39634 41258 39990 41318
rect 37557 41255 37624 41256
rect 39989 41256 39990 41258
rect 40055 41256 40056 41320
rect 39989 41255 40056 41256
rect 42066 41318 42126 41633
rect 42421 41320 42488 41321
rect 42421 41318 42422 41320
rect 42066 41258 42422 41318
rect 426 40814 782 40874
rect 426 40812 427 40814
rect 360 40811 427 40812
rect 722 40499 782 40814
rect 41704 40876 41771 40877
rect 41704 40812 41705 40876
rect 41770 40874 41771 40876
rect 42066 40874 42126 41258
rect 42421 41256 42422 41258
rect 42487 41256 42488 41320
rect 42421 41255 42488 41256
rect 41770 40814 42126 40874
rect 41770 40812 41771 40814
rect 41704 40811 41771 40812
rect 1713 40241 1779 40242
rect 1713 40176 1714 40241
rect 1778 40176 1779 40241
rect 1713 40175 1779 40176
rect 1716 39880 1776 40175
rect 3154 39880 3214 40603
rect 5586 39880 5646 40603
rect 8018 39880 8078 40603
rect 10450 39880 10510 40603
rect 12882 39880 12942 40603
rect 15314 39880 15374 40603
rect 17746 39880 17806 40603
rect 20178 39880 20238 40603
rect 22610 39880 22670 40603
rect 25042 39880 25102 40603
rect 27474 39880 27534 40603
rect 29906 39880 29966 40603
rect 32338 39880 32398 40603
rect 34770 39880 34830 40603
rect 37202 39880 37262 40603
rect 39634 39880 39694 40603
rect -272 39820 103 39880
rect 1401 39820 1776 39880
rect 2432 39820 40416 39880
rect 41072 39820 41447 39880
rect -272 39525 -212 39820
rect -275 39524 -209 39525
rect -275 39459 -274 39524
rect -210 39459 -209 39524
rect -275 39458 -209 39459
rect 722 38886 782 39201
rect 1077 38888 1144 38889
rect 1077 38886 1078 38888
rect 722 38826 1078 38886
rect 360 38444 427 38445
rect 360 38380 361 38444
rect 426 38442 427 38444
rect 722 38442 782 38826
rect 1077 38824 1078 38826
rect 1143 38824 1144 38888
rect 1077 38823 1144 38824
rect 2793 38759 2859 38760
rect 2793 38695 2794 38759
rect 2858 38695 2859 38759
rect 2793 38694 2859 38695
rect 2796 38445 2856 38694
rect 426 38382 782 38442
rect 426 38380 427 38382
rect 360 38379 427 38380
rect 722 38067 782 38382
rect 2793 38444 2859 38445
rect 2793 38380 2794 38444
rect 2858 38380 2859 38444
rect 2793 38379 2859 38380
rect 1713 37809 1779 37810
rect 1713 37744 1714 37809
rect 1778 37744 1779 37809
rect 1713 37743 1779 37744
rect 1716 37448 1776 37743
rect 3154 37448 3214 39820
rect 5586 37448 5646 39820
rect 7657 38759 7723 38760
rect 7657 38695 7658 38759
rect 7722 38695 7723 38759
rect 7657 38694 7723 38695
rect 7660 38445 7720 38694
rect 7657 38444 7723 38445
rect 7657 38380 7658 38444
rect 7722 38380 7723 38444
rect 7657 38379 7723 38380
rect 8018 37448 8078 39820
rect 10450 37448 10510 39820
rect 12521 38759 12587 38760
rect 12521 38695 12522 38759
rect 12586 38695 12587 38759
rect 12521 38694 12587 38695
rect 12524 38445 12584 38694
rect 12521 38444 12587 38445
rect 12521 38380 12522 38444
rect 12586 38380 12587 38444
rect 12521 38379 12587 38380
rect 12882 37448 12942 39820
rect 15314 37448 15374 39820
rect 17385 38759 17451 38760
rect 17385 38695 17386 38759
rect 17450 38695 17451 38759
rect 17385 38694 17451 38695
rect 17388 38445 17448 38694
rect 17385 38444 17451 38445
rect 17385 38380 17386 38444
rect 17450 38380 17451 38444
rect 17385 38379 17451 38380
rect 17746 37448 17806 39820
rect 20178 37448 20238 39820
rect 22249 38759 22315 38760
rect 22249 38695 22250 38759
rect 22314 38695 22315 38759
rect 22249 38694 22315 38695
rect 22252 38445 22312 38694
rect 22249 38444 22315 38445
rect 22249 38380 22250 38444
rect 22314 38380 22315 38444
rect 22249 38379 22315 38380
rect 22610 37448 22670 39820
rect 25042 37448 25102 39820
rect 27113 38759 27179 38760
rect 27113 38695 27114 38759
rect 27178 38695 27179 38759
rect 27113 38694 27179 38695
rect 27116 38445 27176 38694
rect 27113 38444 27179 38445
rect 27113 38380 27114 38444
rect 27178 38380 27179 38444
rect 27113 38379 27179 38380
rect 27474 37448 27534 39820
rect 29906 37448 29966 39820
rect 31977 38759 32043 38760
rect 31977 38695 31978 38759
rect 32042 38695 32043 38759
rect 31977 38694 32043 38695
rect 31980 38445 32040 38694
rect 31977 38444 32043 38445
rect 31977 38380 31978 38444
rect 32042 38380 32043 38444
rect 31977 38379 32043 38380
rect 32338 37448 32398 39820
rect 34770 37448 34830 39820
rect 36841 38759 36907 38760
rect 36841 38695 36842 38759
rect 36906 38695 36907 38759
rect 36841 38694 36907 38695
rect 36844 38445 36904 38694
rect 36841 38444 36907 38445
rect 36841 38380 36842 38444
rect 36906 38380 36907 38444
rect 36841 38379 36907 38380
rect 37202 37448 37262 39820
rect 39634 37448 39694 39820
rect 41072 39525 41132 39820
rect 41069 39524 41135 39525
rect 41069 39459 41070 39524
rect 41134 39459 41135 39524
rect 41069 39458 41135 39459
rect 42066 38886 42126 40814
rect 43057 40241 43123 40242
rect 43057 40176 43058 40241
rect 43122 40176 43123 40241
rect 43057 40175 43123 40176
rect 43060 39880 43120 40175
rect 42745 39820 43120 39880
rect 42421 38888 42488 38889
rect 42421 38886 42422 38888
rect 42066 38826 42422 38886
rect 41704 38444 41771 38445
rect 41704 38380 41705 38444
rect 41770 38442 41771 38444
rect 42066 38442 42126 38826
rect 42421 38824 42422 38826
rect 42487 38824 42488 38888
rect 42421 38823 42488 38824
rect 43412 38760 43472 43862
rect 43409 38759 43475 38760
rect 43409 38695 43410 38759
rect 43474 38695 43475 38759
rect 43409 38694 43475 38695
rect 41770 38382 42126 38442
rect 41770 38380 41771 38382
rect 41704 38379 41771 38380
rect -272 37388 103 37448
rect 1401 37388 1776 37448
rect 2432 37388 40416 37448
rect 41072 37388 41447 37448
rect -272 37093 -212 37388
rect -275 37092 -209 37093
rect -275 37027 -274 37092
rect -210 37027 -209 37092
rect -275 37026 -209 37027
rect 722 36454 782 36769
rect 1077 36456 1144 36457
rect 1077 36454 1078 36456
rect 722 36394 1078 36454
rect -627 36141 -561 36142
rect -627 36077 -626 36141
rect -562 36077 -561 36141
rect -627 36076 -561 36077
rect -624 31278 -564 36076
rect 360 36012 427 36013
rect 360 35948 361 36012
rect 426 36010 427 36012
rect 722 36010 782 36394
rect 1077 36392 1078 36394
rect 1143 36392 1144 36456
rect 1077 36391 1144 36392
rect 426 35950 782 36010
rect 426 35948 427 35950
rect 360 35947 427 35948
rect 722 35635 782 35950
rect 1713 35377 1779 35378
rect 1713 35312 1714 35377
rect 1778 35312 1779 35377
rect 1713 35311 1779 35312
rect 1716 35016 1776 35311
rect 3154 35016 3214 37388
rect 5586 35016 5646 37388
rect 8018 35016 8078 37388
rect 10450 35016 10510 37388
rect 12882 35016 12942 37388
rect 15314 35016 15374 37388
rect 17746 35016 17806 37388
rect 20178 35016 20238 37388
rect 22610 35016 22670 37388
rect 25042 35016 25102 37388
rect 27474 35016 27534 37388
rect 29906 35016 29966 37388
rect 32338 35016 32398 37388
rect 34770 35016 34830 37388
rect 37202 35016 37262 37388
rect 39634 35016 39694 37388
rect 41072 37093 41132 37388
rect 41069 37092 41135 37093
rect 41069 37027 41070 37092
rect 41134 37027 41135 37092
rect 41069 37026 41135 37027
rect 42066 36454 42126 38382
rect 43057 37809 43123 37810
rect 43057 37744 43058 37809
rect 43122 37744 43123 37809
rect 43057 37743 43123 37744
rect 43060 37448 43120 37743
rect 42745 37388 43120 37448
rect 42421 36456 42488 36457
rect 42421 36454 42422 36456
rect 42066 36394 42422 36454
rect 41704 36012 41771 36013
rect 41704 35948 41705 36012
rect 41770 36010 41771 36012
rect 42066 36010 42126 36394
rect 42421 36392 42422 36394
rect 42487 36392 42488 36456
rect 42421 36391 42488 36392
rect 41770 35950 42126 36010
rect 41770 35948 41771 35950
rect 41704 35947 41771 35948
rect -272 34956 103 35016
rect 1401 34956 1776 35016
rect 2432 34956 40416 35016
rect 41072 34956 41447 35016
rect -272 34661 -212 34956
rect -275 34660 -209 34661
rect -275 34595 -274 34660
rect -210 34595 -209 34660
rect -275 34594 -209 34595
rect 722 34022 782 34337
rect 1077 34024 1144 34025
rect 1077 34022 1078 34024
rect 722 33962 1078 34022
rect 360 33580 427 33581
rect 360 33516 361 33580
rect 426 33578 427 33580
rect 722 33578 782 33962
rect 1077 33960 1078 33962
rect 1143 33960 1144 34024
rect 1077 33959 1144 33960
rect 2793 33895 2859 33896
rect 2793 33831 2794 33895
rect 2858 33831 2859 33895
rect 2793 33830 2859 33831
rect 2796 33581 2856 33830
rect 426 33518 782 33578
rect 426 33516 427 33518
rect 360 33515 427 33516
rect 722 33203 782 33518
rect 2793 33580 2859 33581
rect 2793 33516 2794 33580
rect 2858 33516 2859 33580
rect 2793 33515 2859 33516
rect 1713 32945 1779 32946
rect 1713 32880 1714 32945
rect 1778 32880 1779 32945
rect 1713 32879 1779 32880
rect 1716 32584 1776 32879
rect 3154 32584 3214 34956
rect 5586 32584 5646 34956
rect 7657 33895 7723 33896
rect 7657 33831 7658 33895
rect 7722 33831 7723 33895
rect 7657 33830 7723 33831
rect 7660 33581 7720 33830
rect 7657 33580 7723 33581
rect 7657 33516 7658 33580
rect 7722 33516 7723 33580
rect 7657 33515 7723 33516
rect 8018 32584 8078 34956
rect 10450 32584 10510 34956
rect 12521 33895 12587 33896
rect 12521 33831 12522 33895
rect 12586 33831 12587 33895
rect 12521 33830 12587 33831
rect 12524 33581 12584 33830
rect 12521 33580 12587 33581
rect 12521 33516 12522 33580
rect 12586 33516 12587 33580
rect 12521 33515 12587 33516
rect 12882 32584 12942 34956
rect 15314 32584 15374 34956
rect 17385 33895 17451 33896
rect 17385 33831 17386 33895
rect 17450 33831 17451 33895
rect 17385 33830 17451 33831
rect 17388 33581 17448 33830
rect 17385 33580 17451 33581
rect 17385 33516 17386 33580
rect 17450 33516 17451 33580
rect 17385 33515 17451 33516
rect 17746 32584 17806 34956
rect 20178 32584 20238 34956
rect 22249 33895 22315 33896
rect 22249 33831 22250 33895
rect 22314 33831 22315 33895
rect 22249 33830 22315 33831
rect 22252 33581 22312 33830
rect 22249 33580 22315 33581
rect 22249 33516 22250 33580
rect 22314 33516 22315 33580
rect 22249 33515 22315 33516
rect 22610 32584 22670 34956
rect 25042 32584 25102 34956
rect 27113 33895 27179 33896
rect 27113 33831 27114 33895
rect 27178 33831 27179 33895
rect 27113 33830 27179 33831
rect 27116 33581 27176 33830
rect 27113 33580 27179 33581
rect 27113 33516 27114 33580
rect 27178 33516 27179 33580
rect 27113 33515 27179 33516
rect 27474 32584 27534 34956
rect 29906 32584 29966 34956
rect 31977 33895 32043 33896
rect 31977 33831 31978 33895
rect 32042 33831 32043 33895
rect 31977 33830 32043 33831
rect 31980 33581 32040 33830
rect 31977 33580 32043 33581
rect 31977 33516 31978 33580
rect 32042 33516 32043 33580
rect 31977 33515 32043 33516
rect 32338 32584 32398 34956
rect 34770 32584 34830 34956
rect 36841 33895 36907 33896
rect 36841 33831 36842 33895
rect 36906 33831 36907 33895
rect 36841 33830 36907 33831
rect 36844 33581 36904 33830
rect 36841 33580 36907 33581
rect 36841 33516 36842 33580
rect 36906 33516 36907 33580
rect 36841 33515 36907 33516
rect 37202 32584 37262 34956
rect 39634 32584 39694 34956
rect 41072 34661 41132 34956
rect 41069 34660 41135 34661
rect 41069 34595 41070 34660
rect 41134 34595 41135 34660
rect 41069 34594 41135 34595
rect 42066 34022 42126 35950
rect 43057 35377 43123 35378
rect 43057 35312 43058 35377
rect 43122 35312 43123 35377
rect 43057 35311 43123 35312
rect 43060 35016 43120 35311
rect 42745 34956 43120 35016
rect 42421 34024 42488 34025
rect 42421 34022 42422 34024
rect 42066 33962 42422 34022
rect 41704 33580 41771 33581
rect 41704 33516 41705 33580
rect 41770 33578 41771 33580
rect 42066 33578 42126 33962
rect 42421 33960 42422 33962
rect 42487 33960 42488 34024
rect 42421 33959 42488 33960
rect 43412 33896 43472 38694
rect 43536 36328 43596 44118
rect 43533 36327 43599 36328
rect 43533 36263 43534 36327
rect 43598 36263 43599 36327
rect 43533 36262 43599 36263
rect 43409 33895 43475 33896
rect 43409 33831 43410 33895
rect 43474 33831 43475 33895
rect 43409 33830 43475 33831
rect 41770 33518 42126 33578
rect 41770 33516 41771 33518
rect 41704 33515 41771 33516
rect -272 32524 103 32584
rect 1401 32524 1776 32584
rect 2432 32524 40416 32584
rect 41072 32524 41447 32584
rect -272 32229 -212 32524
rect -275 32228 -209 32229
rect -275 32163 -274 32228
rect -210 32163 -209 32228
rect -275 32162 -209 32163
rect 722 31590 782 31905
rect 1077 31592 1144 31593
rect 1077 31590 1078 31592
rect 722 31530 1078 31590
rect -627 31277 -561 31278
rect -627 31213 -626 31277
rect -562 31213 -561 31277
rect -627 31212 -561 31213
rect -751 26599 -685 26600
rect -751 26535 -750 26599
rect -686 26535 -685 26599
rect -751 26534 -685 26535
rect -748 23982 -688 26534
rect -624 26414 -564 31212
rect 360 31148 427 31149
rect 360 31084 361 31148
rect 426 31146 427 31148
rect 722 31146 782 31530
rect 1077 31528 1078 31530
rect 1143 31528 1144 31592
rect 1077 31527 1144 31528
rect 426 31086 782 31146
rect 426 31084 427 31086
rect 360 31083 427 31084
rect 722 30771 782 31086
rect 1713 30513 1779 30514
rect 1713 30448 1714 30513
rect 1778 30448 1779 30513
rect 1713 30447 1779 30448
rect 1716 30152 1776 30447
rect 3154 30152 3214 32524
rect 5586 30152 5646 32524
rect 8018 30152 8078 32524
rect 10450 30152 10510 32524
rect 12882 30152 12942 32524
rect 15314 30152 15374 32524
rect 17746 30152 17806 32524
rect 20178 30152 20238 32524
rect 22610 30152 22670 32524
rect 25042 30152 25102 32524
rect 27474 30152 27534 32524
rect 29906 30152 29966 32524
rect 32338 30152 32398 32524
rect 34770 30152 34830 32524
rect 37202 30152 37262 32524
rect 39634 30152 39694 32524
rect 41072 32229 41132 32524
rect 41069 32228 41135 32229
rect 41069 32163 41070 32228
rect 41134 32163 41135 32228
rect 41069 32162 41135 32163
rect 42066 31590 42126 33518
rect 43057 32945 43123 32946
rect 43057 32880 43058 32945
rect 43122 32880 43123 32945
rect 43057 32879 43123 32880
rect 43060 32584 43120 32879
rect 42745 32524 43120 32584
rect 42421 31592 42488 31593
rect 42421 31590 42422 31592
rect 42066 31530 42422 31590
rect 41704 31148 41771 31149
rect 41704 31084 41705 31148
rect 41770 31146 41771 31148
rect 42066 31146 42126 31530
rect 42421 31528 42422 31530
rect 42487 31528 42488 31592
rect 42421 31527 42488 31528
rect 41770 31086 42126 31146
rect 41770 31084 41771 31086
rect 41704 31083 41771 31084
rect -272 30092 103 30152
rect 1401 30092 1776 30152
rect 2432 30092 40416 30152
rect 41072 30092 41447 30152
rect -272 29797 -212 30092
rect -275 29796 -209 29797
rect -275 29731 -274 29796
rect -210 29731 -209 29796
rect -275 29730 -209 29731
rect 722 29158 782 29473
rect 1077 29160 1144 29161
rect 1077 29158 1078 29160
rect 722 29098 1078 29158
rect 360 28716 427 28717
rect 360 28652 361 28716
rect 426 28714 427 28716
rect 722 28714 782 29098
rect 1077 29096 1078 29098
rect 1143 29096 1144 29160
rect 1077 29095 1144 29096
rect 2793 29031 2859 29032
rect 2793 28967 2794 29031
rect 2858 28967 2859 29031
rect 2793 28966 2859 28967
rect 2796 28717 2856 28966
rect 426 28654 782 28714
rect 426 28652 427 28654
rect 360 28651 427 28652
rect 722 28339 782 28654
rect 2793 28716 2859 28717
rect 2793 28652 2794 28716
rect 2858 28652 2859 28716
rect 2793 28651 2859 28652
rect 1713 28081 1779 28082
rect 1713 28016 1714 28081
rect 1778 28016 1779 28081
rect 1713 28015 1779 28016
rect 1716 27720 1776 28015
rect 3154 27720 3214 30092
rect 5586 27720 5646 30092
rect 7657 29031 7723 29032
rect 7657 28967 7658 29031
rect 7722 28967 7723 29031
rect 7657 28966 7723 28967
rect 7660 28717 7720 28966
rect 7657 28716 7723 28717
rect 7657 28652 7658 28716
rect 7722 28652 7723 28716
rect 7657 28651 7723 28652
rect 8018 27720 8078 30092
rect 10450 27720 10510 30092
rect 12521 29031 12587 29032
rect 12521 28967 12522 29031
rect 12586 28967 12587 29031
rect 12521 28966 12587 28967
rect 12524 28717 12584 28966
rect 12521 28716 12587 28717
rect 12521 28652 12522 28716
rect 12586 28652 12587 28716
rect 12521 28651 12587 28652
rect 12882 27720 12942 30092
rect 15314 27720 15374 30092
rect 17385 29031 17451 29032
rect 17385 28967 17386 29031
rect 17450 28967 17451 29031
rect 17385 28966 17451 28967
rect 17388 28717 17448 28966
rect 17385 28716 17451 28717
rect 17385 28652 17386 28716
rect 17450 28652 17451 28716
rect 17385 28651 17451 28652
rect 17746 27720 17806 30092
rect 20178 27720 20238 30092
rect 22249 29031 22315 29032
rect 22249 28967 22250 29031
rect 22314 28967 22315 29031
rect 22249 28966 22315 28967
rect 22252 28717 22312 28966
rect 22249 28716 22315 28717
rect 22249 28652 22250 28716
rect 22314 28652 22315 28716
rect 22249 28651 22315 28652
rect 22610 27720 22670 30092
rect 25042 27720 25102 30092
rect 27113 29031 27179 29032
rect 27113 28967 27114 29031
rect 27178 28967 27179 29031
rect 27113 28966 27179 28967
rect 27116 28717 27176 28966
rect 27113 28716 27179 28717
rect 27113 28652 27114 28716
rect 27178 28652 27179 28716
rect 27113 28651 27179 28652
rect 27474 27720 27534 30092
rect 29906 27720 29966 30092
rect 31977 29031 32043 29032
rect 31977 28967 31978 29031
rect 32042 28967 32043 29031
rect 31977 28966 32043 28967
rect 31980 28717 32040 28966
rect 31977 28716 32043 28717
rect 31977 28652 31978 28716
rect 32042 28652 32043 28716
rect 31977 28651 32043 28652
rect 32338 27720 32398 30092
rect 34770 27720 34830 30092
rect 36841 29031 36907 29032
rect 36841 28967 36842 29031
rect 36906 28967 36907 29031
rect 36841 28966 36907 28967
rect 36844 28717 36904 28966
rect 36841 28716 36907 28717
rect 36841 28652 36842 28716
rect 36906 28652 36907 28716
rect 36841 28651 36907 28652
rect 37202 27720 37262 30092
rect 39634 27720 39694 30092
rect 41072 29797 41132 30092
rect 41069 29796 41135 29797
rect 41069 29731 41070 29796
rect 41134 29731 41135 29796
rect 41069 29730 41135 29731
rect 42066 29158 42126 31086
rect 43057 30513 43123 30514
rect 43057 30448 43058 30513
rect 43122 30448 43123 30513
rect 43057 30447 43123 30448
rect 43060 30152 43120 30447
rect 42745 30092 43120 30152
rect 42421 29160 42488 29161
rect 42421 29158 42422 29160
rect 42066 29098 42422 29158
rect 41704 28716 41771 28717
rect 41704 28652 41705 28716
rect 41770 28714 41771 28716
rect 42066 28714 42126 29098
rect 42421 29096 42422 29098
rect 42487 29096 42488 29160
rect 42421 29095 42488 29096
rect 43412 29032 43472 33830
rect 43536 31464 43596 36262
rect 43533 31463 43599 31464
rect 43533 31399 43534 31463
rect 43598 31399 43599 31463
rect 43533 31398 43599 31399
rect 43409 29031 43475 29032
rect 43409 28967 43410 29031
rect 43474 28967 43475 29031
rect 43409 28966 43475 28967
rect 41770 28654 42126 28714
rect 41770 28652 41771 28654
rect 41704 28651 41771 28652
rect -272 27660 103 27720
rect 1401 27660 1776 27720
rect 2432 27660 40416 27720
rect 41072 27660 41447 27720
rect -272 27365 -212 27660
rect -275 27364 -209 27365
rect -275 27299 -274 27364
rect -210 27299 -209 27364
rect -275 27298 -209 27299
rect 722 26726 782 27041
rect 1077 26728 1144 26729
rect 1077 26726 1078 26728
rect 722 26666 1078 26726
rect -627 26413 -561 26414
rect -627 26349 -626 26413
rect -562 26349 -561 26413
rect -627 26348 -561 26349
rect -751 23981 -685 23982
rect -751 23917 -750 23981
rect -686 23917 -685 23981
rect -751 23916 -685 23917
rect -875 21363 -809 21364
rect -875 21299 -874 21363
rect -810 21299 -809 21363
rect -875 21298 -809 21299
rect -872 16488 -812 21298
rect -748 19118 -688 23916
rect -751 19117 -685 19118
rect -751 19053 -750 19117
rect -686 19053 -685 19117
rect -751 19052 -685 19053
rect -748 16500 -688 19052
rect -624 16686 -564 26348
rect 360 26284 427 26285
rect 360 26220 361 26284
rect 426 26282 427 26284
rect 722 26282 782 26666
rect 1077 26664 1078 26666
rect 1143 26664 1144 26728
rect 1077 26663 1144 26664
rect 426 26222 782 26282
rect 426 26220 427 26222
rect 360 26219 427 26220
rect 722 25907 782 26222
rect 1713 25649 1779 25650
rect 1713 25584 1714 25649
rect 1778 25584 1779 25649
rect 1713 25583 1779 25584
rect 1716 25288 1776 25583
rect 3154 25288 3214 27660
rect 5586 25288 5646 27660
rect 8018 25288 8078 27660
rect 10450 25288 10510 27660
rect 12882 25288 12942 27660
rect 15314 25288 15374 27660
rect 17746 25288 17806 27660
rect 20178 25288 20238 27660
rect 22610 25288 22670 27660
rect 25042 25288 25102 27660
rect 27474 25288 27534 27660
rect 29906 25288 29966 27660
rect 32338 25288 32398 27660
rect 34770 25288 34830 27660
rect 37202 25288 37262 27660
rect 39634 25288 39694 27660
rect 41072 27365 41132 27660
rect 41069 27364 41135 27365
rect 41069 27299 41070 27364
rect 41134 27299 41135 27364
rect 41069 27298 41135 27299
rect 42066 26726 42126 28654
rect 43057 28081 43123 28082
rect 43057 28016 43058 28081
rect 43122 28016 43123 28081
rect 43057 28015 43123 28016
rect 43060 27720 43120 28015
rect 42745 27660 43120 27720
rect 42421 26728 42488 26729
rect 42421 26726 42422 26728
rect 42066 26666 42422 26726
rect 41704 26284 41771 26285
rect 41704 26220 41705 26284
rect 41770 26282 41771 26284
rect 42066 26282 42126 26666
rect 42421 26664 42422 26666
rect 42487 26664 42488 26728
rect 42421 26663 42488 26664
rect 41770 26222 42126 26282
rect 41770 26220 41771 26222
rect 41704 26219 41771 26220
rect -272 25228 103 25288
rect 1401 25228 1776 25288
rect 2432 25228 40416 25288
rect 41072 25228 41447 25288
rect -272 24933 -212 25228
rect -275 24932 -209 24933
rect -275 24867 -274 24932
rect -210 24867 -209 24932
rect -275 24866 -209 24867
rect 722 24294 782 24609
rect 1077 24296 1144 24297
rect 1077 24294 1078 24296
rect 722 24234 1078 24294
rect 360 23852 427 23853
rect 360 23788 361 23852
rect 426 23850 427 23852
rect 722 23850 782 24234
rect 1077 24232 1078 24234
rect 1143 24232 1144 24296
rect 1077 24231 1144 24232
rect 2793 24167 2859 24168
rect 2793 24103 2794 24167
rect 2858 24103 2859 24167
rect 2793 24102 2859 24103
rect 2796 23853 2856 24102
rect 426 23790 782 23850
rect 426 23788 427 23790
rect 360 23787 427 23788
rect 722 23475 782 23790
rect 2793 23852 2859 23853
rect 2793 23788 2794 23852
rect 2858 23788 2859 23852
rect 2793 23787 2859 23788
rect 1713 23217 1779 23218
rect 1713 23152 1714 23217
rect 1778 23152 1779 23217
rect 1713 23151 1779 23152
rect 1716 22856 1776 23151
rect 3154 22856 3214 25228
rect 5586 22856 5646 25228
rect 7657 24167 7723 24168
rect 7657 24103 7658 24167
rect 7722 24103 7723 24167
rect 7657 24102 7723 24103
rect 7660 23853 7720 24102
rect 7657 23852 7723 23853
rect 7657 23788 7658 23852
rect 7722 23788 7723 23852
rect 7657 23787 7723 23788
rect 8018 22856 8078 25228
rect 10450 22856 10510 25228
rect 12521 24167 12587 24168
rect 12521 24103 12522 24167
rect 12586 24103 12587 24167
rect 12521 24102 12587 24103
rect 12524 23853 12584 24102
rect 12521 23852 12587 23853
rect 12521 23788 12522 23852
rect 12586 23788 12587 23852
rect 12521 23787 12587 23788
rect 12882 22856 12942 25228
rect 15314 22856 15374 25228
rect 17385 24167 17451 24168
rect 17385 24103 17386 24167
rect 17450 24103 17451 24167
rect 17385 24102 17451 24103
rect 17388 23853 17448 24102
rect 17385 23852 17451 23853
rect 17385 23788 17386 23852
rect 17450 23788 17451 23852
rect 17385 23787 17451 23788
rect 17746 22856 17806 25228
rect 20178 22856 20238 25228
rect 22249 24167 22315 24168
rect 22249 24103 22250 24167
rect 22314 24103 22315 24167
rect 22249 24102 22315 24103
rect 22252 23853 22312 24102
rect 22249 23852 22315 23853
rect 22249 23788 22250 23852
rect 22314 23788 22315 23852
rect 22249 23787 22315 23788
rect 22610 22856 22670 25228
rect 25042 22856 25102 25228
rect 27113 24167 27179 24168
rect 27113 24103 27114 24167
rect 27178 24103 27179 24167
rect 27113 24102 27179 24103
rect 27116 23853 27176 24102
rect 27113 23852 27179 23853
rect 27113 23788 27114 23852
rect 27178 23788 27179 23852
rect 27113 23787 27179 23788
rect 27474 22856 27534 25228
rect 29906 22856 29966 25228
rect 31977 24167 32043 24168
rect 31977 24103 31978 24167
rect 32042 24103 32043 24167
rect 31977 24102 32043 24103
rect 31980 23853 32040 24102
rect 31977 23852 32043 23853
rect 31977 23788 31978 23852
rect 32042 23788 32043 23852
rect 31977 23787 32043 23788
rect 32338 22856 32398 25228
rect 34770 22856 34830 25228
rect 36841 24167 36907 24168
rect 36841 24103 36842 24167
rect 36906 24103 36907 24167
rect 36841 24102 36907 24103
rect 36844 23853 36904 24102
rect 36841 23852 36907 23853
rect 36841 23788 36842 23852
rect 36906 23788 36907 23852
rect 36841 23787 36907 23788
rect 37202 22856 37262 25228
rect 39634 22856 39694 25228
rect 41072 24933 41132 25228
rect 41069 24932 41135 24933
rect 41069 24867 41070 24932
rect 41134 24867 41135 24932
rect 41069 24866 41135 24867
rect 42066 24294 42126 26222
rect 43057 25649 43123 25650
rect 43057 25584 43058 25649
rect 43122 25584 43123 25649
rect 43057 25583 43123 25584
rect 43060 25288 43120 25583
rect 42745 25228 43120 25288
rect 42421 24296 42488 24297
rect 42421 24294 42422 24296
rect 42066 24234 42422 24294
rect 41704 23852 41771 23853
rect 41704 23788 41705 23852
rect 41770 23850 41771 23852
rect 42066 23850 42126 24234
rect 42421 24232 42422 24234
rect 42487 24232 42488 24296
rect 42421 24231 42488 24232
rect 43412 24168 43472 28966
rect 43409 24167 43475 24168
rect 43409 24103 43410 24167
rect 43474 24103 43475 24167
rect 43409 24102 43475 24103
rect 41770 23790 42126 23850
rect 41770 23788 41771 23790
rect 41704 23787 41771 23788
rect -272 22796 103 22856
rect 1401 22796 1776 22856
rect 2432 22796 40416 22856
rect 41072 22796 41447 22856
rect -272 22501 -212 22796
rect -275 22500 -209 22501
rect -275 22435 -274 22500
rect -210 22435 -209 22500
rect -275 22434 -209 22435
rect 722 21862 782 22177
rect 1077 21864 1144 21865
rect 1077 21862 1078 21864
rect 722 21802 1078 21862
rect 360 21234 427 21235
rect 360 21170 361 21234
rect 426 21232 427 21234
rect 722 21232 782 21802
rect 1077 21800 1078 21802
rect 1143 21800 1144 21864
rect 1077 21799 1144 21800
rect 426 21172 782 21232
rect 426 21170 427 21172
rect 360 21169 427 21170
rect 722 20857 782 21172
rect 1713 20599 1779 20600
rect 1713 20534 1714 20599
rect 1778 20534 1779 20599
rect 1713 20533 1779 20534
rect 1716 20238 1776 20533
rect 3154 20238 3214 22796
rect 5586 20238 5646 22796
rect 8018 20238 8078 22796
rect 10450 20238 10510 22796
rect 10805 21864 10871 21865
rect 10805 21799 10806 21864
rect 10870 21799 10871 21864
rect 10805 21798 10871 21799
rect 10808 21365 10868 21798
rect 12521 21735 12587 21736
rect 12521 21671 12522 21735
rect 12586 21671 12587 21735
rect 12521 21670 12587 21671
rect 10805 21364 10871 21365
rect 10805 21299 10806 21364
rect 10870 21299 10871 21364
rect 10805 21298 10871 21299
rect 12524 21235 12584 21670
rect 12521 21234 12587 21235
rect 12521 21170 12522 21234
rect 12586 21170 12587 21234
rect 12521 21169 12587 21170
rect 12882 20238 12942 22796
rect 15314 20238 15374 22796
rect 17746 20238 17806 22796
rect 20178 20238 20238 22796
rect 22249 21549 22315 21550
rect 22249 21485 22250 21549
rect 22314 21485 22315 21549
rect 22249 21484 22315 21485
rect 22252 21235 22312 21484
rect 22249 21234 22315 21235
rect 22249 21170 22250 21234
rect 22314 21170 22315 21234
rect 22249 21169 22315 21170
rect 22610 20238 22670 22796
rect 25042 20238 25102 22796
rect 27474 20238 27534 22796
rect 29906 20238 29966 22796
rect 32338 20238 32398 22796
rect 34770 20238 34830 22796
rect 37202 20238 37262 22796
rect 39634 20238 39694 22796
rect 41072 22501 41132 22796
rect 41069 22500 41135 22501
rect 41069 22435 41070 22500
rect 41134 22435 41135 22500
rect 41069 22434 41135 22435
rect 39989 21864 40055 21865
rect 39989 21799 39990 21864
rect 40054 21799 40055 21864
rect 39989 21798 40055 21799
rect 42066 21862 42126 23790
rect 43057 23217 43123 23218
rect 43057 23152 43058 23217
rect 43122 23152 43123 23217
rect 43057 23151 43123 23152
rect 43060 22856 43120 23151
rect 42745 22796 43120 22856
rect 42421 21864 42488 21865
rect 42421 21862 42422 21864
rect 42066 21802 42422 21862
rect 39992 21365 40052 21798
rect 39989 21364 40055 21365
rect 39989 21299 39990 21364
rect 40054 21299 40055 21364
rect 39989 21298 40055 21299
rect 41704 21234 41771 21235
rect 41704 21170 41705 21234
rect 41770 21232 41771 21234
rect 42066 21232 42126 21802
rect 42421 21800 42422 21802
rect 42487 21800 42488 21864
rect 42421 21799 42488 21800
rect 41770 21172 42126 21232
rect 41770 21170 41771 21172
rect 41704 21169 41771 21170
rect -272 20178 103 20238
rect 1401 20178 1776 20238
rect 2432 20178 40416 20238
rect 41072 20178 41447 20238
rect -272 19883 -212 20178
rect -275 19882 -209 19883
rect -275 19817 -274 19882
rect -210 19817 -209 19882
rect -275 19816 -209 19817
rect 722 19244 782 19559
rect 1077 19246 1144 19247
rect 1077 19244 1078 19246
rect 722 19184 1078 19244
rect 360 18802 427 18803
rect 360 18738 361 18802
rect 426 18800 427 18802
rect 722 18800 782 19184
rect 1077 19182 1078 19184
rect 1143 19182 1144 19246
rect 1077 19181 1144 19182
rect 426 18740 782 18800
rect 426 18738 427 18740
rect 360 18737 427 18738
rect 722 18425 782 18740
rect 1713 18167 1779 18168
rect 1713 18102 1714 18167
rect 1778 18102 1779 18167
rect 1713 18101 1779 18102
rect 1716 17806 1776 18101
rect 3154 17806 3214 20178
rect 5586 17806 5646 20178
rect 5941 19246 6007 19247
rect 5941 19181 5942 19246
rect 6006 19181 6007 19246
rect 5941 19180 6007 19181
rect 5944 18933 6004 19180
rect 5941 18932 6007 18933
rect 5941 18867 5942 18932
rect 6006 18867 6007 18932
rect 5941 18866 6007 18867
rect 8018 17806 8078 20178
rect 10450 17806 10510 20178
rect 10805 19246 10871 19247
rect 10805 19181 10806 19246
rect 10870 19181 10871 19246
rect 10805 19180 10871 19181
rect 10808 18933 10868 19180
rect 10805 18932 10871 18933
rect 10805 18867 10806 18932
rect 10870 18867 10871 18932
rect 10805 18866 10871 18867
rect 12882 17806 12942 20178
rect 15314 17806 15374 20178
rect 15669 19246 15735 19247
rect 15669 19181 15670 19246
rect 15734 19181 15735 19246
rect 15669 19180 15735 19181
rect 15672 18933 15732 19180
rect 15669 18932 15735 18933
rect 15669 18867 15670 18932
rect 15734 18867 15735 18932
rect 15669 18866 15735 18867
rect 17746 17806 17806 20178
rect 20178 17806 20238 20178
rect 20533 19246 20599 19247
rect 20533 19181 20534 19246
rect 20598 19181 20599 19246
rect 20533 19180 20599 19181
rect 20536 18933 20596 19180
rect 20533 18932 20599 18933
rect 20533 18867 20534 18932
rect 20598 18867 20599 18932
rect 20533 18866 20599 18867
rect 22610 17806 22670 20178
rect 25042 17806 25102 20178
rect 25397 19246 25463 19247
rect 25397 19181 25398 19246
rect 25462 19181 25463 19246
rect 25397 19180 25463 19181
rect 25400 18933 25460 19180
rect 25397 18932 25463 18933
rect 25397 18867 25398 18932
rect 25462 18867 25463 18932
rect 25397 18866 25463 18867
rect 27474 17806 27534 20178
rect 29906 17806 29966 20178
rect 30261 19246 30327 19247
rect 30261 19181 30262 19246
rect 30326 19181 30327 19246
rect 30261 19180 30327 19181
rect 30264 18933 30324 19180
rect 30261 18932 30327 18933
rect 30261 18867 30262 18932
rect 30326 18867 30327 18932
rect 30261 18866 30327 18867
rect 32338 17806 32398 20178
rect 34770 17806 34830 20178
rect 35125 19246 35191 19247
rect 35125 19181 35126 19246
rect 35190 19181 35191 19246
rect 35125 19180 35191 19181
rect 35128 18933 35188 19180
rect 35125 18932 35191 18933
rect 35125 18867 35126 18932
rect 35190 18867 35191 18932
rect 35125 18866 35191 18867
rect 37202 17806 37262 20178
rect 39634 17806 39694 20178
rect 41072 19883 41132 20178
rect 41069 19882 41135 19883
rect 41069 19817 41070 19882
rect 41134 19817 41135 19882
rect 41069 19816 41135 19817
rect 39989 19246 40055 19247
rect 39989 19181 39990 19246
rect 40054 19181 40055 19246
rect 39989 19180 40055 19181
rect 42066 19244 42126 21172
rect 43057 20599 43123 20600
rect 43057 20534 43058 20599
rect 43122 20534 43123 20599
rect 43057 20533 43123 20534
rect 43060 20238 43120 20533
rect 42745 20178 43120 20238
rect 42421 19246 42488 19247
rect 42421 19244 42422 19246
rect 42066 19184 42422 19244
rect 39992 18933 40052 19180
rect 39989 18932 40055 18933
rect 39989 18867 39990 18932
rect 40054 18867 40055 18932
rect 39989 18866 40055 18867
rect 41704 18802 41771 18803
rect 41704 18738 41705 18802
rect 41770 18800 41771 18802
rect 42066 18800 42126 19184
rect 42421 19182 42422 19184
rect 42487 19182 42488 19246
rect 42421 19181 42488 19182
rect 43412 18932 43472 24102
rect 43409 18931 43475 18932
rect 43409 18867 43410 18931
rect 43474 18867 43475 18931
rect 43409 18866 43475 18867
rect 41770 18740 42126 18800
rect 41770 18738 41771 18740
rect 41704 18737 41771 18738
rect -272 17746 103 17806
rect 1401 17746 1776 17806
rect 2432 17746 40416 17806
rect 41072 17746 41447 17806
rect -272 17451 -212 17746
rect -275 17450 -209 17451
rect -275 17385 -274 17450
rect -210 17385 -209 17450
rect -275 17384 -209 17385
rect 722 16812 782 17127
rect 1077 16814 1144 16815
rect 1077 16812 1078 16814
rect 722 16752 1078 16812
rect -627 16685 -561 16686
rect -627 16621 -626 16685
rect -562 16621 -561 16685
rect -627 16620 -561 16621
rect -751 16499 -685 16500
rect -751 16435 -750 16499
rect -686 16435 -685 16499
rect -751 16434 -685 16435
rect -624 11822 -564 16620
rect 360 16370 427 16371
rect 360 16306 361 16370
rect 426 16368 427 16370
rect 722 16368 782 16752
rect 1077 16750 1078 16752
rect 1143 16750 1144 16814
rect 1077 16749 1144 16750
rect 426 16308 782 16368
rect 426 16306 427 16308
rect 360 16305 427 16306
rect 722 15993 782 16308
rect 1713 15735 1779 15736
rect 1713 15670 1714 15735
rect 1778 15670 1779 15735
rect 1713 15669 1779 15670
rect 1716 15374 1776 15669
rect 3154 15374 3214 17746
rect 5586 15374 5646 17746
rect 8018 15374 8078 17746
rect 10450 15374 10510 17746
rect 12882 15374 12942 17746
rect 15314 15374 15374 17746
rect 17746 15374 17806 17746
rect 20178 15374 20238 17746
rect 22610 15374 22670 17746
rect 25042 15374 25102 17746
rect 27474 15374 27534 17746
rect 29906 15374 29966 17746
rect 32338 15374 32398 17746
rect 34770 15374 34830 17746
rect 37202 15374 37262 17746
rect 39634 15374 39694 17746
rect 41072 17451 41132 17746
rect 41069 17450 41135 17451
rect 41069 17385 41070 17450
rect 41134 17385 41135 17450
rect 41069 17384 41135 17385
rect 42066 16812 42126 18740
rect 43057 18167 43123 18168
rect 43057 18102 43058 18167
rect 43122 18102 43123 18167
rect 43057 18101 43123 18102
rect 43060 17806 43120 18101
rect 42745 17746 43120 17806
rect 42421 16814 42488 16815
rect 42421 16812 42422 16814
rect 42066 16752 42422 16812
rect 41704 16370 41771 16371
rect 41704 16306 41705 16370
rect 41770 16368 41771 16370
rect 42066 16368 42126 16752
rect 42421 16750 42422 16752
rect 42487 16750 42488 16814
rect 42421 16749 42488 16750
rect 41770 16308 42126 16368
rect 41770 16306 41771 16308
rect 41704 16305 41771 16306
rect -272 15314 103 15374
rect 1401 15314 1776 15374
rect 2432 15314 40416 15374
rect 41072 15314 41447 15374
rect -272 15019 -212 15314
rect -275 15018 -209 15019
rect -275 14953 -274 15018
rect -210 14953 -209 15018
rect -275 14952 -209 14953
rect 722 14380 782 14695
rect 1077 14382 1144 14383
rect 1077 14380 1078 14382
rect 722 14320 1078 14380
rect 360 13938 427 13939
rect 360 13874 361 13938
rect 426 13936 427 13938
rect 722 13936 782 14320
rect 1077 14318 1078 14320
rect 1143 14318 1144 14382
rect 1077 14317 1144 14318
rect 426 13876 782 13936
rect 426 13874 427 13876
rect 360 13873 427 13874
rect 722 13561 782 13876
rect 1713 13303 1779 13304
rect 1713 13238 1714 13303
rect 1778 13238 1779 13303
rect 1713 13237 1779 13238
rect 1716 12942 1776 13237
rect 3154 12942 3214 15314
rect 5586 12942 5646 15314
rect 5941 14382 6007 14383
rect 5941 14317 5942 14382
rect 6006 14317 6007 14382
rect 5941 14316 6007 14317
rect 5944 14069 6004 14316
rect 5941 14068 6007 14069
rect 5941 14003 5942 14068
rect 6006 14003 6007 14068
rect 5941 14002 6007 14003
rect 8018 12942 8078 15314
rect 10450 12942 10510 15314
rect 10805 14382 10871 14383
rect 10805 14317 10806 14382
rect 10870 14317 10871 14382
rect 10805 14316 10871 14317
rect 10808 14069 10868 14316
rect 10805 14068 10871 14069
rect 10805 14003 10806 14068
rect 10870 14003 10871 14068
rect 10805 14002 10871 14003
rect 12882 12942 12942 15314
rect 15314 12942 15374 15314
rect 15669 14382 15735 14383
rect 15669 14317 15670 14382
rect 15734 14317 15735 14382
rect 15669 14316 15735 14317
rect 15672 14069 15732 14316
rect 15669 14068 15735 14069
rect 15669 14003 15670 14068
rect 15734 14003 15735 14068
rect 15669 14002 15735 14003
rect 17746 12942 17806 15314
rect 20178 12942 20238 15314
rect 20533 14382 20599 14383
rect 20533 14317 20534 14382
rect 20598 14317 20599 14382
rect 20533 14316 20599 14317
rect 20536 14069 20596 14316
rect 20533 14068 20599 14069
rect 20533 14003 20534 14068
rect 20598 14003 20599 14068
rect 20533 14002 20599 14003
rect 22610 12942 22670 15314
rect 25042 12942 25102 15314
rect 25397 14382 25463 14383
rect 25397 14317 25398 14382
rect 25462 14317 25463 14382
rect 25397 14316 25463 14317
rect 25400 14069 25460 14316
rect 25397 14068 25463 14069
rect 25397 14003 25398 14068
rect 25462 14003 25463 14068
rect 25397 14002 25463 14003
rect 27474 12942 27534 15314
rect 29906 12942 29966 15314
rect 30261 14382 30327 14383
rect 30261 14317 30262 14382
rect 30326 14317 30327 14382
rect 30261 14316 30327 14317
rect 30264 14069 30324 14316
rect 30261 14068 30327 14069
rect 30261 14003 30262 14068
rect 30326 14003 30327 14068
rect 30261 14002 30327 14003
rect 32338 12942 32398 15314
rect 34770 12942 34830 15314
rect 35125 14382 35191 14383
rect 35125 14317 35126 14382
rect 35190 14317 35191 14382
rect 35125 14316 35191 14317
rect 35128 14069 35188 14316
rect 35125 14068 35191 14069
rect 35125 14003 35126 14068
rect 35190 14003 35191 14068
rect 35125 14002 35191 14003
rect 37202 12942 37262 15314
rect 39634 12942 39694 15314
rect 41072 15019 41132 15314
rect 41069 15018 41135 15019
rect 41069 14953 41070 15018
rect 41134 14953 41135 15018
rect 41069 14952 41135 14953
rect 39989 14382 40055 14383
rect 39989 14317 39990 14382
rect 40054 14317 40055 14382
rect 39989 14316 40055 14317
rect 42066 14380 42126 16308
rect 43057 15735 43123 15736
rect 43057 15670 43058 15735
rect 43122 15670 43123 15735
rect 43057 15669 43123 15670
rect 43060 15374 43120 15669
rect 42745 15314 43120 15374
rect 42421 14382 42488 14383
rect 42421 14380 42422 14382
rect 42066 14320 42422 14380
rect 39992 14069 40052 14316
rect 39989 14068 40055 14069
rect 39989 14003 39990 14068
rect 40054 14003 40055 14068
rect 39989 14002 40055 14003
rect 41704 13938 41771 13939
rect 41704 13874 41705 13938
rect 41770 13936 41771 13938
rect 42066 13936 42126 14320
rect 42421 14318 42422 14320
rect 42487 14318 42488 14382
rect 42421 14317 42488 14318
rect 43412 14068 43472 18866
rect 43409 14067 43475 14068
rect 43409 14003 43410 14067
rect 43474 14003 43475 14067
rect 43409 14002 43475 14003
rect 41770 13876 42126 13936
rect 41770 13874 41771 13876
rect 41704 13873 41771 13874
rect -272 12882 103 12942
rect 1401 12882 1776 12942
rect 2432 12882 40416 12942
rect 41072 12882 41447 12942
rect -272 12587 -212 12882
rect -275 12586 -209 12587
rect -275 12521 -274 12586
rect -210 12521 -209 12586
rect -275 12520 -209 12521
rect 722 11948 782 12263
rect 1077 11950 1144 11951
rect 1077 11948 1078 11950
rect 722 11888 1078 11948
rect -627 11821 -561 11822
rect -627 11757 -626 11821
rect -562 11757 -561 11821
rect -627 11756 -561 11757
rect -624 6958 -564 11756
rect 360 11506 427 11507
rect 360 11442 361 11506
rect 426 11504 427 11506
rect 722 11504 782 11888
rect 1077 11886 1078 11888
rect 1143 11886 1144 11950
rect 1077 11885 1144 11886
rect 426 11444 782 11504
rect 426 11442 427 11444
rect 360 11441 427 11442
rect 722 11129 782 11444
rect 1713 10871 1779 10872
rect 1713 10806 1714 10871
rect 1778 10806 1779 10871
rect 1713 10805 1779 10806
rect 1716 10510 1776 10805
rect 3154 10510 3214 12882
rect 5586 10510 5646 12882
rect 8018 10510 8078 12882
rect 10450 10510 10510 12882
rect 12882 10510 12942 12882
rect 15314 10510 15374 12882
rect 17746 10510 17806 12882
rect 20178 10510 20238 12882
rect 22610 10510 22670 12882
rect 25042 10510 25102 12882
rect 27474 10510 27534 12882
rect 29906 10510 29966 12882
rect 32338 10510 32398 12882
rect 34770 10510 34830 12882
rect 37202 10510 37262 12882
rect 39634 10510 39694 12882
rect 41072 12587 41132 12882
rect 41069 12586 41135 12587
rect 41069 12521 41070 12586
rect 41134 12521 41135 12586
rect 41069 12520 41135 12521
rect 42066 11948 42126 13876
rect 43057 13303 43123 13304
rect 43057 13238 43058 13303
rect 43122 13238 43123 13303
rect 43057 13237 43123 13238
rect 43060 12942 43120 13237
rect 42745 12882 43120 12942
rect 42421 11950 42488 11951
rect 42421 11948 42422 11950
rect 42066 11888 42422 11948
rect 41704 11506 41771 11507
rect 41704 11442 41705 11506
rect 41770 11504 41771 11506
rect 42066 11504 42126 11888
rect 42421 11886 42422 11888
rect 42487 11886 42488 11950
rect 42421 11885 42488 11886
rect 41770 11444 42126 11504
rect 41770 11442 41771 11444
rect 41704 11441 41771 11442
rect -272 10450 103 10510
rect 1401 10450 1776 10510
rect 2432 10450 40416 10510
rect 41072 10450 41447 10510
rect -272 10155 -212 10450
rect -275 10154 -209 10155
rect -275 10089 -274 10154
rect -210 10089 -209 10154
rect -275 10088 -209 10089
rect 722 9516 782 9831
rect 1077 9518 1144 9519
rect 1077 9516 1078 9518
rect 722 9456 1078 9516
rect 360 9074 427 9075
rect 360 9010 361 9074
rect 426 9072 427 9074
rect 722 9072 782 9456
rect 1077 9454 1078 9456
rect 1143 9454 1144 9518
rect 1077 9453 1144 9454
rect 426 9012 782 9072
rect 426 9010 427 9012
rect 360 9009 427 9010
rect 722 8697 782 9012
rect 1713 8439 1779 8440
rect 1713 8374 1714 8439
rect 1778 8374 1779 8439
rect 1713 8373 1779 8374
rect 1716 8078 1776 8373
rect 3154 8078 3214 10450
rect 5586 8078 5646 10450
rect 5941 9518 6007 9519
rect 5941 9453 5942 9518
rect 6006 9453 6007 9518
rect 5941 9452 6007 9453
rect 5944 9205 6004 9452
rect 5941 9204 6007 9205
rect 5941 9139 5942 9204
rect 6006 9139 6007 9204
rect 5941 9138 6007 9139
rect 8018 8078 8078 10450
rect 10450 8078 10510 10450
rect 10805 9518 10871 9519
rect 10805 9453 10806 9518
rect 10870 9453 10871 9518
rect 10805 9452 10871 9453
rect 10808 9205 10868 9452
rect 10805 9204 10871 9205
rect 10805 9139 10806 9204
rect 10870 9139 10871 9204
rect 10805 9138 10871 9139
rect 12882 8078 12942 10450
rect 15314 8078 15374 10450
rect 15669 9518 15735 9519
rect 15669 9453 15670 9518
rect 15734 9453 15735 9518
rect 15669 9452 15735 9453
rect 15672 9205 15732 9452
rect 15669 9204 15735 9205
rect 15669 9139 15670 9204
rect 15734 9139 15735 9204
rect 15669 9138 15735 9139
rect 17746 8078 17806 10450
rect 20178 8078 20238 10450
rect 20533 9518 20599 9519
rect 20533 9453 20534 9518
rect 20598 9453 20599 9518
rect 20533 9452 20599 9453
rect 20536 9205 20596 9452
rect 20533 9204 20599 9205
rect 20533 9139 20534 9204
rect 20598 9139 20599 9204
rect 20533 9138 20599 9139
rect 22610 8078 22670 10450
rect 25042 8078 25102 10450
rect 25397 9518 25463 9519
rect 25397 9453 25398 9518
rect 25462 9453 25463 9518
rect 25397 9452 25463 9453
rect 25400 9205 25460 9452
rect 25397 9204 25463 9205
rect 25397 9139 25398 9204
rect 25462 9139 25463 9204
rect 25397 9138 25463 9139
rect 27474 8078 27534 10450
rect 29906 8078 29966 10450
rect 30261 9518 30327 9519
rect 30261 9453 30262 9518
rect 30326 9453 30327 9518
rect 30261 9452 30327 9453
rect 30264 9205 30324 9452
rect 30261 9204 30327 9205
rect 30261 9139 30262 9204
rect 30326 9139 30327 9204
rect 30261 9138 30327 9139
rect 32338 8078 32398 10450
rect 34770 8078 34830 10450
rect 35125 9518 35191 9519
rect 35125 9453 35126 9518
rect 35190 9453 35191 9518
rect 35125 9452 35191 9453
rect 35128 9205 35188 9452
rect 35125 9204 35191 9205
rect 35125 9139 35126 9204
rect 35190 9139 35191 9204
rect 35125 9138 35191 9139
rect 37202 8078 37262 10450
rect 39634 8078 39694 10450
rect 41072 10155 41132 10450
rect 41069 10154 41135 10155
rect 41069 10089 41070 10154
rect 41134 10089 41135 10154
rect 41069 10088 41135 10089
rect 39989 9518 40055 9519
rect 39989 9453 39990 9518
rect 40054 9453 40055 9518
rect 39989 9452 40055 9453
rect 42066 9516 42126 11444
rect 43057 10871 43123 10872
rect 43057 10806 43058 10871
rect 43122 10806 43123 10871
rect 43057 10805 43123 10806
rect 43060 10510 43120 10805
rect 42745 10450 43120 10510
rect 42421 9518 42488 9519
rect 42421 9516 42422 9518
rect 42066 9456 42422 9516
rect 39992 9205 40052 9452
rect 39989 9204 40055 9205
rect 39989 9139 39990 9204
rect 40054 9139 40055 9204
rect 39989 9138 40055 9139
rect 41704 9074 41771 9075
rect 41704 9010 41705 9074
rect 41770 9072 41771 9074
rect 42066 9072 42126 9456
rect 42421 9454 42422 9456
rect 42487 9454 42488 9518
rect 42421 9453 42488 9454
rect 43412 9204 43472 14002
rect 43536 11636 43596 31398
rect 43660 28846 43720 44374
rect 43657 28845 43723 28846
rect 43657 28781 43658 28845
rect 43722 28781 43723 28845
rect 43657 28780 43723 28781
rect 43660 14254 43720 28780
rect 43784 21736 43844 44630
rect 43781 21735 43847 21736
rect 43781 21671 43782 21735
rect 43846 21671 43847 21735
rect 43781 21670 43847 21671
rect 43657 14253 43723 14254
rect 43657 14189 43658 14253
rect 43722 14189 43723 14253
rect 43657 14188 43723 14189
rect 43533 11635 43599 11636
rect 43533 11571 43534 11635
rect 43598 11571 43599 11635
rect 43533 11570 43599 11571
rect 43409 9203 43475 9204
rect 43409 9139 43410 9203
rect 43474 9139 43475 9203
rect 43409 9138 43475 9139
rect 41770 9012 42126 9072
rect 41770 9010 41771 9012
rect 41704 9009 41771 9010
rect -272 8018 103 8078
rect 1401 8018 1776 8078
rect 2432 8018 40416 8078
rect 41072 8018 41447 8078
rect -272 7723 -212 8018
rect -275 7722 -209 7723
rect -275 7657 -274 7722
rect -210 7657 -209 7722
rect -275 7656 -209 7657
rect 722 7084 782 7399
rect 1077 7086 1144 7087
rect 1077 7084 1078 7086
rect 722 7024 1078 7084
rect -627 6957 -561 6958
rect -627 6893 -626 6957
rect -562 6893 -561 6957
rect -627 6892 -561 6893
rect -624 2094 -564 6892
rect 360 6642 427 6643
rect 360 6578 361 6642
rect 426 6640 427 6642
rect 722 6640 782 7024
rect 1077 7022 1078 7024
rect 1143 7022 1144 7086
rect 1077 7021 1144 7022
rect 426 6580 782 6640
rect 426 6578 427 6580
rect 360 6577 427 6578
rect 722 6265 782 6580
rect 1713 6007 1779 6008
rect 1713 5942 1714 6007
rect 1778 5942 1779 6007
rect 1713 5941 1779 5942
rect 1716 5646 1776 5941
rect 3154 5646 3214 8018
rect 5586 5646 5646 8018
rect 8018 5646 8078 8018
rect 10450 5646 10510 8018
rect 12882 5646 12942 8018
rect 15314 5646 15374 8018
rect 17746 5646 17806 8018
rect 20178 5646 20238 8018
rect 22610 5646 22670 8018
rect 25042 5646 25102 8018
rect 27474 5646 27534 8018
rect 29906 5646 29966 8018
rect 32338 5646 32398 8018
rect 34770 5646 34830 8018
rect 37202 5646 37262 8018
rect 39634 5646 39694 8018
rect 41072 7723 41132 8018
rect 41069 7722 41135 7723
rect 41069 7657 41070 7722
rect 41134 7657 41135 7722
rect 41069 7656 41135 7657
rect 42066 7084 42126 9012
rect 43057 8439 43123 8440
rect 43057 8374 43058 8439
rect 43122 8374 43123 8439
rect 43057 8373 43123 8374
rect 43060 8078 43120 8373
rect 42745 8018 43120 8078
rect 42421 7086 42488 7087
rect 42421 7084 42422 7086
rect 42066 7024 42422 7084
rect 41704 6642 41771 6643
rect 41704 6578 41705 6642
rect 41770 6640 41771 6642
rect 42066 6640 42126 7024
rect 42421 7022 42422 7024
rect 42487 7022 42488 7086
rect 42421 7021 42488 7022
rect 41770 6580 42126 6640
rect 41770 6578 41771 6580
rect 41704 6577 41771 6578
rect -272 5586 103 5646
rect 1401 5586 1776 5646
rect 2432 5586 40416 5646
rect 41072 5586 41447 5646
rect -272 5291 -212 5586
rect -275 5290 -209 5291
rect -275 5225 -274 5290
rect -210 5225 -209 5290
rect -275 5224 -209 5225
rect 722 4652 782 4967
rect 1077 4654 1144 4655
rect 1077 4652 1078 4654
rect 722 4592 1078 4652
rect 360 4210 427 4211
rect 360 4146 361 4210
rect 426 4208 427 4210
rect 722 4208 782 4592
rect 1077 4590 1078 4592
rect 1143 4590 1144 4654
rect 1077 4589 1144 4590
rect 426 4148 782 4208
rect 426 4146 427 4148
rect 360 4145 427 4146
rect 722 3833 782 4148
rect 1713 3575 1779 3576
rect 1713 3510 1714 3575
rect 1778 3510 1779 3575
rect 1713 3509 1779 3510
rect 1716 3214 1776 3509
rect 3154 3214 3214 5586
rect 5586 3214 5646 5586
rect 5941 4654 6007 4655
rect 5941 4589 5942 4654
rect 6006 4589 6007 4654
rect 5941 4588 6007 4589
rect 5944 4341 6004 4588
rect 5941 4340 6007 4341
rect 5941 4275 5942 4340
rect 6006 4275 6007 4340
rect 5941 4274 6007 4275
rect 8018 3214 8078 5586
rect 10450 3214 10510 5586
rect 10805 4654 10871 4655
rect 10805 4589 10806 4654
rect 10870 4589 10871 4654
rect 10805 4588 10871 4589
rect 10808 4341 10868 4588
rect 10805 4340 10871 4341
rect 10805 4275 10806 4340
rect 10870 4275 10871 4340
rect 10805 4274 10871 4275
rect 12882 3214 12942 5586
rect 15314 3214 15374 5586
rect 15669 4654 15735 4655
rect 15669 4589 15670 4654
rect 15734 4589 15735 4654
rect 15669 4588 15735 4589
rect 15672 4341 15732 4588
rect 15669 4340 15735 4341
rect 15669 4275 15670 4340
rect 15734 4275 15735 4340
rect 15669 4274 15735 4275
rect 17746 3214 17806 5586
rect 20178 3214 20238 5586
rect 20533 4654 20599 4655
rect 20533 4589 20534 4654
rect 20598 4589 20599 4654
rect 20533 4588 20599 4589
rect 20536 4341 20596 4588
rect 20533 4340 20599 4341
rect 20533 4275 20534 4340
rect 20598 4275 20599 4340
rect 20533 4274 20599 4275
rect 22610 3214 22670 5586
rect 25042 3214 25102 5586
rect 25397 4654 25463 4655
rect 25397 4589 25398 4654
rect 25462 4589 25463 4654
rect 25397 4588 25463 4589
rect 25400 4341 25460 4588
rect 25397 4340 25463 4341
rect 25397 4275 25398 4340
rect 25462 4275 25463 4340
rect 25397 4274 25463 4275
rect 27474 3214 27534 5586
rect 29906 3214 29966 5586
rect 30261 4654 30327 4655
rect 30261 4589 30262 4654
rect 30326 4589 30327 4654
rect 30261 4588 30327 4589
rect 30264 4341 30324 4588
rect 30261 4340 30327 4341
rect 30261 4275 30262 4340
rect 30326 4275 30327 4340
rect 30261 4274 30327 4275
rect 32338 3214 32398 5586
rect 34770 3214 34830 5586
rect 35125 4654 35191 4655
rect 35125 4589 35126 4654
rect 35190 4589 35191 4654
rect 35125 4588 35191 4589
rect 35128 4341 35188 4588
rect 35125 4340 35191 4341
rect 35125 4275 35126 4340
rect 35190 4275 35191 4340
rect 35125 4274 35191 4275
rect 37202 3214 37262 5586
rect 39634 3214 39694 5586
rect 41072 5291 41132 5586
rect 41069 5290 41135 5291
rect 41069 5225 41070 5290
rect 41134 5225 41135 5290
rect 41069 5224 41135 5225
rect 39989 4654 40055 4655
rect 39989 4589 39990 4654
rect 40054 4589 40055 4654
rect 39989 4588 40055 4589
rect 42066 4652 42126 6580
rect 43057 6007 43123 6008
rect 43057 5942 43058 6007
rect 43122 5942 43123 6007
rect 43057 5941 43123 5942
rect 43060 5646 43120 5941
rect 42745 5586 43120 5646
rect 42421 4654 42488 4655
rect 42421 4652 42422 4654
rect 42066 4592 42422 4652
rect 39992 4341 40052 4588
rect 39989 4340 40055 4341
rect 39989 4275 39990 4340
rect 40054 4275 40055 4340
rect 39989 4274 40055 4275
rect 41704 4210 41771 4211
rect 41704 4146 41705 4210
rect 41770 4208 41771 4210
rect 42066 4208 42126 4592
rect 42421 4590 42422 4592
rect 42487 4590 42488 4654
rect 42421 4589 42488 4590
rect 43412 4341 43472 9138
rect 43536 6772 43596 11570
rect 43533 6771 43599 6772
rect 43533 6707 43534 6771
rect 43598 6707 43599 6771
rect 43533 6706 43599 6707
rect 43409 4340 43475 4341
rect 43409 4275 43410 4340
rect 43474 4275 43475 4340
rect 43409 4274 43475 4275
rect 41770 4148 42126 4208
rect 41770 4146 41771 4148
rect 41704 4145 41771 4146
rect -272 3154 103 3214
rect 1401 3154 1776 3214
rect 2432 3154 40416 3214
rect 41072 3154 41447 3214
rect -272 2859 -212 3154
rect -275 2858 -209 2859
rect -275 2793 -274 2858
rect -210 2793 -209 2858
rect -275 2792 -209 2793
rect 722 2220 782 2535
rect 3154 2431 3214 3154
rect 5586 2431 5646 3154
rect 8018 2431 8078 3154
rect 10450 2431 10510 3154
rect 12882 2431 12942 3154
rect 15314 2431 15374 3154
rect 17746 2431 17806 3154
rect 20178 2431 20238 3154
rect 22610 2431 22670 3154
rect 25042 2431 25102 3154
rect 27474 2431 27534 3154
rect 29906 2431 29966 3154
rect 32338 2431 32398 3154
rect 34770 2431 34830 3154
rect 37202 2431 37262 3154
rect 39634 2431 39694 3154
rect 41072 2859 41132 3154
rect 41069 2858 41135 2859
rect 41069 2793 41070 2858
rect 41134 2793 41135 2858
rect 41069 2792 41135 2793
rect 1077 2222 1144 2223
rect 1077 2220 1078 2222
rect 722 2160 1078 2220
rect -627 2093 -561 2094
rect -627 2029 -626 2093
rect -562 2029 -561 2093
rect -627 2028 -561 2029
rect 360 1778 427 1779
rect 360 1714 361 1778
rect 426 1776 427 1778
rect 722 1776 782 2160
rect 1077 2158 1078 2160
rect 1143 2158 1144 2222
rect 1077 2157 1144 2158
rect 42066 2220 42126 4148
rect 43057 3575 43123 3576
rect 43057 3510 43058 3575
rect 43122 3510 43123 3575
rect 43057 3509 43123 3510
rect 43060 3214 43120 3509
rect 42745 3154 43120 3214
rect 42421 2222 42488 2223
rect 42421 2220 42422 2222
rect 42066 2160 42422 2220
rect 426 1716 782 1776
rect 426 1714 427 1716
rect 360 1713 427 1714
rect 722 782 782 1716
rect 2792 1778 2859 1779
rect 2792 1714 2793 1778
rect 2858 1776 2859 1778
rect 5224 1778 5291 1779
rect 2858 1716 3214 1776
rect 2858 1714 2859 1716
rect 2792 1713 2859 1714
rect 3154 1468 3214 1716
rect 5224 1714 5225 1778
rect 5290 1776 5291 1778
rect 7656 1778 7723 1779
rect 5290 1716 5646 1776
rect 5290 1714 5291 1716
rect 5224 1713 5291 1714
rect 5586 1401 5646 1716
rect 7656 1714 7657 1778
rect 7722 1776 7723 1778
rect 10088 1778 10155 1779
rect 7722 1716 8078 1776
rect 7722 1714 7723 1716
rect 7656 1713 7723 1714
rect 8018 1401 8078 1716
rect 10088 1714 10089 1778
rect 10154 1776 10155 1778
rect 12520 1778 12587 1779
rect 10154 1716 10510 1776
rect 10154 1714 10155 1716
rect 10088 1713 10155 1714
rect 10450 1401 10510 1716
rect 12520 1714 12521 1778
rect 12586 1776 12587 1778
rect 14952 1778 15019 1779
rect 12586 1716 12942 1776
rect 12586 1714 12587 1716
rect 12520 1713 12587 1714
rect 12882 1401 12942 1716
rect 14952 1714 14953 1778
rect 15018 1776 15019 1778
rect 17384 1778 17451 1779
rect 15018 1716 15374 1776
rect 15018 1714 15019 1716
rect 14952 1713 15019 1714
rect 15314 1401 15374 1716
rect 17384 1714 17385 1778
rect 17450 1776 17451 1778
rect 19816 1778 19883 1779
rect 17450 1716 17806 1776
rect 17450 1714 17451 1716
rect 17384 1713 17451 1714
rect 17746 1401 17806 1716
rect 19816 1714 19817 1778
rect 19882 1776 19883 1778
rect 22248 1778 22315 1779
rect 19882 1716 20238 1776
rect 19882 1714 19883 1716
rect 19816 1713 19883 1714
rect 20178 1401 20238 1716
rect 22248 1714 22249 1778
rect 22314 1776 22315 1778
rect 24680 1778 24747 1779
rect 22314 1716 22670 1776
rect 22314 1714 22315 1716
rect 22248 1713 22315 1714
rect 22610 1401 22670 1716
rect 24680 1714 24681 1778
rect 24746 1776 24747 1778
rect 27112 1778 27179 1779
rect 24746 1716 25102 1776
rect 24746 1714 24747 1716
rect 24680 1713 24747 1714
rect 25042 1401 25102 1716
rect 27112 1714 27113 1778
rect 27178 1776 27179 1778
rect 29544 1778 29611 1779
rect 27178 1716 27534 1776
rect 27178 1714 27179 1716
rect 27112 1713 27179 1714
rect 27474 1401 27534 1716
rect 29544 1714 29545 1778
rect 29610 1776 29611 1778
rect 31976 1778 32043 1779
rect 29610 1716 29966 1776
rect 29610 1714 29611 1716
rect 29544 1713 29611 1714
rect 29906 1401 29966 1716
rect 31976 1714 31977 1778
rect 32042 1776 32043 1778
rect 34408 1778 34475 1779
rect 32042 1716 32398 1776
rect 32042 1714 32043 1716
rect 31976 1713 32043 1714
rect 32338 1401 32398 1716
rect 34408 1714 34409 1778
rect 34474 1776 34475 1778
rect 36840 1778 36907 1779
rect 34474 1716 34830 1776
rect 34474 1714 34475 1716
rect 34408 1713 34475 1714
rect 34770 1401 34830 1716
rect 36840 1714 36841 1778
rect 36906 1776 36907 1778
rect 39272 1778 39339 1779
rect 36906 1716 37262 1776
rect 36906 1714 36907 1716
rect 36840 1713 36907 1714
rect 37202 1401 37262 1716
rect 39272 1714 39273 1778
rect 39338 1776 39339 1778
rect 41704 1778 41771 1779
rect 39338 1716 39694 1776
rect 39338 1714 39339 1716
rect 39272 1713 39339 1714
rect 39634 1401 39694 1716
rect 41704 1714 41705 1778
rect 41770 1776 41771 1778
rect 42066 1776 42126 2160
rect 42421 2158 42422 2160
rect 42487 2158 42488 2222
rect 42421 2157 42488 2158
rect 41770 1716 42126 1776
rect 41770 1714 41771 1716
rect 41704 1713 41771 1714
rect 1713 1143 1779 1144
rect 1713 1078 1714 1143
rect 1778 1078 1779 1143
rect 1713 1077 1779 1078
rect 4145 1143 4211 1144
rect 4145 1078 4146 1143
rect 4210 1078 4211 1143
rect 4145 1077 4211 1078
rect 6577 1143 6643 1144
rect 6577 1078 6578 1143
rect 6642 1078 6643 1143
rect 6577 1077 6643 1078
rect 9009 1143 9075 1144
rect 9009 1078 9010 1143
rect 9074 1078 9075 1143
rect 9009 1077 9075 1078
rect 11441 1143 11507 1144
rect 11441 1078 11442 1143
rect 11506 1078 11507 1143
rect 11441 1077 11507 1078
rect 13873 1143 13939 1144
rect 13873 1078 13874 1143
rect 13938 1078 13939 1143
rect 13873 1077 13939 1078
rect 16305 1143 16371 1144
rect 16305 1078 16306 1143
rect 16370 1078 16371 1143
rect 16305 1077 16371 1078
rect 18737 1143 18803 1144
rect 18737 1078 18738 1143
rect 18802 1078 18803 1143
rect 18737 1077 18803 1078
rect 21169 1143 21235 1144
rect 21169 1078 21170 1143
rect 21234 1078 21235 1143
rect 21169 1077 21235 1078
rect 23601 1143 23667 1144
rect 23601 1078 23602 1143
rect 23666 1078 23667 1143
rect 23601 1077 23667 1078
rect 26033 1143 26099 1144
rect 26033 1078 26034 1143
rect 26098 1078 26099 1143
rect 26033 1077 26099 1078
rect 28465 1143 28531 1144
rect 28465 1078 28466 1143
rect 28530 1078 28531 1143
rect 28465 1077 28531 1078
rect 30897 1143 30963 1144
rect 30897 1078 30898 1143
rect 30962 1078 30963 1143
rect 30897 1077 30963 1078
rect 33329 1143 33395 1144
rect 33329 1078 33330 1143
rect 33394 1078 33395 1143
rect 33329 1077 33395 1078
rect 35761 1143 35827 1144
rect 35761 1078 35762 1143
rect 35826 1078 35827 1143
rect 35761 1077 35827 1078
rect 38193 1143 38259 1144
rect 38193 1078 38194 1143
rect 38258 1078 38259 1143
rect 38193 1077 38259 1078
rect 40625 1143 40691 1144
rect 40625 1078 40626 1143
rect 40690 1078 40691 1143
rect 40625 1077 40691 1078
rect 1716 782 1776 1077
rect 4148 782 4208 1077
rect 6580 782 6640 1077
rect 9012 782 9072 1077
rect 11444 782 11504 1077
rect 13876 782 13936 1077
rect 16308 782 16368 1077
rect 18740 782 18800 1077
rect 21172 782 21232 1077
rect 23604 782 23664 1077
rect 26036 782 26096 1077
rect 28468 782 28528 1077
rect 30900 782 30960 1077
rect 33332 782 33392 1077
rect 35764 782 35824 1077
rect 38196 782 38256 1077
rect 40628 782 40688 1077
rect 42066 782 42126 1716
rect 43057 1143 43123 1144
rect 43057 1078 43058 1143
rect 43122 1078 43123 1143
rect 43057 1077 43123 1078
rect 43060 782 43120 1077
rect -272 722 43120 782
rect -272 427 -212 722
rect -275 426 -209 427
rect -275 361 -274 426
rect -210 361 -209 426
rect -275 360 -209 361
rect 722 -212 782 722
rect 2160 427 2220 722
rect 4592 427 4652 722
rect 7024 427 7084 722
rect 9456 427 9516 722
rect 11888 427 11948 722
rect 14320 427 14380 722
rect 16752 427 16812 722
rect 19184 427 19244 722
rect 21616 427 21676 722
rect 24048 427 24108 722
rect 26480 427 26540 722
rect 28912 427 28972 722
rect 31344 427 31404 722
rect 33776 427 33836 722
rect 36208 427 36268 722
rect 38640 427 38700 722
rect 41072 427 41132 722
rect 2157 426 2223 427
rect 2157 361 2158 426
rect 2222 361 2223 426
rect 2157 360 2223 361
rect 4589 426 4655 427
rect 4589 361 4590 426
rect 4654 361 4655 426
rect 4589 360 4655 361
rect 7021 426 7087 427
rect 7021 361 7022 426
rect 7086 361 7087 426
rect 7021 360 7087 361
rect 9453 426 9519 427
rect 9453 361 9454 426
rect 9518 361 9519 426
rect 9453 360 9519 361
rect 11885 426 11951 427
rect 11885 361 11886 426
rect 11950 361 11951 426
rect 11885 360 11951 361
rect 14317 426 14383 427
rect 14317 361 14318 426
rect 14382 361 14383 426
rect 14317 360 14383 361
rect 16749 426 16815 427
rect 16749 361 16750 426
rect 16814 361 16815 426
rect 16749 360 16815 361
rect 19181 426 19247 427
rect 19181 361 19182 426
rect 19246 361 19247 426
rect 19181 360 19247 361
rect 21613 426 21679 427
rect 21613 361 21614 426
rect 21678 361 21679 426
rect 21613 360 21679 361
rect 24045 426 24111 427
rect 24045 361 24046 426
rect 24110 361 24111 426
rect 24045 360 24111 361
rect 26477 426 26543 427
rect 26477 361 26478 426
rect 26542 361 26543 426
rect 26477 360 26543 361
rect 28909 426 28975 427
rect 28909 361 28910 426
rect 28974 361 28975 426
rect 28909 360 28975 361
rect 31341 426 31407 427
rect 31341 361 31342 426
rect 31406 361 31407 426
rect 31341 360 31407 361
rect 33773 426 33839 427
rect 33773 361 33774 426
rect 33838 361 33839 426
rect 33773 360 33839 361
rect 36205 426 36271 427
rect 36205 361 36206 426
rect 36270 361 36271 426
rect 36205 360 36271 361
rect 38637 426 38703 427
rect 38637 361 38638 426
rect 38702 361 38703 426
rect 38637 360 38703 361
rect 41069 426 41135 427
rect 41069 361 41070 426
rect 41134 361 41135 426
rect 41069 360 41135 361
rect 1077 -210 1144 -209
rect 1077 -212 1078 -210
rect 722 -272 1078 -212
rect 1077 -274 1078 -272
rect 1143 -274 1144 -210
rect 3154 -212 3214 36
rect 3509 -210 3576 -209
rect 3509 -212 3510 -210
rect 3154 -272 3510 -212
rect 1077 -275 1144 -274
rect 3509 -274 3510 -272
rect 3575 -274 3576 -210
rect 5586 -212 5646 103
rect 5941 -210 6008 -209
rect 5941 -212 5942 -210
rect 5586 -272 5942 -212
rect 3509 -275 3576 -274
rect 5941 -274 5942 -272
rect 6007 -274 6008 -210
rect 8018 -212 8078 103
rect 8373 -210 8440 -209
rect 8373 -212 8374 -210
rect 8018 -272 8374 -212
rect 5941 -275 6008 -274
rect 8373 -274 8374 -272
rect 8439 -274 8440 -210
rect 10450 -212 10510 103
rect 10805 -210 10872 -209
rect 10805 -212 10806 -210
rect 10450 -272 10806 -212
rect 8373 -275 8440 -274
rect 10805 -274 10806 -272
rect 10871 -274 10872 -210
rect 12882 -212 12942 103
rect 13237 -210 13304 -209
rect 13237 -212 13238 -210
rect 12882 -272 13238 -212
rect 10805 -275 10872 -274
rect 13237 -274 13238 -272
rect 13303 -274 13304 -210
rect 15314 -212 15374 103
rect 15669 -210 15736 -209
rect 15669 -212 15670 -210
rect 15314 -272 15670 -212
rect 13237 -275 13304 -274
rect 15669 -274 15670 -272
rect 15735 -274 15736 -210
rect 17746 -212 17806 103
rect 18101 -210 18168 -209
rect 18101 -212 18102 -210
rect 17746 -272 18102 -212
rect 15669 -275 15736 -274
rect 18101 -274 18102 -272
rect 18167 -274 18168 -210
rect 20178 -212 20238 103
rect 20533 -210 20600 -209
rect 20533 -212 20534 -210
rect 20178 -272 20534 -212
rect 18101 -275 18168 -274
rect 20533 -274 20534 -272
rect 20599 -274 20600 -210
rect 22610 -212 22670 103
rect 22965 -210 23032 -209
rect 22965 -212 22966 -210
rect 22610 -272 22966 -212
rect 20533 -275 20600 -274
rect 22965 -274 22966 -272
rect 23031 -274 23032 -210
rect 25042 -212 25102 103
rect 25397 -210 25464 -209
rect 25397 -212 25398 -210
rect 25042 -272 25398 -212
rect 22965 -275 23032 -274
rect 25397 -274 25398 -272
rect 25463 -274 25464 -210
rect 27474 -212 27534 103
rect 27829 -210 27896 -209
rect 27829 -212 27830 -210
rect 27474 -272 27830 -212
rect 25397 -275 25464 -274
rect 27829 -274 27830 -272
rect 27895 -274 27896 -210
rect 29906 -212 29966 103
rect 30261 -210 30328 -209
rect 30261 -212 30262 -210
rect 29906 -272 30262 -212
rect 27829 -275 27896 -274
rect 30261 -274 30262 -272
rect 30327 -274 30328 -210
rect 32338 -212 32398 103
rect 32693 -210 32760 -209
rect 32693 -212 32694 -210
rect 32338 -272 32694 -212
rect 30261 -275 30328 -274
rect 32693 -274 32694 -272
rect 32759 -274 32760 -210
rect 34770 -212 34830 103
rect 35125 -210 35192 -209
rect 35125 -212 35126 -210
rect 34770 -272 35126 -212
rect 32693 -275 32760 -274
rect 35125 -274 35126 -272
rect 35191 -274 35192 -210
rect 37202 -212 37262 103
rect 37557 -210 37624 -209
rect 37557 -212 37558 -210
rect 37202 -272 37558 -212
rect 35125 -275 35192 -274
rect 37557 -274 37558 -272
rect 37623 -274 37624 -210
rect 39634 -212 39694 103
rect 39989 -210 40056 -209
rect 39989 -212 39990 -210
rect 39634 -272 39990 -212
rect 37557 -275 37624 -274
rect 39989 -274 39990 -272
rect 40055 -274 40056 -210
rect 42066 -212 42126 722
rect 42421 -210 42488 -209
rect 42421 -212 42422 -210
rect 42066 -272 42422 -212
rect 39989 -275 40056 -274
rect 42421 -274 42422 -272
rect 42487 -274 42488 -210
rect 42421 -275 42488 -274
use switch  switch_0
timestamp 1757220954
transform 1 0 9282 0 1 46477
box 1296 -1584 3268 244
use switch  switch_2
timestamp 1757220954
transform 1 0 13226 0 1 46477
box 1296 -1584 3268 244
use switch  switch_3
timestamp 1757220954
transform 1 0 17170 0 1 46477
box 1296 -1584 3268 244
use switch  switch_4
timestamp 1757220954
transform 1 0 21114 0 1 46477
box 1296 -1584 3268 244
use switch  switch_5
timestamp 1757220954
transform 1 0 25058 0 1 46477
box 1296 -1584 3268 244
use switch  switch_6
timestamp 1757220954
transform 1 0 32946 0 1 46477
box 1296 -1584 3268 244
use switch  switch_7
timestamp 1757220954
transform 1 0 29002 0 1 46477
box 1296 -1584 3268 244
use switch  switch_8
timestamp 1757220954
transform 1 0 5338 0 1 46477
box 1296 -1584 3268 244
use unit_cap  unit_cap_0
timestamp 1757220954
transform 1 0 90 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_1
timestamp 1757220954
transform 1 0 90 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_2
timestamp 1757220954
transform 1 0 90 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_3
timestamp 1757220954
transform 1 0 90 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_4
timestamp 1757220954
transform 1 0 90 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_5
timestamp 1757220954
transform 1 0 90 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_6
timestamp 1757220954
transform 1 0 90 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_7
timestamp 1757220954
transform 1 0 90 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_8
timestamp 1757220954
transform 1 0 90 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_9
timestamp 1757220954
transform 1 0 90 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_10
timestamp 1757220954
transform 1 0 90 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_11
timestamp 1757220954
transform 1 0 90 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_12
timestamp 1757220954
transform 1 0 90 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_13
timestamp 1757220954
transform 1 0 90 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_14
timestamp 1757220954
transform 1 0 90 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_15
timestamp 1757220954
transform 1 0 90 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_16
timestamp 1757220954
transform 1 0 90 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_17
timestamp 1757220954
transform 1 0 90 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_18
timestamp 1757220954
transform 1 0 2522 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_19
timestamp 1757220954
transform 1 0 2522 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_20
timestamp 1757220954
transform 1 0 2522 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_21
timestamp 1757220954
transform 1 0 2522 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_22
timestamp 1757220954
transform 1 0 2522 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_23
timestamp 1757220954
transform 1 0 2522 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_24
timestamp 1757220954
transform 1 0 2522 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_25
timestamp 1757220954
transform 1 0 2522 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_26
timestamp 1757220954
transform 1 0 2522 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_27
timestamp 1757220954
transform 1 0 2522 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_28
timestamp 1757220954
transform 1 0 2522 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_29
timestamp 1757220954
transform 1 0 2522 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_30
timestamp 1757220954
transform 1 0 2522 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_31
timestamp 1757220954
transform 1 0 2522 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_32
timestamp 1757220954
transform 1 0 2522 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_33
timestamp 1757220954
transform 1 0 2522 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_34
timestamp 1757220954
transform 1 0 2522 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_35
timestamp 1757220954
transform 1 0 2522 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_36
timestamp 1757220954
transform 1 0 4954 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_37
timestamp 1757220954
transform 1 0 4954 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_38
timestamp 1757220954
transform 1 0 4954 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_39
timestamp 1757220954
transform 1 0 4954 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_40
timestamp 1757220954
transform 1 0 4954 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_41
timestamp 1757220954
transform 1 0 4954 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_42
timestamp 1757220954
transform 1 0 4954 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_43
timestamp 1757220954
transform 1 0 4954 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_44
timestamp 1757220954
transform 1 0 4954 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_45
timestamp 1757220954
transform 1 0 4954 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_46
timestamp 1757220954
transform 1 0 4954 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_47
timestamp 1757220954
transform 1 0 4954 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_48
timestamp 1757220954
transform 1 0 4954 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_49
timestamp 1757220954
transform 1 0 4954 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_50
timestamp 1757220954
transform 1 0 4954 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_51
timestamp 1757220954
transform 1 0 4954 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_52
timestamp 1757220954
transform 1 0 4954 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_53
timestamp 1757220954
transform 1 0 4954 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_54
timestamp 1757220954
transform 1 0 7386 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_55
timestamp 1757220954
transform 1 0 7386 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_56
timestamp 1757220954
transform 1 0 7386 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_57
timestamp 1757220954
transform 1 0 7386 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_58
timestamp 1757220954
transform 1 0 7386 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_59
timestamp 1757220954
transform 1 0 7386 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_60
timestamp 1757220954
transform 1 0 7386 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_61
timestamp 1757220954
transform 1 0 7386 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_62
timestamp 1757220954
transform 1 0 7386 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_63
timestamp 1757220954
transform 1 0 7386 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_64
timestamp 1757220954
transform 1 0 7386 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_65
timestamp 1757220954
transform 1 0 7386 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_66
timestamp 1757220954
transform 1 0 7386 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_67
timestamp 1757220954
transform 1 0 7386 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_68
timestamp 1757220954
transform 1 0 7386 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_69
timestamp 1757220954
transform 1 0 7386 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_70
timestamp 1757220954
transform 1 0 7386 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_71
timestamp 1757220954
transform 1 0 7386 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_72
timestamp 1757220954
transform 1 0 9818 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_73
timestamp 1757220954
transform 1 0 9818 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_74
timestamp 1757220954
transform 1 0 9818 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_75
timestamp 1757220954
transform 1 0 9818 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_76
timestamp 1757220954
transform 1 0 9818 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_77
timestamp 1757220954
transform 1 0 9818 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_78
timestamp 1757220954
transform 1 0 9818 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_79
timestamp 1757220954
transform 1 0 9818 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_80
timestamp 1757220954
transform 1 0 9818 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_81
timestamp 1757220954
transform 1 0 9818 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_82
timestamp 1757220954
transform 1 0 9818 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_83
timestamp 1757220954
transform 1 0 9818 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_84
timestamp 1757220954
transform 1 0 9818 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_85
timestamp 1757220954
transform 1 0 9818 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_86
timestamp 1757220954
transform 1 0 9818 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_87
timestamp 1757220954
transform 1 0 9818 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_88
timestamp 1757220954
transform 1 0 9818 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_89
timestamp 1757220954
transform 1 0 9818 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_90
timestamp 1757220954
transform 1 0 12250 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_91
timestamp 1757220954
transform 1 0 12250 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_92
timestamp 1757220954
transform 1 0 12250 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_93
timestamp 1757220954
transform 1 0 12250 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_94
timestamp 1757220954
transform 1 0 12250 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_95
timestamp 1757220954
transform 1 0 12250 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_96
timestamp 1757220954
transform 1 0 12250 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_97
timestamp 1757220954
transform 1 0 12250 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_98
timestamp 1757220954
transform 1 0 12250 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_99
timestamp 1757220954
transform 1 0 12250 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_100
timestamp 1757220954
transform 1 0 12250 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_101
timestamp 1757220954
transform 1 0 12250 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_102
timestamp 1757220954
transform 1 0 12250 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_103
timestamp 1757220954
transform 1 0 12250 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_104
timestamp 1757220954
transform 1 0 12250 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_105
timestamp 1757220954
transform 1 0 12250 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_106
timestamp 1757220954
transform 1 0 12250 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_107
timestamp 1757220954
transform 1 0 12250 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_108
timestamp 1757220954
transform 1 0 14682 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_109
timestamp 1757220954
transform 1 0 14682 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_110
timestamp 1757220954
transform 1 0 14682 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_111
timestamp 1757220954
transform 1 0 14682 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_112
timestamp 1757220954
transform 1 0 14682 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_113
timestamp 1757220954
transform 1 0 14682 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_114
timestamp 1757220954
transform 1 0 14682 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_115
timestamp 1757220954
transform 1 0 14682 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_116
timestamp 1757220954
transform 1 0 14682 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_117
timestamp 1757220954
transform 1 0 14682 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_118
timestamp 1757220954
transform 1 0 14682 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_119
timestamp 1757220954
transform 1 0 14682 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_120
timestamp 1757220954
transform 1 0 14682 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_121
timestamp 1757220954
transform 1 0 14682 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_122
timestamp 1757220954
transform 1 0 14682 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_123
timestamp 1757220954
transform 1 0 14682 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_124
timestamp 1757220954
transform 1 0 14682 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_125
timestamp 1757220954
transform 1 0 14682 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_126
timestamp 1757220954
transform 1 0 17114 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_127
timestamp 1757220954
transform 1 0 17114 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_128
timestamp 1757220954
transform 1 0 17114 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_129
timestamp 1757220954
transform 1 0 17114 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_130
timestamp 1757220954
transform 1 0 17114 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_131
timestamp 1757220954
transform 1 0 17114 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_132
timestamp 1757220954
transform 1 0 17114 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_133
timestamp 1757220954
transform 1 0 17114 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_134
timestamp 1757220954
transform 1 0 17114 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_135
timestamp 1757220954
transform 1 0 17114 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_136
timestamp 1757220954
transform 1 0 17114 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_137
timestamp 1757220954
transform 1 0 17114 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_138
timestamp 1757220954
transform 1 0 17114 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_139
timestamp 1757220954
transform 1 0 17114 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_140
timestamp 1757220954
transform 1 0 17114 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_141
timestamp 1757220954
transform 1 0 17114 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_142
timestamp 1757220954
transform 1 0 17114 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_143
timestamp 1757220954
transform 1 0 17114 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_144
timestamp 1757220954
transform 1 0 19546 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_145
timestamp 1757220954
transform 1 0 19546 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_146
timestamp 1757220954
transform 1 0 19546 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_147
timestamp 1757220954
transform 1 0 19546 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_148
timestamp 1757220954
transform 1 0 19546 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_149
timestamp 1757220954
transform 1 0 19546 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_150
timestamp 1757220954
transform 1 0 19546 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_151
timestamp 1757220954
transform 1 0 19546 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_152
timestamp 1757220954
transform 1 0 19546 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_154
timestamp 1757220954
transform 1 0 19546 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_155
timestamp 1757220954
transform 1 0 19546 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_156
timestamp 1757220954
transform 1 0 19546 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_157
timestamp 1757220954
transform 1 0 19546 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_158
timestamp 1757220954
transform 1 0 19546 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_159
timestamp 1757220954
transform 1 0 19546 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_160
timestamp 1757220954
transform 1 0 19546 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_161
timestamp 1757220954
transform 1 0 19546 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_162
timestamp 1757220954
transform 1 0 21978 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_163
timestamp 1757220954
transform 1 0 21978 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_164
timestamp 1757220954
transform 1 0 21978 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_165
timestamp 1757220954
transform 1 0 21978 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_166
timestamp 1757220954
transform 1 0 21978 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_167
timestamp 1757220954
transform 1 0 21978 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_168
timestamp 1757220954
transform 1 0 21978 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_169
timestamp 1757220954
transform 1 0 21978 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_170
timestamp 1757220954
transform 1 0 21978 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_171
timestamp 1757220954
transform 1 0 21978 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_172
timestamp 1757220954
transform 1 0 21978 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_173
timestamp 1757220954
transform 1 0 21978 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_174
timestamp 1757220954
transform 1 0 21978 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_175
timestamp 1757220954
transform 1 0 21978 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_176
timestamp 1757220954
transform 1 0 21978 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_177
timestamp 1757220954
transform 1 0 21978 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_178
timestamp 1757220954
transform 1 0 21978 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_179
timestamp 1757220954
transform 1 0 21978 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_180
timestamp 1757220954
transform 1 0 24410 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_181
timestamp 1757220954
transform 1 0 24410 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_182
timestamp 1757220954
transform 1 0 24410 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_183
timestamp 1757220954
transform 1 0 24410 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_184
timestamp 1757220954
transform 1 0 24410 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_185
timestamp 1757220954
transform 1 0 24410 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_186
timestamp 1757220954
transform 1 0 24410 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_187
timestamp 1757220954
transform 1 0 24410 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_188
timestamp 1757220954
transform 1 0 24410 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_189
timestamp 1757220954
transform 1 0 24410 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_190
timestamp 1757220954
transform 1 0 24410 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_191
timestamp 1757220954
transform 1 0 24410 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_192
timestamp 1757220954
transform 1 0 24410 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_193
timestamp 1757220954
transform 1 0 24410 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_194
timestamp 1757220954
transform 1 0 24410 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_195
timestamp 1757220954
transform 1 0 24410 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_196
timestamp 1757220954
transform 1 0 24410 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_197
timestamp 1757220954
transform 1 0 24410 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_198
timestamp 1757220954
transform 1 0 26842 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_199
timestamp 1757220954
transform 1 0 26842 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_200
timestamp 1757220954
transform 1 0 26842 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_201
timestamp 1757220954
transform 1 0 26842 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_202
timestamp 1757220954
transform 1 0 26842 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_203
timestamp 1757220954
transform 1 0 26842 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_204
timestamp 1757220954
transform 1 0 26842 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_205
timestamp 1757220954
transform 1 0 26842 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_206
timestamp 1757220954
transform 1 0 26842 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_207
timestamp 1757220954
transform 1 0 26842 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_208
timestamp 1757220954
transform 1 0 26842 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_209
timestamp 1757220954
transform 1 0 26842 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_210
timestamp 1757220954
transform 1 0 26842 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_211
timestamp 1757220954
transform 1 0 26842 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_212
timestamp 1757220954
transform 1 0 26842 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_213
timestamp 1757220954
transform 1 0 26842 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_214
timestamp 1757220954
transform 1 0 26842 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_215
timestamp 1757220954
transform 1 0 26842 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_216
timestamp 1757220954
transform 1 0 29274 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_217
timestamp 1757220954
transform 1 0 29274 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_218
timestamp 1757220954
transform 1 0 29274 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_219
timestamp 1757220954
transform 1 0 29274 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_220
timestamp 1757220954
transform 1 0 29274 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_221
timestamp 1757220954
transform 1 0 29274 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_222
timestamp 1757220954
transform 1 0 29274 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_223
timestamp 1757220954
transform 1 0 29274 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_224
timestamp 1757220954
transform 1 0 29274 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_225
timestamp 1757220954
transform 1 0 29274 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_226
timestamp 1757220954
transform 1 0 29274 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_227
timestamp 1757220954
transform 1 0 29274 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_228
timestamp 1757220954
transform 1 0 29274 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_229
timestamp 1757220954
transform 1 0 29274 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_230
timestamp 1757220954
transform 1 0 29274 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_231
timestamp 1757220954
transform 1 0 29274 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_232
timestamp 1757220954
transform 1 0 29274 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_233
timestamp 1757220954
transform 1 0 29274 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_234
timestamp 1757220954
transform 1 0 31706 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_235
timestamp 1757220954
transform 1 0 31706 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_236
timestamp 1757220954
transform 1 0 31706 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_237
timestamp 1757220954
transform 1 0 31706 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_238
timestamp 1757220954
transform 1 0 31706 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_239
timestamp 1757220954
transform 1 0 31706 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_240
timestamp 1757220954
transform 1 0 31706 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_241
timestamp 1757220954
transform 1 0 31706 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_242
timestamp 1757220954
transform 1 0 31706 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_243
timestamp 1757220954
transform 1 0 31706 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_244
timestamp 1757220954
transform 1 0 31706 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_245
timestamp 1757220954
transform 1 0 31706 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_246
timestamp 1757220954
transform 1 0 31706 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_247
timestamp 1757220954
transform 1 0 31706 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_248
timestamp 1757220954
transform 1 0 31706 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_249
timestamp 1757220954
transform 1 0 31706 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_250
timestamp 1757220954
transform 1 0 31706 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_251
timestamp 1757220954
transform 1 0 31706 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_252
timestamp 1757220954
transform 1 0 34138 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_253
timestamp 1757220954
transform 1 0 34138 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_254
timestamp 1757220954
transform 1 0 34138 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_255
timestamp 1757220954
transform 1 0 34138 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_256
timestamp 1757220954
transform 1 0 34138 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_257
timestamp 1757220954
transform 1 0 34138 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_258
timestamp 1757220954
transform 1 0 34138 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_259
timestamp 1757220954
transform 1 0 34138 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_260
timestamp 1757220954
transform 1 0 34138 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_261
timestamp 1757220954
transform 1 0 34138 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_262
timestamp 1757220954
transform 1 0 34138 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_263
timestamp 1757220954
transform 1 0 34138 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_264
timestamp 1757220954
transform 1 0 34138 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_265
timestamp 1757220954
transform 1 0 34138 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_266
timestamp 1757220954
transform 1 0 34138 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_267
timestamp 1757220954
transform 1 0 34138 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_268
timestamp 1757220954
transform 1 0 34138 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_269
timestamp 1757220954
transform 1 0 34138 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_270
timestamp 1757220954
transform 1 0 36570 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_271
timestamp 1757220954
transform 1 0 36570 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_272
timestamp 1757220954
transform 1 0 36570 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_273
timestamp 1757220954
transform 1 0 36570 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_274
timestamp 1757220954
transform 1 0 36570 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_275
timestamp 1757220954
transform 1 0 36570 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_276
timestamp 1757220954
transform 1 0 36570 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_277
timestamp 1757220954
transform 1 0 36570 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_278
timestamp 1757220954
transform 1 0 36570 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_279
timestamp 1757220954
transform 1 0 36570 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_280
timestamp 1757220954
transform 1 0 36570 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_281
timestamp 1757220954
transform 1 0 36570 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_282
timestamp 1757220954
transform 1 0 36570 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_283
timestamp 1757220954
transform 1 0 36570 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_284
timestamp 1757220954
transform 1 0 36570 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_285
timestamp 1757220954
transform 1 0 36570 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_286
timestamp 1757220954
transform 1 0 36570 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_287
timestamp 1757220954
transform 1 0 36570 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_288
timestamp 1757220954
transform 1 0 39002 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_289
timestamp 1757220954
transform 1 0 39002 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_290
timestamp 1757220954
transform 1 0 39002 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_291
timestamp 1757220954
transform 1 0 39002 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_292
timestamp 1757220954
transform 1 0 39002 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_293
timestamp 1757220954
transform 1 0 39002 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_294
timestamp 1757220954
transform 1 0 39002 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_295
timestamp 1757220954
transform 1 0 39002 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_296
timestamp 1757220954
transform 1 0 39002 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_297
timestamp 1757220954
transform 1 0 39002 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_298
timestamp 1757220954
transform 1 0 39002 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_299
timestamp 1757220954
transform 1 0 39002 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_300
timestamp 1757220954
transform 1 0 39002 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_301
timestamp 1757220954
transform 1 0 39002 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_302
timestamp 1757220954
transform 1 0 39002 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_303
timestamp 1757220954
transform 1 0 39002 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_304
timestamp 1757220954
transform 1 0 39002 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_305
timestamp 1757220954
transform 1 0 39002 0 1 43433
box -90 -1904 1414 -398
use unit_cap  unit_cap_306
timestamp 1757220954
transform 1 0 41434 0 1 1903
box -90 -1904 1414 -398
use unit_cap  unit_cap_307
timestamp 1757220954
transform 1 0 41434 0 1 4335
box -90 -1904 1414 -398
use unit_cap  unit_cap_308
timestamp 1757220954
transform 1 0 41434 0 1 6767
box -90 -1904 1414 -398
use unit_cap  unit_cap_309
timestamp 1757220954
transform 1 0 41434 0 1 9199
box -90 -1904 1414 -398
use unit_cap  unit_cap_310
timestamp 1757220954
transform 1 0 41434 0 1 11631
box -90 -1904 1414 -398
use unit_cap  unit_cap_311
timestamp 1757220954
transform 1 0 41434 0 1 14063
box -90 -1904 1414 -398
use unit_cap  unit_cap_312
timestamp 1757220954
transform 1 0 41434 0 1 16495
box -90 -1904 1414 -398
use unit_cap  unit_cap_313
timestamp 1757220954
transform 1 0 41434 0 1 18927
box -90 -1904 1414 -398
use unit_cap  unit_cap_314
timestamp 1757220954
transform 1 0 41434 0 1 21359
box -90 -1904 1414 -398
use unit_cap  unit_cap_315
timestamp 1757220954
transform 1 0 41434 0 1 23977
box -90 -1904 1414 -398
use unit_cap  unit_cap_316
timestamp 1757220954
transform 1 0 41434 0 1 26409
box -90 -1904 1414 -398
use unit_cap  unit_cap_317
timestamp 1757220954
transform 1 0 41434 0 1 28841
box -90 -1904 1414 -398
use unit_cap  unit_cap_318
timestamp 1757220954
transform 1 0 41434 0 1 31273
box -90 -1904 1414 -398
use unit_cap  unit_cap_319
timestamp 1757220954
transform 1 0 41434 0 1 33705
box -90 -1904 1414 -398
use unit_cap  unit_cap_320
timestamp 1757220954
transform 1 0 41434 0 1 36137
box -90 -1904 1414 -398
use unit_cap  unit_cap_321
timestamp 1757220954
transform 1 0 41434 0 1 38569
box -90 -1904 1414 -398
use unit_cap  unit_cap_322
timestamp 1757220954
transform 1 0 41434 0 1 41001
box -90 -1904 1414 -398
use unit_cap  unit_cap_323
timestamp 1757220954
transform 1 0 41434 0 1 43433
box -90 -1904 1414 -398
<< labels >>
flabel space 2468 2468 3900 3900 0 FreeSans 8000 0 0 0 7
flabel space 2468 7332 3900 8764 0 FreeSans 8000 0 0 0 7
flabel space 2468 12196 3900 13628 0 FreeSans 8000 0 0 0 7
flabel space 2468 17060 3900 18492 0 FreeSans 8000 0 0 0 7
flabel space 4900 2468 6332 3900 0 FreeSans 8000 0 0 0 6
flabel space 2468 4900 3900 6332 0 FreeSans 8000 0 0 0 5
flabel space 2468 9764 3900 11196 0 FreeSans 8000 0 0 0 5
flabel space 2468 14628 3900 16060 0 FreeSans 8000 0 0 0 3
flabel space 2468 19492 3900 20924 0 FreeSans 8000 0 0 0 2
flabel space 7332 19492 8764 20924 0 FreeSans 8000 0 0 0 4
flabel space 17060 19492 18492 20924 0 FreeSans 8000 0 0 0 4
flabel space 7332 14628 8764 16060 0 FreeSans 8000 0 0 0 4
flabel space 17024 14592 18528 16096 0 FreeSans 8000 0 0 0 4
flabel space 26788 19492 28220 20924 0 FreeSans 8000 0 0 0 4
flabel space 26788 14628 28220 16060 0 FreeSans 8000 0 0 0 4
flabel space 36516 19492 37948 20924 0 FreeSans 8000 0 0 0 4
flabel space 36516 14628 37948 16060 0 FreeSans 8000 0 0 0 4
flabel space 12196 14628 13628 16060 0 FreeSans 8000 0 0 0 3
flabel space 21924 14628 23356 16060 0 FreeSans 8000 0 0 0 3
flabel space 31652 14628 33084 16060 0 FreeSans 8000 0 0 0 3
flabel space 31652 19492 33084 20924 0 FreeSans 8000 0 0 0 2
flabel space 12196 19492 13628 20924 0 FreeSans 8000 0 0 0 1
flabel space 21924 19492 23356 20924 0 FreeSans 8000 0 0 0 0
flabel space 38948 19492 40380 20924 0 FreeSans 8000 0 0 0 7
flabel space 36516 17060 37948 18492 0 FreeSans 8000 0 0 0 7
flabel space 38948 14628 40380 16060 0 FreeSans 8000 0 0 0 7
flabel space 34084 14628 35516 16060 0 FreeSans 8000 0 0 0 7
flabel space 34084 19492 35516 20924 0 FreeSans 8000 0 0 0 7
flabel space 31652 17060 33084 18492 0 FreeSans 8000 0 0 0 7
flabel space 29220 14628 30652 16060 0 FreeSans 8000 0 0 0 7
flabel space 29220 19492 30652 20924 0 FreeSans 8000 0 0 0 7
flabel space 26788 17060 28220 18492 0 FreeSans 8000 0 0 0 7
flabel space 24356 14628 25788 16060 0 FreeSans 8000 0 0 0 7
flabel space 24356 19492 25788 20924 0 FreeSans 8000 0 0 0 7
flabel space 21924 17060 23356 18492 0 FreeSans 8000 0 0 0 7
flabel space 19492 19492 20924 20924 0 FreeSans 8000 0 0 0 7
flabel space 14628 19492 16060 20924 0 FreeSans 8000 0 0 0 7
flabel space 9764 19492 11196 20924 0 FreeSans 8000 0 0 0 7
flabel space 4900 19492 6332 20924 0 FreeSans 8000 0 0 0 7
flabel space 7332 17060 8764 18492 0 FreeSans 8000 0 0 0 7
flabel space 12196 17060 13628 18492 0 FreeSans 8000 0 0 0 7
flabel space 17060 17060 18492 18492 0 FreeSans 8000 0 0 0 7
flabel space 19492 14628 20924 16060 0 FreeSans 8000 0 0 0 7
flabel space 14628 14628 16060 16060 0 FreeSans 8000 0 0 0 7
flabel space 9764 14628 11196 16060 0 FreeSans 8000 0 0 0 7
flabel space 4900 14628 6332 16060 0 FreeSans 8000 0 0 0 7
flabel space 7332 12196 8764 13628 0 FreeSans 8000 0 0 0 7
flabel space 4900 9764 6332 11196 0 FreeSans 8000 0 0 0 7
flabel space 7332 7332 8764 8764 0 FreeSans 8000 0 0 0 7
flabel space 9764 9764 11196 11196 0 FreeSans 8000 0 0 0 7
flabel space 12196 12196 13628 13628 0 FreeSans 8000 0 0 0 7
flabel space 17060 12196 18492 13628 0 FreeSans 8000 0 0 0 7
flabel space 21924 12196 23356 13628 0 FreeSans 8000 0 0 0 7
flabel space 24356 9764 25788 11196 0 FreeSans 8000 0 0 0 7
flabel space 19492 9764 20924 11196 0 FreeSans 8000 0 0 0 7
flabel space 14628 9764 16060 11196 0 FreeSans 8000 0 0 0 7
flabel space 17060 7332 18492 8764 0 FreeSans 8000 0 0 0 7
flabel space 12196 7332 13628 8764 0 FreeSans 8000 0 0 0 7
flabel space 26788 12196 28220 13628 0 FreeSans 8000 0 0 0 7
flabel space 31652 12196 33084 13628 0 FreeSans 8000 0 0 0 7
flabel space 29220 9764 30652 11196 0 FreeSans 8000 0 0 0 7
flabel space 36516 12196 37948 13628 0 FreeSans 8000 0 0 0 7
flabel space 38948 9764 40380 11196 0 FreeSans 8000 0 0 0 7
flabel space 34084 9764 35516 11196 0 FreeSans 8000 0 0 0 7
flabel space 36516 7332 37948 8764 0 FreeSans 8000 0 0 0 7
flabel space 38948 4900 40380 6332 0 FreeSans 8000 0 0 0 7
flabel space 34084 4900 35516 6332 0 FreeSans 8000 0 0 0 7
flabel space 29220 4900 30652 6332 0 FreeSans 8000 0 0 0 7
flabel space 31652 7332 33084 8764 0 FreeSans 8000 0 0 0 7
flabel space 26788 7332 28220 8764 0 FreeSans 8000 0 0 0 7
flabel space 24356 4900 25788 6332 0 FreeSans 8000 0 0 0 7
flabel space 21924 7332 23356 8764 0 FreeSans 8000 0 0 0 7
flabel space 19492 4900 20924 6332 0 FreeSans 8000 0 0 0 7
flabel space 14628 4900 16060 6332 0 FreeSans 8000 0 0 0 7
flabel space 9764 4900 11196 6332 0 FreeSans 8000 0 0 0 7
flabel space 4900 4900 6332 6332 0 FreeSans 8000 0 0 0 7
flabel space 7332 2468 8764 3900 0 FreeSans 8000 0 0 0 7
flabel space 12196 2468 13628 3900 0 FreeSans 8000 0 0 0 7
flabel space 17060 2468 18492 3900 0 FreeSans 8000 0 0 0 7
flabel space 21924 2468 23356 3900 0 FreeSans 8000 0 0 0 7
flabel space 26788 2468 28220 3900 0 FreeSans 8000 0 0 0 7
flabel space 31652 2468 33084 3900 0 FreeSans 8000 0 0 0 7
flabel space 36516 2468 37948 3900 0 FreeSans 8000 0 0 0 7
flabel space 38948 2468 40380 3900 0 FreeSans 8000 0 0 0 6
flabel space 38948 7332 40380 8764 0 FreeSans 8000 0 0 0 6
flabel space 38948 12196 40380 13628 0 FreeSans 8000 0 0 0 6
flabel space 38948 17060 40380 18492 0 FreeSans 8000 0 0 0 6
flabel space 34084 17060 35516 18492 0 FreeSans 8000 0 0 0 6
flabel space 29220 17060 30652 18492 0 FreeSans 8000 0 0 0 6
flabel space 24356 17060 25788 18492 0 FreeSans 8000 0 0 0 6
flabel space 19492 17060 20924 18492 0 FreeSans 8000 0 0 0 6
flabel space 14628 17060 16060 18492 0 FreeSans 8000 0 0 0 6
flabel space 9764 17060 11196 18492 0 FreeSans 8000 0 0 0 6
flabel space 4900 17060 6332 18492 0 FreeSans 8000 0 0 0 6
flabel space 4900 12196 6332 13628 0 FreeSans 8000 0 0 0 6
flabel space 9764 12196 11196 13628 0 FreeSans 8000 0 0 0 6
flabel space 14628 12196 16060 13628 0 FreeSans 8000 0 0 0 6
flabel space 19492 12196 20924 13628 0 FreeSans 8000 0 0 0 6
flabel space 24356 12196 25788 13628 0 FreeSans 8000 0 0 0 6
flabel space 29220 12196 30652 13628 0 FreeSans 8000 0 0 0 6
flabel space 34084 12196 35516 13628 0 FreeSans 8000 0 0 0 6
flabel space 34084 7332 35516 8764 0 FreeSans 8000 0 0 0 6
flabel space 34084 2468 35516 3900 0 FreeSans 8000 0 0 0 6
flabel space 29220 2468 30652 3900 0 FreeSans 8000 0 0 0 6
flabel space 29220 7332 30652 8764 0 FreeSans 8000 0 0 0 6
flabel space 24356 2468 25788 3900 0 FreeSans 8000 0 0 0 6
flabel space 24356 7332 25788 8764 0 FreeSans 8000 0 0 0 6
flabel space 19492 7332 20924 8764 0 FreeSans 8000 0 0 0 6
flabel space 19492 2468 20924 3900 0 FreeSans 8000 0 0 0 6
flabel space 14628 2468 16060 3900 0 FreeSans 8000 0 0 0 6
flabel space 14628 7332 16060 8764 0 FreeSans 8000 0 0 0 6
flabel space 9728 2432 11232 3936 0 FreeSans 8000 0 0 0 6
flabel space 9764 7332 11196 8764 0 FreeSans 8000 0 0 0 6
flabel space 4900 7332 6332 8764 0 FreeSans 8000 0 0 0 6
flabel space 7332 9764 8764 11196 0 FreeSans 8000 0 0 0 5
flabel space 7332 4900 8764 6332 0 FreeSans 8000 0 0 0 5
flabel space 12196 4900 13628 6332 0 FreeSans 8000 0 0 0 5
flabel space 12196 9764 13628 11196 0 FreeSans 8000 0 0 0 5
flabel space 17060 9764 18492 11196 0 FreeSans 8000 0 0 0 5
flabel space 21924 9764 23356 11196 0 FreeSans 8000 0 0 0 5
flabel space 26788 9764 28220 11196 0 FreeSans 8000 0 0 0 5
flabel space 31652 9764 33084 11196 0 FreeSans 8000 0 0 0 5
flabel space 36516 9764 37948 11196 0 FreeSans 8000 0 0 0 5
flabel space 36516 4900 37948 6332 0 FreeSans 8000 0 0 0 5
flabel space 31652 4900 33084 6332 0 FreeSans 8000 0 0 0 5
flabel space 26788 4900 28220 6332 0 FreeSans 8000 0 0 0 5
flabel space 21924 4900 23356 6332 0 FreeSans 8000 0 0 0 5
flabel space 17060 4900 18492 6332 0 FreeSans 8000 0 0 0 5
flabel space 2468 22110 3900 23542 0 FreeSans 8000 0 0 0 7
flabel space 2468 26974 3900 28406 0 FreeSans 8000 0 0 0 7
flabel space 2468 31838 3900 33270 0 FreeSans 8000 0 0 0 7
flabel space 2468 36702 3900 38134 0 FreeSans 8000 0 0 0 7
flabel space 2468 39134 3900 40566 0 FreeSans 8000 0 0 0 6
flabel space 4900 36702 6332 38134 0 FreeSans 8000 0 0 0 5
flabel space 2468 34270 3900 35702 0 FreeSans 8000 0 0 0 6
flabel space 4900 31838 6332 33270 0 FreeSans 8000 0 0 0 5
flabel space 2468 29406 3900 30838 0 FreeSans 8000 0 0 0 6
flabel space 2468 24542 3900 25974 0 FreeSans 8000 0 0 0 6
flabel space 9764 36702 11196 38134 0 FreeSans 8000 0 0 0 5
flabel space 9764 31838 11196 33270 0 FreeSans 8000 0 0 0 5
flabel space 14628 31838 16060 33270 0 FreeSans 8000 0 0 0 5
flabel space 19492 31838 20924 33270 0 FreeSans 8000 0 0 0 5
flabel space 19492 36702 20924 38134 0 FreeSans 8000 0 0 0 5
flabel space 14628 36702 16060 38134 0 FreeSans 8000 0 0 0 5
flabel space 24356 31838 25788 33270 0 FreeSans 8000 0 0 0 5
flabel space 24356 36702 25788 38134 0 FreeSans 8000 0 0 0 5
flabel space 29220 36702 30652 38134 0 FreeSans 8000 0 0 0 5
flabel space 34084 36702 35516 38134 0 FreeSans 8000 0 0 0 5
flabel space 38948 36702 40380 38134 0 FreeSans 8000 0 0 0 5
flabel space 38948 31838 40380 33270 0 FreeSans 8000 0 0 0 5
flabel space 34084 31838 35516 33270 0 FreeSans 8000 0 0 0 5
flabel space 29220 31838 30652 33270 0 FreeSans 8000 0 0 0 5
flabel space 4900 39134 6332 40566 0 FreeSans 8000 0 0 0 7
flabel space 9764 39134 11196 40566 0 FreeSans 8000 0 0 0 7
flabel space 14628 39134 16060 40566 0 FreeSans 8000 0 0 0 7
flabel space 19492 39134 20924 40566 0 FreeSans 8000 0 0 0 7
flabel space 24356 39134 25788 40566 0 FreeSans 8000 0 0 0 7
flabel space 29220 39134 30652 40566 0 FreeSans 8000 0 0 0 7
flabel space 34084 39134 35516 40566 0 FreeSans 8000 0 0 0 7
flabel space 38948 39134 40380 40566 0 FreeSans 8000 0 0 0 7
flabel space 36516 36702 37948 38134 0 FreeSans 8000 0 0 0 7
flabel space 38948 34270 40380 35702 0 FreeSans 8000 0 0 0 7
flabel space 34084 34270 35516 35702 0 FreeSans 8000 0 0 0 7
flabel space 31652 36702 33084 38134 0 FreeSans 8000 0 0 0 7
flabel space 29220 34270 30652 35702 0 FreeSans 8000 0 0 0 7
flabel space 26788 36702 28220 38134 0 FreeSans 8000 0 0 0 7
flabel space 24356 34270 25788 35702 0 FreeSans 8000 0 0 0 7
flabel space 21924 36702 23356 38134 0 FreeSans 8000 0 0 0 7
flabel space 19492 34270 20924 35702 0 FreeSans 8000 0 0 0 7
flabel space 17060 36702 18492 38134 0 FreeSans 8000 0 0 0 7
flabel space 14628 34270 16060 35702 0 FreeSans 8000 0 0 0 7
flabel space 12196 36702 13628 38134 0 FreeSans 8000 0 0 0 7
flabel space 7332 36702 8764 38134 0 FreeSans 8000 0 0 0 7
flabel space 4900 34270 6332 35702 0 FreeSans 8000 0 0 0 7
flabel space 7332 31838 8764 33270 0 FreeSans 8000 0 0 0 7
flabel space 12196 31838 13628 33270 0 FreeSans 8000 0 0 0 7
flabel space 9764 34270 11196 35702 0 FreeSans 8000 0 0 0 7
flabel space 17060 31838 18492 33270 0 FreeSans 8000 0 0 0 7
flabel space 21924 31838 23356 33270 0 FreeSans 8000 0 0 0 7
flabel space 26788 31838 28220 33270 0 FreeSans 8000 0 0 0 7
flabel space 36516 31838 37948 33270 0 FreeSans 8000 0 0 0 7
flabel space 31652 31838 33084 33270 0 FreeSans 8000 0 0 0 7
flabel space 4900 26974 6332 28406 0 FreeSans 8000 0 0 0 4
flabel space 14628 26974 16060 28406 0 FreeSans 8000 0 0 0 4
flabel space 4900 22110 6332 23542 0 FreeSans 8000 0 0 0 4
flabel space 14628 22110 16060 23542 0 FreeSans 8000 0 0 0 4
flabel space 24356 22110 25788 23542 0 FreeSans 8000 0 0 0 4
flabel space 24356 26974 25788 28406 0 FreeSans 8000 0 0 0 4
flabel space 34084 26974 35516 28406 0 FreeSans 8000 0 0 0 4
flabel space 34084 22110 35516 23542 0 FreeSans 8000 0 0 0 4
flabel space 29220 26974 30652 28406 0 FreeSans 8000 0 0 0 3
flabel space 38948 26974 40380 28406 0 FreeSans 8000 0 0 0 3
flabel space 19492 26974 20924 28406 0 FreeSans 8000 0 0 0 3
flabel space 9764 26974 11196 28406 0 FreeSans 8000 0 0 0 3
flabel space 9764 22110 11196 23542 0 FreeSans 8000 0 0 0 2
flabel space 38948 22110 40380 23542 0 FreeSans 8000 0 0 0 2
flabel space 29220 22110 30652 23542 0 FreeSans 8000 0 0 0 1
flabel space 19492 22110 20924 23542 0 FreeSans 8000 0 0 0 D
flabel space 4900 29406 6332 30838 0 FreeSans 8000 0 0 0 7
flabel space 9764 29406 11196 30838 0 FreeSans 8000 0 0 0 7
flabel space 7332 26974 8764 28406 0 FreeSans 8000 0 0 0 7
flabel space 12196 26974 13628 28406 0 FreeSans 8000 0 0 0 7
flabel space 14628 29406 16060 30838 0 FreeSans 8000 0 0 0 7
flabel space 17060 26974 18492 28406 0 FreeSans 8000 0 0 0 7
flabel space 19492 29406 20924 30838 0 FreeSans 8000 0 0 0 7
flabel space 21924 26974 23356 28406 0 FreeSans 8000 0 0 0 7
flabel space 24356 29406 25788 30838 0 FreeSans 8000 0 0 0 7
flabel space 26788 26974 28220 28406 0 FreeSans 8000 0 0 0 7
flabel space 31652 26974 33084 28406 0 FreeSans 8000 0 0 0 7
flabel space 36516 26974 37948 28406 0 FreeSans 8000 0 0 0 7
flabel space 38948 29406 40380 30838 0 FreeSans 8000 0 0 0 7
flabel space 34084 29406 35516 30838 0 FreeSans 8000 0 0 0 7
flabel space 29220 29406 30652 30838 0 FreeSans 8000 0 0 0 7
flabel space 4900 24542 6332 25974 0 FreeSans 8000 0 0 0 7
flabel space 9764 24542 11196 25974 0 FreeSans 8000 0 0 0 7
flabel space 14628 24542 16060 25974 0 FreeSans 8000 0 0 0 7
flabel space 19492 24542 20924 25974 0 FreeSans 8000 0 0 0 7
flabel space 24356 24542 25788 25974 0 FreeSans 8000 0 0 0 7
flabel space 21924 22110 23356 23542 0 FreeSans 8000 0 0 0 7
flabel space 26788 22110 28220 23542 0 FreeSans 8000 0 0 0 7
flabel space 29220 24542 30652 25974 0 FreeSans 8000 0 0 0 7
flabel space 31652 22110 33084 23542 0 FreeSans 8000 0 0 0 7
flabel space 34084 24542 35516 25974 0 FreeSans 8000 0 0 0 7
flabel space 36516 22110 37948 23542 0 FreeSans 8000 0 0 0 7
flabel space 38948 24542 40380 25974 0 FreeSans 8000 0 0 0 7
flabel space 17060 22110 18492 23542 0 FreeSans 8000 0 0 0 7
flabel space 12196 22110 13628 23542 0 FreeSans 8000 0 0 0 7
flabel space 7332 22110 8764 23542 0 FreeSans 8000 0 0 0 7
flabel space 7332 39134 8764 40566 0 FreeSans 8000 0 0 0 6
flabel space 12196 39134 13628 40566 0 FreeSans 8000 0 0 0 6
flabel space 7332 34270 8764 35702 0 FreeSans 8000 0 0 0 6
flabel space 7332 29406 8764 30838 0 FreeSans 8000 0 0 0 6
flabel space 7332 24542 8764 25974 0 FreeSans 8000 0 0 0 6
flabel space 12196 24542 13628 25974 0 FreeSans 8000 0 0 0 6
flabel space 17060 24542 18492 25974 0 FreeSans 8000 0 0 0 6
flabel space 21924 24542 23356 25974 0 FreeSans 8000 0 0 0 6
flabel space 26788 24542 28220 25974 0 FreeSans 8000 0 0 0 6
flabel space 36516 24542 37948 25974 0 FreeSans 8000 0 0 0 6
flabel space 31652 24542 33084 25974 0 FreeSans 8000 0 0 0 6
flabel space 36516 29406 37948 30838 0 FreeSans 8000 0 0 0 6
flabel space 36516 34270 37948 35702 0 FreeSans 8000 0 0 0 6
flabel space 36516 39134 37948 40566 0 FreeSans 8000 0 0 0 6
flabel space 31652 39134 33084 40566 0 FreeSans 8000 0 0 0 6
flabel space 31652 34270 33084 35702 0 FreeSans 8000 0 0 0 6
flabel space 31652 29406 33084 30838 0 FreeSans 8000 0 0 0 6
flabel space 26788 29406 28220 30838 0 FreeSans 8000 0 0 0 6
flabel space 26788 34270 28220 35702 0 FreeSans 8000 0 0 0 6
flabel space 26788 39134 28220 40566 0 FreeSans 8000 0 0 0 6
flabel space 21924 39134 23356 40566 0 FreeSans 8000 0 0 0 6
flabel space 21888 34234 23392 35738 0 FreeSans 8000 0 0 0 6
flabel space 21924 29406 23356 30838 0 FreeSans 8000 0 0 0 6
flabel space 17060 29406 18492 30838 0 FreeSans 8000 0 0 0 6
flabel space 12196 29406 13628 30838 0 FreeSans 8000 0 0 0 6
flabel space 12196 34270 13628 35702 0 FreeSans 8000 0 0 0 6
flabel space 17060 34270 18492 35702 0 FreeSans 8000 0 0 0 6
flabel space 17060 39134 18492 40566 0 FreeSans 8000 0 0 0 6
flabel metal4 2432 39820 40416 39880 0 FreeSans 160 0 0 0 OUT
port 8 nsew
flabel metal1 420 44893 41706 44939 0 FreeSans 160 0 0 0 GND
port 9 nsew
flabel metal1 6634 46675 36214 46721 0 FreeSans 160 0 0 0 VDD
port 10 nsew
flabel metal1 7597 45865 8257 45911 0 FreeSans 160 0 0 0 b0
port 11 nsew
flabel metal1 11541 45865 12201 45911 0 FreeSans 160 0 0 0 b1
port 12 nsew
flabel metal1 15485 45865 16145 45911 0 FreeSans 160 0 0 0 b2
port 13 nsew
flabel metal1 19429 45865 20089 45911 0 FreeSans 160 0 0 0 b3
port 14 nsew
flabel metal1 23373 45865 24033 45911 0 FreeSans 160 0 0 0 b4
port 15 nsew
flabel metal1 27317 45865 27977 45911 0 FreeSans 160 0 0 0 b5
port 16 nsew
flabel metal1 31261 45865 31921 45911 0 FreeSans 160 0 0 0 b6
port 17 nsew
flabel metal1 35205 45865 35865 45911 0 FreeSans 160 0 0 0 b7
port 18 nsew
<< end >>
