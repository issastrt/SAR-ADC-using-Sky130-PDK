** sch_path: /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_21-28-41/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.697058823500 8.5u 0.697058823500 8.500001u 0.698823529375 17u 0.698823529375 17.000001u 0.700588235250 25.5u
+ 0.700588235250 25.500001u 0.702352941125 34u 0.702352941125 34.000001u 0.704117647000 42.5u 0.704117647000 42.500001u 0.705882352875 51u
+ 0.705882352875 51.000001u 0.707647058750 59.5u 0.707647058750 59.500001u 0.709411764625 68u 0.709411764625 68.000001u 0.711176470500 76.5u
+ 0.711176470500 76.500001u 0.712941176375 85u 0.712941176375 85.000001u 0.714705882250 93.5u 0.714705882250 93.500001u 0.716470588125 102u
+ 0.716470588125 102.000001u 0.718235294000 110.5u 0.718235294000 110.500001u 0.720000000000 119u 0.720000000000 119.000001u 0.721764705875 127.5u
+ 0.721764705875 127.500001u 0.723529411750 136u 0.723529411750 136.000001u 0.725294117625 144.5u 0.725294117625 144.500001u 0.727058823500 153u
+ 0.727058823500 153.000001u 0.728823529375 161.5u 0.728823529375 161.500001u 0.730588235250 170u 0.730588235250 170.000001u 0.732352941125 178.5u
+ 0.732352941125 178.500001u 0.734117647000 187u 0.734117647000 187.000001u 0.735882352875 195.5u 0.735882352875 195.500001u 0.737647058750 204u
+ 0.737647058750 204.000001u 0.739411764625 212.5u 0.739411764625 212.500001u 0.741176470500 221u 0.741176470500 221.000001u 0.742941176375 229.5u
+ 0.742941176375 229.500001u 0.744705882250 238u 0.744705882250 238.000001u 0.746470588125 246.5u 0.746470588125 246.500001u 0.748235294000 255u
+ 0.748235294000 255.000001u 0.750000000000 263.5u 0.750000000000 263.500001u 0.751764705875 272u 0.751764705875 272.000001u 0.753529411750 280.5u
+ 0.753529411750 280.500001u 0.755294117625 289u 0.755294117625 289.000001u 0.757058823500 297.5u 0.757058823500 297.500001u 0.758823529375 306u
+ 0.758823529375 306.000001u 0.760588235250 314.5u 0.760588235250 314.500001u 0.762352941125 323u 0.762352941125 323.000001u 0.764117647000 331.5u
+ 0.764117647000 331.500001u 0.765882352875 340u 0.765882352875 340.000001u 0.767647058750 348.5u 0.767647058750 348.500001u 0.769411764625 357u
+ 0.769411764625 357.000001u 0.771176470500 365.5u 0.771176470500 365.500001u 0.772941176375 374u 0.772941176375 374.000001u 0.774705882250 382.5u
+ 0.774705882250 382.500001u 0.776470588125 391u 0.776470588125 391.000001u 0.778235294000 399.5u 0.778235294000 399.500001u 0.780000000000 408u
+ 0.780000000000 408.000001u 0.781764705875 416.5u 0.781764705875 416.500001u 0.783529411750 425u 0.783529411750 425.000001u 0.785294117625 433.5u
+ 0.785294117625 433.500001u 0.787058823500 442u 0.787058823500 442.000001u 0.788823529375 450.5u 0.788823529375 450.500001u 0.790588235250 459u
+ 0.790588235250 459.000001u 0.792352941125 467.5u 0.792352941125 467.500001u 0.794117647000 476u 0.794117647000 476.000001u 0.795882352875 484.5u
+ 0.795882352875 484.500001u 0.797647058750 493u 0.797647058750 493.000001u 0.799411764625 501.5u 0.799411764625 501.500001u 0.801176470500 510u
+ 0.801176470500 510.000001u 0.802941176375 518.5u 0.802941176375 518.500001u 0.804705882250 527u 0.804705882250 527.000001u 0.806470588125 535.5u
+ 0.806470588125 535.500001u 0.808235294000 544u 0.808235294000 544.000001u 0.810000000000 552.5u 0.810000000000 552.500001u 0.811764705875 561u
+ 0.811764705875 561.000001u 0.813529411750 569.5u 0.813529411750 569.500001u 0.815294117625 578u 0.815294117625 578.000001u 0.817058823500 586.5u
+ 0.817058823500 586.500001u 0.818823529375 595u 0.818823529375 595.000001u 0.820588235250 603.5u 0.820588235250 603.500001u 0.822352941125 612u
+ 0.822352941125 612.000001u 0.824117647000 620.5u 0.824117647000 620.500001u 0.825882352875 629u 0.825882352875 629.000001u 0.827647058750 637.5u
+ 0.827647058750 637.500001u 0.829411764625 646u 0.829411764625 646.000001u 0.831176470500 654.5u 0.831176470500 654.500001u 0.832941176375 663u
+ 0.832941176375 663.000001u 0.834705882250 671.5u 0.834705882250 671.500001u 0.836470588125 680u 0.836470588125)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/samantha/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 680u uic
  wrdata /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_21-28-41/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
