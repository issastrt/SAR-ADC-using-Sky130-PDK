magic
tech sky130A
magscale 1 2
timestamp 1761401228
<< metal1 >>
rect 1861 -9936 1925 -9930
rect 1861 -9988 1867 -9936
rect 1919 -9988 1925 -9936
rect 1861 -9994 1925 -9988
rect 2304 -11927 2368 -11921
rect 2304 -11979 2310 -11927
rect 2362 -11979 2368 -11927
rect 2304 -11985 2368 -11979
rect 2010 -13500 2074 -13494
rect 2010 -13503 2016 -13500
rect 2005 -13549 2016 -13503
rect 2010 -13552 2016 -13549
rect 2068 -13503 2074 -13500
rect 2068 -13549 2079 -13503
rect 2068 -13552 2074 -13549
rect 2010 -13558 2074 -13552
rect 2304 -15491 2368 -15485
rect 2304 -15543 2310 -15491
rect 2362 -15543 2368 -15491
rect 2304 -15549 2368 -15543
rect 2010 -17064 2074 -17058
rect 2010 -17067 2016 -17064
rect 2005 -17113 2016 -17067
rect 2010 -17116 2016 -17113
rect 2068 -17067 2074 -17064
rect 2068 -17113 2079 -17067
rect 2068 -17116 2074 -17113
rect 2010 -17122 2074 -17116
rect 2304 -19055 2368 -19049
rect 2304 -19107 2310 -19055
rect 2362 -19107 2368 -19055
rect 2304 -19113 2368 -19107
rect 2010 -20628 2074 -20622
rect 2010 -20631 2016 -20628
rect 2005 -20677 2016 -20631
rect 2010 -20680 2016 -20677
rect 2068 -20631 2074 -20628
rect 2068 -20677 2079 -20631
rect 2068 -20680 2074 -20677
rect 2010 -20686 2074 -20680
rect 2304 -22619 2368 -22613
rect 2304 -22671 2310 -22619
rect 2362 -22671 2368 -22619
rect 2304 -22677 2368 -22671
rect 2010 -24192 2074 -24186
rect 2010 -24195 2016 -24192
rect 2005 -24241 2016 -24195
rect 2010 -24244 2016 -24241
rect 2068 -24195 2074 -24192
rect 2068 -24241 2079 -24195
rect 2068 -24244 2074 -24241
rect 2010 -24250 2074 -24244
rect 2304 -26183 2368 -26177
rect 2304 -26235 2310 -26183
rect 2362 -26235 2368 -26183
rect 2304 -26241 2368 -26235
rect 2010 -27756 2074 -27750
rect 2010 -27759 2016 -27756
rect 2005 -27805 2016 -27759
rect 2010 -27808 2016 -27805
rect 2068 -27759 2074 -27756
rect 2068 -27805 2079 -27759
rect 2068 -27808 2074 -27805
rect 2010 -27814 2074 -27808
rect 2304 -29747 2368 -29741
rect 2304 -29799 2310 -29747
rect 2362 -29799 2368 -29747
rect 2304 -29805 2368 -29799
rect 2010 -31320 2074 -31314
rect 2010 -31323 2016 -31320
rect 2005 -31369 2016 -31323
rect 2010 -31372 2016 -31369
rect 2068 -31323 2074 -31320
rect 2068 -31369 2079 -31323
rect 2068 -31372 2074 -31369
rect 2010 -31378 2074 -31372
rect 2304 -33311 2368 -33305
rect 2304 -33363 2310 -33311
rect 2362 -33363 2368 -33311
rect 2304 -33369 2368 -33363
rect 2010 -34884 2074 -34878
rect 2010 -34887 2016 -34884
rect 2005 -34933 2016 -34887
rect 2010 -34936 2016 -34933
rect 2068 -34887 2074 -34884
rect 2068 -34933 2079 -34887
rect 2068 -34936 2074 -34933
rect 2010 -34942 2074 -34936
rect 2304 -36875 2368 -36869
rect 2304 -36927 2310 -36875
rect 2362 -36927 2368 -36875
rect 2304 -36933 2368 -36927
rect 2010 -38448 2074 -38442
rect 2010 -38451 2016 -38448
rect 2005 -38497 2016 -38451
rect 2010 -38500 2016 -38497
rect 2068 -38451 2074 -38448
rect 2068 -38497 2079 -38451
rect 2068 -38500 2074 -38497
rect 2010 -38506 2074 -38500
rect 2304 -40439 2368 -40433
rect 2304 -40491 2310 -40439
rect 2362 -40491 2368 -40439
rect 2304 -40497 2368 -40491
rect 2010 -42012 2074 -42006
rect 2010 -42015 2016 -42012
rect 2005 -42061 2016 -42015
rect 2010 -42064 2016 -42061
rect 2068 -42015 2074 -42012
rect 2068 -42061 2079 -42015
rect 2068 -42064 2074 -42061
rect 2010 -42070 2074 -42064
rect 2304 -44003 2368 -43997
rect 2304 -44055 2310 -44003
rect 2362 -44055 2368 -44003
rect 2304 -44061 2368 -44055
rect 2010 -45576 2074 -45570
rect 2010 -45579 2016 -45576
rect 2005 -45625 2016 -45579
rect 2010 -45628 2016 -45625
rect 2068 -45579 2074 -45576
rect 2068 -45625 2079 -45579
rect 2068 -45628 2074 -45625
rect 2010 -45634 2074 -45628
rect 2304 -47567 2368 -47561
rect 2304 -47619 2310 -47567
rect 2362 -47619 2368 -47567
rect 2304 -47625 2368 -47619
rect 2010 -49140 2074 -49134
rect 2010 -49143 2016 -49140
rect 2005 -49189 2016 -49143
rect 2010 -49192 2016 -49189
rect 2068 -49143 2074 -49140
rect 2068 -49189 2079 -49143
rect 2068 -49192 2074 -49189
rect 2010 -49198 2074 -49192
rect 2304 -51131 2368 -51125
rect 2304 -51183 2310 -51131
rect 2362 -51183 2368 -51131
rect 2304 -51189 2368 -51183
rect 2010 -52704 2074 -52698
rect 2010 -52707 2016 -52704
rect 2005 -52753 2016 -52707
rect 2010 -52756 2016 -52753
rect 2068 -52707 2074 -52704
rect 2068 -52753 2079 -52707
rect 2068 -52756 2074 -52753
rect 2010 -52762 2074 -52756
rect 2304 -54695 2368 -54689
rect 2304 -54747 2310 -54695
rect 2362 -54747 2368 -54695
rect 2304 -54753 2368 -54747
rect 2010 -56268 2074 -56262
rect 2010 -56271 2016 -56268
rect 2005 -56317 2016 -56271
rect 2010 -56320 2016 -56317
rect 2068 -56271 2074 -56268
rect 2068 -56317 2079 -56271
rect 2068 -56320 2074 -56317
rect 2010 -56326 2074 -56320
rect 2304 -58259 2368 -58253
rect 2304 -58311 2310 -58259
rect 2362 -58311 2368 -58259
rect 2304 -58317 2368 -58311
rect 2010 -59832 2074 -59826
rect 2010 -59835 2016 -59832
rect 2005 -59881 2016 -59835
rect 2010 -59884 2016 -59881
rect 2068 -59835 2074 -59832
rect 2068 -59881 2079 -59835
rect 2068 -59884 2074 -59881
rect 2010 -59890 2074 -59884
rect 2304 -61823 2368 -61817
rect 2304 -61875 2310 -61823
rect 2362 -61875 2368 -61823
rect 2304 -61881 2368 -61875
rect 2002 -63396 2082 -63382
rect 2002 -63448 2016 -63396
rect 2068 -63448 2082 -63396
rect 2002 -63462 2082 -63448
rect 2304 -65387 2368 -65381
rect 2304 -65439 2310 -65387
rect 2362 -65439 2368 -65387
rect 2304 -65445 2368 -65439
rect 2002 -66960 2082 -66946
rect 2002 -67012 2016 -66960
rect 2068 -67012 2082 -66960
rect 2002 -67026 2082 -67012
<< via1 >>
rect 1867 -9988 1919 -9936
rect 2310 -11979 2362 -11927
rect 2016 -13552 2068 -13500
rect 2310 -15543 2362 -15491
rect 2016 -17116 2068 -17064
rect 2310 -19107 2362 -19055
rect 2016 -20680 2068 -20628
rect 2310 -22671 2362 -22619
rect 2016 -24244 2068 -24192
rect 2310 -26235 2362 -26183
rect 2016 -27808 2068 -27756
rect 2310 -29799 2362 -29747
rect 2016 -31372 2068 -31320
rect 2310 -33363 2362 -33311
rect 2016 -34936 2068 -34884
rect 2310 -36927 2362 -36875
rect 2016 -38500 2068 -38448
rect 2310 -40491 2362 -40439
rect 2016 -42064 2068 -42012
rect 2310 -44055 2362 -44003
rect 2016 -45628 2068 -45576
rect 2310 -47619 2362 -47567
rect 2016 -49192 2068 -49140
rect 2310 -51183 2362 -51131
rect 2016 -52756 2068 -52704
rect 2310 -54747 2362 -54695
rect 2016 -56320 2068 -56268
rect 2310 -58311 2362 -58259
rect 2016 -59884 2068 -59832
rect 2310 -61875 2362 -61823
rect 2016 -63448 2068 -63396
rect 2310 -65439 2362 -65387
rect 2016 -67012 2068 -66960
<< metal2 >>
rect 2299 -9004 2373 -8995
rect 2299 -9060 2308 -9004
rect 2364 -9060 2373 -9004
rect 2299 -9069 2373 -9060
rect 1853 -9934 1933 -9922
rect 1853 -9990 1865 -9934
rect 1921 -9990 1933 -9934
rect 1853 -10002 1933 -9990
rect 1720 -10173 1794 -10164
rect 1720 -10229 1729 -10173
rect 1785 -10229 1794 -10173
rect 1720 -10238 1794 -10229
rect 2296 -11925 9154 -11913
rect 2296 -11927 9086 -11925
rect 2296 -11979 2310 -11927
rect 2362 -11979 9086 -11927
rect 2296 -11981 9086 -11979
rect 9142 -11981 9154 -11925
rect 2296 -11993 9154 -11981
rect 2005 -12688 2079 -12679
rect 2005 -12744 2014 -12688
rect 2070 -12744 2079 -12688
rect 2005 -12753 2079 -12744
rect 1720 -13259 1794 -13250
rect 1720 -13315 1729 -13259
rect 1785 -13315 1794 -13259
rect 1720 -13324 1794 -13315
rect 2002 -13498 2082 -13486
rect 2002 -13554 2014 -13498
rect 2070 -13554 2082 -13498
rect 2002 -13566 2082 -13554
rect 2296 -15489 9154 -15477
rect 2296 -15491 9086 -15489
rect 2296 -15543 2310 -15491
rect 2362 -15543 9086 -15491
rect 2296 -15545 9086 -15543
rect 9142 -15545 9154 -15489
rect 2296 -15557 9154 -15545
rect 2002 -17062 2082 -17050
rect 2002 -17118 2014 -17062
rect 2070 -17118 2082 -17062
rect 2002 -17130 2082 -17118
rect 2296 -19053 9154 -19041
rect 2296 -19055 9086 -19053
rect 2296 -19107 2310 -19055
rect 2362 -19107 9086 -19055
rect 2296 -19109 9086 -19107
rect 9142 -19109 9154 -19053
rect 2296 -19121 9154 -19109
rect 2002 -20626 2082 -20614
rect 2002 -20682 2014 -20626
rect 2070 -20682 2082 -20626
rect 2002 -20694 2082 -20682
rect 2296 -22617 9154 -22605
rect 2296 -22619 9086 -22617
rect 2296 -22671 2310 -22619
rect 2362 -22671 9086 -22619
rect 2296 -22673 9086 -22671
rect 9142 -22673 9154 -22617
rect 2296 -22685 9154 -22673
rect 2002 -24190 2082 -24178
rect 2002 -24246 2014 -24190
rect 2070 -24246 2082 -24190
rect 2002 -24258 2082 -24246
rect 2296 -26181 9154 -26169
rect 2296 -26183 9086 -26181
rect 2296 -26235 2310 -26183
rect 2362 -26235 9086 -26183
rect 2296 -26237 9086 -26235
rect 9142 -26237 9154 -26181
rect 2296 -26249 9154 -26237
rect 2002 -27754 2082 -27742
rect 2002 -27810 2014 -27754
rect 2070 -27810 2082 -27754
rect 2002 -27822 2082 -27810
rect 2296 -29745 9154 -29733
rect 2296 -29747 9086 -29745
rect 2296 -29799 2310 -29747
rect 2362 -29799 9086 -29747
rect 2296 -29801 9086 -29799
rect 9142 -29801 9154 -29745
rect 2296 -29813 9154 -29801
rect 2002 -31318 2082 -31306
rect 2002 -31374 2014 -31318
rect 2070 -31374 2082 -31318
rect 2002 -31386 2082 -31374
rect 2296 -33309 9154 -33297
rect 2296 -33311 9086 -33309
rect 2296 -33363 2310 -33311
rect 2362 -33363 9086 -33311
rect 2296 -33365 9086 -33363
rect 9142 -33365 9154 -33309
rect 2296 -33377 9154 -33365
rect 2002 -34882 2082 -34870
rect 2002 -34938 2014 -34882
rect 2070 -34938 2082 -34882
rect 2002 -34950 2082 -34938
rect 2296 -36873 9154 -36861
rect 2296 -36875 9086 -36873
rect 2296 -36927 2310 -36875
rect 2362 -36927 9086 -36875
rect 2296 -36929 9086 -36927
rect 9142 -36929 9154 -36873
rect 2296 -36941 9154 -36929
rect 2002 -38446 2082 -38434
rect 2002 -38502 2014 -38446
rect 2070 -38502 2082 -38446
rect 2002 -38514 2082 -38502
rect 2296 -40437 9154 -40425
rect 2296 -40439 9086 -40437
rect 2296 -40491 2310 -40439
rect 2362 -40491 9086 -40439
rect 2296 -40493 9086 -40491
rect 9142 -40493 9154 -40437
rect 2296 -40505 9154 -40493
rect 2002 -42010 2082 -41998
rect 2002 -42066 2014 -42010
rect 2070 -42066 2082 -42010
rect 2002 -42078 2082 -42066
rect 2296 -44001 9154 -43989
rect 2296 -44003 9086 -44001
rect 2296 -44055 2310 -44003
rect 2362 -44055 9086 -44003
rect 2296 -44057 9086 -44055
rect 9142 -44057 9154 -44001
rect 2296 -44069 9154 -44057
rect 2002 -45574 2082 -45562
rect 2002 -45630 2014 -45574
rect 2070 -45630 2082 -45574
rect 2002 -45642 2082 -45630
rect 2296 -47565 9154 -47553
rect 2296 -47567 9086 -47565
rect 2296 -47619 2310 -47567
rect 2362 -47619 9086 -47567
rect 2296 -47621 9086 -47619
rect 9142 -47621 9154 -47565
rect 2296 -47633 9154 -47621
rect 2002 -49138 2082 -49126
rect 2002 -49194 2014 -49138
rect 2070 -49194 2082 -49138
rect 2002 -49206 2082 -49194
rect 2296 -51129 9154 -51117
rect 2296 -51131 9086 -51129
rect 2296 -51183 2310 -51131
rect 2362 -51183 9086 -51131
rect 2296 -51185 9086 -51183
rect 9142 -51185 9154 -51129
rect 2296 -51197 9154 -51185
rect 2002 -52702 2082 -52690
rect 2002 -52758 2014 -52702
rect 2070 -52758 2082 -52702
rect 2002 -52770 2082 -52758
rect 2296 -54693 9154 -54681
rect 2296 -54695 9086 -54693
rect 2296 -54747 2310 -54695
rect 2362 -54747 9086 -54695
rect 2296 -54749 9086 -54747
rect 9142 -54749 9154 -54693
rect 2296 -54761 9154 -54749
rect 2002 -56266 2082 -56254
rect 2002 -56322 2014 -56266
rect 2070 -56322 2082 -56266
rect 2002 -56334 2082 -56322
rect 2296 -58257 9154 -58245
rect 2296 -58259 9086 -58257
rect 2296 -58311 2310 -58259
rect 2362 -58311 9086 -58259
rect 2296 -58313 9086 -58311
rect 9142 -58313 9154 -58257
rect 2296 -58325 9154 -58313
rect 2002 -59830 2082 -59818
rect 2002 -59886 2014 -59830
rect 2070 -59886 2082 -59830
rect 2002 -59898 2082 -59886
rect 2296 -61821 9154 -61809
rect 2296 -61823 9086 -61821
rect 2296 -61875 2310 -61823
rect 2362 -61875 9086 -61823
rect 2296 -61877 9086 -61875
rect 9142 -61877 9154 -61821
rect 2296 -61889 9154 -61877
rect 2002 -63394 2082 -63382
rect 2002 -63450 2014 -63394
rect 2070 -63450 2082 -63394
rect 2002 -63462 2082 -63450
rect 2296 -65385 9154 -65373
rect 2296 -65387 9086 -65385
rect 2296 -65439 2310 -65387
rect 2362 -65439 9086 -65387
rect 2296 -65441 9086 -65439
rect 9142 -65441 9154 -65385
rect 2296 -65453 9154 -65441
rect 2002 -66958 2082 -66946
rect 2002 -67014 2014 -66958
rect 2070 -67014 2082 -66958
rect 2002 -67026 2082 -67014
rect 2296 -66958 9154 -66946
rect 2296 -67014 2308 -66958
rect 2364 -67014 9086 -66958
rect 9142 -67014 9154 -66958
rect 2296 -67026 9154 -67014
<< via2 >>
rect 2308 -9060 2364 -9004
rect 1865 -9936 1921 -9934
rect 1865 -9988 1867 -9936
rect 1867 -9988 1919 -9936
rect 1919 -9988 1921 -9936
rect 1865 -9990 1921 -9988
rect 1729 -10229 1785 -10173
rect 9086 -11981 9142 -11925
rect 2014 -12744 2070 -12688
rect 1729 -13315 1785 -13259
rect 2014 -13500 2070 -13498
rect 2014 -13552 2016 -13500
rect 2016 -13552 2068 -13500
rect 2068 -13552 2070 -13500
rect 2014 -13554 2070 -13552
rect 9086 -15545 9142 -15489
rect 2014 -17064 2070 -17062
rect 2014 -17116 2016 -17064
rect 2016 -17116 2068 -17064
rect 2068 -17116 2070 -17064
rect 2014 -17118 2070 -17116
rect 9086 -19109 9142 -19053
rect 2014 -20628 2070 -20626
rect 2014 -20680 2016 -20628
rect 2016 -20680 2068 -20628
rect 2068 -20680 2070 -20628
rect 2014 -20682 2070 -20680
rect 9086 -22673 9142 -22617
rect 2014 -24192 2070 -24190
rect 2014 -24244 2016 -24192
rect 2016 -24244 2068 -24192
rect 2068 -24244 2070 -24192
rect 2014 -24246 2070 -24244
rect 9086 -26237 9142 -26181
rect 2014 -27756 2070 -27754
rect 2014 -27808 2016 -27756
rect 2016 -27808 2068 -27756
rect 2068 -27808 2070 -27756
rect 2014 -27810 2070 -27808
rect 9086 -29801 9142 -29745
rect 2014 -31320 2070 -31318
rect 2014 -31372 2016 -31320
rect 2016 -31372 2068 -31320
rect 2068 -31372 2070 -31320
rect 2014 -31374 2070 -31372
rect 9086 -33365 9142 -33309
rect 2014 -34884 2070 -34882
rect 2014 -34936 2016 -34884
rect 2016 -34936 2068 -34884
rect 2068 -34936 2070 -34884
rect 2014 -34938 2070 -34936
rect 9086 -36929 9142 -36873
rect 2014 -38448 2070 -38446
rect 2014 -38500 2016 -38448
rect 2016 -38500 2068 -38448
rect 2068 -38500 2070 -38448
rect 2014 -38502 2070 -38500
rect 9086 -40493 9142 -40437
rect 2014 -42012 2070 -42010
rect 2014 -42064 2016 -42012
rect 2016 -42064 2068 -42012
rect 2068 -42064 2070 -42012
rect 2014 -42066 2070 -42064
rect 9086 -44057 9142 -44001
rect 2014 -45576 2070 -45574
rect 2014 -45628 2016 -45576
rect 2016 -45628 2068 -45576
rect 2068 -45628 2070 -45576
rect 2014 -45630 2070 -45628
rect 9086 -47621 9142 -47565
rect 2014 -49140 2070 -49138
rect 2014 -49192 2016 -49140
rect 2016 -49192 2068 -49140
rect 2068 -49192 2070 -49140
rect 2014 -49194 2070 -49192
rect 9086 -51185 9142 -51129
rect 2014 -52704 2070 -52702
rect 2014 -52756 2016 -52704
rect 2016 -52756 2068 -52704
rect 2068 -52756 2070 -52704
rect 2014 -52758 2070 -52756
rect 9086 -54749 9142 -54693
rect 2014 -56268 2070 -56266
rect 2014 -56320 2016 -56268
rect 2016 -56320 2068 -56268
rect 2068 -56320 2070 -56268
rect 2014 -56322 2070 -56320
rect 9086 -58313 9142 -58257
rect 2014 -59832 2070 -59830
rect 2014 -59884 2016 -59832
rect 2016 -59884 2068 -59832
rect 2068 -59884 2070 -59832
rect 2014 -59886 2070 -59884
rect 9086 -61877 9142 -61821
rect 2014 -63396 2070 -63394
rect 2014 -63448 2016 -63396
rect 2016 -63448 2068 -63396
rect 2068 -63448 2070 -63396
rect 2014 -63450 2070 -63448
rect 9086 -65441 9142 -65385
rect 2014 -66960 2070 -66958
rect 2014 -67012 2016 -66960
rect 2016 -67012 2068 -66960
rect 2068 -67012 2070 -66960
rect 2014 -67014 2070 -67012
rect 2308 -67014 2364 -66958
rect 9086 -67014 9142 -66958
<< metal3 >>
rect 635 -68740 695 -8212
rect 2303 -9004 2369 -8999
rect 2303 -9060 2308 -9004
rect 2364 -9060 2369 -9004
rect 2303 -9065 2369 -9060
rect 1860 -9934 1926 -9929
rect 1860 -9990 1865 -9934
rect 1921 -9990 1926 -9934
rect 1860 -9995 1926 -9990
rect 1724 -10173 1790 -10168
rect 1724 -10229 1729 -10173
rect 1785 -10229 1790 -10173
rect 1724 -10234 1790 -10229
rect 1727 -13254 1787 -10234
rect 2012 -12683 2072 -10742
rect 1724 -13259 1790 -13254
rect 1724 -13315 1729 -13259
rect 1785 -13315 1790 -13259
rect 1724 -13320 1790 -13315
rect 1863 -67272 1923 -12686
rect 2009 -12688 2075 -12683
rect 2009 -12744 2014 -12688
rect 2070 -12744 2075 -12688
rect 2009 -12749 2075 -12744
rect 2012 -13493 2072 -13310
rect 2009 -13498 2075 -13493
rect 2009 -13554 2014 -13498
rect 2070 -13554 2075 -13498
rect 2009 -13559 2075 -13554
rect 2012 -17057 2072 -13559
rect 2009 -17062 2075 -17057
rect 2009 -17118 2014 -17062
rect 2070 -17118 2075 -17062
rect 2009 -17123 2075 -17118
rect 2012 -20621 2072 -17123
rect 2009 -20626 2075 -20621
rect 2009 -20682 2014 -20626
rect 2070 -20682 2075 -20626
rect 2009 -20687 2075 -20682
rect 2012 -24185 2072 -20687
rect 2009 -24190 2075 -24185
rect 2009 -24246 2014 -24190
rect 2070 -24246 2075 -24190
rect 2009 -24251 2075 -24246
rect 2012 -27749 2072 -24251
rect 2009 -27754 2075 -27749
rect 2009 -27810 2014 -27754
rect 2070 -27810 2075 -27754
rect 2009 -27815 2075 -27810
rect 2012 -31313 2072 -27815
rect 2009 -31318 2075 -31313
rect 2009 -31374 2014 -31318
rect 2070 -31374 2075 -31318
rect 2009 -31379 2075 -31374
rect 2012 -34877 2072 -31379
rect 2009 -34882 2075 -34877
rect 2009 -34938 2014 -34882
rect 2070 -34938 2075 -34882
rect 2009 -34943 2075 -34938
rect 2012 -38441 2072 -34943
rect 2009 -38446 2075 -38441
rect 2009 -38502 2014 -38446
rect 2070 -38502 2075 -38446
rect 2009 -38507 2075 -38502
rect 2012 -42005 2072 -38507
rect 2009 -42010 2075 -42005
rect 2009 -42066 2014 -42010
rect 2070 -42066 2075 -42010
rect 2009 -42071 2075 -42066
rect 2012 -45569 2072 -42071
rect 2009 -45574 2075 -45569
rect 2009 -45630 2014 -45574
rect 2070 -45630 2075 -45574
rect 2009 -45635 2075 -45630
rect 2012 -49133 2072 -45635
rect 2009 -49138 2075 -49133
rect 2009 -49194 2014 -49138
rect 2070 -49194 2075 -49138
rect 2009 -49199 2075 -49194
rect 2012 -52697 2072 -49199
rect 2009 -52702 2075 -52697
rect 2009 -52758 2014 -52702
rect 2070 -52758 2075 -52702
rect 2009 -52763 2075 -52758
rect 2012 -56261 2072 -52763
rect 2009 -56266 2075 -56261
rect 2009 -56322 2014 -56266
rect 2070 -56322 2075 -56266
rect 2009 -56327 2075 -56322
rect 2012 -59825 2072 -56327
rect 2009 -59830 2075 -59825
rect 2009 -59886 2014 -59830
rect 2070 -59886 2075 -59830
rect 2009 -59891 2075 -59886
rect 2012 -63389 2072 -59891
rect 2009 -63394 2075 -63389
rect 2009 -63450 2014 -63394
rect 2070 -63450 2075 -63394
rect 2009 -63455 2075 -63450
rect 2012 -66953 2072 -63455
rect 2306 -66953 2366 -9065
rect 2009 -66958 2075 -66953
rect 2009 -67014 2014 -66958
rect 2070 -67014 2075 -66958
rect 2009 -67019 2075 -67014
rect 2303 -66958 2369 -66953
rect 2303 -67014 2308 -66958
rect 2364 -67014 2369 -66958
rect 2303 -67019 2369 -67014
rect 2012 -67826 2072 -67019
rect 2920 -67272 2980 -9690
rect 9084 -11920 9144 -9580
rect 9081 -11925 9147 -11920
rect 9081 -11981 9086 -11925
rect 9142 -11981 9147 -11925
rect 9081 -11986 9147 -11981
rect 9084 -15484 9144 -13144
rect 9081 -15489 9147 -15484
rect 9081 -15545 9086 -15489
rect 9142 -15545 9147 -15489
rect 9081 -15550 9147 -15545
rect 9084 -19048 9144 -16708
rect 9081 -19053 9147 -19048
rect 9081 -19109 9086 -19053
rect 9142 -19109 9147 -19053
rect 9081 -19114 9147 -19109
rect 9084 -22612 9144 -20272
rect 9081 -22617 9147 -22612
rect 9081 -22673 9086 -22617
rect 9142 -22673 9147 -22617
rect 9081 -22678 9147 -22673
rect 9084 -26176 9144 -23836
rect 9081 -26181 9147 -26176
rect 9081 -26237 9086 -26181
rect 9142 -26237 9147 -26181
rect 9081 -26242 9147 -26237
rect 9084 -29740 9144 -27400
rect 9081 -29745 9147 -29740
rect 9081 -29801 9086 -29745
rect 9142 -29801 9147 -29745
rect 9081 -29806 9147 -29801
rect 9084 -33304 9144 -30964
rect 9081 -33309 9147 -33304
rect 9081 -33365 9086 -33309
rect 9142 -33365 9147 -33309
rect 9081 -33370 9147 -33365
rect 9084 -36868 9144 -34528
rect 9081 -36873 9147 -36868
rect 9081 -36929 9086 -36873
rect 9142 -36929 9147 -36873
rect 9081 -36934 9147 -36929
rect 9084 -40432 9144 -38092
rect 9081 -40437 9147 -40432
rect 9081 -40493 9086 -40437
rect 9142 -40493 9147 -40437
rect 9081 -40498 9147 -40493
rect 9084 -43996 9144 -41656
rect 9081 -44001 9147 -43996
rect 9081 -44057 9086 -44001
rect 9142 -44057 9147 -44001
rect 9081 -44062 9147 -44057
rect 9084 -47560 9144 -45220
rect 9081 -47565 9147 -47560
rect 9081 -47621 9086 -47565
rect 9142 -47621 9147 -47565
rect 9081 -47626 9147 -47621
rect 9084 -51124 9144 -48784
rect 9081 -51129 9147 -51124
rect 9081 -51185 9086 -51129
rect 9142 -51185 9147 -51129
rect 9081 -51190 9147 -51185
rect 9084 -54688 9144 -52348
rect 9081 -54693 9147 -54688
rect 9081 -54749 9086 -54693
rect 9142 -54749 9147 -54693
rect 9081 -54754 9147 -54749
rect 9084 -58252 9144 -55912
rect 9081 -58257 9147 -58252
rect 9081 -58313 9086 -58257
rect 9142 -58313 9147 -58257
rect 9081 -58318 9147 -58313
rect 9084 -61816 9144 -59476
rect 9081 -61821 9147 -61816
rect 9081 -61877 9086 -61821
rect 9142 -61877 9147 -61821
rect 9081 -61882 9147 -61877
rect 9084 -65380 9144 -63040
rect 9081 -65385 9147 -65380
rect 9081 -65441 9086 -65385
rect 9142 -65441 9147 -65385
rect 9081 -65446 9147 -65441
rect 9081 -66958 9147 -66953
rect 9081 -67014 9086 -66958
rect 9142 -67014 9147 -66958
rect 9081 -67019 9147 -67014
use D_FlipFlop  D_FlipFlop_0
timestamp 1761392116
transform 1 0 606 0 1 -9985
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_1
timestamp 1761392116
transform 1 0 606 0 1 -13549
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_2
timestamp 1761392116
transform 1 0 606 0 1 -17113
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_3
timestamp 1761392116
transform 1 0 606 0 1 -20677
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_4
timestamp 1761392116
transform 1 0 606 0 1 -24241
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_5
timestamp 1761392116
transform 1 0 606 0 1 -27805
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_6
timestamp 1761392116
transform 1 0 606 0 1 -31369
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_7
timestamp 1761392116
transform 1 0 606 0 1 -34933
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_8
timestamp 1761392116
transform 1 0 606 0 1 -38497
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_9
timestamp 1761392116
transform 1 0 606 0 1 -42061
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_10
timestamp 1761392116
transform 1 0 606 0 1 -45625
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_11
timestamp 1761392116
transform 1 0 606 0 1 -49189
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_12
timestamp 1761392116
transform 1 0 606 0 1 -52753
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_13
timestamp 1761392116
transform 1 0 606 0 1 -56317
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_14
timestamp 1761392116
transform 1 0 606 0 1 -59881
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_15
timestamp 1761392116
transform 1 0 606 0 1 -63445
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_16
timestamp 1761392116
transform 1 0 606 0 1 -67009
box 0 -1799 8762 1845
<< labels >>
flabel metal3 2920 -67272 2980 -9690 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 1863 -67272 1923 -12686 0 FreeSans 160 90 0 0 EN
port 1 nsew
flabel metal3 635 -68740 695 -8212 0 FreeSans 160 90 0 0 GND
port 2 nsew
flabel metal3 9084 -11942 9144 -9580 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal3 9084 -15506 9144 -13144 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal3 9084 -19070 9144 -16708 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal3 9084 -22634 9144 -20272 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal3 9084 -26198 9144 -23836 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal3 9084 -29762 9144 -27400 0 FreeSans 160 0 0 0 Q5
port 8 nsew
flabel metal3 9084 -33326 9144 -30964 0 FreeSans 160 0 0 0 Q6
port 9 nsew
flabel metal3 9084 -36890 9144 -34528 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal3 9084 -40454 9144 -38092 0 FreeSans 160 0 0 0 Q8
port 11 nsew
flabel metal3 9084 -44018 9144 -41656 0 FreeSans 160 0 0 0 Q9
port 12 nsew
flabel metal3 9084 -47582 9144 -45220 0 FreeSans 160 0 0 0 Q10
port 13 nsew
flabel metal3 9084 -51146 9144 -48784 0 FreeSans 160 0 0 0 Q11
port 14 nsew
flabel metal3 9084 -54710 9144 -52348 0 FreeSans 160 0 0 0 Q12
port 15 nsew
flabel metal3 9084 -58274 9144 -55912 0 FreeSans 160 0 0 0 Q13
port 16 nsew
flabel metal3 9084 -61838 9144 -59476 0 FreeSans 160 0 0 0 Q14
port 17 nsew
flabel metal3 9084 -65402 9144 -63040 0 FreeSans 160 0 0 0 Q15
port 18 nsew
flabel metal3 2012 -67826 2072 -13310 0 FreeSans 160 0 0 0 VDD
port 19 nsew
<< end >>
