magic
tech sky130A
magscale 1 2
timestamp 1761291873
<< dnwell >>
rect 24583 14110 26613 29565
rect 24583 -1560 30792 14110
rect 24560 -2160 30792 -1560
rect 24583 -2191 30792 -2160
rect 24583 -2197 26613 -2191
<< nwell >>
rect 24473 29359 26723 29675
rect 24473 -1985 24795 29359
rect 26407 14220 26723 29359
rect 28818 19081 29237 29675
rect 29235 17354 29951 19081
rect 29235 17337 29560 17354
rect 29633 17337 29951 17354
rect 29235 17081 29951 17337
rect 26407 13904 30902 14220
rect 30586 -1985 30902 13904
rect 24473 -2307 30902 -1985
<< pwell >>
rect 24850 12337 26328 29265
rect 24850 617 28850 12337
rect 24850 -1964 29969 617
rect 27899 -1985 27965 -1964
rect 28952 -1985 29018 -1964
<< mvnsubdiff >>
rect 24540 29588 26656 29608
rect 24540 29554 24634 29588
rect 26576 29554 26656 29588
rect 24540 29534 26656 29554
rect 24540 29528 24620 29534
rect 24540 -2146 24560 29528
rect 24600 -2146 24620 29528
rect 26582 29528 26656 29534
rect 26582 14157 26602 29528
rect 26636 14157 26656 29528
rect 26582 14153 26656 14157
rect 26582 14133 30835 14153
rect 26582 14099 26672 14133
rect 30755 14099 30835 14133
rect 26582 14079 30835 14099
rect 24540 -2160 24620 -2146
rect 30761 14073 30835 14079
rect 30761 -2154 30781 14073
rect 30815 -2154 30835 14073
rect 30761 -2160 30835 -2154
rect 24540 -2180 30835 -2160
rect 24540 -2220 24620 -2180
rect 30755 -2220 30835 -2180
rect 24540 -2240 30835 -2220
<< mvnsubdiffcont >>
rect 24634 29554 26576 29588
rect 24560 -2146 24600 29528
rect 26602 14157 26636 29528
rect 26672 14099 30755 14133
rect 30781 -2154 30815 14073
rect 24620 -2220 30755 -2180
<< locali >>
rect 24634 29715 26576 29721
rect 24634 29681 24640 29715
rect 26570 29681 26576 29715
rect 24634 29588 26576 29681
rect 27657 29715 28743 29721
rect 27657 29681 27663 29715
rect 28737 29681 28743 29715
rect 24560 29554 24634 29588
rect 26576 29554 26636 29588
rect 27657 29563 28743 29681
rect 29313 29715 29873 29721
rect 29313 29681 29319 29715
rect 29867 29681 29873 29715
rect 29313 29563 29873 29681
rect 24560 29528 24600 29554
rect 26602 29528 26636 29554
rect 26602 14133 26636 14157
rect 26602 14099 26672 14133
rect 30755 14099 30815 14133
rect 30781 14073 30815 14099
rect 24982 -1970 26196 -1829
rect 24982 -2004 24988 -1970
rect 26190 -2004 26196 -1970
rect 24982 -2010 26196 -2004
rect 27426 -1970 28438 -1817
rect 27426 -2004 27432 -1970
rect 28432 -2004 28438 -1970
rect 27426 -2010 28438 -2004
rect 29457 -1970 29825 -1817
rect 29457 -2004 29463 -1970
rect 29819 -2004 29825 -1970
rect 29457 -2010 29825 -2004
rect 24560 -2180 24600 -2146
rect 30781 -2180 30815 -2154
rect 24560 -2220 24620 -2180
rect 30755 -2220 30815 -2180
<< viali >>
rect 24640 29681 26570 29715
rect 27663 29681 28737 29715
rect 29319 29681 29867 29715
rect 24988 -2004 26190 -1970
rect 27432 -2004 28432 -1970
rect 29463 -2004 29819 -1970
<< metal1 >>
rect 24473 29715 29951 29738
rect 24473 29681 24640 29715
rect 26570 29681 27663 29715
rect 28737 29681 29319 29715
rect 29867 29681 29951 29715
rect 24473 29658 29951 29681
rect 25016 28667 26162 29658
rect 27837 29419 28037 29499
rect 28162 29378 28238 29658
rect 28363 29419 28563 29499
rect 29327 29378 29403 29658
rect 29493 29419 29693 29499
rect 27755 19337 27831 29378
rect 28043 29298 28357 29378
rect 28043 19378 28119 29298
rect 28281 19378 28357 29298
rect 28569 19458 28645 29378
rect 29327 29298 29487 29378
rect 28569 19444 28708 19458
rect 28569 19392 28642 19444
rect 28694 19392 28708 19444
rect 28569 19378 28708 19392
rect 27695 19323 28559 19337
rect 27695 19271 27709 19323
rect 27761 19271 28559 19323
rect 27695 19257 28559 19271
rect 29407 17378 29487 29298
rect 29699 17444 29779 29378
rect 29699 17392 29713 17444
rect 29765 17392 29779 17444
rect 29699 17378 29779 17392
rect 29493 17320 29560 17337
rect 29561 17323 29625 17329
rect 29561 17320 29567 17323
rect 29493 17271 29567 17320
rect 29619 17320 29625 17323
rect 29633 17320 29693 17337
rect 29619 17271 29693 17320
rect 29493 17257 29693 17271
rect 27778 12163 27978 12177
rect 27778 12111 27911 12163
rect 27963 12111 27978 12163
rect 27778 12100 27978 12111
rect 27778 12097 27897 12100
rect 27899 12097 27978 12100
rect 28422 12097 28622 12177
rect 27700 12055 27764 12057
rect 27692 12051 27768 12055
rect 27692 11999 27706 12051
rect 27758 11999 27768 12051
rect 27692 11995 27768 11999
rect 27692 9065 27772 11995
rect 27984 9133 28064 12065
rect 27984 9081 27998 9133
rect 28050 9081 28064 9133
rect 27984 9065 28064 9081
rect 28336 9133 28416 12065
rect 28336 9081 28350 9133
rect 28402 9081 28416 9133
rect 28336 9065 28416 9081
rect 28628 12051 28708 12065
rect 28628 11999 28642 12051
rect 28694 11999 28708 12051
rect 28628 9065 28708 11999
rect 27778 8953 27978 9033
rect 28422 9020 28495 9033
rect 28499 9020 28622 9033
rect 28422 9019 28622 9020
rect 28422 8967 28509 9019
rect 28561 8967 28622 9019
rect 28422 8953 28622 8967
rect 27510 2391 27710 2471
rect 28154 2391 28354 2471
rect 25981 -1587 26045 -1581
rect 25981 -1639 25987 -1587
rect 26039 -1639 26045 -1587
rect 25981 -1645 26045 -1639
rect 27424 -1587 27504 2359
rect 27424 -1639 27438 -1587
rect 27490 -1639 27504 -1587
rect 27424 -1673 27504 -1639
rect 27716 -1575 27796 2359
rect 27716 -1627 27730 -1575
rect 27782 -1627 27796 -1575
rect 27716 -1641 27796 -1627
rect 28068 2336 28148 2359
rect 28068 2284 28082 2336
rect 28134 2284 28148 2336
rect 28068 -1641 28148 2284
rect 28360 -1575 28440 2359
rect 29541 391 29741 471
rect 28360 -1627 28374 -1575
rect 28426 -1627 28440 -1575
rect 28360 -1641 28440 -1627
rect 29455 -1575 29535 359
rect 29455 -1627 29469 -1575
rect 29521 -1627 29535 -1575
rect 29455 -1641 29535 -1627
rect 29747 292 29827 359
rect 29747 240 29761 292
rect 29813 240 29827 292
rect 29747 -1641 29827 240
rect 27424 -1753 29737 -1673
rect 24850 -1961 29969 -1947
rect 24850 -1970 27906 -1961
rect 27958 -1970 28959 -1961
rect 24850 -2004 24988 -1970
rect 26190 -2004 27432 -1970
rect 28432 -2004 28959 -1970
rect 24850 -2013 27906 -2004
rect 27958 -2013 28959 -2004
rect 29011 -1970 29969 -1961
rect 29011 -2004 29463 -1970
rect 29819 -2004 29969 -1970
rect 29011 -2013 29969 -2004
rect 24850 -2027 29969 -2013
<< via1 >>
rect 28642 19392 28694 19444
rect 27709 19271 27761 19323
rect 29713 17392 29765 17444
rect 29567 17271 29619 17323
rect 27911 12111 27963 12163
rect 27706 11999 27758 12051
rect 27998 9081 28050 9133
rect 28350 9081 28402 9133
rect 28642 11999 28694 12051
rect 28509 8967 28561 9019
rect 25987 -1639 26039 -1587
rect 27438 -1639 27490 -1587
rect 27730 -1627 27782 -1575
rect 28082 2284 28134 2336
rect 28374 -1627 28426 -1575
rect 29469 -1627 29521 -1575
rect 29761 240 29813 292
rect 27906 -1970 27958 -1961
rect 27906 -2004 27958 -1970
rect 27906 -2013 27958 -2004
rect 28959 -2013 29011 -1961
<< metal2 >>
rect 28628 19446 28708 19458
rect 28628 19390 28640 19446
rect 28696 19390 28708 19446
rect 28628 19378 28708 19390
rect 27695 19325 27775 19337
rect 27695 19269 27707 19325
rect 27763 19269 27775 19325
rect 27695 19257 27775 19269
rect 29699 17446 30238 17458
rect 29699 17444 30173 17446
rect 29699 17392 29713 17444
rect 29765 17392 30173 17444
rect 29699 17390 30173 17392
rect 30229 17390 30238 17446
rect 29699 17378 30238 17390
rect 28628 17325 29633 17337
rect 28628 17269 28640 17325
rect 28696 17269 29565 17325
rect 29621 17269 29633 17325
rect 28628 17257 29633 17269
rect 27897 12165 27977 12177
rect 27897 12109 27909 12165
rect 27965 12109 27977 12165
rect 27897 12097 27977 12109
rect 27692 12053 27772 12065
rect 27692 11997 27704 12053
rect 27760 11997 27772 12053
rect 27692 11985 27772 11997
rect 28628 12053 28708 12065
rect 28628 11997 28640 12053
rect 28696 11997 28708 12053
rect 28628 11985 28708 11997
rect 27984 9135 28416 9147
rect 27984 9133 28172 9135
rect 27984 9081 27998 9133
rect 28050 9081 28172 9133
rect 27984 9079 28172 9081
rect 28228 9133 28416 9135
rect 28228 9081 28350 9133
rect 28402 9081 28416 9133
rect 28228 9079 28416 9081
rect 27984 9067 28416 9079
rect 28495 9021 28575 9033
rect 28495 8965 28507 9021
rect 28563 8965 28575 9021
rect 28495 8953 28575 8965
rect 28068 2338 28148 2350
rect 28068 2282 28080 2338
rect 28136 2282 28148 2338
rect 28068 2270 28148 2282
rect 29747 294 30238 306
rect 29747 292 30173 294
rect 29747 240 29761 292
rect 29813 240 30173 292
rect 29747 238 30173 240
rect 30229 238 30238 294
rect 29747 226 30238 238
rect 27716 -1573 29535 -1561
rect 25981 -1587 27504 -1573
rect 25981 -1639 25987 -1587
rect 26039 -1639 27438 -1587
rect 27490 -1639 27504 -1587
rect 25981 -1653 27504 -1639
rect 27716 -1575 27904 -1573
rect 27716 -1627 27730 -1575
rect 27782 -1627 27904 -1575
rect 27716 -1629 27904 -1627
rect 27960 -1575 28957 -1573
rect 27960 -1627 28374 -1575
rect 28426 -1627 28957 -1575
rect 27960 -1629 28957 -1627
rect 29013 -1575 29535 -1573
rect 29013 -1627 29469 -1575
rect 29521 -1627 29535 -1575
rect 29013 -1629 29535 -1627
rect 27716 -1641 29535 -1629
rect 27892 -1959 27972 -1947
rect 27892 -2015 27904 -1959
rect 27960 -2015 27972 -1959
rect 27892 -2027 27972 -2015
rect 28945 -1959 29025 -1947
rect 28945 -2015 28957 -1959
rect 29013 -2015 29025 -1959
rect 28945 -2027 29025 -2015
<< via2 >>
rect 28640 19444 28696 19446
rect 28640 19392 28642 19444
rect 28642 19392 28694 19444
rect 28694 19392 28696 19444
rect 28640 19390 28696 19392
rect 27707 19323 27763 19325
rect 27707 19271 27709 19323
rect 27709 19271 27761 19323
rect 27761 19271 27763 19323
rect 27707 19269 27763 19271
rect 30173 17390 30229 17446
rect 28640 17269 28696 17325
rect 29565 17323 29621 17325
rect 29565 17271 29567 17323
rect 29567 17271 29619 17323
rect 29619 17271 29621 17323
rect 29565 17269 29621 17271
rect 27909 12163 27965 12165
rect 27909 12111 27911 12163
rect 27911 12111 27963 12163
rect 27963 12111 27965 12163
rect 27909 12109 27965 12111
rect 27704 12051 27760 12053
rect 27704 11999 27706 12051
rect 27706 11999 27758 12051
rect 27758 11999 27760 12051
rect 27704 11997 27760 11999
rect 28640 12051 28696 12053
rect 28640 11999 28642 12051
rect 28642 11999 28694 12051
rect 28694 11999 28696 12051
rect 28640 11997 28696 11999
rect 28172 9079 28228 9135
rect 28507 9019 28563 9021
rect 28507 8967 28509 9019
rect 28509 8967 28561 9019
rect 28561 8967 28563 9019
rect 28507 8965 28563 8967
rect 28080 2336 28136 2338
rect 28080 2284 28082 2336
rect 28082 2284 28134 2336
rect 28134 2284 28136 2336
rect 28080 2282 28136 2284
rect 30173 238 30229 294
rect 27904 -1629 27960 -1573
rect 28957 -1629 29013 -1573
rect 27904 -1961 27960 -1959
rect 27904 -2013 27906 -1961
rect 27906 -2013 27958 -1961
rect 27958 -2013 27960 -1961
rect 27904 -2015 27960 -2013
rect 28957 -1961 29013 -1959
rect 28957 -2013 28959 -1961
rect 28959 -2013 29011 -1961
rect 29011 -2013 29013 -1961
rect 28957 -2015 29013 -2013
<< metal3 >>
rect 28635 19446 28701 19451
rect 28635 19390 28640 19446
rect 28696 19390 28701 19446
rect 28635 19385 28701 19390
rect 27702 19325 27768 19330
rect 27702 19269 27707 19325
rect 27763 19269 27768 19325
rect 27702 19257 27768 19269
rect 27702 12058 27762 19257
rect 28638 17330 28698 19385
rect 30168 17446 30234 17451
rect 30168 17390 30173 17446
rect 30229 17390 30234 17446
rect 30168 17385 30234 17390
rect 28635 17325 28701 17330
rect 28635 17269 28640 17325
rect 28696 17269 28701 17325
rect 28635 17264 28701 17269
rect 29560 17325 29626 17330
rect 29560 17269 29565 17325
rect 29621 17269 29626 17325
rect 29560 17264 29626 17269
rect 27899 12475 27975 12481
rect 27899 12411 27905 12475
rect 27969 12411 27975 12475
rect 27899 12405 27975 12411
rect 27907 12170 27967 12405
rect 27904 12165 27970 12170
rect 27904 12109 27909 12165
rect 27965 12109 27970 12165
rect 27904 12104 27970 12109
rect 28638 12058 28698 17264
rect 29563 13429 29623 17264
rect 29555 13423 29631 13429
rect 29555 13359 29561 13423
rect 29625 13359 29631 13423
rect 29555 13353 29631 13359
rect 27699 12053 27765 12058
rect 27699 11997 27704 12053
rect 27760 11997 27765 12053
rect 27699 11992 27765 11997
rect 28635 12053 28701 12058
rect 28635 11997 28640 12053
rect 28696 11997 28701 12053
rect 28635 11992 28701 11997
rect 30171 11311 30231 17385
rect 30163 11305 30239 11311
rect 30163 11241 30169 11305
rect 30233 11241 30239 11305
rect 30163 11235 30239 11241
rect 28167 9135 28233 9140
rect 28167 9079 28172 9135
rect 28228 9079 28233 9135
rect 28167 9074 28233 9079
rect 28170 2692 28230 9074
rect 28502 9021 28568 9026
rect 28502 8965 28507 9021
rect 28563 8965 28568 9021
rect 28502 8960 28568 8965
rect 28505 8735 28565 8960
rect 28497 8729 28573 8735
rect 28497 8665 28503 8729
rect 28567 8665 28573 8729
rect 28497 8659 28573 8665
rect 28947 5357 29023 5363
rect 28947 5293 28953 5357
rect 29017 5293 29023 5357
rect 28947 5287 29023 5293
rect 28079 2632 28230 2692
rect 28079 2343 28139 2632
rect 28075 2338 28141 2343
rect 28075 2282 28080 2338
rect 28136 2282 28141 2338
rect 28075 2277 28141 2282
rect 28955 -1568 29015 5287
rect 30171 299 30231 11235
rect 30168 294 30234 299
rect 30168 238 30173 294
rect 30229 238 30234 294
rect 30168 233 30234 238
rect 27899 -1573 27965 -1568
rect 27899 -1629 27904 -1573
rect 27960 -1629 27965 -1573
rect 27899 -1634 27965 -1629
rect 28952 -1573 29018 -1568
rect 28952 -1629 28957 -1573
rect 29013 -1629 29018 -1573
rect 28952 -1634 29018 -1629
rect 27902 -1954 27962 -1634
rect 28955 -1954 29015 -1634
rect 27899 -1959 27965 -1954
rect 27899 -2015 27904 -1959
rect 27960 -2015 27965 -1959
rect 27899 -2020 27965 -2015
rect 28952 -1959 29018 -1954
rect 28952 -2015 28957 -1959
rect 29013 -2015 29018 -1959
rect 28952 -2020 29018 -2015
<< via3 >>
rect 27905 12411 27969 12475
rect 29561 13359 29625 13423
rect 30169 11241 30233 11305
rect 28503 8665 28567 8729
rect 28953 5293 29017 5357
<< via4 >>
rect 29475 13423 29711 13509
rect 29475 13359 29561 13423
rect 29561 13359 29625 13423
rect 29625 13359 29711 13423
rect 29475 13273 29711 13359
rect 27819 12475 28055 12561
rect 27819 12411 27905 12475
rect 27905 12411 27969 12475
rect 27969 12411 28055 12475
rect 27819 12325 28055 12411
rect 30083 11305 30319 11391
rect 30083 11241 30169 11305
rect 30169 11241 30233 11305
rect 30233 11241 30319 11305
rect 30083 11155 30319 11241
rect 28417 8729 28653 8815
rect 28417 8665 28503 8729
rect 28503 8665 28567 8729
rect 28567 8665 28653 8729
rect 28417 8579 28653 8665
rect 28867 5357 29103 5443
rect 28867 5293 28953 5357
rect 28953 5293 29017 5357
rect 29017 5293 29103 5357
rect 28867 5207 29103 5293
<< metal5 >>
rect 29433 13509 29753 13533
rect 29433 13273 29475 13509
rect 29711 13273 29753 13509
rect 27777 12561 28097 12881
rect 27777 12325 27819 12561
rect 28055 12325 28097 12561
rect 27777 12301 28097 12325
rect 29433 12128 29753 13273
rect 29103 11391 30343 11433
rect 29103 11155 30083 11391
rect 30319 11155 30343 11391
rect 29103 11113 30343 11155
rect 28375 8815 28695 8839
rect 28375 8579 28417 8815
rect 28653 8579 28695 8815
rect 28375 8259 28695 8579
rect 29433 6180 29753 11113
rect 28835 5443 30165 5485
rect 28835 5207 28867 5443
rect 29103 5207 30165 5443
rect 28835 5165 30165 5207
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_0
timestamp 1756481424
transform 0 1 29593 -1 0 6071
box -884 -281 906 281
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_1
timestamp 1756481424
transform 0 1 29593 -1 0 12019
box -884 -281 906 281
use sky130_fd_pr__nfet_g5v0d10v5_94KJBV  sky130_fd_pr__nfet_g5v0d10v5_94KJBV_0
timestamp 1756538730
transform 1 0 27878 0 1 10565
box -328 -1758 328 1758
use sky130_fd_pr__nfet_g5v0d10v5_94KJBV  sky130_fd_pr__nfet_g5v0d10v5_94KJBV_1
timestamp 1756538730
transform 1 0 28522 0 1 10565
box -328 -1758 328 1758
use sky130_fd_pr__nfet_g5v0d10v5_DTGLBV  sky130_fd_pr__nfet_g5v0d10v5_DTGLBV_1
timestamp 1756538730
transform 1 0 28254 0 1 359
box -328 -2258 328 2258
use sky130_fd_pr__nfet_g5v0d10v5_DTGLBV  sky130_fd_pr__nfet_g5v0d10v5_DTGLBV_2
timestamp 1756538730
transform 1 0 27610 0 1 359
box -328 -2258 328 2258
use sky130_fd_pr__res_xhigh_po_5p73_2WP2GG  sky130_fd_pr__res_xhigh_po_5p73_2WP2GG_0
timestamp 1756481424
transform 1 0 25589 0 1 13683
box -739 -15582 739 15582
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM3
timestamp 1756481424
transform 1 0 27937 0 1 24378
box -358 -5297 358 5297
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM4
timestamp 1756481424
transform 1 0 28463 0 1 24378
box -358 -5297 358 5297
use sky130_fd_pr__nfet_g5v0d10v5_Q3M7H8  XM6
timestamp 1756481424
transform 1 0 29641 0 1 -641
box -328 -1258 328 1258
use sky130_fd_pr__pfet_g5v0d10v5_UX3D7Q  XM9
timestamp 1756481424
transform 1 0 29593 0 1 23378
box -358 -6297 358 6297
<< labels >>
flabel metal5 27777 12561 28097 12881 0 FreeSans 800 0 0 0 Vinm
port 3 nsew
flabel metal5 29433 6180 29753 10857 0 FreeSans 800 0 0 0 Vout
port 5 nsew
flabel metal1 25175 -2010 27906 -1964 0 FreeSans 160 0 0 0 VSS
port 6 nsew
flabel metal5 28375 8259 28695 8579 0 FreeSans 800 0 0 0 Vinp
port 4 nsew
flabel metal1 26570 29658 27663 29738 0 FreeSans 160 0 0 0 VDD
port 7 nsew
<< end >>
