magic
tech sky130A
magscale 1 2
timestamp 1753263907
<< nwell >>
rect 1906 370 1948 1252
rect 3222 370 3264 1252
<< locali >>
rect 2122 1292 2434 1298
rect 2122 1258 2128 1292
rect 2428 1258 2434 1292
rect 2122 1140 2434 1258
rect 2736 1292 3048 1298
rect 2736 1258 2742 1292
rect 3042 1258 3048 1292
rect 2736 1140 3048 1258
rect 2050 -490 2506 -402
rect 2050 -524 2056 -490
rect 2500 -524 2506 -490
rect 2050 -530 2506 -524
rect 2664 -490 3120 -402
rect 2664 -524 2670 -490
rect 3114 -524 3120 -490
rect 2664 -530 3120 -524
<< viali >>
rect 2128 1258 2428 1292
rect 2742 1258 3042 1292
rect 2056 -524 2500 -490
rect 2670 -524 3114 -490
<< metal1 >>
rect 1906 1292 3264 1298
rect 1906 1258 2128 1292
rect 2428 1258 2742 1292
rect 3042 1258 3264 1292
rect 1906 1252 3264 1258
rect 2562 955 2608 1252
rect 2356 909 2814 955
rect 2145 725 2209 731
rect 2145 673 2151 725
rect 2203 673 2209 725
rect 2145 667 2209 673
rect 2961 725 3025 731
rect 2961 673 2967 725
rect 3019 713 3025 725
rect 3019 673 3138 713
rect 2961 667 3138 673
rect 2255 94 2301 626
rect 2869 94 2915 626
rect 3092 62 3138 667
rect 3042 16 3138 62
rect 2032 -226 2128 -180
rect 2428 -226 2742 -180
rect 2032 -484 2078 -226
rect 1906 -490 3264 -484
rect 1906 -524 2056 -490
rect 2500 -524 2670 -490
rect 3114 -524 3264 -490
rect 1906 -530 3264 -524
<< via1 >>
rect 2151 673 2203 725
rect 2967 673 3019 725
<< metal2 >>
rect 2145 725 2209 731
rect 2145 673 2151 725
rect 2203 722 2209 725
rect 2961 725 3025 731
rect 2961 722 2967 725
rect 2203 676 2967 722
rect 2203 673 2209 676
rect 2145 667 2209 673
rect 2961 673 2967 676
rect 3019 673 3025 725
rect 2961 667 3025 673
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1753016136
transform 1 0 2892 0 1 811
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM2
timestamp 1753016136
transform 1 0 2278 0 1 811
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM3
timestamp 1753016136
transform 1 0 2892 0 1 -82
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4
timestamp 1753016136
transform 1 0 2278 0 1 -82
box -372 -402 372 402
<< labels >>
flabel metal1 1906 -530 3264 -484 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 1906 1252 3264 1298 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 2255 94 2301 626 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 2869 94 2915 626 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal1 3092 16 3138 713 0 FreeSans 160 90 0 0 Vout
port 4 nsew
<< end >>
