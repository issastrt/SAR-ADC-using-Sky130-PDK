magic
tech sky130A
magscale 1 2
timestamp 1761392116
<< nwell >>
rect 1906 370 1948 1252
rect 3222 370 3264 1252
<< mvpsubdiff >>
rect 1954 238 2014 272
rect 3156 238 3216 272
rect 1954 212 1988 238
rect 1954 -402 1988 -376
rect 3182 212 3216 238
rect 3182 -402 3216 -376
rect 1954 -436 2014 -402
rect 3156 -436 3216 -402
<< mvpsubdiffcont >>
rect 2014 238 3156 272
rect 1954 -376 1988 212
rect 3182 -376 3216 212
rect 2014 -436 3156 -402
<< locali >>
rect 2122 1292 2434 1298
rect 2122 1258 2128 1292
rect 2428 1258 2434 1292
rect 2122 1140 2434 1258
rect 2736 1292 3048 1298
rect 2736 1258 2742 1292
rect 3042 1258 3048 1292
rect 2736 1140 3048 1258
rect 1954 238 2014 272
rect 3156 238 3216 272
rect 1954 212 1988 238
rect 1954 -402 1988 -376
rect 3182 212 3216 238
rect 3182 -402 3216 -376
rect 1954 -436 2014 -402
rect 3156 -436 3216 -402
rect 2050 -490 2506 -436
rect 2050 -524 2056 -490
rect 2500 -524 2506 -490
rect 2050 -530 2506 -524
rect 2664 -490 3120 -436
rect 2664 -524 2670 -490
rect 3114 -524 3120 -490
rect 2664 -530 3120 -524
<< viali >>
rect 2128 1258 2428 1292
rect 2742 1258 3042 1292
rect 2056 -524 2500 -490
rect 2670 -524 3114 -490
<< metal1 >>
rect 1906 1292 3264 1315
rect 1906 1258 2128 1292
rect 2428 1258 2742 1292
rect 3042 1258 3264 1292
rect 1906 1235 3264 1258
rect 2206 996 2350 1076
rect 2545 955 2625 1235
rect 2820 996 2964 1076
rect 2120 733 2200 955
rect 2120 681 2134 733
rect 2186 681 2200 733
rect 2120 667 2200 681
rect 2356 875 2814 955
rect 2356 667 2436 875
rect 2734 667 2814 875
rect 2970 747 3050 955
rect 2970 733 3206 747
rect 2970 681 2984 733
rect 3036 681 3206 733
rect 2970 667 3206 681
rect 2206 546 2350 626
rect 2820 546 2964 626
rect 2238 174 2318 546
rect 2852 174 2932 546
rect 2134 94 2422 174
rect 2748 94 3036 174
rect 3126 62 3206 667
rect 2048 -146 2128 62
rect 1964 -226 2128 -146
rect 2428 -146 2508 62
rect 2662 -146 2742 62
rect 2428 -226 2742 -146
rect 3042 -18 3206 62
rect 3042 -226 3122 -18
rect 1964 -467 2044 -226
rect 2134 -338 2422 -258
rect 2748 -338 3036 -258
rect 1906 -490 3264 -467
rect 1906 -524 2056 -490
rect 2500 -524 2670 -490
rect 3114 -524 3264 -490
rect 1906 -547 3264 -524
<< via1 >>
rect 2134 681 2186 733
rect 2984 681 3036 733
<< metal2 >>
rect 2120 733 3050 747
rect 2120 681 2134 733
rect 2186 681 2984 733
rect 3036 681 3050 733
rect 2120 667 3050 681
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1757220954
transform 1 0 2892 0 1 811
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM2
timestamp 1757220954
transform 1 0 2278 0 1 811
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM3
timestamp 1757220954
transform 1 0 2892 0 1 -82
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4
timestamp 1757220954
transform 1 0 2278 0 1 -82
box -372 -402 372 402
<< labels >>
flabel metal1 1906 -530 3264 -484 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 1906 1252 3264 1298 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 3126 -18 3206 747 0 FreeSans 160 0 0 0 Vout
port 4 nsew
flabel metal1 2852 94 2932 626 0 FreeSans 160 0 0 0 B
port 6 nsew
flabel metal1 2238 94 2318 626 0 FreeSans 160 0 0 0 A
port 2 nsew
<< end >>
