magic
tech sky130A
magscale 1 2
timestamp 1761375837
<< nwell >>
rect 2023 -528 2065 354
rect 3953 -528 3995 354
<< mvpsubdiff >>
rect 2071 -660 2131 -626
rect 3887 -660 3947 -626
rect 2071 -686 2105 -660
rect 2071 -1300 2105 -1274
rect 3913 -686 3947 -660
rect 3913 -1300 3947 -1274
rect 2071 -1334 2131 -1300
rect 3887 -1334 3947 -1300
<< mvpsubdiffcont >>
rect 2131 -660 3887 -626
rect 2071 -1274 2105 -686
rect 3913 -1274 3947 -686
rect 2131 -1334 3887 -1300
<< locali >>
rect 2239 394 2551 400
rect 2239 360 2245 394
rect 2545 360 2551 394
rect 2239 242 2551 360
rect 2853 394 3165 400
rect 2853 360 2859 394
rect 3159 360 3165 394
rect 2853 242 3165 360
rect 3467 394 3779 400
rect 3467 360 3473 394
rect 3773 360 3779 394
rect 3467 242 3779 360
rect 2071 -660 2131 -626
rect 3887 -660 3947 -626
rect 2071 -686 2105 -660
rect 2071 -1300 2105 -1274
rect 3913 -686 3947 -660
rect 3913 -1300 3947 -1274
rect 2071 -1334 2131 -1300
rect 3887 -1334 3947 -1300
rect 2167 -1388 2623 -1334
rect 2167 -1422 2173 -1388
rect 2617 -1422 2623 -1388
rect 2167 -1428 2623 -1422
rect 2781 -1388 3237 -1334
rect 2781 -1422 2787 -1388
rect 3231 -1422 3237 -1388
rect 2781 -1428 3237 -1422
rect 3395 -1388 3851 -1334
rect 3395 -1422 3401 -1388
rect 3845 -1422 3851 -1388
rect 3395 -1428 3851 -1422
<< viali >>
rect 2245 360 2545 394
rect 2859 360 3159 394
rect 3473 360 3773 394
rect 2173 -1422 2617 -1388
rect 2787 -1422 3231 -1388
rect 3401 -1422 3845 -1388
<< metal1 >>
rect 2023 394 3995 417
rect 2023 360 2245 394
rect 2545 360 2859 394
rect 3159 360 3473 394
rect 3773 360 3995 394
rect 2023 337 3995 360
rect 2153 57 2233 337
rect 2323 98 2467 178
rect 2937 98 3081 178
rect 3276 57 3356 337
rect 3551 98 3695 178
rect 2153 -23 2317 57
rect 2237 -231 2317 -23
rect 2473 -23 2931 57
rect 2473 -231 2553 -23
rect 2851 -165 2931 -23
rect 2851 -217 2865 -165
rect 2917 -217 2931 -165
rect 2851 -231 2931 -217
rect 3087 -23 3545 57
rect 3087 -231 3167 -23
rect 3465 -231 3545 -23
rect 3701 -151 3781 57
rect 3701 -165 3937 -151
rect 3701 -217 3715 -165
rect 3767 -217 3937 -165
rect 3701 -231 3937 -217
rect 2323 -352 2467 -272
rect 2937 -352 3081 -272
rect 3551 -352 3695 -272
rect 2355 -724 2435 -352
rect 2969 -724 3049 -352
rect 3583 -724 3663 -352
rect 2251 -804 2539 -724
rect 2865 -804 3153 -724
rect 3479 -804 3767 -724
rect 3857 -836 3937 -231
rect 2165 -1044 2245 -836
rect 2081 -1124 2245 -1044
rect 2545 -1044 2625 -836
rect 2779 -1044 2859 -836
rect 2545 -1124 2859 -1044
rect 3159 -1044 3239 -836
rect 3393 -1044 3473 -836
rect 3159 -1124 3473 -1044
rect 3773 -916 3937 -836
rect 3773 -1124 3853 -916
rect 2081 -1365 2161 -1124
rect 2251 -1236 2539 -1156
rect 2865 -1236 3153 -1156
rect 3479 -1236 3767 -1156
rect 2023 -1388 3995 -1365
rect 2023 -1422 2173 -1388
rect 2617 -1422 2787 -1388
rect 3231 -1422 3401 -1388
rect 3845 -1422 3995 -1388
rect 2023 -1445 3995 -1422
<< via1 >>
rect 2865 -217 2917 -165
rect 3715 -217 3767 -165
<< metal2 >>
rect 2851 -165 3781 -151
rect 2851 -217 2865 -165
rect 2917 -217 3715 -165
rect 3767 -217 3781 -165
rect 2851 -231 3781 -217
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1757220954
transform 1 0 3623 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM2
timestamp 1757220954
transform 1 0 3009 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM3
timestamp 1757220954
transform 1 0 2395 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4
timestamp 1757220954
transform 1 0 3623 0 1 -980
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM5
timestamp 1757220954
transform 1 0 3009 0 1 -980
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM6
timestamp 1757220954
transform 1 0 2395 0 1 -980
box -372 -402 372 402
<< labels >>
flabel metal1 2023 -1428 3995 -1382 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 2023 354 3995 400 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 2372 -804 2418 -272 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 2986 -804 3032 -272 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal1 3600 -804 3646 -272 0 FreeSans 160 0 0 0 C
port 4 nsew
flabel metal1 3857 -916 3937 -151 0 FreeSans 160 0 0 0 Vout
port 5 nsew
<< end >>
