** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/SAR-ADC-using-Sky130-PDK.sch
.subckt SAR-ADC-using-Sky130-PDK VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 GND
*.PININFO EN:I CLK:I VDD:I Vin:I Q0:O Q2:O Q3:O Q4:O Q5:O Q6:O Q7:O Q1:O Vbias:I GND:I
x2 net23 Compout Q0 net1 net32 FFCLR GND VDD D_FlipFlop_for_Ring
x4 net19 Compout Q2 net2 net33 FFCLR GND VDD D_FlipFlop_for_Ring
x5 net17 Compout Q3 net3 net34 FFCLR GND VDD D_FlipFlop_for_Ring
x6 net15 Compout Q4 net4 net35 FFCLR GND VDD D_FlipFlop_for_Ring
x7 net13 Compout Q5 net5 net36 FFCLR GND VDD D_FlipFlop_for_Ring
x8 net11 Compout Q6 net6 net37 FFCLR GND VDD D_FlipFlop_for_Ring
x9 FFCLR Compout Q7 net7 net38 EN GND VDD D_FlipFlop_for_Ring
x3 net21 Compout Q1 net8 net39 FFCLR GND VDD D_FlipFlop_for_Ring
x18 net9 net23 net30 GND VDD Nand_Gate
x19 net22 net21 net31 GND VDD Nand_Gate
x20 net20 net19 net25 GND VDD Nand_Gate
x21 net18 net17 net26 GND VDD Nand_Gate
x10 net30 CLK net1 GND VDD And_Gate
x27 DACout Q7 Q6 Q5 Q4 Q3 Q2 Q1 Q0 GND VDD CDAC8_v2
x1 Compout DACout Vin VDD Vbias comparator
x26 VDD net11 net9 net13 net14 net15 net16 net10 net18 net19 net20 net21 net22 net23 FFCLR net12 net17 CLK EN GND
+ RING_COUNTER_FINAL
* noconn #net32
* noconn #net39
* noconn #net33
* noconn #net34
* noconn #net36
* noconn #net35
* noconn #net37
* noconn #net38
x22 net16 net15 net27 GND VDD Nand_Gate
x23 net14 net13 net28 GND VDD Nand_Gate
x24 net12 net11 net29 GND VDD Nand_Gate
x25 net10 FFCLR net24 GND VDD Nand_Gate
x11 net31 CLK net8 GND VDD And_Gate
x12 net25 CLK net2 GND VDD And_Gate
x13 net26 CLK net3 GND VDD And_Gate
x14 net27 CLK net4 GND VDD And_Gate
x15 net28 CLK net5 GND VDD And_Gate
x16 net29 CLK net6 GND VDD And_Gate
x17 net24 CLK net7 GND VDD And_Gate
.ends

* expanding   symbol:  D_FlipFlop_for_Ring.sym # of pins=8
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/D_FlipFlop_for_Ring.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/D_FlipFlop_for_Ring.sch
.subckt D_FlipFlop_for_Ring nPRE D Q CLK Qbar nCLR GND VDD
*.PININFO D:I CLK:I nPRE:I nCLR:I Q:O Qbar:O VDD:I GND:I
x1 CLK net6 GND VDD Inverter
x2 CLK D nCLR net1 GND VDD 3-input-nand
x3 net4 net6 net7 GND VDD Nand_Gate
x4 CLK net5 nPRE net2 GND VDD 3-input-nand
x5 Q net8 nCLR Qbar GND VDD 3-input-nand
x6 Qbar net7 nPRE Q GND VDD 3-input-nand
x7 net3 net6 net8 GND VDD Nand_Gate
x8 net3 net1 nPRE net4 GND VDD 3-input-nand
x9 net4 net2 nCLR net3 GND VDD 3-input-nand
x10 D net5 GND VDD Inverter
.ends


* expanding   symbol:  Nand_Gate.sym # of pins=5
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/Nand_Gate.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/Nand_Gate.sch
.subckt Nand_Gate A B Vout GND VDD
*.PININFO A:I B:I VDD:I GND:I Vout:O
XM1 Vout B VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout A VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout B net1 GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 A GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  And_Gate.sym # of pins=5
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/And_Gate.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/And_Gate.sch
.subckt And_Gate A B Vout GND VDD
*.PININFO Vout:O A:I B:I VDD:I GND:I
XM1 net1 B VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 A VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 B net2 GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 A GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vout net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout net1 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CDAC8_v2.sym # of pins=11
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/CDAC8_v2.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/CDAC8_v2.sch
.subckt CDAC8_v2 OUT b7 b6 b5 b4 b3 b2 b1 b0 GND VDD
*.PININFO b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I VDD:I GND:I OUT:O
x1 VDD GND net1 b0 VDD GND switch_symbol
x2 VDD GND net2 b1 VDD GND switch_symbol
x3 VDD GND net3 b2 VDD GND switch_symbol
x4 VDD GND net4 b3 VDD GND switch_symbol
x5 VDD GND net5 b4 VDD GND switch_symbol
x6 VDD GND net6 b5 VDD GND switch_symbol
x7 VDD GND net7 b6 VDD GND switch_symbol
x8 VDD GND net8 b7 VDD GND switch_symbol
XC0 OUT net1 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=1 m=1
XC1 OUT net2 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=2 m=2
XC2 OUT net3 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=4 m=4
XC3 OUT net4 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=8 m=8
XC4 OUT net5 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=16 m=16
XC5 OUT net6 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=32 m=32
XC6 OUT net7 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=64 m=64
XC7 OUT net8 sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=128 m=128
XC8 GND GND sky130_fd_pr__cap_mim_m3_1 W=6.88 L=6.88 MF=68 m=68
.ends


* expanding   symbol:  comparator.sym # of pins=5
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/comparator.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/comparator.sch
.subckt comparator Vout Vinm Vinp VDD VSS
*.PININFO Vout:O Vinp:I Vinm:I VDD:I VSS:I
XM9 Vout net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=60 nf=1 ad=17.4 as=17.4 pd=120.58 ps=120.58 nrd=0.00483333333333333
+ nrs=0.00483333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058 nrs=0.0058 sa=0
+ sb=0 sd=0 mult=1 m=1
XM4 net2 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=1 ad=14.5 as=14.5 pd=100.58 ps=100.58 nrd=0.0058 nrs=0.0058 sa=0
+ sb=0 sd=0 mult=1 m=1
XM1 net1 Vinm net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=15 nf=1 ad=4.35 as=4.35 pd=30.58 ps=30.58 nrd=0.0193333333333333
+ nrs=0.0193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 Vinp net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=15 nf=1 ad=4.35 as=4.35 pd=30.58 ps=30.58 nrd=0.0193333333333333
+ nrs=0.0193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad=2.9 as=2.9 pd=20.58 ps=20.58 nrd=0.029 nrs=0.029 sa=0 sb=0
+ sd=0 mult=1 m=1
XM5 net3 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=1 ad=5.8 as=5.8 pd=40.58 ps=40.58 nrd=0.0145 nrs=0.0145 sa=0 sb=0
+ sd=0 mult=1 m=1
XM7 net4 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=20 nf=1 ad=5.8 as=5.8 pd=40.58 ps=40.58 nrd=0.0145 nrs=0.0145 sa=0 sb=0
+ sd=0 mult=1 m=1
XR1 net4 VDD VSS sky130_fd_pr__res_xhigh_po_5p73 L=150 mult=1 m=1
XC3 net2 Vout sky130_fd_pr__cap_mim_m3_2 W=5.35 L=2 MF=1 m=1
XC1 Vout VSS sky130_fd_pr__cap_mim_m3_2 W=5.35 L=2 MF=1 m=1
.ends


* expanding   symbol:  RING_COUNTER_FINAL.sym # of pins=20
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/RING_COUNTER_FINAL.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/RING_COUNTER_FINAL.sch
.subckt RING_COUNTER_FINAL VDD Q2 Q15 Q4 Q5 Q6 Q7 Q1 Q9 Q10 Q11 Q12 Q13 Q14 Q0 Q3 Q8 CLK EN GND
*.PININFO Q0:O Q1:O Q2:O Q3:O Q4:O Q5:O Q6:O Q7:O Q8:O Q9:O Q10:O Q11:O Q12:O Q13:O Q14:O Q15:O CLK:I EN:I VDD:I GND:I
x1 VDD net1 Q0 CLK net2 EN GND VDD D_FlipFlop_for_Ring
x2 EN Q0 Q1 CLK net3 VDD GND VDD D_FlipFlop_for_Ring
x3 EN Q1 Q2 CLK net4 VDD GND VDD D_FlipFlop_for_Ring
x4 EN Q2 Q3 CLK net5 VDD GND VDD D_FlipFlop_for_Ring
x5 EN Q3 Q4 CLK net6 VDD GND VDD D_FlipFlop_for_Ring
x6 EN Q4 Q5 CLK net7 VDD GND VDD D_FlipFlop_for_Ring
x7 EN Q5 Q6 CLK net8 VDD GND VDD D_FlipFlop_for_Ring
x8 EN Q6 Q7 CLK net9 VDD GND VDD D_FlipFlop_for_Ring
x9 EN Q7 Q8 CLK net10 VDD GND VDD D_FlipFlop_for_Ring
x10 EN Q8 Q9 CLK net11 VDD GND VDD D_FlipFlop_for_Ring
x11 EN Q9 Q10 CLK net12 VDD GND VDD D_FlipFlop_for_Ring
x12 EN Q10 Q11 CLK net13 VDD GND VDD D_FlipFlop_for_Ring
x13 EN Q11 Q12 CLK net14 VDD GND VDD D_FlipFlop_for_Ring
x14 EN Q12 Q13 CLK net15 VDD GND VDD D_FlipFlop_for_Ring
x15 EN Q13 Q14 CLK net16 VDD GND VDD D_FlipFlop_for_Ring
x16 EN Q14 Q15 CLK net17 VDD GND VDD D_FlipFlop_for_Ring
x17 EN Q15 net1 CLK net18 VDD GND VDD D_FlipFlop_for_Ring
* noconn #net2
* noconn #net3
* noconn #net4
* noconn #net5
* noconn #net6
* noconn #net7
* noconn #net8
* noconn #net9
* noconn #net10
* noconn #net11
* noconn #net12
* noconn #net13
* noconn #net14
* noconn #net18
* noconn #net17
* noconn #net16
* noconn #net15
.ends


* expanding   symbol:  Inverter.sym # of pins=4
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/Inverter.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/Inverter.sch
.subckt Inverter Vin Vout GND VDD
*.PININFO Vout:O Vin:I VDD:I GND:I
XM1 Vout Vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  3-input-nand.sym # of pins=6
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/3-input-nand.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/3-input-nand.sch
.subckt 3-input-nand C B A Vout GND VDD
*.PININFO A:I B:I Vout:O C:I VDD:I GND:I
XM1 Vout C VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout B VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout A VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vout C net1 GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 B net2 GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 A GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  switch_symbol.sym # of pins=6
** sym_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/switch_symbol.sym
** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/xschem/switch_symbol.sch
.subckt switch_symbol B A Z Vref VDD GND
*.PININFO Vref:I Z:B A:B B:B VDD:I GND:I
XM2 Z Vref B GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM1 B net1 Z VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM3 A Vref Z VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 Vref VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.720 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM4 Z net1 A GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 Vref GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1.44 W=1.44 nf=1 ad=0.4176 as=0.4176 pd=3.46 ps=3.46 nrd=0.201388888888889
+ nrs=0.201388888888889 sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
