magic
tech sky130A
magscale 1 2
timestamp 1757220954
<< nwell >>
rect 1296 -684 1338 198
rect 1961 -503 1989 -3
rect 3226 -684 3268 198
<< mvpsubdiff >>
rect 1344 -816 1404 -782
rect 3160 -816 3220 -782
rect 1344 -842 1378 -816
rect 1344 -1456 1378 -1430
rect 3186 -842 3220 -816
rect 3186 -1456 3220 -1430
rect 1344 -1490 1404 -1456
rect 3160 -1490 3220 -1456
<< mvpsubdiffcont >>
rect 1404 -816 3160 -782
rect 1344 -1430 1378 -842
rect 3186 -1430 3220 -842
rect 1404 -1490 3160 -1456
<< locali >>
rect 1512 238 1824 244
rect 1512 204 1518 238
rect 1818 204 1824 238
rect 1512 86 1824 204
rect 2126 238 2438 244
rect 2126 204 2132 238
rect 2432 204 2438 238
rect 2126 86 2438 204
rect 2740 238 3052 244
rect 2740 204 2746 238
rect 3046 204 3052 238
rect 2740 86 3052 204
rect 1344 -816 1404 -782
rect 3160 -816 3220 -782
rect 1344 -842 1378 -816
rect 1344 -1456 1378 -1430
rect 3186 -842 3220 -816
rect 3186 -1456 3220 -1430
rect 1344 -1490 1404 -1456
rect 3160 -1490 3220 -1456
rect 1440 -1544 1896 -1490
rect 1440 -1578 1446 -1544
rect 1890 -1578 1896 -1544
rect 1440 -1584 1896 -1578
rect 2054 -1544 2510 -1490
rect 2054 -1578 2060 -1544
rect 2504 -1578 2510 -1544
rect 2054 -1584 2510 -1578
rect 2668 -1544 3124 -1490
rect 2668 -1578 2674 -1544
rect 3118 -1578 3124 -1544
rect 2668 -1584 3124 -1578
<< viali >>
rect 1518 204 1818 238
rect 2132 204 2432 238
rect 2746 204 3046 238
rect 1446 -1578 1890 -1544
rect 2060 -1578 2504 -1544
rect 2674 -1578 3118 -1544
<< metal1 >>
rect 1296 238 3268 244
rect 1296 204 1518 238
rect 1818 204 2132 238
rect 2432 204 2746 238
rect 3046 204 3268 238
rect 1296 198 3268 204
rect 2724 -99 2770 198
rect 2351 -105 2415 -99
rect 2351 -157 2357 -105
rect 2409 -157 2415 -105
rect 2724 -145 2772 -99
rect 2351 -163 2415 -157
rect 1535 -329 1599 -323
rect 1535 -381 1541 -329
rect 1593 -381 1599 -329
rect 1535 -387 1599 -381
rect 1791 -387 2190 -341
rect 3014 -387 3140 -341
rect 1645 -767 1691 -448
rect 1636 -773 1700 -767
rect 1636 -825 1642 -773
rect 1694 -825 1700 -773
rect 1636 -831 1700 -825
rect 1645 -948 1691 -831
rect 1463 -994 1527 -988
rect 1952 -992 1998 -387
rect 2259 -566 2305 -440
rect 2873 -566 2919 -442
rect 2259 -612 2919 -566
rect 2259 -940 2305 -612
rect 2873 -942 2919 -612
rect 3094 -767 3140 -387
rect 3085 -773 3149 -767
rect 3085 -825 3091 -773
rect 3143 -825 3149 -773
rect 3085 -831 3149 -825
rect 3094 -992 3140 -831
rect 1463 -1046 1469 -994
rect 1521 -1046 1527 -994
rect 1863 -1020 2092 -992
rect 1864 -1038 2092 -1020
rect 3086 -1038 3140 -992
rect 1463 -1052 1527 -1046
rect 2423 -1222 2487 -1216
rect 2423 -1274 2429 -1222
rect 2481 -1274 2487 -1222
rect 2423 -1280 2487 -1274
rect 2652 -1280 2700 -1234
rect 2652 -1538 2698 -1280
rect 1296 -1544 3268 -1538
rect 1296 -1578 1446 -1544
rect 1890 -1578 2060 -1544
rect 2504 -1578 2674 -1544
rect 3118 -1578 3268 -1544
rect 1296 -1584 3268 -1578
<< via1 >>
rect 2357 -157 2409 -105
rect 1541 -381 1593 -329
rect 1642 -825 1694 -773
rect 3091 -825 3143 -773
rect 1469 -1046 1521 -994
rect 2429 -1274 2481 -1222
<< metal2 >>
rect 2083 -103 2157 -94
rect 2083 -159 2092 -103
rect 2148 -108 2157 -103
rect 2351 -105 2415 -99
rect 2351 -108 2357 -105
rect 2148 -154 2357 -108
rect 2148 -159 2157 -154
rect 2083 -168 2157 -159
rect 2351 -157 2357 -154
rect 2409 -157 2415 -105
rect 2351 -163 2415 -157
rect 1535 -329 1599 -323
rect 1535 -381 1541 -329
rect 1593 -332 1599 -329
rect 1793 -327 1867 -318
rect 1793 -332 1802 -327
rect 1593 -378 1802 -332
rect 1593 -381 1599 -378
rect 1535 -387 1599 -381
rect 1793 -383 1802 -378
rect 1858 -383 1867 -327
rect 1793 -392 1867 -383
rect 1636 -773 1700 -767
rect 1636 -825 1642 -773
rect 1694 -776 1700 -773
rect 3085 -773 3149 -767
rect 3085 -776 3091 -773
rect 1694 -822 3091 -776
rect 1694 -825 1700 -822
rect 1636 -831 1700 -825
rect 3085 -825 3091 -822
rect 3143 -825 3149 -773
rect 3085 -831 3149 -825
rect 1463 -994 1527 -988
rect 1463 -1046 1469 -994
rect 1521 -997 1527 -994
rect 2083 -992 2157 -983
rect 2083 -997 2092 -992
rect 1521 -1043 2092 -997
rect 1521 -1046 1527 -1043
rect 1463 -1052 1527 -1046
rect 2083 -1048 2092 -1043
rect 2148 -1048 2157 -992
rect 2083 -1057 2157 -1048
rect 1793 -1220 1867 -1211
rect 1793 -1276 1802 -1220
rect 1858 -1225 1867 -1220
rect 2423 -1222 2487 -1216
rect 2423 -1225 2429 -1222
rect 1858 -1271 2429 -1225
rect 1858 -1276 1867 -1271
rect 1793 -1285 1867 -1276
rect 2423 -1274 2429 -1271
rect 2481 -1274 2487 -1222
rect 2423 -1280 2487 -1274
<< via2 >>
rect 2092 -159 2148 -103
rect 1802 -383 1858 -327
rect 2092 -1048 2148 -992
rect 1802 -1276 1858 -1220
<< metal3 >>
rect 2087 -103 2153 -98
rect 2087 -159 2092 -103
rect 2148 -159 2153 -103
rect 2087 -164 2153 -159
rect 1797 -327 1863 -322
rect 1797 -383 1802 -327
rect 1858 -383 1863 -327
rect 1797 -388 1863 -383
rect 1800 -1215 1860 -388
rect 2090 -987 2150 -164
rect 2087 -992 2153 -987
rect 2087 -1048 2092 -992
rect 2148 -1048 2153 -992
rect 2087 -1053 2153 -1048
rect 1797 -1220 1863 -1215
rect 1797 -1276 1802 -1220
rect 1858 -1276 1863 -1220
rect 1797 -1281 1863 -1276
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1757220954
transform 1 0 1668 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM2
timestamp 1757220954
transform 1 0 2282 0 1 -1136
box -372 -402 372 402
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM3
timestamp 1757220954
transform 1 0 2282 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4
timestamp 1757220954
transform 1 0 1668 0 1 -1136
box -372 -402 372 402
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM5
timestamp 1757220954
transform 1 0 2896 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM6
timestamp 1757220954
transform 1 0 2896 0 1 -1136
box -372 -402 372 402
<< labels >>
flabel metal1 1296 -1584 3268 -1538 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 1296 198 3268 244 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 2259 -612 2919 -566 0 FreeSans 160 0 0 0 Vref
port 6 nsew
flabel metal1 1952 -1038 1998 -341 0 FreeSans 160 0 0 0 Z
port 2 nsew
flabel metal3 2090 -992 2150 -159 0 FreeSans 160 0 0 0 A
port 3 nsew
flabel metal3 1800 -1220 1860 -383 0 FreeSans 160 0 0 0 B
port 4 nsew
<< end >>
