magic
tech sky130A
magscale 1 2
timestamp 1757047045
<< nwell >>
rect 61005 48259 61079 48271
rect 83085 48259 83159 48271
<< pwell >>
rect 61005 48197 61079 48209
rect 83085 48197 83159 48209
<< metal1 >>
rect 127370 49190 127434 49196
rect 127370 49187 127376 49190
rect 48421 49141 127376 49187
rect 127370 49138 127376 49141
rect 127428 49138 127434 49190
rect 127370 49132 127434 49138
rect 49375 48518 49439 48524
rect 49375 48466 49381 48518
rect 49433 48466 49439 48518
rect 49375 48460 49439 48466
rect 71455 48518 71519 48524
rect 71455 48466 71461 48518
rect 71513 48466 71519 48518
rect 71455 48460 71519 48466
rect 93535 48518 93599 48524
rect 93535 48466 93541 48518
rect 93593 48466 93599 48518
rect 93535 48460 93599 48466
rect 115615 48518 115679 48524
rect 115615 48466 115621 48518
rect 115673 48466 115679 48518
rect 115615 48460 115679 48466
rect 61019 48266 61065 48271
rect 83099 48266 83145 48271
rect 48761 48260 48825 48266
rect 48761 48208 48767 48260
rect 48819 48208 48825 48260
rect 48761 48202 48825 48208
rect 49598 48260 49662 48266
rect 49598 48208 49604 48260
rect 49656 48208 49662 48260
rect 49598 48202 49662 48208
rect 59429 48260 59493 48266
rect 59429 48208 59435 48260
rect 59487 48208 59493 48260
rect 59429 48202 59493 48208
rect 61010 48260 61074 48266
rect 61010 48208 61016 48260
rect 61068 48208 61074 48260
rect 61010 48202 61074 48208
rect 70841 48260 70905 48266
rect 70841 48208 70847 48260
rect 70899 48208 70905 48260
rect 70841 48202 70905 48208
rect 71678 48260 71742 48266
rect 71678 48208 71684 48260
rect 71736 48208 71742 48260
rect 71678 48202 71742 48208
rect 81509 48260 81573 48266
rect 81509 48208 81515 48260
rect 81567 48208 81573 48260
rect 81509 48202 81573 48208
rect 83090 48260 83154 48266
rect 83090 48208 83096 48260
rect 83148 48208 83154 48260
rect 83090 48202 83154 48208
rect 92921 48260 92985 48266
rect 92921 48208 92927 48260
rect 92979 48208 92985 48260
rect 92921 48202 92985 48208
rect 93758 48260 93822 48266
rect 93758 48208 93764 48260
rect 93816 48208 93822 48260
rect 93758 48202 93822 48208
rect 103589 48260 103653 48266
rect 103589 48208 103595 48260
rect 103647 48208 103653 48260
rect 103589 48202 103653 48208
rect 105170 48260 105234 48266
rect 105170 48208 105176 48260
rect 105228 48208 105234 48260
rect 105170 48202 105234 48208
rect 115001 48260 115065 48266
rect 115001 48208 115007 48260
rect 115059 48208 115065 48260
rect 115001 48202 115065 48208
rect 115838 48260 115902 48266
rect 115838 48208 115844 48260
rect 115896 48208 115902 48260
rect 115838 48202 115902 48208
rect 125669 48260 125733 48266
rect 125669 48208 125675 48260
rect 125727 48208 125733 48260
rect 125669 48202 125733 48208
rect 61019 48197 61065 48202
rect 83099 48197 83145 48202
rect 60043 48032 60107 48038
rect 60043 47980 60049 48032
rect 60101 47980 60107 48032
rect 60043 47974 60107 47980
rect 82123 48032 82187 48038
rect 82123 47980 82129 48032
rect 82181 47980 82187 48032
rect 82123 47974 82187 47980
rect 104203 48032 104267 48038
rect 104203 47980 104209 48032
rect 104261 47980 104267 48032
rect 104203 47974 104267 47980
rect 126283 48032 126347 48038
rect 126283 47980 126289 48032
rect 126341 47980 126347 48032
rect 126283 47974 126347 47980
rect 127250 47954 127314 47960
rect 127250 47902 127256 47954
rect 127308 47902 127314 47954
rect 127250 47896 127314 47902
rect 138272 47860 138336 47866
rect 138272 47808 138278 47860
rect 138330 47808 138336 47860
rect 138272 47802 138336 47808
rect 116382 47408 116446 47414
rect 116382 47405 116388 47408
rect 29386 47359 116388 47405
rect 116381 47356 116388 47359
rect 116440 47405 116446 47408
rect 127627 47405 127721 47441
rect 116440 47359 125339 47405
rect 127431 47395 127721 47405
rect 127431 47359 127673 47395
rect 116440 47356 116447 47359
rect 116381 47349 116447 47356
rect 77238 45668 77302 45674
rect 77238 45616 77244 45668
rect 77296 45616 77302 45668
rect 136643 45662 136707 45668
rect 136643 45659 136649 45662
rect 77238 45610 77302 45616
rect 127721 45613 136649 45659
rect 136643 45610 136649 45613
rect 136701 45610 136707 45662
rect 136643 45604 136707 45610
rect 77581 44996 77645 45002
rect 77581 44944 77587 44996
rect 77639 44944 77645 44996
rect 77581 44938 77645 44944
rect 77238 42121 77302 42127
rect 77238 42069 77244 42121
rect 77296 42069 77302 42121
rect 136643 42098 136707 42104
rect 136643 42095 136649 42098
rect 77238 42063 77302 42069
rect 127721 42049 136649 42095
rect 136643 42046 136649 42049
rect 136701 42046 136707 42098
rect 136643 42040 136707 42046
rect 77581 41865 77645 41871
rect 77581 41813 77587 41865
rect 77639 41813 77645 41865
rect 77581 41807 77645 41813
rect 77238 38549 77302 38555
rect 77238 38497 77244 38549
rect 77296 38497 77302 38549
rect 136643 38534 136707 38540
rect 136643 38531 136649 38534
rect 77238 38491 77302 38497
rect 127721 38485 136649 38531
rect 136643 38482 136649 38485
rect 136701 38482 136707 38534
rect 136643 38476 136707 38482
rect 77581 38293 77645 38299
rect 77581 38241 77587 38293
rect 77639 38241 77645 38293
rect 77581 38235 77645 38241
rect 77238 34977 77302 34983
rect 77238 34925 77244 34977
rect 77296 34925 77302 34977
rect 136643 34970 136707 34976
rect 136643 34967 136649 34970
rect 77238 34919 77302 34925
rect 136483 34921 136649 34967
rect 136643 34918 136649 34921
rect 136701 34918 136707 34970
rect 136643 34912 136707 34918
rect 77581 34721 77645 34727
rect 77581 34669 77587 34721
rect 77639 34669 77645 34721
rect 77581 34663 77645 34669
rect 136643 29291 136707 29297
rect 136643 29288 136649 29291
rect 136483 29242 136649 29288
rect 136643 29239 136649 29242
rect 136701 29239 136707 29291
rect 136643 29233 136707 29239
rect 77238 29133 77302 29139
rect 77238 29081 77244 29133
rect 77296 29081 77302 29133
rect 77238 29075 77302 29081
rect 77581 27577 77645 27583
rect 77581 27525 77587 27577
rect 77639 27525 77645 27577
rect 77581 27519 77645 27525
rect 136643 25727 136707 25733
rect 136643 25724 136649 25727
rect 127721 25678 136649 25724
rect 136643 25675 136649 25678
rect 136701 25675 136707 25727
rect 136643 25669 136707 25675
rect 77238 25561 77302 25567
rect 77238 25509 77244 25561
rect 77296 25509 77302 25561
rect 77238 25503 77302 25509
rect 77581 24005 77645 24011
rect 77581 23953 77587 24005
rect 77639 23953 77645 24005
rect 77581 23947 77645 23953
rect 136643 22163 136707 22169
rect 136643 22160 136649 22163
rect 127721 22114 136649 22160
rect 136643 22111 136649 22114
rect 136701 22111 136707 22163
rect 136643 22105 136707 22111
rect 77238 21985 77302 21991
rect 77238 21933 77244 21985
rect 77296 21933 77302 21985
rect 77238 21927 77302 21933
rect 77581 20429 77645 20435
rect 77581 20377 77587 20429
rect 77639 20377 77645 20429
rect 77581 20371 77645 20377
rect 136088 19222 136134 19754
rect 77238 18873 77302 18879
rect 77238 18821 77244 18873
rect 77296 18821 77302 18873
rect 77238 18815 77302 18821
rect 77679 18647 77743 18653
rect 77679 18595 77685 18647
rect 77737 18595 77743 18647
rect 136643 18599 136707 18605
rect 136643 18596 136649 18599
rect 77679 18589 77743 18595
rect 127721 18550 136649 18596
rect 136643 18547 136649 18550
rect 136701 18547 136707 18599
rect 136643 18541 136707 18547
rect 115620 18502 115684 18508
rect 115620 18499 115626 18502
rect 37381 18453 115626 18499
rect 115620 18450 115626 18453
rect 115678 18499 115684 18502
rect 115678 18453 116391 18499
rect 115678 18450 115684 18453
rect 115620 18444 115684 18450
rect 49970 17917 50034 17923
rect 49970 17865 49976 17917
rect 50028 17865 50034 17917
rect 49970 17859 50034 17865
rect 72050 17917 72114 17923
rect 72050 17865 72056 17917
rect 72108 17865 72114 17917
rect 72050 17859 72114 17865
rect 94130 17917 94194 17923
rect 94130 17865 94136 17917
rect 94188 17865 94194 17917
rect 94130 17859 94194 17865
rect 116210 17917 116274 17923
rect 116210 17865 116216 17917
rect 116268 17865 116274 17917
rect 116210 17859 116274 17865
rect 48389 17830 48453 17836
rect 48389 17778 48395 17830
rect 48447 17778 48453 17830
rect 48389 17772 48453 17778
rect 70469 17830 70533 17836
rect 70469 17778 70475 17830
rect 70527 17778 70533 17830
rect 70469 17772 70533 17778
rect 92549 17830 92613 17836
rect 92549 17778 92555 17830
rect 92607 17778 92613 17830
rect 92549 17772 92613 17778
rect 114629 17830 114693 17836
rect 114629 17778 114635 17830
rect 114687 17778 114693 17830
rect 114629 17772 114693 17778
rect 37721 17572 37785 17578
rect 37721 17520 37727 17572
rect 37779 17520 37785 17572
rect 37721 17514 37785 17520
rect 38558 17572 38622 17578
rect 38558 17520 38564 17572
rect 38616 17520 38622 17572
rect 38558 17514 38622 17520
rect 49003 17572 49067 17578
rect 49003 17520 49009 17572
rect 49061 17520 49067 17572
rect 49003 17514 49067 17520
rect 59801 17572 59865 17578
rect 59801 17520 59807 17572
rect 59859 17520 59865 17572
rect 59801 17514 59865 17520
rect 60638 17572 60702 17578
rect 60638 17520 60644 17572
rect 60696 17520 60702 17572
rect 60638 17514 60702 17520
rect 71083 17572 71147 17578
rect 71083 17520 71089 17572
rect 71141 17520 71147 17572
rect 71083 17514 71147 17520
rect 81881 17572 81945 17578
rect 81881 17520 81887 17572
rect 81939 17520 81945 17572
rect 81881 17514 81945 17520
rect 82718 17572 82782 17578
rect 82718 17520 82724 17572
rect 82776 17520 82782 17572
rect 82718 17514 82782 17520
rect 93163 17572 93227 17578
rect 93163 17520 93169 17572
rect 93221 17520 93227 17572
rect 93163 17514 93227 17520
rect 103961 17572 104025 17578
rect 103961 17520 103967 17572
rect 104019 17520 104025 17572
rect 103961 17514 104025 17520
rect 104798 17572 104862 17578
rect 104798 17520 104804 17572
rect 104856 17520 104862 17572
rect 104798 17514 104862 17520
rect 115243 17572 115307 17578
rect 115243 17520 115249 17572
rect 115301 17520 115307 17572
rect 115243 17514 115307 17520
rect 38335 17344 38399 17350
rect 38335 17292 38341 17344
rect 38393 17292 38399 17344
rect 38335 17286 38399 17292
rect 60415 17344 60479 17350
rect 60415 17292 60421 17344
rect 60473 17292 60479 17344
rect 60415 17286 60479 17292
rect 82495 17344 82559 17350
rect 82495 17292 82501 17344
rect 82553 17292 82559 17344
rect 82495 17286 82559 17292
rect 104575 17344 104639 17350
rect 104575 17292 104581 17344
rect 104633 17292 104639 17344
rect 104575 17286 104639 17292
rect 77679 16720 77743 16726
rect 77679 16717 77685 16720
rect 37381 16671 77685 16717
rect 77679 16668 77685 16671
rect 77737 16717 77743 16720
rect 114836 16720 114900 16726
rect 114836 16717 114842 16720
rect 77737 16671 114842 16717
rect 77737 16668 77743 16671
rect 77679 16662 77743 16668
rect 114836 16668 114842 16671
rect 114894 16717 114900 16720
rect 114894 16671 116391 16717
rect 114894 16668 114900 16671
rect 114836 16662 114900 16668
rect 140592 16601 140991 16647
rect 142718 16601 142802 16647
rect 125180 14610 125244 14616
rect 125180 14558 125186 14610
rect 125238 14558 125244 14610
rect 125180 14552 125244 14558
<< via1 >>
rect 127376 49138 127428 49190
rect 49381 48466 49433 48518
rect 71461 48466 71513 48518
rect 93541 48466 93593 48518
rect 115621 48466 115673 48518
rect 48767 48208 48819 48260
rect 49604 48208 49656 48260
rect 59435 48208 59487 48260
rect 61016 48208 61068 48260
rect 70847 48208 70899 48260
rect 71684 48208 71736 48260
rect 81515 48208 81567 48260
rect 83096 48208 83148 48260
rect 92927 48208 92979 48260
rect 93764 48208 93816 48260
rect 103595 48208 103647 48260
rect 105176 48208 105228 48260
rect 115007 48208 115059 48260
rect 115844 48208 115896 48260
rect 125675 48208 125727 48260
rect 60049 47980 60101 48032
rect 82129 47980 82181 48032
rect 104209 47980 104261 48032
rect 126289 47980 126341 48032
rect 127256 47902 127308 47954
rect 138278 47808 138330 47860
rect 116388 47356 116440 47408
rect 77244 45616 77296 45668
rect 136649 45610 136701 45662
rect 77587 44944 77639 44996
rect 77244 42069 77296 42121
rect 136649 42046 136701 42098
rect 77587 41813 77639 41865
rect 77244 38497 77296 38549
rect 136649 38482 136701 38534
rect 77587 38241 77639 38293
rect 77244 34925 77296 34977
rect 136649 34918 136701 34970
rect 77587 34669 77639 34721
rect 136649 29239 136701 29291
rect 77244 29081 77296 29133
rect 77587 27525 77639 27577
rect 136649 25675 136701 25727
rect 77244 25509 77296 25561
rect 77587 23953 77639 24005
rect 136649 22111 136701 22163
rect 77244 21933 77296 21985
rect 77587 20377 77639 20429
rect 77244 18821 77296 18873
rect 77685 18595 77737 18647
rect 136649 18547 136701 18599
rect 115626 18450 115678 18502
rect 49976 17865 50028 17917
rect 72056 17865 72108 17917
rect 94136 17865 94188 17917
rect 116216 17865 116268 17917
rect 48395 17778 48447 17830
rect 70475 17778 70527 17830
rect 92555 17778 92607 17830
rect 114635 17778 114687 17830
rect 37727 17520 37779 17572
rect 38564 17520 38616 17572
rect 49009 17520 49061 17572
rect 59807 17520 59859 17572
rect 60644 17520 60696 17572
rect 71089 17520 71141 17572
rect 81887 17520 81939 17572
rect 82724 17520 82776 17572
rect 93169 17520 93221 17572
rect 103967 17520 104019 17572
rect 104804 17520 104856 17572
rect 115249 17520 115301 17572
rect 38341 17292 38393 17344
rect 60421 17292 60473 17344
rect 82501 17292 82553 17344
rect 104581 17292 104633 17344
rect 77685 16668 77737 16720
rect 114842 16668 114894 16720
rect 125186 14558 125238 14610
<< metal2 >>
rect 48122 52317 48196 52326
rect 48122 52261 48131 52317
rect 48187 52261 48196 52317
rect 48122 52252 48196 52261
rect 59162 52317 59236 52326
rect 59162 52261 59171 52317
rect 59227 52261 59236 52317
rect 59162 52252 59236 52261
rect 70202 52317 70276 52326
rect 70202 52261 70211 52317
rect 70267 52261 70276 52317
rect 70202 52252 70276 52261
rect 81242 52317 81316 52326
rect 81242 52261 81251 52317
rect 81307 52261 81316 52317
rect 81242 52252 81316 52261
rect 92282 52317 92356 52326
rect 92282 52261 92291 52317
rect 92347 52261 92356 52317
rect 92282 52252 92356 52261
rect 103322 52317 103396 52326
rect 103322 52261 103331 52317
rect 103387 52261 103396 52317
rect 103322 52252 103396 52261
rect 114362 52317 114436 52326
rect 114362 52261 114371 52317
rect 114427 52261 114436 52317
rect 114362 52252 114436 52261
rect 127370 49190 127434 49196
rect 127370 49138 127376 49190
rect 127428 49187 127434 49190
rect 136638 49192 136712 49201
rect 136638 49187 136647 49192
rect 127428 49141 136647 49187
rect 127428 49138 127434 49141
rect 127370 49132 127434 49138
rect 136638 49136 136647 49141
rect 136703 49136 136712 49192
rect 136638 49127 136712 49136
rect 49375 48518 49439 48524
rect 49375 48466 49381 48518
rect 49433 48515 49439 48518
rect 59162 48520 59236 48529
rect 59162 48515 59171 48520
rect 49433 48469 59171 48515
rect 49433 48466 49439 48469
rect 49375 48460 49439 48466
rect 59162 48464 59171 48469
rect 59227 48464 59236 48520
rect 59162 48455 59236 48464
rect 71455 48518 71519 48524
rect 71455 48466 71461 48518
rect 71513 48515 71519 48518
rect 81242 48520 81316 48529
rect 81242 48515 81251 48520
rect 71513 48469 81251 48515
rect 71513 48466 71519 48469
rect 71455 48460 71519 48466
rect 81242 48464 81251 48469
rect 81307 48464 81316 48520
rect 81242 48455 81316 48464
rect 93535 48518 93599 48524
rect 93535 48466 93541 48518
rect 93593 48515 93599 48518
rect 103322 48520 103396 48529
rect 103322 48515 103331 48520
rect 93593 48469 103331 48515
rect 93593 48466 93599 48469
rect 93535 48460 93599 48466
rect 103322 48464 103331 48469
rect 103387 48464 103396 48520
rect 103322 48455 103396 48464
rect 115615 48518 115679 48524
rect 115615 48466 115621 48518
rect 115673 48515 115679 48518
rect 124832 48520 124906 48529
rect 124832 48515 124841 48520
rect 115673 48469 124841 48515
rect 115673 48466 115679 48469
rect 115615 48460 115679 48466
rect 124832 48464 124841 48469
rect 124897 48464 124906 48520
rect 124832 48455 124906 48464
rect 48122 48262 48196 48271
rect 48122 48206 48131 48262
rect 48187 48257 48196 48262
rect 48761 48260 48825 48266
rect 48761 48257 48767 48260
rect 48187 48211 48767 48257
rect 48187 48206 48196 48211
rect 48122 48197 48196 48206
rect 48761 48208 48767 48211
rect 48819 48208 48825 48260
rect 48761 48202 48825 48208
rect 49598 48260 49662 48266
rect 49598 48208 49604 48260
rect 49656 48257 49662 48260
rect 59429 48260 59493 48266
rect 59429 48257 59435 48260
rect 49656 48211 59435 48257
rect 49656 48208 49662 48211
rect 49598 48202 49662 48208
rect 59429 48208 59435 48211
rect 59487 48208 59493 48260
rect 59429 48202 59493 48208
rect 61005 48262 61079 48271
rect 61005 48206 61014 48262
rect 61070 48206 61079 48262
rect 61005 48197 61079 48206
rect 70202 48262 70276 48271
rect 70202 48206 70211 48262
rect 70267 48257 70276 48262
rect 70841 48260 70905 48266
rect 70841 48257 70847 48260
rect 70267 48211 70847 48257
rect 70267 48206 70276 48211
rect 70202 48197 70276 48206
rect 70841 48208 70847 48211
rect 70899 48208 70905 48260
rect 70841 48202 70905 48208
rect 71678 48260 71742 48266
rect 71678 48208 71684 48260
rect 71736 48257 71742 48260
rect 81509 48260 81573 48266
rect 81509 48257 81515 48260
rect 71736 48211 81515 48257
rect 71736 48208 71742 48211
rect 71678 48202 71742 48208
rect 81509 48208 81515 48211
rect 81567 48208 81573 48260
rect 81509 48202 81573 48208
rect 83085 48262 83159 48271
rect 83085 48206 83094 48262
rect 83150 48206 83159 48262
rect 83085 48197 83159 48206
rect 92282 48262 92356 48271
rect 92282 48206 92291 48262
rect 92347 48257 92356 48262
rect 92921 48260 92985 48266
rect 92921 48257 92927 48260
rect 92347 48211 92927 48257
rect 92347 48206 92356 48211
rect 92282 48197 92356 48206
rect 92921 48208 92927 48211
rect 92979 48208 92985 48260
rect 92921 48202 92985 48208
rect 93758 48260 93822 48266
rect 93758 48208 93764 48260
rect 93816 48257 93822 48260
rect 103589 48260 103653 48266
rect 103589 48257 103595 48260
rect 93816 48211 103595 48257
rect 93816 48208 93822 48211
rect 93758 48202 93822 48208
rect 103589 48208 103595 48211
rect 103647 48208 103653 48260
rect 103589 48202 103653 48208
rect 105165 48262 105239 48271
rect 105165 48206 105174 48262
rect 105230 48206 105239 48262
rect 105165 48197 105239 48206
rect 114362 48262 114436 48271
rect 114362 48206 114371 48262
rect 114427 48257 114436 48262
rect 115001 48260 115065 48266
rect 115001 48257 115007 48260
rect 114427 48211 115007 48257
rect 114427 48206 114436 48211
rect 114362 48197 114436 48206
rect 115001 48208 115007 48211
rect 115059 48208 115065 48260
rect 115001 48202 115065 48208
rect 115838 48260 115902 48266
rect 115838 48208 115844 48260
rect 115896 48257 115902 48260
rect 125669 48260 125733 48266
rect 125669 48257 125675 48260
rect 115896 48211 125675 48257
rect 115896 48208 115902 48211
rect 115838 48202 115902 48208
rect 125669 48208 125675 48211
rect 125727 48208 125733 48260
rect 125669 48202 125733 48208
rect 60043 48032 60107 48038
rect 60043 48029 60049 48032
rect 59935 47983 60049 48029
rect 60043 47980 60049 47983
rect 60101 48029 60107 48032
rect 78587 48034 78661 48043
rect 78587 48029 78596 48034
rect 60101 47983 78596 48029
rect 60101 47980 60107 47983
rect 60043 47974 60107 47980
rect 78587 47978 78596 47983
rect 78652 48029 78661 48034
rect 82123 48032 82187 48038
rect 82123 48029 82129 48032
rect 78652 47983 82129 48029
rect 78652 47978 78661 47983
rect 78587 47969 78661 47978
rect 82123 47980 82129 47983
rect 82181 48029 82187 48032
rect 104203 48032 104267 48038
rect 104203 48029 104209 48032
rect 82181 47983 104209 48029
rect 82181 47980 82187 47983
rect 82123 47974 82187 47980
rect 104203 47980 104209 47983
rect 104261 48029 104267 48032
rect 115196 48034 115270 48043
rect 115196 48029 115205 48034
rect 104261 47983 115205 48029
rect 104261 47980 104267 47983
rect 104203 47974 104267 47980
rect 115196 47978 115205 47983
rect 115261 48029 115270 48034
rect 126283 48032 126347 48038
rect 126283 48029 126289 48032
rect 115261 47983 126289 48029
rect 115261 47978 115270 47983
rect 115196 47969 115270 47978
rect 126283 47980 126289 47983
rect 126341 48029 126347 48032
rect 126341 47983 126455 48029
rect 126341 47980 126347 47983
rect 126283 47974 126347 47980
rect 127245 47956 127319 47965
rect 127245 47900 127254 47956
rect 127310 47900 127319 47956
rect 127245 47891 127319 47900
rect 136638 47862 136712 47871
rect 136638 47806 136647 47862
rect 136703 47857 136712 47862
rect 138272 47860 138336 47866
rect 138272 47857 138278 47860
rect 136703 47811 138278 47857
rect 136703 47806 136712 47811
rect 136638 47797 136712 47806
rect 138272 47808 138278 47811
rect 138330 47808 138336 47860
rect 138272 47802 138336 47808
rect 116377 47410 116451 47419
rect 116377 47354 116386 47410
rect 116442 47354 116451 47410
rect 116377 47345 116451 47354
rect 136074 46594 136148 46603
rect 136074 46538 136083 46594
rect 136139 46538 136148 46594
rect 136074 46529 136148 46538
rect 77238 45668 77302 45674
rect 77238 45616 77244 45668
rect 77296 45665 77302 45668
rect 127955 45670 128029 45679
rect 127955 45665 127964 45670
rect 77296 45619 127964 45665
rect 77296 45616 77302 45619
rect 77238 45610 77302 45616
rect 127955 45614 127964 45619
rect 128020 45614 128029 45670
rect 127955 45605 128029 45614
rect 136638 45664 136712 45673
rect 136638 45608 136647 45664
rect 136703 45608 136712 45664
rect 136638 45599 136712 45608
rect 77581 44996 77645 45002
rect 77581 44944 77587 44996
rect 77639 44993 77645 44996
rect 77956 44998 78030 45007
rect 77956 44993 77965 44998
rect 77639 44947 77965 44993
rect 77639 44944 77645 44947
rect 77581 44938 77645 44944
rect 77956 44942 77965 44947
rect 78021 44942 78030 44998
rect 77956 44933 78030 44942
rect 136074 43030 136148 43039
rect 136074 42974 136083 43030
rect 136139 42974 136148 43030
rect 136074 42965 136148 42974
rect 77238 42121 77302 42127
rect 77238 42069 77244 42121
rect 77296 42118 77302 42121
rect 127955 42123 128029 42132
rect 127955 42118 127964 42123
rect 77296 42072 127964 42118
rect 77296 42069 77302 42072
rect 77238 42063 77302 42069
rect 127955 42067 127964 42072
rect 128020 42067 128029 42123
rect 127955 42058 128029 42067
rect 136638 42100 136712 42109
rect 136638 42044 136647 42100
rect 136703 42044 136712 42100
rect 136638 42035 136712 42044
rect 77581 41865 77645 41871
rect 77581 41813 77587 41865
rect 77639 41862 77645 41865
rect 77956 41867 78030 41876
rect 77956 41862 77965 41867
rect 77639 41816 77965 41862
rect 77639 41813 77645 41816
rect 77581 41807 77645 41813
rect 77956 41811 77965 41816
rect 78021 41811 78030 41867
rect 77956 41802 78030 41811
rect 136074 39466 136148 39475
rect 136074 39410 136083 39466
rect 136139 39410 136148 39466
rect 136074 39401 136148 39410
rect 77238 38549 77302 38555
rect 77238 38497 77244 38549
rect 77296 38546 77302 38549
rect 127955 38551 128029 38560
rect 127955 38546 127964 38551
rect 77296 38500 127964 38546
rect 77296 38497 77302 38500
rect 77238 38491 77302 38497
rect 127955 38495 127964 38500
rect 128020 38495 128029 38551
rect 127955 38486 128029 38495
rect 136638 38536 136712 38545
rect 136638 38480 136647 38536
rect 136703 38480 136712 38536
rect 136638 38471 136712 38480
rect 77581 38293 77645 38299
rect 77581 38241 77587 38293
rect 77639 38290 77645 38293
rect 77956 38295 78030 38304
rect 77956 38290 77965 38295
rect 77639 38244 77965 38290
rect 77639 38241 77645 38244
rect 77581 38235 77645 38241
rect 77956 38239 77965 38244
rect 78021 38239 78030 38295
rect 77956 38230 78030 38239
rect 136074 35902 136148 35911
rect 136074 35846 136083 35902
rect 136139 35846 136148 35902
rect 136074 35837 136148 35846
rect 134744 35425 134818 35434
rect 134744 35369 134753 35425
rect 134809 35420 134818 35425
rect 135010 35425 135084 35434
rect 135010 35420 135019 35425
rect 134809 35374 135019 35420
rect 134809 35369 134818 35374
rect 134744 35360 134818 35369
rect 135010 35369 135019 35374
rect 135075 35369 135084 35425
rect 135010 35360 135084 35369
rect 77238 34977 77302 34983
rect 77238 34925 77244 34977
rect 77296 34974 77302 34977
rect 127955 34974 128029 34981
rect 77296 34972 128029 34974
rect 77296 34928 127964 34972
rect 77296 34925 77302 34928
rect 77238 34919 77302 34925
rect 127955 34916 127964 34928
rect 128020 34916 128029 34972
rect 127955 34907 128029 34916
rect 136638 34972 136712 34981
rect 136638 34916 136647 34972
rect 136703 34916 136712 34972
rect 136638 34907 136712 34916
rect 77581 34721 77645 34727
rect 77581 34669 77587 34721
rect 77639 34718 77645 34721
rect 77956 34723 78030 34732
rect 77956 34718 77965 34723
rect 77639 34672 77965 34718
rect 77639 34669 77645 34672
rect 77581 34663 77645 34669
rect 77956 34667 77965 34672
rect 78021 34667 78030 34723
rect 77956 34658 78030 34667
rect 134744 32501 134818 32510
rect 134744 32445 134753 32501
rect 134809 32496 134818 32501
rect 135010 32501 135084 32510
rect 135010 32496 135019 32501
rect 134809 32450 135019 32496
rect 134809 32445 134818 32450
rect 134744 32436 134818 32445
rect 135010 32445 135019 32450
rect 135075 32445 135084 32501
rect 135010 32436 135084 32445
rect 136074 30223 136148 30232
rect 136074 30167 136083 30223
rect 136139 30167 136148 30223
rect 136074 30158 136148 30167
rect 136638 29293 136712 29302
rect 136638 29237 136647 29293
rect 136703 29237 136712 29293
rect 136638 29228 136712 29237
rect 77238 29133 77302 29139
rect 77238 29081 77244 29133
rect 77296 29130 77302 29133
rect 127955 29135 128029 29144
rect 127955 29130 127964 29135
rect 77296 29084 127964 29130
rect 77296 29081 77302 29084
rect 77238 29075 77302 29081
rect 127955 29079 127964 29084
rect 128020 29079 128029 29135
rect 127955 29046 128029 29079
rect 77581 27577 77645 27583
rect 77581 27525 77587 27577
rect 77639 27574 77645 27577
rect 77956 27579 78030 27588
rect 77956 27574 77965 27579
rect 77639 27528 77965 27574
rect 77639 27525 77645 27528
rect 77581 27519 77645 27525
rect 77956 27523 77965 27528
rect 78021 27523 78030 27579
rect 77956 27514 78030 27523
rect 136074 26659 136148 26668
rect 136074 26603 136083 26659
rect 136139 26603 136148 26659
rect 136074 26594 136148 26603
rect 136638 25729 136712 25738
rect 136638 25673 136647 25729
rect 136703 25673 136712 25729
rect 136638 25664 136712 25673
rect 77238 25561 77302 25567
rect 77238 25509 77244 25561
rect 77296 25557 77302 25561
rect 127955 25562 128029 25571
rect 127955 25557 127964 25562
rect 77296 25511 127964 25557
rect 77296 25509 77302 25511
rect 77238 25503 77302 25509
rect 127955 25506 127964 25511
rect 128020 25506 128029 25562
rect 127955 25482 128029 25506
rect 77581 24005 77645 24011
rect 77581 23953 77587 24005
rect 77639 24002 77645 24005
rect 77956 24007 78030 24016
rect 77956 24002 77965 24007
rect 77639 23956 77965 24002
rect 77639 23953 77645 23956
rect 77581 23947 77645 23953
rect 77956 23951 77965 23956
rect 78021 23951 78030 24007
rect 77956 23942 78030 23951
rect 136074 23095 136148 23104
rect 136074 23039 136083 23095
rect 136139 23039 136148 23095
rect 136074 23030 136148 23039
rect 136638 22165 136712 22174
rect 136638 22109 136647 22165
rect 136703 22109 136712 22165
rect 136638 22100 136712 22109
rect 77238 21985 77302 21991
rect 77238 21933 77244 21985
rect 77296 21982 77302 21985
rect 127955 21989 128029 21998
rect 127955 21982 127964 21989
rect 77296 21936 127964 21982
rect 77296 21933 77302 21936
rect 77238 21927 77302 21933
rect 127955 21933 127964 21936
rect 128020 21933 128029 21989
rect 127955 21918 128029 21933
rect 77581 20429 77645 20435
rect 77581 20377 77587 20429
rect 77639 20426 77645 20429
rect 77956 20431 78030 20440
rect 77956 20426 77965 20431
rect 77639 20380 77965 20426
rect 77639 20377 77645 20380
rect 77581 20371 77645 20377
rect 77956 20375 77965 20380
rect 78021 20375 78030 20431
rect 77956 20366 78030 20375
rect 136074 19531 136148 19540
rect 136074 19475 136083 19531
rect 136139 19475 136148 19531
rect 136074 19466 136148 19475
rect 77238 18873 77302 18879
rect 77238 18821 77244 18873
rect 77296 18870 77302 18873
rect 127955 18873 128029 18891
rect 127955 18870 127964 18873
rect 77296 18824 127964 18870
rect 77296 18821 77302 18824
rect 77238 18815 77302 18821
rect 127955 18817 127964 18824
rect 128020 18817 128029 18873
rect 127955 18808 128029 18817
rect 77674 18649 77748 18658
rect 77674 18593 77683 18649
rect 77739 18593 77748 18649
rect 77674 18584 77748 18593
rect 136638 18601 136712 18610
rect 136638 18545 136647 18601
rect 136703 18545 136712 18601
rect 136638 18536 136712 18545
rect 115615 18504 115689 18513
rect 115615 18448 115624 18504
rect 115680 18448 115689 18504
rect 115615 18439 115689 18448
rect 49965 17920 50039 17929
rect 49965 17864 49974 17920
rect 50030 17864 50039 17920
rect 49965 17855 50039 17864
rect 72045 17919 72119 17928
rect 72045 17863 72054 17919
rect 72110 17863 72119 17919
rect 72045 17855 72119 17863
rect 94125 17919 94199 17928
rect 94125 17863 94134 17919
rect 94190 17863 94199 17919
rect 94125 17855 94199 17863
rect 116205 17919 116279 17928
rect 116205 17863 116214 17919
rect 116270 17863 116279 17919
rect 116205 17854 116279 17863
rect 48389 17830 48453 17836
rect 48389 17827 48395 17830
rect 48353 17781 48395 17827
rect 48389 17778 48395 17781
rect 48447 17827 48453 17830
rect 70469 17830 70533 17836
rect 70469 17827 70475 17830
rect 48447 17781 70475 17827
rect 48447 17778 48453 17781
rect 48389 17772 48453 17778
rect 70469 17778 70475 17781
rect 70527 17827 70533 17830
rect 78587 17832 78661 17841
rect 78587 17827 78596 17832
rect 70527 17781 78596 17827
rect 70527 17778 70533 17781
rect 70469 17772 70533 17778
rect 78587 17776 78596 17781
rect 78652 17827 78661 17832
rect 92549 17830 92613 17836
rect 92549 17827 92555 17830
rect 78652 17781 92555 17827
rect 78652 17776 78661 17781
rect 78587 17767 78661 17776
rect 92549 17778 92555 17781
rect 92607 17827 92613 17830
rect 114629 17830 114693 17836
rect 114629 17827 114635 17830
rect 92607 17781 114635 17827
rect 92607 17778 92613 17781
rect 92549 17772 92613 17778
rect 114629 17778 114635 17781
rect 114687 17827 114693 17830
rect 115196 17832 115270 17841
rect 115196 17827 115205 17832
rect 114687 17781 115205 17827
rect 114687 17778 114693 17781
rect 114629 17772 114693 17778
rect 115196 17776 115205 17781
rect 115261 17776 115270 17832
rect 115196 17767 115270 17776
rect 37177 17574 37251 17583
rect 37177 17518 37186 17574
rect 37242 17569 37251 17574
rect 37721 17572 37785 17578
rect 37721 17569 37727 17572
rect 37242 17523 37727 17569
rect 37242 17518 37251 17523
rect 37177 17509 37251 17518
rect 37721 17520 37727 17523
rect 37779 17520 37785 17572
rect 37721 17514 37785 17520
rect 38558 17572 38622 17578
rect 38558 17520 38564 17572
rect 38616 17569 38622 17572
rect 49003 17572 49067 17578
rect 49003 17569 49009 17572
rect 38616 17523 49009 17569
rect 38616 17520 38622 17523
rect 38558 17514 38622 17520
rect 49003 17520 49009 17523
rect 49061 17520 49067 17572
rect 49003 17514 49067 17520
rect 59257 17574 59331 17583
rect 59257 17518 59266 17574
rect 59322 17569 59331 17574
rect 59801 17572 59865 17578
rect 59801 17569 59807 17572
rect 59322 17523 59807 17569
rect 59322 17518 59331 17523
rect 59257 17509 59331 17518
rect 59801 17520 59807 17523
rect 59859 17520 59865 17572
rect 59801 17514 59865 17520
rect 60638 17572 60702 17578
rect 60638 17520 60644 17572
rect 60696 17569 60702 17572
rect 71083 17572 71147 17578
rect 71083 17569 71089 17572
rect 60696 17523 71089 17569
rect 60696 17520 60702 17523
rect 60638 17514 60702 17520
rect 71083 17520 71089 17523
rect 71141 17520 71147 17572
rect 71083 17514 71147 17520
rect 81337 17574 81411 17583
rect 81337 17518 81346 17574
rect 81402 17569 81411 17574
rect 81881 17572 81945 17578
rect 81881 17569 81887 17572
rect 81402 17523 81887 17569
rect 81402 17518 81411 17523
rect 81337 17509 81411 17518
rect 81881 17520 81887 17523
rect 81939 17520 81945 17572
rect 81881 17514 81945 17520
rect 82718 17572 82782 17578
rect 82718 17520 82724 17572
rect 82776 17569 82782 17572
rect 93163 17572 93227 17578
rect 93163 17569 93169 17572
rect 82776 17523 93169 17569
rect 82776 17520 82782 17523
rect 82718 17514 82782 17520
rect 93163 17520 93169 17523
rect 93221 17520 93227 17572
rect 93163 17514 93227 17520
rect 103417 17574 103491 17583
rect 103417 17518 103426 17574
rect 103482 17569 103491 17574
rect 103961 17572 104025 17578
rect 103961 17569 103967 17572
rect 103482 17523 103967 17569
rect 103482 17518 103491 17523
rect 103417 17509 103491 17518
rect 103961 17520 103967 17523
rect 104019 17520 104025 17572
rect 103961 17514 104025 17520
rect 104798 17572 104862 17578
rect 104798 17520 104804 17572
rect 104856 17569 104862 17572
rect 115243 17572 115307 17578
rect 115243 17569 115249 17572
rect 104856 17523 115249 17569
rect 104856 17520 104862 17523
rect 104798 17514 104862 17520
rect 115243 17520 115249 17523
rect 115301 17520 115307 17572
rect 115243 17514 115307 17520
rect 38335 17344 38399 17350
rect 38335 17341 38341 17344
rect 38227 17295 38341 17341
rect 38335 17292 38341 17295
rect 38393 17341 38399 17344
rect 48217 17346 48291 17355
rect 48217 17341 48226 17346
rect 38393 17295 48226 17341
rect 38393 17292 38399 17295
rect 38335 17286 38399 17292
rect 48217 17290 48226 17295
rect 48282 17290 48291 17346
rect 48217 17281 48291 17290
rect 60415 17344 60479 17350
rect 60415 17292 60421 17344
rect 60473 17341 60479 17344
rect 70297 17346 70371 17355
rect 70297 17341 70306 17346
rect 60473 17295 70306 17341
rect 60473 17292 60479 17295
rect 60415 17286 60479 17292
rect 70297 17290 70306 17295
rect 70362 17290 70371 17346
rect 70297 17281 70371 17290
rect 82495 17344 82559 17350
rect 82495 17292 82501 17344
rect 82553 17341 82559 17344
rect 92377 17346 92451 17355
rect 92377 17341 92386 17346
rect 82553 17295 92386 17341
rect 82553 17292 82559 17295
rect 82495 17286 82559 17292
rect 92377 17290 92386 17295
rect 92442 17290 92451 17346
rect 92377 17281 92451 17290
rect 104575 17344 104639 17350
rect 104575 17292 104581 17344
rect 104633 17341 104639 17344
rect 114457 17346 114531 17355
rect 114457 17341 114466 17346
rect 104633 17295 114466 17341
rect 104633 17292 104639 17295
rect 104575 17286 104639 17292
rect 114457 17290 114466 17295
rect 114522 17290 114531 17346
rect 114457 17281 114531 17290
rect 77674 16722 77748 16731
rect 77674 16666 77683 16722
rect 77739 16666 77748 16722
rect 77674 16657 77748 16666
rect 114831 16722 114905 16731
rect 114831 16666 114840 16722
rect 114896 16666 114905 16722
rect 114831 16657 114905 16666
rect 37177 15542 37251 15551
rect 37177 15486 37186 15542
rect 37242 15486 37251 15542
rect 37177 15477 37251 15486
rect 48217 15542 48291 15551
rect 48217 15486 48226 15542
rect 48282 15486 48291 15542
rect 48217 15477 48291 15486
rect 59257 15542 59331 15551
rect 59257 15486 59266 15542
rect 59322 15486 59331 15542
rect 59257 15477 59331 15486
rect 70297 15542 70371 15551
rect 70297 15486 70306 15542
rect 70362 15486 70371 15542
rect 70297 15477 70371 15486
rect 81337 15542 81411 15551
rect 81337 15486 81346 15542
rect 81402 15486 81411 15542
rect 81337 15477 81411 15486
rect 92377 15542 92451 15551
rect 92377 15486 92386 15542
rect 92442 15486 92451 15542
rect 92377 15477 92451 15486
rect 103417 15542 103491 15551
rect 103417 15486 103426 15542
rect 103482 15486 103491 15542
rect 103417 15477 103491 15486
rect 114457 15542 114531 15551
rect 114457 15486 114466 15542
rect 114522 15486 114531 15542
rect 114457 15477 114531 15486
rect 125180 14610 125244 14616
rect 125180 14558 125186 14610
rect 125238 14607 125244 14610
rect 136638 14612 136712 14621
rect 136638 14607 136647 14612
rect 125238 14561 136647 14607
rect 125238 14558 125244 14561
rect 125180 14552 125244 14558
rect 136638 14556 136647 14561
rect 136703 14556 136712 14612
rect 136638 14547 136712 14556
<< via2 >>
rect 48131 52261 48187 52317
rect 59171 52261 59227 52317
rect 70211 52261 70267 52317
rect 81251 52261 81307 52317
rect 92291 52261 92347 52317
rect 103331 52261 103387 52317
rect 114371 52261 114427 52317
rect 136647 49136 136703 49192
rect 59171 48464 59227 48520
rect 81251 48464 81307 48520
rect 103331 48464 103387 48520
rect 124841 48464 124897 48520
rect 48131 48206 48187 48262
rect 61014 48260 61070 48262
rect 61014 48208 61016 48260
rect 61016 48208 61068 48260
rect 61068 48208 61070 48260
rect 61014 48206 61070 48208
rect 70211 48206 70267 48262
rect 83094 48260 83150 48262
rect 83094 48208 83096 48260
rect 83096 48208 83148 48260
rect 83148 48208 83150 48260
rect 83094 48206 83150 48208
rect 92291 48206 92347 48262
rect 105174 48260 105230 48262
rect 105174 48208 105176 48260
rect 105176 48208 105228 48260
rect 105228 48208 105230 48260
rect 105174 48206 105230 48208
rect 114371 48206 114427 48262
rect 78596 47978 78652 48034
rect 115205 47978 115261 48034
rect 127254 47954 127310 47956
rect 127254 47902 127256 47954
rect 127256 47902 127308 47954
rect 127308 47902 127310 47954
rect 127254 47900 127310 47902
rect 136647 47806 136703 47862
rect 116386 47408 116442 47410
rect 116386 47356 116388 47408
rect 116388 47356 116440 47408
rect 116440 47356 116442 47408
rect 116386 47354 116442 47356
rect 136083 46538 136139 46594
rect 127964 45614 128020 45670
rect 136647 45662 136703 45664
rect 136647 45610 136649 45662
rect 136649 45610 136701 45662
rect 136701 45610 136703 45662
rect 136647 45608 136703 45610
rect 77965 44942 78021 44998
rect 136083 42974 136139 43030
rect 127964 42067 128020 42123
rect 136647 42098 136703 42100
rect 136647 42046 136649 42098
rect 136649 42046 136701 42098
rect 136701 42046 136703 42098
rect 136647 42044 136703 42046
rect 77965 41811 78021 41867
rect 136083 39410 136139 39466
rect 127964 38495 128020 38551
rect 136647 38534 136703 38536
rect 136647 38482 136649 38534
rect 136649 38482 136701 38534
rect 136701 38482 136703 38534
rect 136647 38480 136703 38482
rect 77965 38239 78021 38295
rect 136083 35846 136139 35902
rect 134753 35369 134809 35425
rect 135019 35369 135075 35425
rect 127964 34916 128020 34972
rect 136647 34970 136703 34972
rect 136647 34918 136649 34970
rect 136649 34918 136701 34970
rect 136701 34918 136703 34970
rect 136647 34916 136703 34918
rect 77965 34667 78021 34723
rect 134753 32445 134809 32501
rect 135019 32445 135075 32501
rect 136083 30167 136139 30223
rect 136647 29291 136703 29293
rect 136647 29239 136649 29291
rect 136649 29239 136701 29291
rect 136701 29239 136703 29291
rect 136647 29237 136703 29239
rect 127964 29079 128020 29135
rect 77965 27523 78021 27579
rect 136083 26603 136139 26659
rect 136647 25727 136703 25729
rect 136647 25675 136649 25727
rect 136649 25675 136701 25727
rect 136701 25675 136703 25727
rect 136647 25673 136703 25675
rect 127964 25506 128020 25562
rect 77965 23951 78021 24007
rect 136083 23039 136139 23095
rect 136647 22163 136703 22165
rect 136647 22111 136649 22163
rect 136649 22111 136701 22163
rect 136701 22111 136703 22163
rect 136647 22109 136703 22111
rect 127964 21933 128020 21989
rect 77965 20375 78021 20431
rect 136083 19475 136139 19531
rect 127964 18817 128020 18873
rect 77683 18647 77739 18649
rect 77683 18595 77685 18647
rect 77685 18595 77737 18647
rect 77737 18595 77739 18647
rect 77683 18593 77739 18595
rect 136647 18599 136703 18601
rect 136647 18547 136649 18599
rect 136649 18547 136701 18599
rect 136701 18547 136703 18599
rect 136647 18545 136703 18547
rect 115624 18502 115680 18504
rect 115624 18450 115626 18502
rect 115626 18450 115678 18502
rect 115678 18450 115680 18502
rect 115624 18448 115680 18450
rect 49974 17917 50030 17920
rect 49974 17865 49976 17917
rect 49976 17865 50028 17917
rect 50028 17865 50030 17917
rect 49974 17864 50030 17865
rect 72054 17917 72110 17919
rect 72054 17865 72056 17917
rect 72056 17865 72108 17917
rect 72108 17865 72110 17917
rect 72054 17863 72110 17865
rect 94134 17917 94190 17919
rect 94134 17865 94136 17917
rect 94136 17865 94188 17917
rect 94188 17865 94190 17917
rect 94134 17863 94190 17865
rect 116214 17917 116270 17919
rect 116214 17865 116216 17917
rect 116216 17865 116268 17917
rect 116268 17865 116270 17917
rect 116214 17863 116270 17865
rect 78596 17776 78652 17832
rect 115205 17776 115261 17832
rect 37186 17518 37242 17574
rect 59266 17518 59322 17574
rect 81346 17518 81402 17574
rect 103426 17518 103482 17574
rect 48226 17290 48282 17346
rect 70306 17290 70362 17346
rect 92386 17290 92442 17346
rect 114466 17290 114522 17346
rect 77683 16720 77739 16722
rect 77683 16668 77685 16720
rect 77685 16668 77737 16720
rect 77737 16668 77739 16720
rect 77683 16666 77739 16668
rect 114840 16720 114896 16722
rect 114840 16668 114842 16720
rect 114842 16668 114894 16720
rect 114894 16668 114896 16720
rect 114840 16666 114896 16668
rect 37186 15486 37242 15542
rect 48226 15486 48282 15542
rect 59266 15486 59322 15542
rect 70306 15486 70362 15542
rect 81346 15486 81402 15542
rect 92386 15486 92442 15542
rect 103426 15486 103482 15542
rect 114466 15486 114522 15542
rect 136647 14556 136703 14612
<< metal3 >>
rect 48126 52317 48192 52322
rect 48126 52261 48131 52317
rect 48187 52261 48192 52317
rect 48126 52256 48192 52261
rect 59166 52317 59232 52322
rect 59166 52261 59171 52317
rect 59227 52261 59232 52317
rect 59166 52256 59232 52261
rect 70206 52317 70272 52322
rect 70206 52261 70211 52317
rect 70267 52261 70272 52317
rect 70206 52256 70272 52261
rect 81246 52317 81312 52322
rect 81246 52261 81251 52317
rect 81307 52261 81312 52317
rect 81246 52256 81312 52261
rect 92286 52317 92352 52322
rect 92286 52261 92291 52317
rect 92347 52261 92352 52317
rect 92286 52256 92352 52261
rect 103326 52317 103392 52322
rect 103326 52261 103331 52317
rect 103387 52261 103392 52317
rect 103326 52256 103392 52261
rect 114366 52317 114432 52322
rect 114366 52261 114371 52317
rect 114427 52261 114432 52317
rect 114366 52256 114432 52261
rect 48129 48267 48189 52256
rect 59169 48525 59229 52256
rect 59166 48520 59232 48525
rect 59166 48464 59171 48520
rect 59227 48464 59232 48520
rect 59166 48459 59232 48464
rect 70209 48267 70269 52256
rect 81249 48525 81309 52256
rect 81246 48520 81312 48525
rect 81246 48464 81251 48520
rect 81307 48464 81312 48520
rect 81246 48459 81312 48464
rect 92289 48267 92349 52256
rect 103329 48525 103389 52256
rect 103326 48520 103392 48525
rect 103326 48464 103331 48520
rect 103387 48464 103392 48520
rect 103326 48459 103392 48464
rect 114369 48267 114429 52256
rect 48126 48262 48192 48267
rect 48126 48206 48131 48262
rect 48187 48206 48192 48262
rect 48126 48201 48192 48206
rect 61009 48262 61075 48267
rect 61009 48206 61014 48262
rect 61070 48206 61075 48262
rect 61009 48201 61075 48206
rect 70206 48262 70272 48267
rect 70206 48206 70211 48262
rect 70267 48206 70272 48262
rect 70206 48201 70272 48206
rect 83089 48262 83155 48267
rect 83089 48206 83094 48262
rect 83150 48206 83155 48262
rect 83089 48201 83155 48206
rect 92286 48262 92352 48267
rect 92286 48206 92291 48262
rect 92347 48206 92352 48262
rect 92286 48201 92352 48206
rect 105169 48262 105235 48267
rect 105169 48206 105174 48262
rect 105230 48206 105235 48262
rect 105169 48201 105235 48206
rect 114366 48262 114432 48267
rect 114366 48206 114371 48262
rect 114427 48206 114432 48262
rect 114366 48201 114432 48206
rect 48129 36806 48189 48201
rect 48121 36800 48197 36806
rect 48121 36736 48127 36800
rect 48191 36736 48197 36800
rect 48121 36730 48197 36736
rect 61012 36625 61072 48201
rect 70209 38575 70269 48201
rect 78591 48034 78657 48039
rect 78591 47978 78596 48034
rect 78652 47978 78657 48034
rect 78591 47973 78657 47978
rect 77960 44998 78026 45003
rect 77960 44942 77965 44998
rect 78021 44942 78026 44998
rect 77960 44937 78026 44942
rect 77963 41872 78023 41876
rect 77960 41867 78026 41872
rect 77960 41811 77965 41867
rect 78021 41811 78026 41867
rect 77960 41806 78026 41811
rect 77963 41802 78023 41806
rect 70201 38569 70277 38575
rect 70201 38505 70207 38569
rect 70271 38505 70277 38569
rect 70201 38499 70277 38505
rect 77963 38300 78023 38304
rect 77960 38295 78026 38300
rect 77960 38239 77965 38295
rect 78021 38239 78026 38295
rect 77960 38234 78026 38239
rect 77963 38230 78023 38234
rect 61004 36619 61080 36625
rect 61004 36555 61010 36619
rect 61074 36555 61080 36619
rect 61004 36549 61080 36555
rect 77963 34728 78023 34732
rect 77960 34723 78026 34728
rect 77960 34667 77965 34723
rect 78021 34667 78026 34723
rect 77960 34662 78026 34667
rect 77963 34658 78023 34662
rect 77963 27584 78023 27588
rect 77960 27579 78026 27584
rect 77960 27523 77965 27579
rect 78021 27523 78026 27579
rect 77960 27518 78026 27523
rect 77963 27514 78023 27518
rect 77963 24012 78023 24016
rect 77960 24007 78026 24012
rect 77960 23951 77965 24007
rect 78021 23951 78026 24007
rect 77960 23946 78026 23951
rect 77963 23942 78023 23946
rect 70296 22517 70372 22523
rect 70296 22453 70302 22517
rect 70366 22453 70372 22517
rect 70296 22447 70372 22453
rect 48216 18865 48292 18871
rect 48216 18801 48222 18865
rect 48286 18801 48292 18865
rect 48216 18795 48292 18801
rect 37181 17574 37247 17579
rect 37181 17518 37186 17574
rect 37242 17518 37247 17574
rect 37181 17513 37247 17518
rect 37184 15547 37244 17513
rect 48224 17351 48284 18795
rect 49964 18658 50040 18664
rect 49964 18594 49970 18658
rect 50034 18594 50040 18658
rect 49964 18588 50040 18594
rect 49972 17925 50032 18588
rect 49969 17920 50035 17925
rect 49969 17864 49974 17920
rect 50030 17864 50035 17920
rect 49969 17859 50035 17864
rect 59261 17574 59327 17579
rect 59261 17518 59266 17574
rect 59322 17518 59327 17574
rect 59261 17513 59327 17518
rect 48221 17346 48287 17351
rect 48221 17290 48226 17346
rect 48282 17290 48287 17346
rect 48221 17285 48287 17290
rect 48224 15547 48284 17285
rect 59264 15547 59324 17513
rect 70304 17351 70364 22447
rect 72044 22297 72120 22303
rect 72044 22233 72050 22297
rect 72114 22233 72120 22297
rect 72044 22227 72120 22233
rect 72052 17924 72112 22227
rect 77963 20436 78023 20440
rect 77960 20431 78026 20436
rect 77960 20375 77965 20431
rect 78021 20375 78026 20431
rect 77960 20370 78026 20375
rect 77963 20366 78023 20370
rect 77678 18649 77744 18654
rect 77678 18593 77683 18649
rect 77739 18593 77744 18649
rect 77678 18588 77744 18593
rect 72049 17919 72115 17924
rect 72049 17863 72054 17919
rect 72110 17863 72115 17919
rect 72049 17858 72115 17863
rect 70301 17346 70367 17351
rect 70301 17290 70306 17346
rect 70362 17290 70367 17346
rect 70301 17285 70367 17290
rect 70304 15547 70364 17285
rect 77681 16727 77741 18588
rect 78594 17837 78654 47973
rect 83092 38355 83152 48201
rect 92289 42148 92349 48201
rect 92281 42142 92357 42148
rect 92281 42078 92287 42142
rect 92351 42078 92357 42142
rect 92281 42072 92357 42078
rect 105172 41920 105232 48201
rect 114369 45716 114429 48201
rect 115200 48034 115266 48039
rect 115200 47978 115205 48034
rect 115261 47978 115266 48034
rect 115200 47973 115266 47978
rect 116384 47415 116444 49628
rect 116381 47410 116447 47415
rect 116381 47354 116386 47410
rect 116442 47354 116447 47410
rect 116381 47349 116447 47354
rect 114361 45710 114437 45716
rect 114361 45646 114367 45710
rect 114431 45646 114437 45710
rect 114361 45640 114437 45646
rect 105164 41914 105240 41920
rect 105164 41850 105170 41914
rect 105234 41850 105240 41914
rect 105164 41844 105240 41850
rect 83084 38349 83160 38355
rect 83084 38285 83090 38349
rect 83154 38285 83160 38349
rect 83084 38279 83160 38285
rect 103809 36800 103885 36806
rect 103809 36736 103815 36800
rect 103879 36736 103885 36800
rect 103809 36730 103885 36736
rect 103817 35000 103877 36730
rect 106094 36619 106170 36625
rect 106094 36555 106100 36619
rect 106164 36555 106170 36619
rect 106094 36549 106170 36555
rect 103809 34994 103885 35000
rect 103809 34930 103815 34994
rect 103879 34930 103885 34994
rect 103809 34924 103885 34930
rect 106102 34806 106162 36549
rect 106094 34800 106170 34806
rect 106094 34736 106100 34800
rect 106164 34736 106170 34800
rect 106094 34730 106170 34736
rect 118049 33118 118109 49365
rect 125329 49141 125389 51309
rect 136642 49192 136708 49197
rect 136642 49136 136647 49192
rect 136703 49136 136708 49192
rect 136642 49131 136708 49136
rect 124836 48520 124902 48525
rect 124836 48464 124841 48520
rect 124897 48464 124902 48520
rect 124836 48459 124902 48464
rect 127249 47956 127315 47961
rect 127249 47900 127254 47956
rect 127310 47900 127315 47956
rect 127249 47895 127315 47900
rect 127252 45579 127312 47895
rect 136645 47867 136705 49131
rect 136642 47862 136708 47867
rect 136642 47806 136647 47862
rect 136703 47806 136708 47862
rect 136642 47801 136708 47806
rect 136073 46594 136149 46604
rect 136073 46538 136083 46594
rect 136139 46538 136149 46594
rect 136073 46528 136149 46538
rect 127959 45670 128025 45675
rect 127959 45614 127964 45670
rect 128020 45614 128025 45670
rect 127959 45609 128025 45614
rect 127244 45573 127320 45579
rect 127244 45509 127250 45573
rect 127314 45509 127320 45573
rect 127244 45503 127320 45509
rect 134101 45573 134177 45579
rect 134101 45509 134107 45573
rect 134171 45509 134177 45573
rect 134101 45503 134177 45509
rect 127959 42123 128025 42128
rect 127959 42067 127964 42123
rect 128020 42067 128025 42123
rect 127959 42062 128025 42067
rect 134101 41914 134177 41920
rect 134101 41850 134107 41914
rect 134171 41850 134177 41914
rect 134101 41844 134177 41850
rect 127959 38551 128025 38556
rect 127959 38495 127964 38551
rect 128020 38495 128025 38551
rect 127959 38490 128025 38495
rect 134101 38349 134177 38355
rect 134101 38285 134107 38349
rect 134171 38285 134177 38349
rect 134101 38279 134177 38285
rect 135017 35430 135077 45925
rect 135158 45710 135234 45716
rect 135158 45646 135164 45710
rect 135228 45646 135234 45710
rect 135158 45640 135234 45646
rect 136081 43040 136141 46528
rect 136645 45669 136705 47801
rect 136642 45664 136708 45669
rect 136642 45608 136647 45664
rect 136703 45608 136708 45664
rect 136642 45603 136708 45608
rect 136073 43030 136149 43040
rect 136073 42974 136083 43030
rect 136139 42974 136149 43030
rect 136073 42964 136149 42974
rect 135158 42142 135234 42148
rect 135158 42078 135164 42142
rect 135228 42078 135234 42142
rect 135158 42072 135234 42078
rect 136081 39476 136141 42964
rect 136645 42105 136705 45603
rect 136642 42100 136708 42105
rect 136642 42044 136647 42100
rect 136703 42044 136708 42100
rect 136642 42039 136708 42044
rect 136073 39466 136149 39476
rect 136073 39410 136083 39466
rect 136139 39410 136149 39466
rect 136073 39400 136149 39410
rect 135158 38569 135234 38575
rect 135158 38505 135164 38569
rect 135228 38505 135234 38569
rect 135158 38499 135234 38505
rect 136081 35912 136141 39400
rect 136645 38541 136705 42039
rect 136642 38536 136708 38541
rect 136642 38480 136647 38536
rect 136703 38480 136708 38536
rect 136642 38475 136708 38480
rect 136073 35902 136149 35912
rect 136073 35846 136083 35902
rect 136139 35846 136149 35902
rect 136073 35836 136149 35846
rect 134748 35425 134814 35430
rect 134748 35369 134753 35425
rect 134809 35369 134814 35425
rect 134748 35364 134814 35369
rect 135014 35425 135080 35430
rect 135014 35369 135019 35425
rect 135075 35369 135080 35425
rect 135014 35364 135080 35369
rect 134751 35000 134811 35364
rect 134743 34994 134819 35000
rect 127959 34972 128025 34977
rect 127959 34916 127964 34972
rect 128020 34916 128025 34972
rect 134743 34930 134749 34994
rect 134813 34930 134819 34994
rect 134743 34924 134819 34930
rect 127959 34911 128025 34916
rect 134101 34800 134177 34806
rect 134101 34736 134107 34800
rect 134171 34736 134177 34800
rect 134101 34730 134177 34736
rect 134106 34721 134172 34730
rect 118041 33112 118117 33118
rect 118041 33048 118047 33112
rect 118111 33048 118117 33112
rect 118041 33042 118117 33048
rect 114456 29653 114532 29659
rect 114456 29589 114462 29653
rect 114526 29589 114532 29653
rect 114456 29583 114532 29589
rect 92376 26085 92452 26091
rect 92376 26021 92382 26085
rect 92446 26021 92452 26085
rect 92376 26015 92452 26021
rect 78591 17832 78657 17837
rect 78591 17776 78596 17832
rect 78652 17776 78657 17832
rect 78591 17771 78657 17776
rect 81341 17574 81407 17579
rect 81341 17518 81346 17574
rect 81402 17518 81407 17574
rect 81341 17513 81407 17518
rect 77678 16722 77744 16727
rect 77678 16666 77683 16722
rect 77739 16666 77744 16722
rect 77678 16661 77744 16666
rect 81344 15547 81404 17513
rect 92384 17351 92444 26015
rect 94124 25886 94200 25892
rect 94124 25822 94130 25886
rect 94194 25822 94200 25886
rect 94124 25816 94200 25822
rect 94132 17924 94192 25816
rect 94129 17919 94195 17924
rect 94129 17863 94134 17919
rect 94190 17863 94195 17919
rect 94129 17858 94195 17863
rect 103421 17574 103487 17579
rect 103421 17518 103426 17574
rect 103482 17518 103487 17574
rect 103421 17513 103487 17518
rect 92381 17346 92447 17351
rect 92381 17290 92386 17346
rect 92442 17290 92447 17346
rect 92381 17285 92447 17290
rect 92384 15547 92444 17285
rect 103424 15547 103484 17513
rect 114464 17351 114524 29583
rect 116204 29455 116280 29461
rect 116204 29391 116210 29455
rect 116274 29391 116280 29455
rect 116204 29385 116280 29391
rect 115619 18504 115685 18509
rect 115619 18448 115624 18504
rect 115680 18448 115685 18504
rect 115619 18443 115685 18448
rect 116212 17924 116272 29385
rect 116209 17919 116275 17924
rect 116209 17863 116214 17919
rect 116270 17863 116275 17919
rect 116209 17858 116275 17863
rect 115200 17832 115266 17837
rect 115200 17776 115205 17832
rect 115261 17776 115266 17832
rect 115200 17771 115266 17776
rect 114461 17346 114527 17351
rect 114461 17290 114466 17346
rect 114522 17290 114527 17346
rect 114461 17285 114527 17290
rect 114464 15547 114524 17285
rect 114835 16722 114901 16727
rect 114835 16666 114840 16722
rect 114896 16666 114901 16722
rect 114835 16661 114901 16666
rect 118049 16578 118109 33042
rect 134751 32506 134811 34924
rect 135017 33118 135077 35233
rect 135158 34994 135234 35000
rect 135158 34930 135164 34994
rect 135228 34930 135234 34994
rect 135158 34924 135234 34930
rect 135009 33112 135085 33118
rect 135009 33048 135015 33112
rect 135079 33048 135085 33112
rect 135009 33042 135085 33048
rect 134748 32501 134814 32506
rect 134748 32445 134753 32501
rect 134809 32445 134814 32501
rect 134748 32440 134814 32445
rect 135014 32501 135080 32506
rect 135014 32445 135019 32501
rect 135075 32445 135080 32501
rect 135014 32440 135080 32445
rect 134106 29461 134172 29490
rect 134101 29455 134177 29461
rect 134101 29391 134107 29455
rect 134171 29391 134177 29455
rect 134101 29385 134177 29391
rect 127959 29135 128025 29140
rect 127959 29079 127964 29135
rect 128020 29079 128025 29135
rect 127959 29042 128025 29079
rect 134106 25892 134172 25924
rect 134101 25886 134177 25892
rect 134101 25822 134107 25886
rect 134171 25822 134177 25886
rect 134101 25816 134177 25822
rect 127959 25562 128025 25567
rect 127959 25506 127964 25562
rect 128020 25506 128025 25562
rect 127959 25478 128025 25506
rect 134106 22303 134172 22364
rect 134101 22297 134177 22303
rect 134101 22233 134107 22297
rect 134171 22233 134177 22297
rect 134101 22227 134177 22233
rect 127959 21989 128025 21994
rect 127959 21933 127964 21989
rect 128020 21933 128025 21989
rect 127959 21914 128025 21933
rect 127959 18873 128025 18892
rect 127959 18817 127964 18873
rect 128020 18817 128025 18873
rect 127959 18812 128025 18817
rect 134101 18658 134177 18664
rect 134101 18594 134107 18658
rect 134171 18594 134177 18658
rect 134101 18588 134177 18594
rect 135017 17402 135077 32440
rect 136081 30233 136141 35836
rect 136645 34977 136705 38475
rect 136642 34972 136708 34977
rect 136642 34916 136647 34972
rect 136703 34916 136708 34972
rect 136642 34911 136708 34916
rect 136518 31014 136578 33195
rect 136073 30223 136149 30233
rect 136073 30167 136083 30223
rect 136139 30167 136149 30223
rect 136073 30157 136149 30167
rect 135158 29653 135234 29659
rect 135158 29589 135164 29653
rect 135228 29589 135234 29653
rect 135158 29583 135234 29589
rect 136081 26669 136141 30157
rect 136645 29298 136705 34911
rect 136642 29293 136708 29298
rect 136642 29237 136647 29293
rect 136703 29237 136708 29293
rect 136642 29232 136708 29237
rect 136073 26663 136149 26669
rect 136073 26599 136079 26663
rect 136143 26599 136149 26663
rect 136073 26593 136149 26599
rect 135158 26085 135234 26091
rect 135158 26021 135164 26085
rect 135228 26021 135234 26085
rect 135158 26015 135234 26021
rect 136081 23105 136141 26593
rect 136645 25734 136705 29232
rect 136642 25729 136708 25734
rect 136642 25673 136647 25729
rect 136703 25673 136708 25729
rect 136642 25668 136708 25673
rect 136073 23095 136149 23105
rect 136073 23039 136083 23095
rect 136139 23039 136149 23095
rect 136073 23029 136149 23039
rect 135158 22517 135234 22523
rect 135158 22453 135164 22517
rect 135228 22453 135234 22517
rect 135158 22447 135234 22453
rect 136081 19541 136141 23029
rect 136645 22170 136705 25668
rect 136642 22165 136708 22170
rect 136642 22109 136647 22165
rect 136703 22109 136708 22165
rect 136642 22104 136708 22109
rect 136073 19531 136149 19541
rect 136073 19475 136083 19531
rect 136139 19475 136149 19531
rect 136073 19465 136149 19475
rect 135158 18865 135234 18871
rect 135158 18801 135164 18865
rect 135228 18801 135234 18865
rect 135158 18795 135234 18801
rect 136518 16824 136578 20327
rect 136645 18606 136705 22104
rect 136642 18601 136708 18606
rect 136642 18545 136647 18601
rect 136703 18545 136708 18601
rect 136642 18540 136708 18545
rect 136515 16758 136581 16824
rect 37181 15542 37247 15547
rect 37181 15486 37186 15542
rect 37242 15486 37247 15542
rect 37181 15481 37247 15486
rect 48221 15542 48287 15547
rect 48221 15486 48226 15542
rect 48282 15486 48287 15542
rect 48221 15481 48287 15486
rect 59261 15542 59327 15547
rect 59261 15486 59266 15542
rect 59322 15486 59327 15542
rect 59261 15481 59327 15486
rect 70301 15542 70367 15547
rect 70301 15486 70306 15542
rect 70362 15486 70367 15542
rect 70301 15481 70367 15486
rect 81341 15542 81407 15547
rect 81341 15486 81346 15542
rect 81402 15486 81407 15542
rect 81341 15481 81407 15486
rect 92381 15542 92447 15547
rect 92381 15486 92386 15542
rect 92442 15486 92447 15542
rect 92381 15481 92447 15486
rect 103421 15542 103487 15547
rect 103421 15486 103426 15542
rect 103482 15486 103487 15542
rect 103421 15481 103487 15486
rect 114461 15542 114527 15547
rect 114461 15486 114466 15542
rect 114522 15486 114527 15542
rect 114461 15481 114527 15486
rect 125276 12835 125336 16338
rect 136645 14617 136705 18540
rect 136642 14612 136708 14617
rect 136642 14556 136647 14612
rect 136703 14556 136708 14612
rect 136642 14551 136708 14556
rect 125273 12830 125339 12835
rect 125273 12769 125276 12830
rect 125336 12769 125339 12830
<< via3 >>
rect 48127 36736 48191 36800
rect 70207 38505 70271 38569
rect 61010 36555 61074 36619
rect 70302 22453 70366 22517
rect 48222 18801 48286 18865
rect 49970 18594 50034 18658
rect 72050 22233 72114 22297
rect 92287 42078 92351 42142
rect 114367 45646 114431 45710
rect 105170 41850 105234 41914
rect 83090 38285 83154 38349
rect 103815 36736 103879 36800
rect 106100 36555 106164 36619
rect 103815 34930 103879 34994
rect 106100 34736 106164 34800
rect 127250 45509 127314 45573
rect 134107 45509 134171 45573
rect 134107 41850 134171 41914
rect 134107 38285 134171 38349
rect 135164 45646 135228 45710
rect 135164 42078 135228 42142
rect 135164 38505 135228 38569
rect 134749 34930 134813 34994
rect 134107 34736 134171 34800
rect 118047 33048 118111 33112
rect 114462 29589 114526 29653
rect 92382 26021 92446 26085
rect 94130 25822 94194 25886
rect 116210 29391 116274 29455
rect 135164 34930 135228 34994
rect 135015 33048 135079 33112
rect 134107 29391 134171 29455
rect 134107 25822 134171 25886
rect 134107 22233 134171 22297
rect 134107 18594 134171 18658
rect 135164 29589 135228 29653
rect 136079 26659 136143 26663
rect 136079 26603 136083 26659
rect 136083 26603 136139 26659
rect 136139 26603 136143 26659
rect 136079 26599 136143 26603
rect 135164 26021 135228 26085
rect 135164 22453 135228 22517
rect 135164 18801 135228 18865
<< metal4 >>
rect 114366 45710 114432 45711
rect 114366 45646 114367 45710
rect 114431 45708 114432 45710
rect 135163 45710 135229 45711
rect 135163 45708 135164 45710
rect 114431 45648 135164 45708
rect 114431 45646 114432 45648
rect 114366 45645 114432 45646
rect 135163 45646 135164 45648
rect 135228 45646 135229 45710
rect 135163 45645 135229 45646
rect 127249 45573 127315 45574
rect 127249 45509 127250 45573
rect 127314 45571 127315 45573
rect 134106 45573 134172 45574
rect 134106 45571 134107 45573
rect 127314 45511 134107 45571
rect 127314 45509 127315 45511
rect 127249 45508 127315 45509
rect 134106 45509 134107 45511
rect 134171 45509 134172 45573
rect 134106 45508 134172 45509
rect 92286 42142 92352 42143
rect 92286 42078 92287 42142
rect 92351 42140 92352 42142
rect 135163 42142 135229 42143
rect 135163 42140 135164 42142
rect 92351 42080 135164 42140
rect 92351 42078 92352 42080
rect 92286 42077 92352 42078
rect 135163 42078 135164 42080
rect 135228 42078 135229 42142
rect 135163 42077 135229 42078
rect 105169 41914 105235 41915
rect 105169 41850 105170 41914
rect 105234 41912 105235 41914
rect 134106 41914 134172 41915
rect 134106 41912 134107 41914
rect 105234 41852 134107 41912
rect 105234 41850 105235 41852
rect 105169 41849 105235 41850
rect 134106 41850 134107 41852
rect 134171 41850 134172 41914
rect 134106 41849 134172 41850
rect 70206 38569 70272 38570
rect 70206 38505 70207 38569
rect 70271 38567 70272 38569
rect 135163 38569 135229 38570
rect 135163 38567 135164 38569
rect 70271 38507 135164 38567
rect 70271 38505 70272 38507
rect 70206 38504 70272 38505
rect 135163 38505 135164 38507
rect 135228 38505 135229 38569
rect 135163 38504 135229 38505
rect 83089 38349 83155 38350
rect 83089 38285 83090 38349
rect 83154 38347 83155 38349
rect 134106 38349 134172 38350
rect 134106 38347 134107 38349
rect 83154 38287 134107 38347
rect 83154 38285 83155 38287
rect 83089 38284 83155 38285
rect 134106 38285 134107 38287
rect 134171 38285 134172 38349
rect 134106 38284 134172 38285
rect 48126 36800 48192 36801
rect 48126 36736 48127 36800
rect 48191 36798 48192 36800
rect 103814 36800 103880 36801
rect 103814 36798 103815 36800
rect 48191 36738 103815 36798
rect 48191 36736 48192 36738
rect 48126 36735 48192 36736
rect 103814 36736 103815 36738
rect 103879 36736 103880 36800
rect 103814 36735 103880 36736
rect 61009 36619 61075 36620
rect 61009 36555 61010 36619
rect 61074 36617 61075 36619
rect 106099 36619 106165 36620
rect 106099 36617 106100 36619
rect 61074 36557 106100 36617
rect 61074 36555 61075 36557
rect 61009 36554 61075 36555
rect 106099 36555 106100 36557
rect 106164 36555 106165 36619
rect 106099 36554 106165 36555
rect 103814 34994 103880 34995
rect 103814 34930 103815 34994
rect 103879 34992 103880 34994
rect 134748 34994 134814 34995
rect 134748 34992 134749 34994
rect 103879 34932 134749 34992
rect 103879 34930 103880 34932
rect 103814 34929 103880 34930
rect 134748 34930 134749 34932
rect 134813 34992 134814 34994
rect 135163 34994 135229 34995
rect 135163 34992 135164 34994
rect 134813 34932 135164 34992
rect 134813 34930 134814 34932
rect 134748 34929 134814 34930
rect 135163 34930 135164 34932
rect 135228 34930 135229 34994
rect 135163 34929 135229 34930
rect 106099 34800 106165 34801
rect 106099 34736 106100 34800
rect 106164 34798 106165 34800
rect 134106 34800 134172 34801
rect 134106 34798 134107 34800
rect 106164 34738 134107 34798
rect 106164 34736 106165 34738
rect 106099 34735 106165 34736
rect 134106 34736 134107 34738
rect 134171 34736 134172 34800
rect 134106 34735 134172 34736
rect 118046 33112 118112 33113
rect 118046 33048 118047 33112
rect 118111 33110 118112 33112
rect 135014 33112 135080 33113
rect 135014 33110 135015 33112
rect 118111 33050 135015 33110
rect 118111 33048 118112 33050
rect 118046 33047 118112 33048
rect 135014 33048 135015 33050
rect 135079 33048 135080 33112
rect 135014 33047 135080 33048
rect 114461 29653 114527 29654
rect 114461 29589 114462 29653
rect 114526 29651 114527 29653
rect 135163 29653 135229 29654
rect 135163 29651 135164 29653
rect 114526 29591 135164 29651
rect 114526 29589 114527 29591
rect 114461 29588 114527 29589
rect 135163 29589 135164 29591
rect 135228 29589 135229 29653
rect 135163 29588 135229 29589
rect 116209 29455 116275 29456
rect 116209 29391 116210 29455
rect 116274 29453 116275 29455
rect 134106 29455 134172 29456
rect 134106 29453 134107 29455
rect 116274 29393 134107 29453
rect 116274 29391 116275 29393
rect 116209 29390 116275 29391
rect 134106 29391 134107 29393
rect 134171 29391 134172 29455
rect 134106 29390 134172 29391
rect 136078 26663 136144 26664
rect 136078 26599 136079 26663
rect 136143 26661 136144 26663
rect 136143 26601 138515 26661
rect 136143 26599 136144 26601
rect 136078 26598 136144 26599
rect 92381 26085 92447 26086
rect 92381 26021 92382 26085
rect 92446 26083 92447 26085
rect 135163 26085 135229 26086
rect 135163 26083 135164 26085
rect 92446 26023 135164 26083
rect 92446 26021 92447 26023
rect 92381 26020 92447 26021
rect 135163 26021 135164 26023
rect 135228 26021 135229 26085
rect 135163 26020 135229 26021
rect 94129 25886 94195 25887
rect 94129 25822 94130 25886
rect 94194 25884 94195 25886
rect 134106 25886 134172 25887
rect 134106 25884 134107 25886
rect 94194 25824 134107 25884
rect 94194 25822 94195 25824
rect 94129 25821 94195 25822
rect 134106 25822 134107 25824
rect 134171 25822 134172 25886
rect 134106 25821 134172 25822
rect 70301 22517 70367 22518
rect 70301 22453 70302 22517
rect 70366 22515 70367 22517
rect 135163 22517 135229 22518
rect 135163 22515 135164 22517
rect 70366 22455 135164 22515
rect 70366 22453 70367 22455
rect 70301 22452 70367 22453
rect 135163 22453 135164 22455
rect 135228 22453 135229 22517
rect 135163 22452 135229 22453
rect 72049 22297 72115 22298
rect 72049 22233 72050 22297
rect 72114 22295 72115 22297
rect 134106 22297 134172 22298
rect 134106 22295 134107 22297
rect 72114 22235 134107 22295
rect 72114 22233 72115 22235
rect 72049 22232 72115 22233
rect 134106 22233 134107 22235
rect 134171 22233 134172 22297
rect 134106 22232 134172 22233
rect 48221 18865 48287 18866
rect 48221 18801 48222 18865
rect 48286 18863 48287 18865
rect 135163 18865 135229 18866
rect 135163 18863 135164 18865
rect 48286 18803 135164 18863
rect 48286 18801 48287 18803
rect 48221 18800 48287 18801
rect 135163 18801 135164 18803
rect 135228 18801 135229 18865
rect 135163 18800 135229 18801
rect 49969 18658 50035 18659
rect 49969 18594 49970 18658
rect 50034 18656 50035 18658
rect 134106 18658 134172 18659
rect 134106 18656 134107 18658
rect 50034 18596 134107 18656
rect 50034 18594 50035 18596
rect 49969 18593 50035 18594
rect 134106 18594 134107 18596
rect 134171 18594 134172 18658
rect 134106 18593 134172 18594
rect 111889 14554 115201 14614
<< via4 >>
rect 138515 26513 138751 26749
<< metal5 >>
rect 121416 32899 140449 33249
rect 140129 31492 140449 32899
rect 140129 31172 140432 31492
rect 139531 26870 139851 27190
use And_Gate  And_Gate_0
timestamp 1756481424
transform 1 0 71687 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_1
timestamp 1756481424
transform 1 0 49607 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_2
timestamp 1756481424
transform 1 0 93767 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_3
timestamp 1756481424
transform 1 0 115847 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_4
timestamp 1756481424
transform 1 0 82727 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_5
timestamp 1756481424
transform 1 0 60647 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_6
timestamp 1756481424
transform 1 0 104807 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_7
timestamp 1756481424
transform 1 0 126887 0 1 47569
box -1558 -210 544 1618
use CDAC8  CDAC8_0
timestamp 1756481424
transform 1 0 68478 0 1 21136
box -39092 -2552 55448 26024
use Comparator  Comparator_0
timestamp 1756559655
transform -1 0 168226 0 1 18611
box 24473 -2307 30902 29735
use D_FlipFlop  D_FlipFlop_0
timestamp 1757042133
transform -1 0 136483 0 1 45613
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_1
timestamp 1757042133
transform -1 0 136483 0 1 34921
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1757042133
transform -1 0 136483 0 1 38485
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1757042133
transform -1 0 136483 0 1 42049
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1757042133
transform -1 0 136483 0 1 29242
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1757042133
transform -1 0 136483 0 1 25678
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1757042133
transform -1 0 136483 0 1 22114
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1757042133
transform -1 0 136483 0 1 18550
box -102 -1796 8762 1842
use Nand_Gate  Nand_Gate_0
timestamp 1756481424
transform 1 0 68595 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_1
timestamp 1756481424
transform 1 0 101715 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_2
timestamp 1756481424
transform 1 0 90675 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_3
timestamp 1756481424
transform 1 0 46515 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_4
timestamp 1756481424
transform 1 0 35475 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_5
timestamp 1756481424
transform 1 0 112755 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_6
timestamp 1756481424
transform 1 0 79635 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_7
timestamp 1756481424
transform 1 0 57555 0 1 17201
box 1906 -530 3264 1298
use RingCounter  RingCounter_0
timestamp 1757042133
transform 1 0 28071 0 1 12779
box 88 -14 97272 40399
<< labels >>
flabel metal3 135017 17402 135077 32496 0 FreeSans 160 90 0 0 FFCLR
flabel metal1 127721 38485 136483 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 38485 135739 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 38485 136483 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 38485 133767 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 38485 131795 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 38485 131051 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 38485 129693 38531 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 42049 136483 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 42049 135739 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 42049 136483 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 42049 133767 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 42049 131795 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 42049 131051 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 42049 129693 42095 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 45613 136483 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 45613 135739 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 45613 136483 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 45613 133767 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 45613 131795 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 45613 131051 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 45613 129693 45659 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 25678 136483 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 25678 135739 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 25678 136483 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 25678 133767 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 25678 131795 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 25678 131051 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 25678 129693 25724 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 22114 136483 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 22114 135739 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 22114 136483 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 22114 133767 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 22114 131795 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 22114 131051 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 22114 129693 22160 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 18550 136483 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 133767 18550 135739 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 135739 18550 136483 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131795 18550 133767 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 131051 18550 131795 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 129693 18550 131051 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal1 127721 18550 129693 18596 0 FreeSans 160 180 0 0 VDD
port 12 nsew
flabel metal4 111889 14554 115201 14614 0 FreeSans 160 0 0 0 CLK
port 0 nsew
flabel metal2 77296 18824 127964 18870 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal2 77296 21936 127964 21982 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal2 77296 25511 127964 25557 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal2 77296 29084 127964 29130 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal2 77295 45619 127963 45665 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal3 118049 16578 118109 49365 0 FreeSans 160 0 0 0 EN
port 14 nsew
flabel metal2 77296 38500 127964 38546 0 FreeSans 160 0 0 0 Q6
port 8 nsew
flabel metal2 77296 42072 127964 42118 0 FreeSans 160 0 0 0 Q5
port 9 nsew
flabel metal2 77296 45619 127964 45665 0 FreeSans 160 0 0 0 Q4
port 15 nsew
flabel metal2 77296 34928 127964 34974 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal3 125276 12830 125336 16338 0 FreeSans 160 90 0 0 GND
port 16 nsew
flabel metal1 140592 16601 140991 16647 0 FreeSans 160 0 0 0 Vbias
port 17 nsew
flabel metal5 139531 26870 139851 27190 0 FreeSans 1600 0 0 0 Vin
port 18 nsew
<< end >>
