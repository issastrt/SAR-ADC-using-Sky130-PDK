magic
tech sky130A
magscale 1 2
timestamp 1755588857
<< nwell >>
rect 7192 -763 9164 -702
<< pwell >>
rect 7841 -1859 7901 -1852
<< metal1 >>
rect 7984 25642 8048 25648
rect 7984 25639 7990 25642
rect 7100 23857 7146 25639
rect 7192 25593 7990 25639
rect 7984 25590 7990 25593
rect 8042 25639 8048 25642
rect 8042 25593 9256 25639
rect 8042 25590 8048 25593
rect 7984 25584 8048 25590
rect 8155 24741 8815 24787
rect 7839 24463 7903 24469
rect 7839 24411 7845 24463
rect 7897 24411 7903 24463
rect 7839 24405 7903 24411
rect 7694 23860 7758 23866
rect 7694 23857 7700 23860
rect 7100 23811 7700 23857
rect 7100 20726 7146 23811
rect 7694 23808 7700 23811
rect 7752 23857 7758 23860
rect 7752 23811 9164 23857
rect 7752 23808 7758 23811
rect 7694 23802 7758 23808
rect 7984 22511 8048 22517
rect 7984 22508 7990 22511
rect 7192 22462 7990 22508
rect 7984 22459 7990 22462
rect 8042 22508 8048 22511
rect 9210 22508 9256 25593
rect 8042 22462 9256 22508
rect 8042 22459 8048 22462
rect 7984 22453 8048 22459
rect 8155 21610 8815 21656
rect 7837 21328 7901 21334
rect 7837 21276 7843 21328
rect 7895 21276 7901 21328
rect 7837 21270 7901 21276
rect 7694 20729 7758 20735
rect 7694 20726 7700 20729
rect 7100 20680 7700 20726
rect 7100 17154 7146 20680
rect 7694 20677 7700 20680
rect 7752 20726 7758 20729
rect 7752 20680 9164 20726
rect 7752 20677 7758 20680
rect 7694 20671 7758 20677
rect 7984 18939 8048 18945
rect 7984 18936 7990 18939
rect 7192 18890 7990 18936
rect 7984 18887 7990 18890
rect 8042 18936 8048 18939
rect 9210 18936 9256 22462
rect 8042 18890 9256 18936
rect 8042 18887 8048 18890
rect 7984 18881 8048 18887
rect 8155 18038 8815 18084
rect 7839 17756 7903 17762
rect 7839 17704 7845 17756
rect 7897 17704 7903 17756
rect 7839 17698 7903 17704
rect 7694 17157 7758 17163
rect 7694 17154 7700 17157
rect 7100 17108 7700 17154
rect 7100 13582 7146 17108
rect 7694 17105 7700 17108
rect 7752 17154 7758 17157
rect 7752 17108 9164 17154
rect 7752 17105 7758 17108
rect 7694 17099 7758 17105
rect 7984 15367 8048 15373
rect 7984 15364 7990 15367
rect 7192 15318 7990 15364
rect 7984 15315 7990 15318
rect 8042 15364 8048 15367
rect 9210 15364 9256 18890
rect 8042 15318 9256 15364
rect 8042 15315 8048 15318
rect 7984 15309 8048 15315
rect 8155 14466 8815 14512
rect 7839 14176 7903 14182
rect 7839 14124 7845 14176
rect 7897 14124 7903 14176
rect 7839 14118 7903 14124
rect 7694 13585 7758 13591
rect 7694 13582 7700 13585
rect 7100 13536 7700 13582
rect 7100 6438 7146 13536
rect 7694 13533 7700 13536
rect 7752 13582 7758 13585
rect 7752 13536 9164 13582
rect 7752 13533 7758 13536
rect 7694 13527 7758 13533
rect 7984 8223 8048 8229
rect 7984 8220 7990 8223
rect 7192 8174 7990 8220
rect 7984 8171 7990 8174
rect 8042 8220 8048 8223
rect 9210 8220 9256 15318
rect 8042 8174 9256 8220
rect 8042 8171 8048 8174
rect 7984 8165 8048 8171
rect 8155 7322 8815 7368
rect 7839 7032 7903 7038
rect 7839 6980 7845 7032
rect 7897 6980 7903 7032
rect 7839 6974 7903 6980
rect 7694 6441 7758 6447
rect 7694 6438 7700 6441
rect 7100 6392 7700 6438
rect 7100 2866 7146 6392
rect 7694 6389 7700 6392
rect 7752 6438 7758 6441
rect 7752 6392 9164 6438
rect 7752 6389 7758 6392
rect 7694 6383 7758 6389
rect 7984 4651 8048 4657
rect 7984 4648 7990 4651
rect 7192 4602 7990 4648
rect 7984 4599 7990 4602
rect 8042 4648 8048 4651
rect 9210 4648 9256 8174
rect 8042 4602 9256 4648
rect 8042 4599 8048 4602
rect 7984 4593 8048 4599
rect 8155 3750 8815 3796
rect 7839 3460 7903 3466
rect 7839 3408 7845 3460
rect 7897 3408 7903 3460
rect 7839 3402 7903 3408
rect 7694 2869 7758 2876
rect 7694 2866 7700 2869
rect 7100 2820 7700 2866
rect 7100 -710 7146 2820
rect 7694 2817 7700 2820
rect 7752 2866 7758 2869
rect 7752 2820 9164 2866
rect 7752 2817 7758 2820
rect 7694 2811 7758 2817
rect 7984 1075 8048 1081
rect 7984 1072 7990 1075
rect 7192 1026 7990 1072
rect 7984 1023 7990 1026
rect 8042 1072 8048 1075
rect 9210 1072 9256 4602
rect 8042 1026 9256 1072
rect 8042 1023 8048 1026
rect 7984 1017 8048 1023
rect 8155 174 8815 220
rect 7839 -112 7903 -106
rect 7839 -164 7845 -112
rect 7897 -164 7903 -112
rect 7839 -170 7903 -164
rect 7694 -707 7758 -701
rect 7694 -710 7700 -707
rect 7100 -756 7700 -710
rect 7100 -2538 7146 -756
rect 7694 -759 7700 -756
rect 7752 -710 7758 -707
rect 7752 -756 9164 -710
rect 7752 -759 7758 -756
rect 7694 -765 7758 -759
rect 8155 -1686 8815 -1640
rect 7839 -1822 7903 -1816
rect 7839 -1874 7845 -1822
rect 7897 -1874 7903 -1822
rect 7839 -1880 7903 -1874
rect 7984 -2489 8048 -2483
rect 7984 -2492 7990 -2489
rect 7192 -2538 7990 -2492
rect 7984 -2541 7990 -2538
rect 8042 -2492 8048 -2489
rect 9210 -2492 9256 1026
rect 8042 -2538 9256 -2492
rect 8042 -2541 8048 -2538
rect 7984 -2547 8048 -2541
<< via1 >>
rect 7990 25590 8042 25642
rect 7845 24411 7897 24463
rect 7700 23808 7752 23860
rect 7990 22459 8042 22511
rect 7843 21276 7895 21328
rect 7700 20677 7752 20729
rect 7990 18887 8042 18939
rect 7845 17704 7897 17756
rect 7700 17105 7752 17157
rect 7990 15315 8042 15367
rect 7845 14124 7897 14176
rect 7700 13533 7752 13585
rect 7990 8171 8042 8223
rect 7845 6980 7897 7032
rect 7700 6389 7752 6441
rect 7990 4599 8042 4651
rect 7845 3408 7897 3460
rect 7700 2817 7752 2869
rect 7990 1023 8042 1075
rect 7845 -164 7897 -112
rect 7700 -759 7752 -707
rect 7845 -1874 7897 -1822
rect 7990 -2541 8042 -2489
<< metal2 >>
rect 7979 25644 8053 25653
rect 7979 25588 7988 25644
rect 8044 25588 8053 25644
rect 7979 25579 8053 25588
rect 7834 24465 7908 24474
rect 7834 24409 7843 24465
rect 7899 24409 7908 24465
rect 7834 24400 7908 24409
rect 7689 23862 7763 23871
rect 7689 23806 7698 23862
rect 7754 23806 7763 23862
rect 7689 23797 7763 23806
rect 7979 22513 8053 22522
rect 7979 22457 7988 22513
rect 8044 22457 8053 22513
rect 7979 22448 8053 22457
rect 7832 21330 7906 21339
rect 7832 21274 7841 21330
rect 7897 21274 7906 21330
rect 7832 21265 7906 21274
rect 7689 20731 7763 20740
rect 7689 20675 7698 20731
rect 7754 20675 7763 20731
rect 7689 20666 7763 20675
rect 7979 18941 8053 18950
rect 7979 18885 7988 18941
rect 8044 18885 8053 18941
rect 7979 18876 8053 18885
rect 7834 17758 7908 17767
rect 7834 17702 7843 17758
rect 7899 17702 7908 17758
rect 7834 17693 7908 17702
rect 7689 17159 7763 17168
rect 7689 17103 7698 17159
rect 7754 17103 7763 17159
rect 7689 17094 7763 17103
rect 7979 15369 8053 15378
rect 7979 15313 7988 15369
rect 8044 15313 8053 15369
rect 7979 15304 8053 15313
rect 7834 14178 7908 14187
rect 7834 14122 7843 14178
rect 7899 14122 7908 14178
rect 7834 14113 7908 14122
rect 7689 13587 7763 13596
rect 7689 13531 7698 13587
rect 7754 13531 7763 13587
rect 7689 13522 7763 13531
rect 7979 8225 8053 8234
rect 7979 8169 7988 8225
rect 8044 8169 8053 8225
rect 7979 8160 8053 8169
rect 7834 7034 7908 7043
rect 7834 6978 7843 7034
rect 7899 6978 7908 7034
rect 7834 6969 7908 6978
rect 7689 6443 7763 6452
rect 7689 6387 7698 6443
rect 7754 6387 7763 6443
rect 7689 6378 7763 6387
rect 7979 4653 8053 4662
rect 7979 4597 7988 4653
rect 8044 4597 8053 4653
rect 7979 4588 8053 4597
rect 7834 3462 7908 3471
rect 7834 3406 7843 3462
rect 7899 3406 7908 3462
rect 7834 3397 7908 3406
rect 7689 2871 7763 2880
rect 7689 2815 7698 2871
rect 7754 2815 7763 2871
rect 7689 2806 7763 2815
rect 7979 1077 8053 1086
rect 7979 1021 7988 1077
rect 8044 1021 8053 1077
rect 7979 1012 8053 1021
rect 7834 -110 7908 -101
rect 7834 -166 7843 -110
rect 7899 -166 7908 -110
rect 7834 -175 7908 -166
rect 7689 -705 7763 -696
rect 7689 -761 7698 -705
rect 7754 -761 7763 -705
rect 7689 -770 7763 -761
rect 7834 -1820 7908 -1811
rect 7834 -1876 7843 -1820
rect 7899 -1876 7908 -1820
rect 7834 -1885 7908 -1876
rect 7979 -2487 8053 -2478
rect 7979 -2543 7988 -2487
rect 8044 -2543 8053 -2487
rect 7979 -2552 8053 -2543
<< via2 >>
rect 7988 25642 8044 25644
rect 7988 25590 7990 25642
rect 7990 25590 8042 25642
rect 8042 25590 8044 25642
rect 7988 25588 8044 25590
rect 7843 24463 7899 24465
rect 7843 24411 7845 24463
rect 7845 24411 7897 24463
rect 7897 24411 7899 24463
rect 7843 24409 7899 24411
rect 7698 23860 7754 23862
rect 7698 23808 7700 23860
rect 7700 23808 7752 23860
rect 7752 23808 7754 23860
rect 7698 23806 7754 23808
rect 7988 22511 8044 22513
rect 7988 22459 7990 22511
rect 7990 22459 8042 22511
rect 8042 22459 8044 22511
rect 7988 22457 8044 22459
rect 7841 21328 7897 21330
rect 7841 21276 7843 21328
rect 7843 21276 7895 21328
rect 7895 21276 7897 21328
rect 7841 21274 7897 21276
rect 7698 20729 7754 20731
rect 7698 20677 7700 20729
rect 7700 20677 7752 20729
rect 7752 20677 7754 20729
rect 7698 20675 7754 20677
rect 7988 18939 8044 18941
rect 7988 18887 7990 18939
rect 7990 18887 8042 18939
rect 8042 18887 8044 18939
rect 7988 18885 8044 18887
rect 7843 17756 7899 17758
rect 7843 17704 7845 17756
rect 7845 17704 7897 17756
rect 7897 17704 7899 17756
rect 7843 17702 7899 17704
rect 7698 17157 7754 17159
rect 7698 17105 7700 17157
rect 7700 17105 7752 17157
rect 7752 17105 7754 17157
rect 7698 17103 7754 17105
rect 7988 15367 8044 15369
rect 7988 15315 7990 15367
rect 7990 15315 8042 15367
rect 8042 15315 8044 15367
rect 7988 15313 8044 15315
rect 7843 14176 7899 14178
rect 7843 14124 7845 14176
rect 7845 14124 7897 14176
rect 7897 14124 7899 14176
rect 7843 14122 7899 14124
rect 7698 13585 7754 13587
rect 7698 13533 7700 13585
rect 7700 13533 7752 13585
rect 7752 13533 7754 13585
rect 7698 13531 7754 13533
rect 7988 8223 8044 8225
rect 7988 8171 7990 8223
rect 7990 8171 8042 8223
rect 8042 8171 8044 8223
rect 7988 8169 8044 8171
rect 7843 7032 7899 7034
rect 7843 6980 7845 7032
rect 7845 6980 7897 7032
rect 7897 6980 7899 7032
rect 7843 6978 7899 6980
rect 7698 6441 7754 6443
rect 7698 6389 7700 6441
rect 7700 6389 7752 6441
rect 7752 6389 7754 6441
rect 7698 6387 7754 6389
rect 7988 4651 8044 4653
rect 7988 4599 7990 4651
rect 7990 4599 8042 4651
rect 8042 4599 8044 4651
rect 7988 4597 8044 4599
rect 7843 3460 7899 3462
rect 7843 3408 7845 3460
rect 7845 3408 7897 3460
rect 7897 3408 7899 3460
rect 7843 3406 7899 3408
rect 7698 2869 7754 2871
rect 7698 2817 7700 2869
rect 7700 2817 7752 2869
rect 7752 2817 7754 2869
rect 7698 2815 7754 2817
rect 7988 1075 8044 1077
rect 7988 1023 7990 1075
rect 7990 1023 8042 1075
rect 8042 1023 8044 1075
rect 7988 1021 8044 1023
rect 7843 -112 7899 -110
rect 7843 -164 7845 -112
rect 7845 -164 7897 -112
rect 7897 -164 7899 -112
rect 7843 -166 7899 -164
rect 7698 -707 7754 -705
rect 7698 -759 7700 -707
rect 7700 -759 7752 -707
rect 7752 -759 7754 -707
rect 7698 -761 7754 -759
rect 7843 -1822 7899 -1820
rect 7843 -1874 7845 -1822
rect 7845 -1874 7897 -1822
rect 7897 -1874 7899 -1822
rect 7843 -1876 7899 -1874
rect 7988 -2489 8044 -2487
rect 7988 -2541 7990 -2489
rect 7990 -2541 8042 -2489
rect 8042 -2541 8044 -2489
rect 7988 -2543 8044 -2541
<< metal3 >>
rect 7983 25644 8049 25649
rect 7696 23867 7756 25639
rect 7983 25588 7988 25644
rect 8044 25588 8049 25644
rect 7983 25583 8049 25588
rect 7841 24475 7901 24509
rect 7833 24469 7909 24475
rect 7833 24405 7839 24469
rect 7903 24405 7909 24469
rect 7833 24399 7909 24405
rect 7841 24365 7901 24399
rect 7693 23862 7759 23867
rect 7693 23806 7698 23862
rect 7754 23806 7759 23862
rect 7693 23801 7759 23806
rect 7696 20736 7756 23801
rect 7986 22518 8046 25583
rect 7983 22513 8049 22518
rect 7983 22457 7988 22513
rect 8044 22457 8049 22513
rect 7983 22452 8049 22457
rect 7836 21330 7902 21335
rect 7836 21274 7841 21330
rect 7897 21274 7902 21330
rect 7836 21264 7902 21274
rect 7831 21258 7907 21264
rect 7831 21194 7837 21258
rect 7901 21194 7907 21258
rect 7831 21188 7907 21194
rect 7693 20731 7759 20736
rect 7693 20675 7698 20731
rect 7754 20675 7759 20731
rect 7693 20670 7759 20675
rect 7696 17164 7756 20670
rect 7986 18947 8046 22452
rect 7983 18941 8049 18947
rect 7983 18885 7988 18941
rect 8044 18885 8049 18941
rect 7983 18880 8049 18885
rect 7838 17758 7904 17763
rect 7838 17702 7843 17758
rect 7899 17702 7904 17758
rect 7838 17692 7904 17702
rect 7833 17686 7909 17692
rect 7833 17622 7839 17686
rect 7903 17622 7909 17686
rect 7833 17616 7909 17622
rect 7693 17159 7759 17164
rect 7693 17103 7698 17159
rect 7754 17103 7759 17159
rect 7693 17098 7759 17103
rect 7696 13592 7756 17098
rect 7986 15374 8046 18880
rect 7983 15369 8049 15374
rect 7983 15313 7988 15369
rect 8044 15313 8049 15369
rect 7983 15308 8049 15313
rect 7841 14188 7901 14222
rect 7833 14182 7909 14188
rect 7833 14118 7839 14182
rect 7903 14118 7909 14182
rect 7833 14112 7909 14118
rect 7841 14078 7901 14112
rect 7693 13587 7759 13592
rect 7693 13531 7698 13587
rect 7754 13531 7759 13587
rect 7693 13526 7759 13531
rect 7696 6448 7756 13526
rect 7986 8230 8046 15308
rect 7983 8225 8049 8230
rect 7983 8169 7988 8225
rect 8044 8169 8049 8225
rect 7983 8164 8049 8169
rect 7841 7044 7901 7078
rect 7833 7038 7909 7044
rect 7833 6974 7839 7038
rect 7903 6974 7909 7038
rect 7833 6968 7909 6974
rect 7841 6934 7901 6968
rect 7693 6443 7759 6448
rect 7693 6387 7698 6443
rect 7754 6387 7759 6443
rect 7693 6382 7759 6387
rect 7696 2877 7756 6382
rect 7986 4658 8046 8164
rect 7983 4653 8049 4658
rect 7983 4597 7988 4653
rect 8044 4597 8049 4653
rect 7983 4592 8049 4597
rect 7841 3472 7901 3506
rect 7833 3466 7909 3472
rect 7833 3402 7839 3466
rect 7903 3402 7909 3466
rect 7833 3396 7909 3402
rect 7841 3362 7901 3396
rect 7693 2871 7759 2877
rect 7693 2815 7698 2871
rect 7754 2815 7759 2871
rect 7693 2810 7759 2815
rect 7696 -700 7756 2810
rect 7986 1082 8046 4592
rect 7983 1077 8049 1082
rect 7983 1021 7988 1077
rect 8044 1021 8049 1077
rect 7983 1016 8049 1021
rect 7841 -100 7901 -66
rect 7833 -106 7909 -100
rect 7833 -170 7839 -106
rect 7903 -170 7909 -106
rect 7833 -176 7909 -170
rect 7840 -210 7900 -176
rect 7693 -705 7759 -700
rect 7693 -761 7698 -705
rect 7754 -761 7759 -705
rect 7693 -766 7759 -761
rect 7696 -2538 7756 -766
rect 7838 -1820 7904 -1815
rect 7838 -1876 7843 -1820
rect 7899 -1876 7904 -1820
rect 7838 -1886 7904 -1876
rect 7833 -1892 7909 -1886
rect 7833 -1956 7839 -1892
rect 7903 -1956 7909 -1892
rect 7833 -1962 7909 -1956
rect 7986 -2482 8046 1016
rect 7983 -2487 8049 -2482
rect 7983 -2543 7988 -2487
rect 8044 -2543 8049 -2487
rect 7983 -2548 8049 -2543
<< via3 >>
rect 7839 24465 7903 24469
rect 7839 24409 7843 24465
rect 7843 24409 7899 24465
rect 7899 24409 7903 24465
rect 7839 24405 7903 24409
rect 7837 21194 7901 21258
rect 7839 17622 7903 17686
rect 7839 14178 7903 14182
rect 7839 14122 7843 14178
rect 7843 14122 7899 14178
rect 7899 14122 7903 14178
rect 7839 14118 7903 14122
rect 7839 7034 7903 7038
rect 7839 6978 7843 7034
rect 7843 6978 7899 7034
rect 7899 6978 7903 7034
rect 7839 6974 7903 6978
rect 7839 3462 7903 3466
rect 7839 3406 7843 3462
rect 7843 3406 7899 3462
rect 7899 3406 7903 3462
rect 7839 3402 7903 3406
rect 7839 -110 7903 -106
rect 7839 -166 7843 -110
rect 7843 -166 7899 -110
rect 7899 -166 7903 -110
rect 7839 -170 7903 -166
rect 7839 -1956 7903 -1892
<< metal4 >>
rect -36624 25852 -31280 25912
rect -31044 25852 -25700 25912
rect -25464 25852 -20120 25912
rect -19884 25852 -14540 25912
rect -14304 25852 -8960 25912
rect -8724 25852 -3380 25912
rect -3144 25852 2200 25912
rect 2436 25852 13920 25912
rect 14156 25852 19500 25912
rect 19736 25852 25080 25912
rect 25316 25852 30660 25912
rect 30896 25852 36240 25912
rect 36476 25852 41820 25912
rect 42056 25852 47400 25912
rect 47636 25852 52980 25912
rect -33874 24748 -28530 24808
rect -28294 24748 -22950 24808
rect -22714 24748 -17370 24808
rect -11554 24748 -6210 24808
rect 22566 24748 27910 24808
rect 33726 24748 39070 24808
rect 39306 24748 44650 24808
rect 44886 24748 50230 24808
rect 7838 24469 7904 24470
rect 7838 24467 7839 24469
rect -17134 24407 7839 24467
rect 7838 24405 7839 24407
rect 7903 24467 7904 24469
rect 7903 24407 33490 24467
rect 7903 24405 7904 24407
rect 7838 24404 7904 24405
rect -36624 24066 -31280 24126
rect -31044 24066 -25700 24126
rect -25464 24066 -20120 24126
rect -19884 24066 -14540 24126
rect -14304 24066 -8960 24126
rect -8724 24066 -3380 24126
rect -3144 24066 2200 24126
rect 2436 24066 13920 24126
rect 14156 24066 19500 24126
rect 19736 24066 25080 24126
rect 25316 24066 30660 24126
rect 30896 24066 36240 24126
rect 36476 24066 41820 24126
rect 42056 24066 47400 24126
rect 47636 24066 52980 24126
rect -33874 22962 -28530 23022
rect -28294 22962 -22950 23022
rect -22714 22962 -17370 23022
rect -11554 22962 -6210 23022
rect 22566 22962 27910 23022
rect 33726 22962 39070 23022
rect 39306 22962 44650 23022
rect 44886 22962 50230 23022
rect -36624 22280 -31280 22340
rect -31044 22280 -25700 22340
rect -25464 22280 -20120 22340
rect -19884 22280 -14540 22340
rect -14304 22280 -8960 22340
rect -8724 22280 -3380 22340
rect -3144 22280 2200 22340
rect 2436 22280 13920 22340
rect 14156 22280 19500 22340
rect 19736 22280 25080 22340
rect 25316 22280 30660 22340
rect 30896 22280 36240 22340
rect 36476 22280 41820 22340
rect 42056 22280 47400 22340
rect 47636 22280 52980 22340
rect -33874 21176 -28530 21236
rect -28294 21176 -22950 21236
rect -22714 21176 -17370 21236
rect -11554 21176 -6210 21236
rect 7836 21258 7902 21259
rect 7836 21256 7837 21258
rect -5974 21196 7837 21256
rect 7836 21194 7837 21196
rect 7901 21256 7902 21258
rect 7901 21196 22330 21256
rect 7901 21194 7902 21196
rect 7836 21193 7902 21194
rect 22566 21176 27910 21256
rect 33726 21176 39070 21236
rect 39306 21176 44650 21236
rect 44886 21176 50230 21236
rect 5186 20835 11170 20895
rect -36624 20494 -31280 20554
rect -31044 20494 -25700 20554
rect -25464 20494 -20120 20554
rect -19884 20494 -14540 20554
rect -14304 20494 -8960 20554
rect -8724 20494 -3380 20554
rect -3144 20494 2200 20554
rect 2436 20494 13920 20554
rect 14156 20494 19500 20554
rect 19736 20494 25080 20554
rect 25316 20494 30660 20554
rect 30896 20494 36240 20554
rect 36476 20494 41820 20554
rect 42056 20494 47400 20554
rect 47636 20494 52980 20554
rect -33874 19390 -28530 19450
rect -28294 19390 -22950 19450
rect -22714 19390 -17370 19450
rect -11554 19390 -6210 19450
rect 22566 19390 27910 19450
rect 33726 19390 39070 19450
rect 39306 19390 44650 19450
rect 44886 19390 50230 19450
rect -36624 18708 -31280 18768
rect -31044 18708 -25700 18768
rect -25464 18708 -20120 18768
rect -19884 18708 -14540 18768
rect -14304 18708 -8960 18768
rect -8724 18708 -3380 18768
rect -3144 18708 2200 18768
rect 2436 18708 13920 18768
rect 14156 18708 19500 18768
rect 19736 18708 25080 18768
rect 25316 18708 30660 18768
rect 30896 18708 36240 18768
rect 36476 18708 41820 18768
rect 42056 18708 47400 18768
rect 47636 18708 52980 18768
rect -33874 17604 -28530 17664
rect -28294 17604 -22950 17664
rect -22714 17604 -17370 17664
rect -11554 17604 -6210 17664
rect 7838 17686 7904 17687
rect 7838 17684 7839 17686
rect -394 17624 7839 17684
rect 7838 17622 7839 17624
rect 7903 17684 7904 17686
rect 7903 17624 16750 17684
rect 7903 17622 7904 17624
rect 7838 17621 7904 17622
rect 22566 17604 27910 17664
rect 33726 17604 39070 17664
rect 39306 17604 44650 17664
rect 44886 17604 50230 17664
rect -36624 16922 -31280 16982
rect -31044 16922 -25700 16982
rect -25464 16922 -20120 16982
rect -19884 16922 -14540 16982
rect -14304 16922 -8960 16982
rect -8724 16922 -3380 16982
rect -3144 16922 2200 16982
rect 2436 16922 13920 16982
rect 14156 16922 19500 16982
rect 19736 16922 25080 16982
rect 25316 16922 30660 16982
rect 30896 16922 36240 16982
rect 36476 16922 41820 16982
rect 42056 16922 47400 16982
rect 47636 16922 52980 16982
rect -33874 15818 -28530 15878
rect -28294 15818 -22950 15878
rect -22714 15818 -17370 15878
rect -11554 15818 -6210 15878
rect 22566 15818 27910 15878
rect 33726 15818 39070 15878
rect 39306 15818 44650 15878
rect 44886 15818 50230 15878
rect -36624 15136 -31280 15196
rect -31044 15136 -25700 15196
rect -25464 15136 -20120 15196
rect -19884 15136 -14540 15196
rect -14304 15136 -8960 15196
rect -8724 15136 -3380 15196
rect -3144 15136 2200 15196
rect 2436 15136 13920 15196
rect 14156 15136 19500 15196
rect 19736 15136 25080 15196
rect 25316 15136 30660 15196
rect 30896 15136 36240 15196
rect 36476 15136 41820 15196
rect 42056 15136 47400 15196
rect 47636 15136 52980 15196
rect 7838 14182 7904 14183
rect 7838 14180 7839 14182
rect -28294 14032 -22950 14092
rect -22714 14032 -17370 14092
rect -11554 14032 -6210 14092
rect 5186 14120 7839 14180
rect 7838 14118 7839 14120
rect 7903 14180 7904 14182
rect 7903 14120 11170 14180
rect 7903 14118 7904 14120
rect 7838 14117 7904 14118
rect 22566 14032 27910 14092
rect 33726 14032 39070 14092
rect 39306 14032 44650 14092
rect 44886 14032 50230 14092
rect -36624 13350 -31280 13410
rect -31044 13350 -25700 13410
rect -25464 13350 -20120 13410
rect -19884 13350 -14540 13410
rect -14304 13350 -8960 13410
rect -8724 13350 -3380 13410
rect -3144 13350 2200 13410
rect 2436 13350 13920 13410
rect 14156 13350 19500 13410
rect 19736 13350 25080 13410
rect 25316 13350 30660 13410
rect 30896 13350 36240 13410
rect 36476 13350 41820 13410
rect 42056 13350 47400 13410
rect 47636 13350 52980 13410
rect -33874 12246 -28530 12306
rect -28294 12246 -22950 12306
rect -22714 12246 -17370 12306
rect -11554 12246 -6210 12306
rect 22566 12246 27910 12306
rect 33726 12246 39070 12306
rect 39306 12246 44650 12306
rect 44886 12246 50230 12306
rect -36624 11564 -31280 11624
rect -31044 11564 -25700 11624
rect -25464 11564 -20120 11624
rect -19884 11564 -14540 11624
rect -14304 11564 -8960 11624
rect -8724 11564 -3380 11624
rect -3144 11564 2200 11624
rect 2436 11564 13920 11624
rect 14156 11564 19500 11624
rect 19736 11564 25080 11624
rect 25316 11564 30660 11624
rect 30896 11564 36240 11624
rect 36476 11564 41820 11624
rect 42056 11564 47400 11624
rect 47636 11564 52980 11624
rect -33874 10460 -28530 10520
rect -28294 10460 -22950 10520
rect -22714 10460 -17370 10520
rect -11554 10460 -6210 10520
rect 5186 10548 11170 10608
rect 22566 10460 27910 10520
rect 33726 10460 39070 10520
rect 39306 10460 44650 10520
rect 44886 10460 50230 10520
rect -17134 10119 33490 10179
rect -36624 9778 -31280 9838
rect -31044 9778 -25700 9838
rect -25464 9778 -20120 9838
rect -19884 9778 -14540 9838
rect -14304 9778 -8960 9838
rect -8724 9778 -3380 9838
rect -3144 9778 2200 9838
rect 2436 9778 13920 9838
rect 14156 9778 19500 9838
rect 19736 9778 25080 9838
rect 25316 9778 30660 9838
rect 30896 9778 36240 9838
rect 36476 9778 41820 9838
rect 42056 9778 47400 9838
rect 47636 9778 52980 9838
rect -33874 8674 -28530 8734
rect -28294 8674 -22950 8734
rect -22714 8674 -17370 8734
rect -11554 8674 -6210 8734
rect 22566 8674 27910 8734
rect 33726 8674 39070 8734
rect 39306 8674 44650 8734
rect 44886 8674 50230 8734
rect -36624 7992 -31280 8052
rect -31044 7992 -25700 8052
rect -25464 7992 -20120 8052
rect -19884 7992 -14540 8052
rect -14304 7992 -8960 8052
rect -8724 7992 -3380 8052
rect -3144 7992 2200 8052
rect 2436 7992 13920 8052
rect 14156 7992 19500 8052
rect 19736 7992 25080 8052
rect 25316 7992 30660 8052
rect 30896 7992 36240 8052
rect 36476 7992 41820 8052
rect 42056 7992 47400 8052
rect 47636 7992 52980 8052
rect 7838 7038 7904 7039
rect 7838 7036 7839 7038
rect -33874 6888 -28530 6948
rect -28294 6888 -22950 6948
rect -22714 6888 -17370 6948
rect -11554 6888 -6210 6948
rect 5186 6976 7839 7036
rect 7838 6974 7839 6976
rect 7903 7036 7904 7038
rect 7903 6976 11170 7036
rect 7903 6974 7904 6976
rect 7838 6973 7904 6974
rect 22566 6888 27910 6948
rect 33726 6888 39070 6948
rect 39306 6888 44650 6948
rect 44886 6888 50230 6948
rect -5974 6547 22330 6607
rect -36624 6206 -31280 6266
rect -31044 6206 -25700 6266
rect -25464 6206 -20120 6266
rect -19884 6206 -14540 6266
rect -14304 6206 -8960 6266
rect -8724 6206 -3380 6266
rect -3144 6206 2200 6266
rect 2436 6206 13920 6266
rect 14156 6206 19500 6266
rect 19736 6206 25080 6266
rect 25316 6206 30660 6266
rect 30896 6206 36240 6266
rect 36476 6206 41820 6266
rect 42056 6206 47400 6266
rect 47636 6206 52980 6266
rect -33874 5102 -28530 5162
rect -28294 5102 -22950 5162
rect -22714 5102 -17370 5162
rect -11554 5102 -6210 5162
rect 22566 5102 27910 5162
rect 33726 5102 39070 5162
rect 39306 5102 44650 5162
rect 44886 5102 50230 5162
rect -36624 4420 -31280 4480
rect -31044 4420 -25700 4480
rect -25464 4420 -20120 4480
rect -19884 4420 -14540 4480
rect -14304 4420 -8960 4480
rect -8724 4420 -3380 4480
rect -3144 4420 2200 4480
rect 2436 4420 13920 4480
rect 14156 4420 19500 4480
rect 19736 4420 25080 4480
rect 25316 4420 30660 4480
rect 30896 4420 36240 4480
rect 36476 4420 41820 4480
rect 42056 4420 47400 4480
rect 47636 4420 52980 4480
rect 7838 3466 7904 3467
rect 7838 3464 7839 3466
rect -33874 3316 -28530 3376
rect -28294 3316 -22950 3376
rect -22714 3316 -17370 3376
rect -11554 3316 -6210 3376
rect 5186 3404 7839 3464
rect 7838 3402 7839 3404
rect 7903 3464 7904 3466
rect 7903 3404 11170 3464
rect 7903 3402 7904 3404
rect 7838 3401 7904 3402
rect 22566 3316 27910 3376
rect 33726 3316 39070 3376
rect 39306 3316 44650 3376
rect 44886 3316 50230 3376
rect -394 2975 16750 3035
rect -36624 2634 -31280 2694
rect -31044 2634 -25700 2694
rect -25464 2634 -20120 2694
rect -19884 2634 -14540 2694
rect -14304 2634 -8960 2694
rect -8724 2634 -3380 2694
rect -3144 2634 2200 2694
rect 2436 2634 13920 2694
rect 14156 2634 19500 2694
rect 19736 2634 25080 2694
rect 25316 2634 30660 2694
rect 30896 2634 36240 2694
rect 36476 2634 41820 2694
rect 42056 2634 47400 2694
rect 47636 2634 52980 2694
rect -33874 1530 -28530 1590
rect -28294 1530 -22950 1590
rect -22714 1530 -17370 1590
rect -11554 1530 -6210 1590
rect 5186 1618 11170 1678
rect 22566 1530 27910 1590
rect 33726 1530 39070 1590
rect 39306 1530 44650 1590
rect 44886 1530 50230 1590
rect -36624 848 -31280 908
rect -31044 848 -25700 908
rect -25464 848 -20120 908
rect -19884 848 -14540 908
rect -14304 848 -8960 908
rect -8724 848 -3380 908
rect -3144 848 2200 908
rect 2436 848 13920 908
rect 14156 848 19500 908
rect 19736 848 25080 908
rect 25316 848 30660 908
rect 30896 848 36240 908
rect 36476 848 41820 908
rect 42056 848 47400 908
rect 47636 848 52980 908
rect 7838 -106 7904 -105
rect 7838 -108 7839 -106
rect -33874 -256 -28530 -196
rect -28294 -256 -22950 -196
rect -22714 -256 -17370 -196
rect -11554 -256 -6210 -196
rect 5186 -168 7839 -108
rect 7838 -170 7839 -168
rect 7903 -108 7904 -106
rect 7903 -168 11170 -108
rect 7903 -170 7904 -168
rect 7838 -171 7904 -170
rect 22566 -256 27910 -196
rect 33726 -256 39070 -196
rect 39306 -256 44650 -196
rect 44886 -256 50230 -196
rect -36624 -938 -31280 -878
rect -31044 -938 -25700 -878
rect -25464 -938 -20120 -878
rect -19884 -938 -14540 -878
rect -14304 -938 -8960 -878
rect -8724 -938 -3380 -878
rect -3144 -938 2200 -878
rect 2436 -938 19500 -878
rect 19736 -938 25080 -878
rect 25316 -938 30660 -878
rect 30896 -938 36240 -878
rect 36476 -938 41820 -878
rect 42056 -938 47400 -878
rect 47636 -938 52980 -878
rect 7838 -1892 7904 -1891
rect 7838 -1894 7839 -1892
rect 5186 -1954 7839 -1894
rect 7838 -1956 7839 -1954
rect 7903 -1956 7904 -1892
rect 7838 -1957 7904 -1956
<< via4 >>
rect -36860 25764 -36624 26000
rect -31280 25764 -31044 26000
rect -25700 25764 -25464 26000
rect -20120 25764 -19884 26000
rect -14540 25764 -14304 26000
rect -8960 25764 -8724 26000
rect -3380 25764 -3144 26000
rect 2200 25764 2436 26000
rect 13920 25764 14156 26000
rect 19500 25764 19736 26000
rect 25080 25764 25316 26000
rect 30660 25764 30896 26000
rect 36240 25764 36476 26000
rect 41820 25764 42056 26000
rect 47400 25764 47636 26000
rect 52980 25764 53216 26000
rect -34110 24660 -33874 24896
rect -28530 24660 -28294 24896
rect -22950 24660 -22714 24896
rect -17370 24660 -17134 24896
rect -11790 24660 -11554 24896
rect -6210 24660 -5974 24896
rect 22330 24660 22566 24896
rect 27910 24660 28146 24896
rect 33490 24660 33726 24896
rect 39070 24660 39306 24896
rect 44650 24660 44886 24896
rect 50230 24660 50466 24896
rect -17370 24319 -17134 24555
rect 33490 24319 33726 24555
rect -36860 23978 -36624 24214
rect -31280 23978 -31044 24214
rect -25700 23978 -25464 24214
rect -20120 23978 -19884 24214
rect -14540 23978 -14304 24214
rect -8960 23978 -8724 24214
rect -3380 23978 -3144 24214
rect 2200 23978 2436 24214
rect 13920 23978 14156 24214
rect 19500 23978 19736 24214
rect 25080 23978 25316 24214
rect 30660 23978 30896 24214
rect 36240 23978 36476 24214
rect 41820 23978 42056 24214
rect 47400 23978 47636 24214
rect 52980 23978 53216 24214
rect -34110 22874 -33874 23110
rect -28530 22874 -28294 23110
rect -22950 22874 -22714 23110
rect -17370 22874 -17134 23110
rect -11790 22874 -11554 23110
rect -6210 22874 -5974 23110
rect 22330 22874 22566 23110
rect 27910 22874 28146 23110
rect 33490 22874 33726 23110
rect 39070 22874 39306 23110
rect 44650 22874 44886 23110
rect 50230 22874 50466 23110
rect -36860 22192 -36624 22428
rect -31280 22192 -31044 22428
rect -25700 22192 -25464 22428
rect -20120 22192 -19884 22428
rect -14540 22192 -14304 22428
rect -8960 22192 -8724 22428
rect -3380 22192 -3144 22428
rect 2200 22192 2436 22428
rect 13920 22192 14156 22428
rect 19500 22192 19736 22428
rect 25080 22192 25316 22428
rect 30660 22192 30896 22428
rect 36240 22192 36476 22428
rect 41820 22192 42056 22428
rect 47400 22192 47636 22428
rect 52980 22192 53216 22428
rect -34110 21088 -33874 21324
rect -28530 21088 -28294 21324
rect -22950 21088 -22714 21324
rect -17370 21088 -17134 21324
rect -11790 21088 -11554 21324
rect -6210 21088 -5974 21324
rect 22330 21088 22566 21324
rect 27910 21088 28146 21324
rect 33490 21088 33726 21324
rect 39070 21088 39306 21324
rect 44650 21088 44886 21324
rect 50230 21088 50466 21324
rect 4950 20747 5186 20983
rect 11170 20747 11406 20983
rect -36860 20406 -36624 20642
rect -31280 20406 -31044 20642
rect -25700 20406 -25464 20642
rect -20120 20406 -19884 20642
rect -14540 20406 -14304 20642
rect -8960 20406 -8724 20642
rect -3380 20406 -3144 20642
rect 2200 20406 2436 20642
rect 13920 20406 14156 20642
rect 19500 20406 19736 20642
rect 25080 20406 25316 20642
rect 30660 20406 30896 20642
rect 36240 20406 36476 20642
rect 41820 20406 42056 20642
rect 47400 20406 47636 20642
rect 52980 20406 53216 20642
rect -34110 19302 -33874 19538
rect -28530 19302 -28294 19538
rect -22950 19302 -22714 19538
rect -17370 19302 -17134 19538
rect -11790 19302 -11554 19538
rect -6210 19302 -5974 19538
rect 22330 19302 22566 19538
rect 27910 19302 28146 19538
rect 33490 19302 33726 19538
rect 39070 19302 39306 19538
rect 44650 19302 44886 19538
rect 50230 19302 50466 19538
rect -36860 18620 -36624 18856
rect -31280 18620 -31044 18856
rect -25700 18620 -25464 18856
rect -20120 18620 -19884 18856
rect -14540 18620 -14304 18856
rect -8960 18620 -8724 18856
rect -3380 18620 -3144 18856
rect 2200 18620 2436 18856
rect 13920 18620 14156 18856
rect 19500 18620 19736 18856
rect 25080 18620 25316 18856
rect 30660 18620 30896 18856
rect 36240 18620 36476 18856
rect 41820 18620 42056 18856
rect 47400 18620 47636 18856
rect 52980 18620 53216 18856
rect -34110 17516 -33874 17752
rect -28530 17516 -28294 17752
rect -22950 17516 -22714 17752
rect -17370 17516 -17134 17752
rect -11790 17516 -11554 17752
rect -6210 17516 -5974 17752
rect -630 17516 -394 17752
rect 16750 17516 16986 17752
rect 22330 17516 22566 17752
rect 27910 17516 28146 17752
rect 33490 17516 33726 17752
rect 39070 17516 39306 17752
rect 44650 17516 44886 17752
rect 50230 17516 50466 17752
rect -36860 16834 -36624 17070
rect -31280 16834 -31044 17070
rect -25700 16834 -25464 17070
rect -20120 16834 -19884 17070
rect -14540 16834 -14304 17070
rect -8960 16834 -8724 17070
rect -3380 16834 -3144 17070
rect 2200 16834 2436 17070
rect 13920 16834 14156 17070
rect 19500 16834 19736 17070
rect 25080 16834 25316 17070
rect 30660 16834 30896 17070
rect 36240 16834 36476 17070
rect 41820 16834 42056 17070
rect 47400 16834 47636 17070
rect 52980 16834 53216 17070
rect -34110 15730 -33874 15966
rect -28530 15730 -28294 15966
rect -22950 15730 -22714 15966
rect -17370 15730 -17134 15966
rect -11790 15730 -11554 15966
rect -6210 15730 -5974 15966
rect 22330 15730 22566 15966
rect 27910 15730 28146 15966
rect 33490 15730 33726 15966
rect 39070 15730 39306 15966
rect 44650 15730 44886 15966
rect 50230 15730 50466 15966
rect -36860 15048 -36624 15284
rect -31280 15048 -31044 15284
rect -25700 15048 -25464 15284
rect -20120 15048 -19884 15284
rect -14540 15048 -14304 15284
rect -8960 15048 -8724 15284
rect -3380 15048 -3144 15284
rect 2200 15048 2436 15284
rect 13920 15048 14156 15284
rect 19500 15048 19736 15284
rect 25080 15048 25316 15284
rect 30660 15048 30896 15284
rect 36240 15048 36476 15284
rect 41820 15048 42056 15284
rect 47400 15048 47636 15284
rect 52980 15048 53216 15284
rect -34110 13944 -33874 14180
rect -28530 13944 -28294 14180
rect -22950 13944 -22714 14180
rect -17370 13944 -17134 14180
rect -11790 13944 -11554 14180
rect -6210 13944 -5974 14180
rect 4950 13944 5186 14180
rect 11170 13944 11406 14180
rect 22330 13944 22566 14180
rect 27910 13944 28146 14180
rect 33490 13944 33726 14180
rect 39070 13944 39306 14180
rect 44650 13944 44886 14180
rect 50230 13944 50466 14180
rect -36860 13262 -36624 13498
rect -31280 13262 -31044 13498
rect -25700 13262 -25464 13498
rect -20120 13262 -19884 13498
rect -14540 13262 -14304 13498
rect -8960 13262 -8724 13498
rect -3380 13262 -3144 13498
rect 2200 13262 2436 13498
rect 13920 13262 14156 13498
rect 19500 13262 19736 13498
rect 25080 13262 25316 13498
rect 30660 13262 30896 13498
rect 36240 13262 36476 13498
rect 41820 13262 42056 13498
rect 47400 13262 47636 13498
rect 52980 13262 53216 13498
rect -34110 12158 -33874 12394
rect -28530 12158 -28294 12394
rect -22950 12158 -22714 12394
rect -17370 12158 -17134 12394
rect -11790 12158 -11554 12394
rect -6210 12158 -5974 12394
rect 22330 12158 22566 12394
rect 27910 12158 28146 12394
rect 33490 12158 33726 12394
rect 39070 12158 39306 12394
rect 44650 12158 44886 12394
rect 50230 12158 50466 12394
rect -36860 11476 -36624 11712
rect -31280 11476 -31044 11712
rect -25700 11476 -25464 11712
rect -20120 11476 -19884 11712
rect -14540 11476 -14304 11712
rect -8960 11476 -8724 11712
rect -3380 11476 -3144 11712
rect 2200 11476 2436 11712
rect 13920 11476 14156 11712
rect 19500 11476 19736 11712
rect 25080 11476 25316 11712
rect 30660 11476 30896 11712
rect 36240 11476 36476 11712
rect 41820 11476 42056 11712
rect 47400 11476 47636 11712
rect 52980 11476 53216 11712
rect -34110 10372 -33874 10608
rect -28530 10372 -28294 10608
rect -22950 10372 -22714 10608
rect -17370 10372 -17134 10608
rect -11790 10372 -11554 10608
rect -6210 10372 -5974 10608
rect 4950 10372 5186 10608
rect 11170 10372 11406 10608
rect 22330 10372 22566 10608
rect 27910 10372 28146 10608
rect 33490 10372 33726 10608
rect 39070 10372 39306 10608
rect 44650 10372 44886 10608
rect 50230 10372 50466 10608
rect -17370 10031 -17134 10267
rect 33490 10031 33726 10267
rect -36860 9690 -36624 9926
rect -31280 9690 -31044 9926
rect -25700 9690 -25464 9926
rect -20120 9690 -19884 9926
rect -14540 9690 -14304 9926
rect -8960 9690 -8724 9926
rect -3380 9690 -3144 9926
rect 2200 9690 2436 9926
rect 13920 9690 14156 9926
rect 19500 9690 19736 9926
rect 25080 9690 25316 9926
rect 30660 9690 30896 9926
rect 36240 9690 36476 9926
rect 41820 9690 42056 9926
rect 47400 9690 47636 9926
rect 52980 9690 53216 9926
rect -34110 8586 -33874 8822
rect -28530 8586 -28294 8822
rect -22950 8586 -22714 8822
rect -17370 8586 -17134 8822
rect -11790 8586 -11554 8822
rect -6210 8586 -5974 8822
rect 22330 8586 22566 8822
rect 27910 8586 28146 8822
rect 33490 8586 33726 8822
rect 39070 8586 39306 8822
rect 44650 8586 44886 8822
rect 50230 8586 50466 8822
rect -36860 7904 -36624 8140
rect -31280 7904 -31044 8140
rect -25700 7904 -25464 8140
rect -20120 7904 -19884 8140
rect -14540 7904 -14304 8140
rect -8960 7904 -8724 8140
rect -3380 7904 -3144 8140
rect 2200 7904 2436 8140
rect 13920 7904 14156 8140
rect 19500 7904 19736 8140
rect 25080 7904 25316 8140
rect 30660 7904 30896 8140
rect 36240 7904 36476 8140
rect 41820 7904 42056 8140
rect 47400 7904 47636 8140
rect 52980 7904 53216 8140
rect -34110 6800 -33874 7036
rect -28530 6800 -28294 7036
rect -22950 6800 -22714 7036
rect -17370 6800 -17134 7036
rect -11790 6800 -11554 7036
rect -6210 6800 -5974 7036
rect 4950 6800 5186 7036
rect 11170 6800 11406 7036
rect 22330 6800 22566 7036
rect 27910 6800 28146 7036
rect 33490 6800 33726 7036
rect 39070 6800 39306 7036
rect 44650 6800 44886 7036
rect 50230 6800 50466 7036
rect -6210 6459 -5974 6695
rect 22330 6459 22566 6695
rect -36860 6118 -36624 6354
rect -31280 6118 -31044 6354
rect -25700 6118 -25464 6354
rect -20120 6118 -19884 6354
rect -14540 6118 -14304 6354
rect -8960 6118 -8724 6354
rect -3380 6118 -3144 6354
rect 2200 6118 2436 6354
rect 13920 6118 14156 6354
rect 19500 6118 19736 6354
rect 25080 6118 25316 6354
rect 30660 6118 30896 6354
rect 36240 6118 36476 6354
rect 41820 6118 42056 6354
rect 47400 6118 47636 6354
rect 52980 6118 53216 6354
rect -34110 5014 -33874 5250
rect -28530 5014 -28294 5250
rect -22950 5014 -22714 5250
rect -17370 5014 -17134 5250
rect -11790 5014 -11554 5250
rect -6210 5014 -5974 5250
rect 22330 5014 22566 5250
rect 27910 5014 28146 5250
rect 33490 5014 33726 5250
rect 39070 5014 39306 5250
rect 44650 5014 44886 5250
rect 50230 5014 50466 5250
rect -36860 4332 -36624 4568
rect -31280 4332 -31044 4568
rect -25700 4332 -25464 4568
rect -20120 4332 -19884 4568
rect -14540 4332 -14304 4568
rect -8960 4332 -8724 4568
rect -3380 4332 -3144 4568
rect 2200 4332 2436 4568
rect 13920 4332 14156 4568
rect 19500 4332 19736 4568
rect 25080 4332 25316 4568
rect 30660 4332 30896 4568
rect 36240 4332 36476 4568
rect 41820 4332 42056 4568
rect 47400 4332 47636 4568
rect 52980 4332 53216 4568
rect -34110 3228 -33874 3464
rect -28530 3228 -28294 3464
rect -22950 3228 -22714 3464
rect -17370 3228 -17134 3464
rect -11790 3228 -11554 3464
rect -6210 3228 -5974 3464
rect 4950 3228 5186 3464
rect 11170 3228 11406 3464
rect 22330 3228 22566 3464
rect 27910 3228 28146 3464
rect 33490 3228 33726 3464
rect 39070 3228 39306 3464
rect 44650 3228 44886 3464
rect 50230 3228 50466 3464
rect -630 2887 -394 3123
rect 16750 2887 16986 3123
rect -36860 2546 -36624 2782
rect -31280 2546 -31044 2782
rect -25700 2546 -25464 2782
rect -20120 2546 -19884 2782
rect -14540 2546 -14304 2782
rect -8960 2546 -8724 2782
rect -3380 2546 -3144 2782
rect 2200 2546 2436 2782
rect 13920 2546 14156 2782
rect 19500 2546 19736 2782
rect 25080 2546 25316 2782
rect 30660 2546 30896 2782
rect 36240 2546 36476 2782
rect 41820 2546 42056 2782
rect 47400 2546 47636 2782
rect 52980 2546 53216 2782
rect -34110 1442 -33874 1678
rect -28530 1442 -28294 1678
rect -22950 1442 -22714 1678
rect -17370 1442 -17134 1678
rect -11790 1442 -11554 1678
rect -6210 1442 -5974 1678
rect 4950 1442 5186 1678
rect 11170 1442 11406 1678
rect 22330 1442 22566 1678
rect 27910 1442 28146 1678
rect 33490 1442 33726 1678
rect 39070 1442 39306 1678
rect 44650 1442 44886 1678
rect 50230 1442 50466 1678
rect -36860 760 -36624 996
rect -31280 760 -31044 996
rect -25700 760 -25464 996
rect -20120 760 -19884 996
rect -14540 760 -14304 996
rect -8960 760 -8724 996
rect -3380 760 -3144 996
rect 2200 760 2436 996
rect 13920 760 14156 996
rect 19500 760 19736 996
rect 25080 760 25316 996
rect 30660 760 30896 996
rect 36240 760 36476 996
rect 41820 760 42056 996
rect 47400 760 47636 996
rect 52980 760 53216 996
rect -34110 -344 -33874 -108
rect -28530 -344 -28294 -108
rect -22950 -344 -22714 -108
rect -17370 -344 -17134 -108
rect -11790 -344 -11554 -108
rect -6210 -344 -5974 -108
rect 4950 -344 5186 -108
rect 11170 -344 11406 -108
rect 22330 -344 22566 -108
rect 27910 -344 28146 -108
rect 33490 -344 33726 -108
rect 39070 -344 39306 -108
rect 44650 -344 44886 -108
rect 50230 -344 50466 -108
rect -36860 -1026 -36624 -790
rect -31280 -1026 -31044 -790
rect -25700 -1026 -25464 -790
rect -20120 -1026 -19884 -790
rect -14540 -1026 -14304 -790
rect -8960 -1026 -8724 -790
rect -3380 -1026 -3144 -790
rect 2200 -1026 2436 -790
rect 19500 -1026 19736 -790
rect 25080 -1026 25316 -790
rect 30660 -1026 30896 -790
rect 36240 -1026 36476 -790
rect 41820 -1026 42056 -790
rect 47400 -1026 47636 -790
rect 52980 -1026 53216 -790
rect -34110 -2130 -33874 -1894
rect -28530 -2130 -28294 -1894
rect -22950 -2130 -22714 -1894
rect -17370 -2130 -17134 -1894
rect -11790 -2130 -11554 -1894
rect -6210 -2130 -5974 -1894
rect -630 -2130 -394 -1894
rect 4950 -2130 5186 -1894
rect 16750 -2130 16986 -1894
rect 22330 -2130 22566 -1894
rect 27910 -2130 28146 -1894
rect 33490 -2130 33726 -1894
rect 39070 -2130 39306 -1894
rect 44650 -2130 44886 -1894
rect 50230 -2130 50466 -1894
<< metal5 >>
rect -36902 26000 -36582 26024
rect -36902 25764 -36860 26000
rect -36624 25764 -36582 26000
rect -36902 24214 -36582 25764
rect -31322 26000 -31002 26024
rect -31322 25764 -31280 26000
rect -31044 25764 -31002 26000
rect -36902 23978 -36860 24214
rect -36624 23978 -36582 24214
rect -36902 22428 -36582 23978
rect -36902 22192 -36860 22428
rect -36624 22192 -36582 22428
rect -36902 20642 -36582 22192
rect -36902 20406 -36860 20642
rect -36624 20406 -36582 20642
rect -36902 18856 -36582 20406
rect -36902 18620 -36860 18856
rect -36624 18620 -36582 18856
rect -36902 17070 -36582 18620
rect -36902 16834 -36860 17070
rect -36624 16834 -36582 17070
rect -36902 15284 -36582 16834
rect -36902 15048 -36860 15284
rect -36624 15048 -36582 15284
rect -36902 13498 -36582 15048
rect -36902 13262 -36860 13498
rect -36624 13262 -36582 13498
rect -36902 11712 -36582 13262
rect -36902 11476 -36860 11712
rect -36624 11476 -36582 11712
rect -36902 9926 -36582 11476
rect -36902 9690 -36860 9926
rect -36624 9690 -36582 9926
rect -36902 8140 -36582 9690
rect -36902 7904 -36860 8140
rect -36624 7904 -36582 8140
rect -36902 6354 -36582 7904
rect -36902 6118 -36860 6354
rect -36624 6118 -36582 6354
rect -36902 4568 -36582 6118
rect -36902 4332 -36860 4568
rect -36624 4332 -36582 4568
rect -36902 2782 -36582 4332
rect -36902 2546 -36860 2782
rect -36624 2546 -36582 2782
rect -36902 996 -36582 2546
rect -36902 760 -36860 996
rect -36624 760 -36582 996
rect -36902 -790 -36582 760
rect -36902 -1026 -36860 -790
rect -36624 -1026 -36582 -790
rect -36902 -1894 -36582 -1026
rect -34152 24896 -33832 25696
rect -34152 24660 -34110 24896
rect -33874 24660 -33832 24896
rect -34152 23110 -33832 24660
rect -34152 22874 -34110 23110
rect -33874 22874 -33832 23110
rect -34152 21324 -33832 22874
rect -34152 21088 -34110 21324
rect -33874 21088 -33832 21324
rect -34152 19538 -33832 21088
rect -34152 19302 -34110 19538
rect -33874 19302 -33832 19538
rect -34152 17752 -33832 19302
rect -34152 17516 -34110 17752
rect -33874 17516 -33832 17752
rect -34152 15966 -33832 17516
rect -34152 15730 -34110 15966
rect -33874 15730 -33832 15966
rect -34152 14180 -33832 15730
rect -34152 13944 -34110 14180
rect -33874 13944 -33832 14180
rect -34152 12394 -33832 13944
rect -34152 12158 -34110 12394
rect -33874 12158 -33832 12394
rect -34152 10608 -33832 12158
rect -34152 10372 -34110 10608
rect -33874 10372 -33832 10608
rect -34152 8822 -33832 10372
rect -34152 8586 -34110 8822
rect -33874 8586 -33832 8822
rect -34152 7036 -33832 8586
rect -34152 6800 -34110 7036
rect -33874 6800 -33832 7036
rect -34152 5250 -33832 6800
rect -34152 5014 -34110 5250
rect -33874 5014 -33832 5250
rect -34152 3464 -33832 5014
rect -34152 3228 -34110 3464
rect -33874 3228 -33832 3464
rect -34152 1678 -33832 3228
rect -34152 1442 -34110 1678
rect -33874 1442 -33832 1678
rect -34152 -108 -33832 1442
rect -34152 -344 -34110 -108
rect -33874 -344 -33832 -108
rect -34152 -1894 -33832 -344
rect -31322 24214 -31002 25764
rect -25742 26000 -25422 26024
rect -25742 25764 -25700 26000
rect -25464 25764 -25422 26000
rect -31322 23978 -31280 24214
rect -31044 23978 -31002 24214
rect -31322 22428 -31002 23978
rect -31322 22192 -31280 22428
rect -31044 22192 -31002 22428
rect -31322 20642 -31002 22192
rect -31322 20406 -31280 20642
rect -31044 20406 -31002 20642
rect -31322 18856 -31002 20406
rect -31322 18620 -31280 18856
rect -31044 18620 -31002 18856
rect -31322 17070 -31002 18620
rect -31322 16834 -31280 17070
rect -31044 16834 -31002 17070
rect -31322 15284 -31002 16834
rect -31322 15048 -31280 15284
rect -31044 15048 -31002 15284
rect -31322 13498 -31002 15048
rect -31322 13262 -31280 13498
rect -31044 13262 -31002 13498
rect -31322 11712 -31002 13262
rect -31322 11476 -31280 11712
rect -31044 11476 -31002 11712
rect -31322 9926 -31002 11476
rect -31322 9690 -31280 9926
rect -31044 9690 -31002 9926
rect -31322 8140 -31002 9690
rect -31322 7904 -31280 8140
rect -31044 7904 -31002 8140
rect -31322 6354 -31002 7904
rect -31322 6118 -31280 6354
rect -31044 6118 -31002 6354
rect -31322 4568 -31002 6118
rect -31322 4332 -31280 4568
rect -31044 4332 -31002 4568
rect -31322 2782 -31002 4332
rect -31322 2546 -31280 2782
rect -31044 2546 -31002 2782
rect -31322 996 -31002 2546
rect -31322 760 -31280 996
rect -31044 760 -31002 996
rect -31322 -790 -31002 760
rect -31322 -1026 -31280 -790
rect -31044 -1026 -31002 -790
rect -31322 -1894 -31002 -1026
rect -28572 24896 -28252 25696
rect -28572 24660 -28530 24896
rect -28294 24660 -28252 24896
rect -28572 23110 -28252 24660
rect -28572 22874 -28530 23110
rect -28294 22874 -28252 23110
rect -28572 21324 -28252 22874
rect -28572 21088 -28530 21324
rect -28294 21088 -28252 21324
rect -28572 19538 -28252 21088
rect -28572 19302 -28530 19538
rect -28294 19302 -28252 19538
rect -28572 17752 -28252 19302
rect -28572 17516 -28530 17752
rect -28294 17516 -28252 17752
rect -28572 15966 -28252 17516
rect -28572 15730 -28530 15966
rect -28294 15730 -28252 15966
rect -28572 14180 -28252 15730
rect -28572 13944 -28530 14180
rect -28294 13944 -28252 14180
rect -28572 12394 -28252 13944
rect -28572 12158 -28530 12394
rect -28294 12158 -28252 12394
rect -28572 10608 -28252 12158
rect -28572 10372 -28530 10608
rect -28294 10372 -28252 10608
rect -28572 8822 -28252 10372
rect -28572 8586 -28530 8822
rect -28294 8586 -28252 8822
rect -28572 7036 -28252 8586
rect -28572 6800 -28530 7036
rect -28294 6800 -28252 7036
rect -28572 5250 -28252 6800
rect -28572 5014 -28530 5250
rect -28294 5014 -28252 5250
rect -28572 3464 -28252 5014
rect -28572 3228 -28530 3464
rect -28294 3228 -28252 3464
rect -28572 1678 -28252 3228
rect -28572 1442 -28530 1678
rect -28294 1442 -28252 1678
rect -28572 -108 -28252 1442
rect -28572 -344 -28530 -108
rect -28294 -344 -28252 -108
rect -28572 -1894 -28252 -344
rect -25742 24214 -25422 25764
rect -20162 26000 -19842 26024
rect -20162 25764 -20120 26000
rect -19884 25764 -19842 26000
rect -25742 23978 -25700 24214
rect -25464 23978 -25422 24214
rect -25742 22428 -25422 23978
rect -25742 22192 -25700 22428
rect -25464 22192 -25422 22428
rect -25742 20642 -25422 22192
rect -25742 20406 -25700 20642
rect -25464 20406 -25422 20642
rect -25742 18856 -25422 20406
rect -25742 18620 -25700 18856
rect -25464 18620 -25422 18856
rect -25742 17070 -25422 18620
rect -25742 16834 -25700 17070
rect -25464 16834 -25422 17070
rect -25742 15284 -25422 16834
rect -25742 15048 -25700 15284
rect -25464 15048 -25422 15284
rect -25742 13498 -25422 15048
rect -25742 13262 -25700 13498
rect -25464 13262 -25422 13498
rect -25742 11712 -25422 13262
rect -25742 11476 -25700 11712
rect -25464 11476 -25422 11712
rect -25742 9926 -25422 11476
rect -25742 9690 -25700 9926
rect -25464 9690 -25422 9926
rect -25742 8140 -25422 9690
rect -25742 7904 -25700 8140
rect -25464 7904 -25422 8140
rect -25742 6354 -25422 7904
rect -25742 6118 -25700 6354
rect -25464 6118 -25422 6354
rect -25742 4568 -25422 6118
rect -25742 4332 -25700 4568
rect -25464 4332 -25422 4568
rect -25742 2782 -25422 4332
rect -25742 2546 -25700 2782
rect -25464 2546 -25422 2782
rect -25742 996 -25422 2546
rect -25742 760 -25700 996
rect -25464 760 -25422 996
rect -25742 -790 -25422 760
rect -25742 -1026 -25700 -790
rect -25464 -1026 -25422 -790
rect -25742 -1894 -25422 -1026
rect -22992 24896 -22672 25696
rect -22992 24660 -22950 24896
rect -22714 24660 -22672 24896
rect -22992 23110 -22672 24660
rect -22992 22874 -22950 23110
rect -22714 22874 -22672 23110
rect -22992 21324 -22672 22874
rect -22992 21088 -22950 21324
rect -22714 21088 -22672 21324
rect -22992 19538 -22672 21088
rect -22992 19302 -22950 19538
rect -22714 19302 -22672 19538
rect -22992 17752 -22672 19302
rect -22992 17516 -22950 17752
rect -22714 17516 -22672 17752
rect -22992 15966 -22672 17516
rect -22992 15730 -22950 15966
rect -22714 15730 -22672 15966
rect -22992 14180 -22672 15730
rect -22992 13944 -22950 14180
rect -22714 13944 -22672 14180
rect -22992 12394 -22672 13944
rect -22992 12158 -22950 12394
rect -22714 12158 -22672 12394
rect -22992 10608 -22672 12158
rect -22992 10372 -22950 10608
rect -22714 10372 -22672 10608
rect -22992 8822 -22672 10372
rect -22992 8586 -22950 8822
rect -22714 8586 -22672 8822
rect -22992 7036 -22672 8586
rect -22992 6800 -22950 7036
rect -22714 6800 -22672 7036
rect -22992 5250 -22672 6800
rect -22992 5014 -22950 5250
rect -22714 5014 -22672 5250
rect -22992 3464 -22672 5014
rect -22992 3228 -22950 3464
rect -22714 3228 -22672 3464
rect -22992 1678 -22672 3228
rect -22992 1442 -22950 1678
rect -22714 1442 -22672 1678
rect -22992 -108 -22672 1442
rect -22992 -344 -22950 -108
rect -22714 -344 -22672 -108
rect -22992 -1894 -22672 -344
rect -20162 24214 -19842 25764
rect -14582 26000 -14262 26024
rect -14582 25764 -14540 26000
rect -14304 25764 -14262 26000
rect -20162 23978 -20120 24214
rect -19884 23978 -19842 24214
rect -20162 22428 -19842 23978
rect -20162 22192 -20120 22428
rect -19884 22192 -19842 22428
rect -20162 20642 -19842 22192
rect -20162 20406 -20120 20642
rect -19884 20406 -19842 20642
rect -20162 18856 -19842 20406
rect -20162 18620 -20120 18856
rect -19884 18620 -19842 18856
rect -20162 17070 -19842 18620
rect -20162 16834 -20120 17070
rect -19884 16834 -19842 17070
rect -20162 15284 -19842 16834
rect -20162 15048 -20120 15284
rect -19884 15048 -19842 15284
rect -20162 13498 -19842 15048
rect -20162 13262 -20120 13498
rect -19884 13262 -19842 13498
rect -20162 11712 -19842 13262
rect -20162 11476 -20120 11712
rect -19884 11476 -19842 11712
rect -20162 9926 -19842 11476
rect -20162 9690 -20120 9926
rect -19884 9690 -19842 9926
rect -20162 8140 -19842 9690
rect -20162 7904 -20120 8140
rect -19884 7904 -19842 8140
rect -20162 6354 -19842 7904
rect -20162 6118 -20120 6354
rect -19884 6118 -19842 6354
rect -20162 4568 -19842 6118
rect -20162 4332 -20120 4568
rect -19884 4332 -19842 4568
rect -20162 2782 -19842 4332
rect -20162 2546 -20120 2782
rect -19884 2546 -19842 2782
rect -20162 996 -19842 2546
rect -20162 760 -20120 996
rect -19884 760 -19842 996
rect -20162 -790 -19842 760
rect -20162 -1026 -20120 -790
rect -19884 -1026 -19842 -790
rect -20162 -1894 -19842 -1026
rect -17412 24896 -17092 25696
rect -17412 24660 -17370 24896
rect -17134 24660 -17092 24896
rect -17412 24555 -17092 24660
rect -17412 24319 -17370 24555
rect -17134 24319 -17092 24555
rect -17412 23110 -17092 24319
rect -17412 22874 -17370 23110
rect -17134 22874 -17092 23110
rect -17412 21324 -17092 22874
rect -17412 21088 -17370 21324
rect -17134 21088 -17092 21324
rect -17412 19538 -17092 21088
rect -17412 19302 -17370 19538
rect -17134 19302 -17092 19538
rect -17412 17752 -17092 19302
rect -17412 17516 -17370 17752
rect -17134 17516 -17092 17752
rect -17412 15966 -17092 17516
rect -17412 15730 -17370 15966
rect -17134 15730 -17092 15966
rect -17412 14180 -17092 15730
rect -17412 13944 -17370 14180
rect -17134 13944 -17092 14180
rect -17412 12394 -17092 13944
rect -17412 12158 -17370 12394
rect -17134 12158 -17092 12394
rect -17412 10608 -17092 12158
rect -17412 10372 -17370 10608
rect -17134 10372 -17092 10608
rect -17412 10267 -17092 10372
rect -17412 10031 -17370 10267
rect -17134 10031 -17092 10267
rect -17412 8822 -17092 10031
rect -17412 8586 -17370 8822
rect -17134 8586 -17092 8822
rect -17412 7036 -17092 8586
rect -17412 6800 -17370 7036
rect -17134 6800 -17092 7036
rect -17412 5250 -17092 6800
rect -17412 5014 -17370 5250
rect -17134 5014 -17092 5250
rect -17412 3464 -17092 5014
rect -17412 3228 -17370 3464
rect -17134 3228 -17092 3464
rect -17412 1678 -17092 3228
rect -17412 1442 -17370 1678
rect -17134 1442 -17092 1678
rect -17412 -108 -17092 1442
rect -17412 -344 -17370 -108
rect -17134 -344 -17092 -108
rect -17412 -1894 -17092 -344
rect -14582 24214 -14262 25764
rect -9002 26000 -8682 26024
rect -9002 25764 -8960 26000
rect -8724 25764 -8682 26000
rect -14582 23978 -14540 24214
rect -14304 23978 -14262 24214
rect -14582 22428 -14262 23978
rect -14582 22192 -14540 22428
rect -14304 22192 -14262 22428
rect -14582 20642 -14262 22192
rect -14582 20406 -14540 20642
rect -14304 20406 -14262 20642
rect -14582 18856 -14262 20406
rect -14582 18620 -14540 18856
rect -14304 18620 -14262 18856
rect -14582 17070 -14262 18620
rect -14582 16834 -14540 17070
rect -14304 16834 -14262 17070
rect -14582 15284 -14262 16834
rect -14582 15048 -14540 15284
rect -14304 15048 -14262 15284
rect -14582 13498 -14262 15048
rect -14582 13262 -14540 13498
rect -14304 13262 -14262 13498
rect -14582 11712 -14262 13262
rect -14582 11476 -14540 11712
rect -14304 11476 -14262 11712
rect -14582 9926 -14262 11476
rect -14582 9690 -14540 9926
rect -14304 9690 -14262 9926
rect -14582 8140 -14262 9690
rect -14582 7904 -14540 8140
rect -14304 7904 -14262 8140
rect -14582 6354 -14262 7904
rect -14582 6118 -14540 6354
rect -14304 6118 -14262 6354
rect -14582 4568 -14262 6118
rect -14582 4332 -14540 4568
rect -14304 4332 -14262 4568
rect -14582 2782 -14262 4332
rect -14582 2546 -14540 2782
rect -14304 2546 -14262 2782
rect -14582 996 -14262 2546
rect -14582 760 -14540 996
rect -14304 760 -14262 996
rect -14582 -790 -14262 760
rect -14582 -1026 -14540 -790
rect -14304 -1026 -14262 -790
rect -14582 -1894 -14262 -1026
rect -11832 24896 -11512 25696
rect -11832 24660 -11790 24896
rect -11554 24660 -11512 24896
rect -11832 23110 -11512 24660
rect -11832 22874 -11790 23110
rect -11554 22874 -11512 23110
rect -11832 21324 -11512 22874
rect -11832 21088 -11790 21324
rect -11554 21088 -11512 21324
rect -11832 19538 -11512 21088
rect -11832 19302 -11790 19538
rect -11554 19302 -11512 19538
rect -11832 17752 -11512 19302
rect -11832 17516 -11790 17752
rect -11554 17516 -11512 17752
rect -11832 15966 -11512 17516
rect -11832 15730 -11790 15966
rect -11554 15730 -11512 15966
rect -11832 14180 -11512 15730
rect -11832 13944 -11790 14180
rect -11554 13944 -11512 14180
rect -11832 12394 -11512 13944
rect -11832 12158 -11790 12394
rect -11554 12158 -11512 12394
rect -11832 10608 -11512 12158
rect -11832 10372 -11790 10608
rect -11554 10372 -11512 10608
rect -11832 8822 -11512 10372
rect -11832 8586 -11790 8822
rect -11554 8586 -11512 8822
rect -11832 7036 -11512 8586
rect -11832 6800 -11790 7036
rect -11554 6800 -11512 7036
rect -11832 5250 -11512 6800
rect -11832 5014 -11790 5250
rect -11554 5014 -11512 5250
rect -11832 3464 -11512 5014
rect -11832 3228 -11790 3464
rect -11554 3228 -11512 3464
rect -11832 1678 -11512 3228
rect -11832 1442 -11790 1678
rect -11554 1442 -11512 1678
rect -11832 -108 -11512 1442
rect -11832 -344 -11790 -108
rect -11554 -344 -11512 -108
rect -11832 -1894 -11512 -344
rect -9002 24214 -8682 25764
rect -3422 26000 -3102 26024
rect -3422 25764 -3380 26000
rect -3144 25764 -3102 26000
rect -9002 23978 -8960 24214
rect -8724 23978 -8682 24214
rect -9002 22428 -8682 23978
rect -9002 22192 -8960 22428
rect -8724 22192 -8682 22428
rect -9002 20642 -8682 22192
rect -9002 20406 -8960 20642
rect -8724 20406 -8682 20642
rect -9002 18856 -8682 20406
rect -9002 18620 -8960 18856
rect -8724 18620 -8682 18856
rect -9002 17070 -8682 18620
rect -9002 16834 -8960 17070
rect -8724 16834 -8682 17070
rect -9002 15284 -8682 16834
rect -9002 15048 -8960 15284
rect -8724 15048 -8682 15284
rect -9002 13498 -8682 15048
rect -9002 13262 -8960 13498
rect -8724 13262 -8682 13498
rect -9002 11712 -8682 13262
rect -9002 11476 -8960 11712
rect -8724 11476 -8682 11712
rect -9002 9926 -8682 11476
rect -9002 9690 -8960 9926
rect -8724 9690 -8682 9926
rect -9002 8140 -8682 9690
rect -9002 7904 -8960 8140
rect -8724 7904 -8682 8140
rect -9002 6354 -8682 7904
rect -9002 6118 -8960 6354
rect -8724 6118 -8682 6354
rect -9002 4568 -8682 6118
rect -9002 4332 -8960 4568
rect -8724 4332 -8682 4568
rect -9002 2782 -8682 4332
rect -9002 2546 -8960 2782
rect -8724 2546 -8682 2782
rect -9002 996 -8682 2546
rect -9002 760 -8960 996
rect -8724 760 -8682 996
rect -9002 -790 -8682 760
rect -9002 -1026 -8960 -790
rect -8724 -1026 -8682 -790
rect -9002 -1894 -8682 -1026
rect -6252 24896 -5932 25696
rect -6252 24660 -6210 24896
rect -5974 24660 -5932 24896
rect -6252 23110 -5932 24660
rect -6252 22874 -6210 23110
rect -5974 22874 -5932 23110
rect -6252 21324 -5932 22874
rect -6252 21088 -6210 21324
rect -5974 21088 -5932 21324
rect -6252 19538 -5932 21088
rect -6252 19302 -6210 19538
rect -5974 19302 -5932 19538
rect -6252 17752 -5932 19302
rect -6252 17516 -6210 17752
rect -5974 17516 -5932 17752
rect -6252 15966 -5932 17516
rect -6252 15730 -6210 15966
rect -5974 15730 -5932 15966
rect -6252 14180 -5932 15730
rect -6252 13944 -6210 14180
rect -5974 13944 -5932 14180
rect -6252 12394 -5932 13944
rect -6252 12158 -6210 12394
rect -5974 12158 -5932 12394
rect -6252 10608 -5932 12158
rect -6252 10372 -6210 10608
rect -5974 10372 -5932 10608
rect -6252 8822 -5932 10372
rect -6252 8586 -6210 8822
rect -5974 8586 -5932 8822
rect -6252 7036 -5932 8586
rect -6252 6800 -6210 7036
rect -5974 6800 -5932 7036
rect -6252 6695 -5932 6800
rect -6252 6459 -6210 6695
rect -5974 6459 -5932 6695
rect -6252 5250 -5932 6459
rect -6252 5014 -6210 5250
rect -5974 5014 -5932 5250
rect -6252 3464 -5932 5014
rect -6252 3228 -6210 3464
rect -5974 3228 -5932 3464
rect -6252 1678 -5932 3228
rect -6252 1442 -6210 1678
rect -5974 1442 -5932 1678
rect -6252 -108 -5932 1442
rect -6252 -344 -6210 -108
rect -5974 -344 -5932 -108
rect -6252 -1894 -5932 -344
rect -3422 24214 -3102 25764
rect 2158 26000 2478 26024
rect 2158 25764 2200 26000
rect 2436 25764 2478 26000
rect -3422 23978 -3380 24214
rect -3144 23978 -3102 24214
rect -3422 22428 -3102 23978
rect -3422 22192 -3380 22428
rect -3144 22192 -3102 22428
rect -3422 20642 -3102 22192
rect -3422 20406 -3380 20642
rect -3144 20406 -3102 20642
rect -3422 18856 -3102 20406
rect -3422 18620 -3380 18856
rect -3144 18620 -3102 18856
rect -3422 17070 -3102 18620
rect -3422 16834 -3380 17070
rect -3144 16834 -3102 17070
rect -3422 15284 -3102 16834
rect -3422 15048 -3380 15284
rect -3144 15048 -3102 15284
rect -3422 13498 -3102 15048
rect -3422 13262 -3380 13498
rect -3144 13262 -3102 13498
rect -3422 11712 -3102 13262
rect -3422 11476 -3380 11712
rect -3144 11476 -3102 11712
rect -3422 9926 -3102 11476
rect -3422 9690 -3380 9926
rect -3144 9690 -3102 9926
rect -3422 8140 -3102 9690
rect -3422 7904 -3380 8140
rect -3144 7904 -3102 8140
rect -3422 6354 -3102 7904
rect -3422 6118 -3380 6354
rect -3144 6118 -3102 6354
rect -3422 4568 -3102 6118
rect -3422 4332 -3380 4568
rect -3144 4332 -3102 4568
rect -3422 2782 -3102 4332
rect -3422 2546 -3380 2782
rect -3144 2546 -3102 2782
rect -3422 996 -3102 2546
rect -3422 760 -3380 996
rect -3144 760 -3102 996
rect -3422 -790 -3102 760
rect -3422 -1026 -3380 -790
rect -3144 -1026 -3102 -790
rect -3422 -1894 -3102 -1026
rect -672 17752 -352 25696
rect -672 17516 -630 17752
rect -394 17516 -352 17752
rect -672 3123 -352 17516
rect -672 2887 -630 3123
rect -394 2887 -352 3123
rect -672 -1894 -352 2887
rect 2158 24214 2478 25764
rect 13878 26000 14198 26024
rect 13878 25764 13920 26000
rect 14156 25764 14198 26000
rect 2158 23978 2200 24214
rect 2436 23978 2478 24214
rect 2158 22428 2478 23978
rect 2158 22192 2200 22428
rect 2436 22192 2478 22428
rect 2158 20642 2478 22192
rect 2158 20406 2200 20642
rect 2436 20406 2478 20642
rect 2158 18856 2478 20406
rect 2158 18620 2200 18856
rect 2436 18620 2478 18856
rect 2158 17070 2478 18620
rect 2158 16834 2200 17070
rect 2436 16834 2478 17070
rect 2158 15284 2478 16834
rect 2158 15048 2200 15284
rect 2436 15048 2478 15284
rect 2158 13498 2478 15048
rect 2158 13262 2200 13498
rect 2436 13262 2478 13498
rect 2158 11712 2478 13262
rect 4908 20983 5228 25696
rect 4908 20747 4950 20983
rect 5186 20747 5228 20983
rect 4908 14180 5228 20747
rect 4908 13944 4950 14180
rect 5186 13944 5228 14180
rect 4908 12394 5228 13944
rect 11128 20983 11448 25696
rect 11128 20747 11170 20983
rect 11406 20747 11448 20983
rect 11128 14180 11448 20747
rect 11128 13944 11170 14180
rect 11406 13944 11448 14180
rect 11128 12394 11448 13944
rect 13878 24214 14198 25764
rect 19458 26000 19778 26024
rect 19458 25764 19500 26000
rect 19736 25764 19778 26000
rect 13878 23978 13920 24214
rect 14156 23978 14198 24214
rect 13878 22428 14198 23978
rect 13878 22192 13920 22428
rect 14156 22192 14198 22428
rect 13878 20642 14198 22192
rect 13878 20406 13920 20642
rect 14156 20406 14198 20642
rect 13878 18856 14198 20406
rect 13878 18620 13920 18856
rect 14156 18620 14198 18856
rect 13878 17070 14198 18620
rect 13878 16834 13920 17070
rect 14156 16834 14198 17070
rect 13878 15284 14198 16834
rect 13878 15048 13920 15284
rect 14156 15048 14198 15284
rect 13878 13498 14198 15048
rect 13878 13262 13920 13498
rect 14156 13262 14198 13498
rect 2158 11476 2200 11712
rect 2436 11476 2478 11712
rect 2158 9926 2478 11476
rect 13878 11712 14198 13262
rect 13878 11476 13920 11712
rect 14156 11476 14198 11712
rect 2158 9690 2200 9926
rect 2436 9690 2478 9926
rect 2158 8140 2478 9690
rect 2158 7904 2200 8140
rect 2436 7904 2478 8140
rect 2158 6354 2478 7904
rect 2158 6118 2200 6354
rect 2436 6118 2478 6354
rect 2158 4568 2478 6118
rect 4908 10608 5228 11408
rect 4908 10372 4950 10608
rect 5186 10372 5228 10608
rect 4908 7036 5228 10372
rect 4908 6800 4950 7036
rect 5186 6800 5228 7036
rect 4908 5250 5228 6800
rect 11128 10608 11448 11408
rect 11128 10372 11170 10608
rect 11406 10372 11448 10608
rect 11128 7036 11448 10372
rect 11128 6800 11170 7036
rect 11406 6800 11448 7036
rect 11128 5250 11448 6800
rect 13878 9926 14198 11476
rect 13878 9690 13920 9926
rect 14156 9690 14198 9926
rect 13878 8140 14198 9690
rect 13878 7904 13920 8140
rect 14156 7904 14198 8140
rect 13878 6354 14198 7904
rect 13878 6118 13920 6354
rect 14156 6118 14198 6354
rect 2158 4332 2200 4568
rect 2436 4332 2478 4568
rect 2158 2782 2478 4332
rect 13878 4568 14198 6118
rect 13878 4332 13920 4568
rect 14156 4332 14198 4568
rect 2158 2546 2200 2782
rect 2436 2546 2478 2782
rect 2158 996 2478 2546
rect 4908 3464 5228 4264
rect 4908 3228 4950 3464
rect 5186 3228 5228 3464
rect 4908 1678 5228 3228
rect 4908 1442 4950 1678
rect 5186 1442 5228 1678
rect 4908 1418 5228 1442
rect 11128 3464 11448 4264
rect 11128 3228 11170 3464
rect 11406 3228 11448 3464
rect 11128 1678 11448 3228
rect 11128 1442 11170 1678
rect 11406 1442 11448 1678
rect 11128 1418 11448 1442
rect 13878 2782 14198 4332
rect 13878 2546 13920 2782
rect 14156 2546 14198 2782
rect 2158 760 2200 996
rect 2436 760 2478 996
rect 2158 -790 2478 760
rect 13878 996 14198 2546
rect 13878 760 13920 996
rect 14156 760 14198 996
rect 4908 -108 5228 692
rect 4908 -344 4950 -108
rect 5186 -344 5228 -108
rect 4908 -368 5228 -344
rect 11128 -108 11448 692
rect 13878 -108 14198 760
rect 16708 17752 17028 25696
rect 16708 17516 16750 17752
rect 16986 17516 17028 17752
rect 16708 3123 17028 17516
rect 16708 2887 16750 3123
rect 16986 2887 17028 3123
rect 11128 -344 11170 -108
rect 11406 -344 11448 -108
rect 11128 -368 11448 -344
rect 2158 -1026 2200 -790
rect 2436 -1026 2478 -790
rect 2158 -1894 2478 -1026
rect 4908 -1894 5228 -1094
rect -34152 -2130 -34110 -1894
rect -33874 -2130 -33832 -1894
rect -34152 -2154 -33832 -2130
rect -28572 -2130 -28530 -1894
rect -28294 -2130 -28252 -1894
rect -28572 -2154 -28252 -2130
rect -22992 -2130 -22950 -1894
rect -22714 -2130 -22672 -1894
rect -22992 -2154 -22672 -2130
rect -17412 -2130 -17370 -1894
rect -17134 -2130 -17092 -1894
rect -17412 -2154 -17092 -2130
rect -11832 -2130 -11790 -1894
rect -11554 -2130 -11512 -1894
rect -11832 -2154 -11512 -2130
rect -6252 -2130 -6210 -1894
rect -5974 -2130 -5932 -1894
rect -6252 -2154 -5932 -2130
rect -672 -2130 -630 -1894
rect -394 -2130 -352 -1894
rect -672 -2154 -352 -2130
rect 4908 -2130 4950 -1894
rect 5186 -2130 5228 -1894
rect 4908 -2154 5228 -2130
rect 16708 -1894 17028 2887
rect 19458 24214 19778 25764
rect 25038 26000 25358 26024
rect 25038 25764 25080 26000
rect 25316 25764 25358 26000
rect 19458 23978 19500 24214
rect 19736 23978 19778 24214
rect 19458 22428 19778 23978
rect 19458 22192 19500 22428
rect 19736 22192 19778 22428
rect 19458 20642 19778 22192
rect 19458 20406 19500 20642
rect 19736 20406 19778 20642
rect 19458 18856 19778 20406
rect 19458 18620 19500 18856
rect 19736 18620 19778 18856
rect 19458 17070 19778 18620
rect 19458 16834 19500 17070
rect 19736 16834 19778 17070
rect 19458 15284 19778 16834
rect 19458 15048 19500 15284
rect 19736 15048 19778 15284
rect 19458 13498 19778 15048
rect 19458 13262 19500 13498
rect 19736 13262 19778 13498
rect 19458 11712 19778 13262
rect 19458 11476 19500 11712
rect 19736 11476 19778 11712
rect 19458 9926 19778 11476
rect 19458 9690 19500 9926
rect 19736 9690 19778 9926
rect 19458 8140 19778 9690
rect 19458 7904 19500 8140
rect 19736 7904 19778 8140
rect 19458 6354 19778 7904
rect 19458 6118 19500 6354
rect 19736 6118 19778 6354
rect 19458 4568 19778 6118
rect 19458 4332 19500 4568
rect 19736 4332 19778 4568
rect 19458 2782 19778 4332
rect 19458 2546 19500 2782
rect 19736 2546 19778 2782
rect 19458 996 19778 2546
rect 19458 760 19500 996
rect 19736 760 19778 996
rect 19458 -790 19778 760
rect 19458 -1026 19500 -790
rect 19736 -1026 19778 -790
rect 19458 -1894 19778 -1026
rect 22288 24896 22608 25696
rect 22288 24660 22330 24896
rect 22566 24660 22608 24896
rect 22288 23110 22608 24660
rect 22288 22874 22330 23110
rect 22566 22874 22608 23110
rect 22288 21324 22608 22874
rect 22288 21088 22330 21324
rect 22566 21088 22608 21324
rect 22288 19538 22608 21088
rect 22288 19302 22330 19538
rect 22566 19302 22608 19538
rect 22288 17752 22608 19302
rect 22288 17516 22330 17752
rect 22566 17516 22608 17752
rect 22288 15966 22608 17516
rect 22288 15730 22330 15966
rect 22566 15730 22608 15966
rect 22288 14180 22608 15730
rect 22288 13944 22330 14180
rect 22566 13944 22608 14180
rect 22288 12394 22608 13944
rect 22288 12158 22330 12394
rect 22566 12158 22608 12394
rect 22288 10608 22608 12158
rect 22288 10372 22330 10608
rect 22566 10372 22608 10608
rect 22288 8822 22608 10372
rect 22288 8586 22330 8822
rect 22566 8586 22608 8822
rect 22288 7036 22608 8586
rect 22288 6800 22330 7036
rect 22566 6800 22608 7036
rect 22288 6695 22608 6800
rect 22288 6459 22330 6695
rect 22566 6459 22608 6695
rect 22288 5250 22608 6459
rect 22288 5014 22330 5250
rect 22566 5014 22608 5250
rect 22288 3464 22608 5014
rect 22288 3228 22330 3464
rect 22566 3228 22608 3464
rect 22288 1678 22608 3228
rect 22288 1442 22330 1678
rect 22566 1442 22608 1678
rect 22288 -108 22608 1442
rect 22288 -344 22330 -108
rect 22566 -344 22608 -108
rect 22288 -1894 22608 -344
rect 25038 24214 25358 25764
rect 30618 26000 30938 26024
rect 30618 25764 30660 26000
rect 30896 25764 30938 26000
rect 25038 23978 25080 24214
rect 25316 23978 25358 24214
rect 25038 22428 25358 23978
rect 25038 22192 25080 22428
rect 25316 22192 25358 22428
rect 25038 20642 25358 22192
rect 25038 20406 25080 20642
rect 25316 20406 25358 20642
rect 25038 18856 25358 20406
rect 25038 18620 25080 18856
rect 25316 18620 25358 18856
rect 25038 17070 25358 18620
rect 25038 16834 25080 17070
rect 25316 16834 25358 17070
rect 25038 15284 25358 16834
rect 25038 15048 25080 15284
rect 25316 15048 25358 15284
rect 25038 13498 25358 15048
rect 25038 13262 25080 13498
rect 25316 13262 25358 13498
rect 25038 11712 25358 13262
rect 25038 11476 25080 11712
rect 25316 11476 25358 11712
rect 25038 9926 25358 11476
rect 25038 9690 25080 9926
rect 25316 9690 25358 9926
rect 25038 8140 25358 9690
rect 25038 7904 25080 8140
rect 25316 7904 25358 8140
rect 25038 6354 25358 7904
rect 25038 6118 25080 6354
rect 25316 6118 25358 6354
rect 25038 4568 25358 6118
rect 25038 4332 25080 4568
rect 25316 4332 25358 4568
rect 25038 2782 25358 4332
rect 25038 2546 25080 2782
rect 25316 2546 25358 2782
rect 25038 996 25358 2546
rect 25038 760 25080 996
rect 25316 760 25358 996
rect 25038 -790 25358 760
rect 25038 -1026 25080 -790
rect 25316 -1026 25358 -790
rect 25038 -1894 25358 -1026
rect 27868 24896 28188 25696
rect 27868 24660 27910 24896
rect 28146 24660 28188 24896
rect 27868 23110 28188 24660
rect 27868 22874 27910 23110
rect 28146 22874 28188 23110
rect 27868 21324 28188 22874
rect 27868 21088 27910 21324
rect 28146 21088 28188 21324
rect 27868 19538 28188 21088
rect 27868 19302 27910 19538
rect 28146 19302 28188 19538
rect 27868 17752 28188 19302
rect 27868 17516 27910 17752
rect 28146 17516 28188 17752
rect 27868 15966 28188 17516
rect 27868 15730 27910 15966
rect 28146 15730 28188 15966
rect 27868 14180 28188 15730
rect 27868 13944 27910 14180
rect 28146 13944 28188 14180
rect 27868 12394 28188 13944
rect 27868 12158 27910 12394
rect 28146 12158 28188 12394
rect 27868 10608 28188 12158
rect 27868 10372 27910 10608
rect 28146 10372 28188 10608
rect 27868 8822 28188 10372
rect 27868 8586 27910 8822
rect 28146 8586 28188 8822
rect 27868 7036 28188 8586
rect 27868 6800 27910 7036
rect 28146 6800 28188 7036
rect 27868 5250 28188 6800
rect 27868 5014 27910 5250
rect 28146 5014 28188 5250
rect 27868 3464 28188 5014
rect 27868 3228 27910 3464
rect 28146 3228 28188 3464
rect 27868 1678 28188 3228
rect 27868 1442 27910 1678
rect 28146 1442 28188 1678
rect 27868 -108 28188 1442
rect 27868 -344 27910 -108
rect 28146 -344 28188 -108
rect 27868 -1894 28188 -344
rect 30618 24214 30938 25764
rect 36198 26000 36518 26024
rect 36198 25764 36240 26000
rect 36476 25764 36518 26000
rect 30618 23978 30660 24214
rect 30896 23978 30938 24214
rect 30618 22428 30938 23978
rect 30618 22192 30660 22428
rect 30896 22192 30938 22428
rect 30618 20642 30938 22192
rect 30618 20406 30660 20642
rect 30896 20406 30938 20642
rect 30618 18856 30938 20406
rect 30618 18620 30660 18856
rect 30896 18620 30938 18856
rect 30618 17070 30938 18620
rect 30618 16834 30660 17070
rect 30896 16834 30938 17070
rect 30618 15284 30938 16834
rect 30618 15048 30660 15284
rect 30896 15048 30938 15284
rect 30618 13498 30938 15048
rect 30618 13262 30660 13498
rect 30896 13262 30938 13498
rect 30618 11712 30938 13262
rect 30618 11476 30660 11712
rect 30896 11476 30938 11712
rect 30618 9926 30938 11476
rect 30618 9690 30660 9926
rect 30896 9690 30938 9926
rect 30618 8140 30938 9690
rect 30618 7904 30660 8140
rect 30896 7904 30938 8140
rect 30618 6354 30938 7904
rect 30618 6118 30660 6354
rect 30896 6118 30938 6354
rect 30618 4568 30938 6118
rect 30618 4332 30660 4568
rect 30896 4332 30938 4568
rect 30618 2782 30938 4332
rect 30618 2546 30660 2782
rect 30896 2546 30938 2782
rect 30618 996 30938 2546
rect 30618 760 30660 996
rect 30896 760 30938 996
rect 30618 -790 30938 760
rect 30618 -1026 30660 -790
rect 30896 -1026 30938 -790
rect 30618 -1894 30938 -1026
rect 33448 24896 33768 25696
rect 33448 24660 33490 24896
rect 33726 24660 33768 24896
rect 33448 24555 33768 24660
rect 33448 24319 33490 24555
rect 33726 24319 33768 24555
rect 33448 23110 33768 24319
rect 33448 22874 33490 23110
rect 33726 22874 33768 23110
rect 33448 21324 33768 22874
rect 33448 21088 33490 21324
rect 33726 21088 33768 21324
rect 33448 19538 33768 21088
rect 33448 19302 33490 19538
rect 33726 19302 33768 19538
rect 33448 17752 33768 19302
rect 33448 17516 33490 17752
rect 33726 17516 33768 17752
rect 33448 15966 33768 17516
rect 33448 15730 33490 15966
rect 33726 15730 33768 15966
rect 33448 14180 33768 15730
rect 33448 13944 33490 14180
rect 33726 13944 33768 14180
rect 33448 12394 33768 13944
rect 33448 12158 33490 12394
rect 33726 12158 33768 12394
rect 33448 10608 33768 12158
rect 33448 10372 33490 10608
rect 33726 10372 33768 10608
rect 33448 10267 33768 10372
rect 33448 10031 33490 10267
rect 33726 10031 33768 10267
rect 33448 8822 33768 10031
rect 33448 8586 33490 8822
rect 33726 8586 33768 8822
rect 33448 7036 33768 8586
rect 33448 6800 33490 7036
rect 33726 6800 33768 7036
rect 33448 5250 33768 6800
rect 33448 5014 33490 5250
rect 33726 5014 33768 5250
rect 33448 3464 33768 5014
rect 33448 3228 33490 3464
rect 33726 3228 33768 3464
rect 33448 1678 33768 3228
rect 33448 1442 33490 1678
rect 33726 1442 33768 1678
rect 33448 -108 33768 1442
rect 33448 -344 33490 -108
rect 33726 -344 33768 -108
rect 33448 -1894 33768 -344
rect 36198 24214 36518 25764
rect 41778 26000 42098 26024
rect 41778 25764 41820 26000
rect 42056 25764 42098 26000
rect 36198 23978 36240 24214
rect 36476 23978 36518 24214
rect 36198 22428 36518 23978
rect 36198 22192 36240 22428
rect 36476 22192 36518 22428
rect 36198 20642 36518 22192
rect 36198 20406 36240 20642
rect 36476 20406 36518 20642
rect 36198 18856 36518 20406
rect 36198 18620 36240 18856
rect 36476 18620 36518 18856
rect 36198 17070 36518 18620
rect 36198 16834 36240 17070
rect 36476 16834 36518 17070
rect 36198 15284 36518 16834
rect 36198 15048 36240 15284
rect 36476 15048 36518 15284
rect 36198 13498 36518 15048
rect 36198 13262 36240 13498
rect 36476 13262 36518 13498
rect 36198 11712 36518 13262
rect 36198 11476 36240 11712
rect 36476 11476 36518 11712
rect 36198 9926 36518 11476
rect 36198 9690 36240 9926
rect 36476 9690 36518 9926
rect 36198 8140 36518 9690
rect 36198 7904 36240 8140
rect 36476 7904 36518 8140
rect 36198 6354 36518 7904
rect 36198 6118 36240 6354
rect 36476 6118 36518 6354
rect 36198 4568 36518 6118
rect 36198 4332 36240 4568
rect 36476 4332 36518 4568
rect 36198 2782 36518 4332
rect 36198 2546 36240 2782
rect 36476 2546 36518 2782
rect 36198 996 36518 2546
rect 36198 760 36240 996
rect 36476 760 36518 996
rect 36198 -790 36518 760
rect 36198 -1026 36240 -790
rect 36476 -1026 36518 -790
rect 36198 -1894 36518 -1026
rect 39028 24896 39348 25696
rect 39028 24660 39070 24896
rect 39306 24660 39348 24896
rect 39028 23110 39348 24660
rect 39028 22874 39070 23110
rect 39306 22874 39348 23110
rect 39028 21324 39348 22874
rect 39028 21088 39070 21324
rect 39306 21088 39348 21324
rect 39028 19538 39348 21088
rect 39028 19302 39070 19538
rect 39306 19302 39348 19538
rect 39028 17752 39348 19302
rect 39028 17516 39070 17752
rect 39306 17516 39348 17752
rect 39028 15966 39348 17516
rect 39028 15730 39070 15966
rect 39306 15730 39348 15966
rect 39028 14180 39348 15730
rect 39028 13944 39070 14180
rect 39306 13944 39348 14180
rect 39028 12394 39348 13944
rect 39028 12158 39070 12394
rect 39306 12158 39348 12394
rect 39028 10608 39348 12158
rect 39028 10372 39070 10608
rect 39306 10372 39348 10608
rect 39028 8822 39348 10372
rect 39028 8586 39070 8822
rect 39306 8586 39348 8822
rect 39028 7036 39348 8586
rect 39028 6800 39070 7036
rect 39306 6800 39348 7036
rect 39028 5250 39348 6800
rect 39028 5014 39070 5250
rect 39306 5014 39348 5250
rect 39028 3464 39348 5014
rect 39028 3228 39070 3464
rect 39306 3228 39348 3464
rect 39028 1678 39348 3228
rect 39028 1442 39070 1678
rect 39306 1442 39348 1678
rect 39028 -108 39348 1442
rect 39028 -344 39070 -108
rect 39306 -344 39348 -108
rect 39028 -1894 39348 -344
rect 41778 24214 42098 25764
rect 47358 26000 47678 26024
rect 47358 25764 47400 26000
rect 47636 25764 47678 26000
rect 41778 23978 41820 24214
rect 42056 23978 42098 24214
rect 41778 22428 42098 23978
rect 41778 22192 41820 22428
rect 42056 22192 42098 22428
rect 41778 20642 42098 22192
rect 41778 20406 41820 20642
rect 42056 20406 42098 20642
rect 41778 18856 42098 20406
rect 41778 18620 41820 18856
rect 42056 18620 42098 18856
rect 41778 17070 42098 18620
rect 41778 16834 41820 17070
rect 42056 16834 42098 17070
rect 41778 15284 42098 16834
rect 41778 15048 41820 15284
rect 42056 15048 42098 15284
rect 41778 13498 42098 15048
rect 41778 13262 41820 13498
rect 42056 13262 42098 13498
rect 41778 11712 42098 13262
rect 41778 11476 41820 11712
rect 42056 11476 42098 11712
rect 41778 9926 42098 11476
rect 41778 9690 41820 9926
rect 42056 9690 42098 9926
rect 41778 8140 42098 9690
rect 41778 7904 41820 8140
rect 42056 7904 42098 8140
rect 41778 6354 42098 7904
rect 41778 6118 41820 6354
rect 42056 6118 42098 6354
rect 41778 4568 42098 6118
rect 41778 4332 41820 4568
rect 42056 4332 42098 4568
rect 41778 2782 42098 4332
rect 41778 2546 41820 2782
rect 42056 2546 42098 2782
rect 41778 996 42098 2546
rect 41778 760 41820 996
rect 42056 760 42098 996
rect 41778 -790 42098 760
rect 41778 -1026 41820 -790
rect 42056 -1026 42098 -790
rect 41778 -1894 42098 -1026
rect 44608 24896 44928 25696
rect 44608 24660 44650 24896
rect 44886 24660 44928 24896
rect 44608 23110 44928 24660
rect 44608 22874 44650 23110
rect 44886 22874 44928 23110
rect 44608 21324 44928 22874
rect 44608 21088 44650 21324
rect 44886 21088 44928 21324
rect 44608 19538 44928 21088
rect 44608 19302 44650 19538
rect 44886 19302 44928 19538
rect 44608 17752 44928 19302
rect 44608 17516 44650 17752
rect 44886 17516 44928 17752
rect 44608 15966 44928 17516
rect 44608 15730 44650 15966
rect 44886 15730 44928 15966
rect 44608 14180 44928 15730
rect 44608 13944 44650 14180
rect 44886 13944 44928 14180
rect 44608 12394 44928 13944
rect 44608 12158 44650 12394
rect 44886 12158 44928 12394
rect 44608 10608 44928 12158
rect 44608 10372 44650 10608
rect 44886 10372 44928 10608
rect 44608 8822 44928 10372
rect 44608 8586 44650 8822
rect 44886 8586 44928 8822
rect 44608 7036 44928 8586
rect 44608 6800 44650 7036
rect 44886 6800 44928 7036
rect 44608 5250 44928 6800
rect 44608 5014 44650 5250
rect 44886 5014 44928 5250
rect 44608 3464 44928 5014
rect 44608 3228 44650 3464
rect 44886 3228 44928 3464
rect 44608 1678 44928 3228
rect 44608 1442 44650 1678
rect 44886 1442 44928 1678
rect 44608 -108 44928 1442
rect 44608 -344 44650 -108
rect 44886 -344 44928 -108
rect 44608 -1894 44928 -344
rect 47358 24214 47678 25764
rect 52938 26000 53258 26024
rect 52938 25764 52980 26000
rect 53216 25764 53258 26000
rect 47358 23978 47400 24214
rect 47636 23978 47678 24214
rect 47358 22428 47678 23978
rect 47358 22192 47400 22428
rect 47636 22192 47678 22428
rect 47358 20642 47678 22192
rect 47358 20406 47400 20642
rect 47636 20406 47678 20642
rect 47358 18856 47678 20406
rect 47358 18620 47400 18856
rect 47636 18620 47678 18856
rect 47358 17070 47678 18620
rect 47358 16834 47400 17070
rect 47636 16834 47678 17070
rect 47358 15284 47678 16834
rect 47358 15048 47400 15284
rect 47636 15048 47678 15284
rect 47358 13498 47678 15048
rect 47358 13262 47400 13498
rect 47636 13262 47678 13498
rect 47358 11712 47678 13262
rect 47358 11476 47400 11712
rect 47636 11476 47678 11712
rect 47358 9926 47678 11476
rect 47358 9690 47400 9926
rect 47636 9690 47678 9926
rect 47358 8140 47678 9690
rect 47358 7904 47400 8140
rect 47636 7904 47678 8140
rect 47358 6354 47678 7904
rect 47358 6118 47400 6354
rect 47636 6118 47678 6354
rect 47358 4568 47678 6118
rect 47358 4332 47400 4568
rect 47636 4332 47678 4568
rect 47358 2782 47678 4332
rect 47358 2546 47400 2782
rect 47636 2546 47678 2782
rect 47358 996 47678 2546
rect 47358 760 47400 996
rect 47636 760 47678 996
rect 47358 -790 47678 760
rect 47358 -1026 47400 -790
rect 47636 -1026 47678 -790
rect 47358 -1894 47678 -1026
rect 50188 24896 50508 25696
rect 50188 24660 50230 24896
rect 50466 24660 50508 24896
rect 50188 23110 50508 24660
rect 50188 22874 50230 23110
rect 50466 22874 50508 23110
rect 50188 21324 50508 22874
rect 50188 21088 50230 21324
rect 50466 21088 50508 21324
rect 50188 19538 50508 21088
rect 50188 19302 50230 19538
rect 50466 19302 50508 19538
rect 50188 17752 50508 19302
rect 50188 17516 50230 17752
rect 50466 17516 50508 17752
rect 50188 15966 50508 17516
rect 50188 15730 50230 15966
rect 50466 15730 50508 15966
rect 50188 14180 50508 15730
rect 50188 13944 50230 14180
rect 50466 13944 50508 14180
rect 50188 12394 50508 13944
rect 50188 12158 50230 12394
rect 50466 12158 50508 12394
rect 50188 10608 50508 12158
rect 50188 10372 50230 10608
rect 50466 10372 50508 10608
rect 50188 8822 50508 10372
rect 50188 8586 50230 8822
rect 50466 8586 50508 8822
rect 50188 7036 50508 8586
rect 50188 6800 50230 7036
rect 50466 6800 50508 7036
rect 50188 5250 50508 6800
rect 50188 5014 50230 5250
rect 50466 5014 50508 5250
rect 50188 3464 50508 5014
rect 50188 3228 50230 3464
rect 50466 3228 50508 3464
rect 50188 1678 50508 3228
rect 50188 1442 50230 1678
rect 50466 1442 50508 1678
rect 50188 -108 50508 1442
rect 50188 -344 50230 -108
rect 50466 -344 50508 -108
rect 50188 -1894 50508 -344
rect 52938 24214 53258 25764
rect 52938 23978 52980 24214
rect 53216 23978 53258 24214
rect 52938 22428 53258 23978
rect 52938 22192 52980 22428
rect 53216 22192 53258 22428
rect 52938 20642 53258 22192
rect 52938 20406 52980 20642
rect 53216 20406 53258 20642
rect 52938 18856 53258 20406
rect 52938 18620 52980 18856
rect 53216 18620 53258 18856
rect 52938 17070 53258 18620
rect 52938 16834 52980 17070
rect 53216 16834 53258 17070
rect 52938 15284 53258 16834
rect 52938 15048 52980 15284
rect 53216 15048 53258 15284
rect 52938 13498 53258 15048
rect 52938 13262 52980 13498
rect 53216 13262 53258 13498
rect 52938 11712 53258 13262
rect 52938 11476 52980 11712
rect 53216 11476 53258 11712
rect 52938 9926 53258 11476
rect 52938 9690 52980 9926
rect 53216 9690 53258 9926
rect 52938 8140 53258 9690
rect 52938 7904 52980 8140
rect 53216 7904 53258 8140
rect 52938 6354 53258 7904
rect 52938 6118 52980 6354
rect 53216 6118 53258 6354
rect 52938 4568 53258 6118
rect 52938 4332 52980 4568
rect 53216 4332 53258 4568
rect 52938 2782 53258 4332
rect 52938 2546 52980 2782
rect 53216 2546 53258 2782
rect 52938 996 53258 2546
rect 52938 760 52980 996
rect 53216 760 53258 996
rect 52938 -790 53258 760
rect 52938 -1026 52980 -790
rect 53216 -1026 53258 -790
rect 52938 -1894 53258 -1026
rect 16708 -2130 16750 -1894
rect 16986 -2130 17028 -1894
rect 16708 -2154 17028 -2130
rect 22288 -2130 22330 -1894
rect 22566 -2130 22608 -1894
rect 22288 -2154 22608 -2130
rect 27868 -2130 27910 -1894
rect 28146 -2130 28188 -1894
rect 27868 -2154 28188 -2130
rect 33448 -2130 33490 -1894
rect 33726 -2130 33768 -1894
rect 33448 -2154 33768 -2130
rect 39028 -2130 39070 -1894
rect 39306 -2130 39348 -1894
rect 39028 -2154 39348 -2130
rect 44608 -2130 44650 -1894
rect 44886 -2130 44928 -1894
rect 44608 -2154 44928 -2130
rect 50188 -2130 50230 -1894
rect 50466 -2130 50508 -1894
rect 50188 -2154 50508 -2130
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_0
timestamp 1755519375
transform 1 0 -8573 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_1
timestamp 1755519375
transform 1 0 -8573 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_2
timestamp 1755519375
transform 1 0 -8573 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_3
timestamp 1755519375
transform 1 0 -8573 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_4
timestamp 1755519375
transform 1 0 -8573 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_5
timestamp 1755519375
transform 1 0 -8573 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_6
timestamp 1755519375
transform 1 0 -8573 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_7
timestamp 1755519375
transform 1 0 -8573 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_8
timestamp 1755519375
transform 1 0 -8573 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_9
timestamp 1755519375
transform 1 0 -8573 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_10
timestamp 1755519375
transform 1 0 -8573 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_11
timestamp 1755519375
transform 1 0 -8573 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_12
timestamp 1755519375
transform 1 0 -8573 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_13
timestamp 1755519375
transform 1 0 -8573 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_14
timestamp 1755519375
transform 1 0 -8573 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_15
timestamp 1755519375
transform 1 0 -30893 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_16
timestamp 1755519375
transform -1 0 19349 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_17
timestamp 1755519375
transform 1 0 2587 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_18
timestamp 1755519375
transform 1 0 2587 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_19
timestamp 1755519375
transform 1 0 2587 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_20
timestamp 1755519375
transform 1 0 2587 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_21
timestamp 1755519375
transform 1 0 2587 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_22
timestamp 1755519375
transform 1 0 2587 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_23
timestamp 1755519375
transform 1 0 2587 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_24
timestamp 1755519375
transform 1 0 2587 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_25
timestamp 1755519375
transform 1 0 2587 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_26
timestamp 1755519375
transform 1 0 2587 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_27
timestamp 1755519375
transform 1 0 2587 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_28
timestamp 1755519375
transform 1 0 2587 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_29
timestamp 1755519375
transform 1 0 2587 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_30
timestamp 1755519375
transform 1 0 2587 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_31
timestamp 1755519375
transform 1 0 2587 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_32
timestamp 1755519375
transform 1 0 -30893 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_33
timestamp 1755519375
transform 1 0 -2993 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_34
timestamp 1755519375
transform 1 0 -2993 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_35
timestamp 1755519375
transform 1 0 -2993 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_36
timestamp 1755519375
transform 1 0 -2993 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_37
timestamp 1755519375
transform 1 0 -2993 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_38
timestamp 1755519375
transform 1 0 -2993 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_39
timestamp 1755519375
transform 1 0 -2993 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_40
timestamp 1755519375
transform 1 0 -2993 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_41
timestamp 1755519375
transform 1 0 -2993 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_42
timestamp 1755519375
transform 1 0 -2993 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_43
timestamp 1755519375
transform 1 0 -2993 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_44
timestamp 1755519375
transform 1 0 -2993 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_45
timestamp 1755519375
transform 1 0 -2993 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_46
timestamp 1755519375
transform 1 0 -2993 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_47
timestamp 1755519375
transform 1 0 -2993 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_48
timestamp 1755519375
transform 1 0 -36473 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_49
timestamp 1755519375
transform 1 0 -14153 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_50
timestamp 1755519375
transform 1 0 -14153 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_51
timestamp 1755519375
transform 1 0 -36473 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_52
timestamp 1755519375
transform 1 0 -14153 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_53
timestamp 1755519375
transform 1 0 -14153 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_54
timestamp 1755519375
transform 1 0 -14153 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_55
timestamp 1755519375
transform 1 0 -14153 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_56
timestamp 1755519375
transform 1 0 -14153 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_57
timestamp 1755519375
transform 1 0 -14153 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_58
timestamp 1755519375
transform 1 0 -14153 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_59
timestamp 1755519375
transform 1 0 -14153 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_60
timestamp 1755519375
transform 1 0 -14153 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_61
timestamp 1755519375
transform 1 0 -14153 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_62
timestamp 1755519375
transform 1 0 -14153 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_63
timestamp 1755519375
transform 1 0 -14153 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_64
timestamp 1755519375
transform 1 0 -14153 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_65
timestamp 1755519375
transform 1 0 2587 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_66
timestamp 1755519375
transform 1 0 -2993 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_67
timestamp 1755519375
transform 1 0 -8573 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_68
timestamp 1755519375
transform 1 0 -14153 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_69
timestamp 1755519375
transform 1 0 -30893 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_70
timestamp 1755519375
transform 1 0 -30893 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_71
timestamp 1755519375
transform 1 0 -36473 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_72
timestamp 1755519375
transform 1 0 -36473 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_73
timestamp 1755519375
transform 1 0 -30893 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_74
timestamp 1755519375
transform 1 0 -30893 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_75
timestamp 1755519375
transform 1 0 -36473 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_76
timestamp 1755519375
transform 1 0 -36473 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_77
timestamp 1755519375
transform 1 0 -30893 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_78
timestamp 1755519375
transform 1 0 -30893 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_79
timestamp 1755519375
transform 1 0 -36473 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_80
timestamp 1755519375
transform 1 0 -36473 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_81
timestamp 1755519375
transform 1 0 -30893 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_82
timestamp 1755519375
transform 1 0 -30893 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_83
timestamp 1755519375
transform 1 0 -36473 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_84
timestamp 1755519375
transform 1 0 -36473 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_85
timestamp 1755519375
transform 1 0 -30893 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_86
timestamp 1755519375
transform 1 0 -30893 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_87
timestamp 1755519375
transform 1 0 -36473 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_88
timestamp 1755519375
transform 1 0 -36473 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_89
timestamp 1755519375
transform 1 0 -30893 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_90
timestamp 1755519375
transform 1 0 -30893 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_91
timestamp 1755519375
transform 1 0 -36473 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_92
timestamp 1755519375
transform 1 0 -36473 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_93
timestamp 1755519375
transform 1 0 -30893 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_94
timestamp 1755519375
transform 1 0 -30893 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_95
timestamp 1755519375
transform 1 0 -36473 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_96
timestamp 1755519375
transform 1 0 -36473 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_97
timestamp 1755519375
transform 1 0 -25313 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_98
timestamp 1755519375
transform 1 0 -25313 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_99
timestamp 1755519375
transform 1 0 -25313 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_100
timestamp 1755519375
transform 1 0 -25313 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_101
timestamp 1755519375
transform 1 0 -19733 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_102
timestamp 1755519375
transform 1 0 -19733 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_103
timestamp 1755519375
transform 1 0 -19733 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_104
timestamp 1755519375
transform 1 0 -19733 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_105
timestamp 1755519375
transform 1 0 -25313 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_106
timestamp 1755519375
transform 1 0 -25313 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_107
timestamp 1755519375
transform 1 0 -25313 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_108
timestamp 1755519375
transform 1 0 -25313 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_109
timestamp 1755519375
transform 1 0 -19733 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_110
timestamp 1755519375
transform 1 0 -19733 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_111
timestamp 1755519375
transform 1 0 -19733 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_112
timestamp 1755519375
transform 1 0 -19733 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_113
timestamp 1755519375
transform 1 0 -25313 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_114
timestamp 1755519375
transform 1 0 -25313 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_115
timestamp 1755519375
transform 1 0 -25313 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_116
timestamp 1755519375
transform 1 0 -19733 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_117
timestamp 1755519375
transform 1 0 -19733 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_118
timestamp 1755519375
transform 1 0 -19733 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_119
timestamp 1755519375
transform 1 0 -25313 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_120
timestamp 1755519375
transform 1 0 -25313 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_121
timestamp 1755519375
transform 1 0 -25313 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_122
timestamp 1755519375
transform 1 0 -25313 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_123
timestamp 1755519375
transform 1 0 -19733 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_124
timestamp 1755519375
transform 1 0 -19733 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_125
timestamp 1755519375
transform 1 0 -19733 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_126
timestamp 1755519375
transform 1 0 -19733 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_127
timestamp 1755519375
transform 1 0 -25313 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_128
timestamp 1755519375
transform 1 0 -19733 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_129
timestamp 1755519375
transform -1 0 52829 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_130
timestamp 1755519375
transform -1 0 47249 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_131
timestamp 1755519375
transform -1 0 41669 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_132
timestamp 1755519375
transform -1 0 36089 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_133
timestamp 1755519375
transform -1 0 30509 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_134
timestamp 1755519375
transform -1 0 24929 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_135
timestamp 1755519375
transform -1 0 19349 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_137
timestamp 1755519375
transform -1 0 52829 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_138
timestamp 1755519375
transform -1 0 47249 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_139
timestamp 1755519375
transform -1 0 41669 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_140
timestamp 1755519375
transform -1 0 36089 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_141
timestamp 1755519375
transform -1 0 30509 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_142
timestamp 1755519375
transform -1 0 24929 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_143
timestamp 1755519375
transform -1 0 19349 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_144
timestamp 1755519375
transform -1 0 13769 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_145
timestamp 1755519375
transform -1 0 52829 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_146
timestamp 1755519375
transform -1 0 47249 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_147
timestamp 1755519375
transform -1 0 41669 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_148
timestamp 1755519375
transform -1 0 36089 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_149
timestamp 1755519375
transform -1 0 30509 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_150
timestamp 1755519375
transform -1 0 24929 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_152
timestamp 1755519375
transform -1 0 13769 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_153
timestamp 1755519375
transform -1 0 52829 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_154
timestamp 1755519375
transform -1 0 47249 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_155
timestamp 1755519375
transform -1 0 41669 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_156
timestamp 1755519375
transform -1 0 36089 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_157
timestamp 1755519375
transform -1 0 30509 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_158
timestamp 1755519375
transform -1 0 24929 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_159
timestamp 1755519375
transform -1 0 19349 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_160
timestamp 1755519375
transform -1 0 13769 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_161
timestamp 1755519375
transform -1 0 52829 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_162
timestamp 1755519375
transform -1 0 47249 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_163
timestamp 1755519375
transform -1 0 41669 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_164
timestamp 1755519375
transform -1 0 36089 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_165
timestamp 1755519375
transform -1 0 30509 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_166
timestamp 1755519375
transform -1 0 24929 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_167
timestamp 1755519375
transform -1 0 19349 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_168
timestamp 1755519375
transform -1 0 13769 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_169
timestamp 1755519375
transform -1 0 52829 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_170
timestamp 1755519375
transform -1 0 47249 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_171
timestamp 1755519375
transform -1 0 41669 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_172
timestamp 1755519375
transform -1 0 36089 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_173
timestamp 1755519375
transform -1 0 30509 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_174
timestamp 1755519375
transform -1 0 24929 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_175
timestamp 1755519375
transform -1 0 19349 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_176
timestamp 1755519375
transform -1 0 13769 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_177
timestamp 1755519375
transform -1 0 52829 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_178
timestamp 1755519375
transform -1 0 47249 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_179
timestamp 1755519375
transform -1 0 41669 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_180
timestamp 1755519375
transform -1 0 36089 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_181
timestamp 1755519375
transform -1 0 30509 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_182
timestamp 1755519375
transform -1 0 24929 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_183
timestamp 1755519375
transform -1 0 19349 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_184
timestamp 1755519375
transform -1 0 13769 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_185
timestamp 1755519375
transform -1 0 52829 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_186
timestamp 1755519375
transform -1 0 47249 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_187
timestamp 1755519375
transform -1 0 41669 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_188
timestamp 1755519375
transform -1 0 36089 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_189
timestamp 1755519375
transform -1 0 30509 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_190
timestamp 1755519375
transform -1 0 24929 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_191
timestamp 1755519375
transform -1 0 19349 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_192
timestamp 1755519375
transform -1 0 13769 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_193
timestamp 1755519375
transform -1 0 52829 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_194
timestamp 1755519375
transform -1 0 47249 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_195
timestamp 1755519375
transform -1 0 41669 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_196
timestamp 1755519375
transform -1 0 36089 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_197
timestamp 1755519375
transform -1 0 30509 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_198
timestamp 1755519375
transform -1 0 24929 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_199
timestamp 1755519375
transform -1 0 19349 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_200
timestamp 1755519375
transform -1 0 13769 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_201
timestamp 1755519375
transform -1 0 52829 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_202
timestamp 1755519375
transform -1 0 47249 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_203
timestamp 1755519375
transform -1 0 41669 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_204
timestamp 1755519375
transform -1 0 36089 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_205
timestamp 1755519375
transform -1 0 30509 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_206
timestamp 1755519375
transform -1 0 24929 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_207
timestamp 1755519375
transform -1 0 19349 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_208
timestamp 1755519375
transform -1 0 13769 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_209
timestamp 1755519375
transform -1 0 52829 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_210
timestamp 1755519375
transform -1 0 47249 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_211
timestamp 1755519375
transform -1 0 41669 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_212
timestamp 1755519375
transform -1 0 36089 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_213
timestamp 1755519375
transform -1 0 30509 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_214
timestamp 1755519375
transform -1 0 24929 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_215
timestamp 1755519375
transform -1 0 19349 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_216
timestamp 1755519375
transform -1 0 13769 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_217
timestamp 1755519375
transform -1 0 52829 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_218
timestamp 1755519375
transform -1 0 47249 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_219
timestamp 1755519375
transform -1 0 41669 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_220
timestamp 1755519375
transform -1 0 36089 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_221
timestamp 1755519375
transform -1 0 30509 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_222
timestamp 1755519375
transform -1 0 24929 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_223
timestamp 1755519375
transform -1 0 19349 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_224
timestamp 1755519375
transform -1 0 13769 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_225
timestamp 1755519375
transform -1 0 52829 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_226
timestamp 1755519375
transform -1 0 47249 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_227
timestamp 1755519375
transform -1 0 41669 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_228
timestamp 1755519375
transform -1 0 36089 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_229
timestamp 1755519375
transform -1 0 30509 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_230
timestamp 1755519375
transform -1 0 24929 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_231
timestamp 1755519375
transform -1 0 19349 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_232
timestamp 1755519375
transform -1 0 13769 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_233
timestamp 1755519375
transform -1 0 52829 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_234
timestamp 1755519375
transform -1 0 47249 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_235
timestamp 1755519375
transform -1 0 41669 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_236
timestamp 1755519375
transform -1 0 36089 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_237
timestamp 1755519375
transform -1 0 30509 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_238
timestamp 1755519375
transform -1 0 24929 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_239
timestamp 1755519375
transform -1 0 19349 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_240
timestamp 1755519375
transform -1 0 13769 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_241
timestamp 1755519375
transform -1 0 52829 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_242
timestamp 1755519375
transform -1 0 47249 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_243
timestamp 1755519375
transform -1 0 41669 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_244
timestamp 1755519375
transform -1 0 36089 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_245
timestamp 1755519375
transform -1 0 30509 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_246
timestamp 1755519375
transform -1 0 24929 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_247
timestamp 1755519375
transform -1 0 19349 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_248
timestamp 1755519375
transform -1 0 13769 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_249
timestamp 1755519375
transform -1 0 13769 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_250
timestamp 1755519375
transform -1 0 19349 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_251
timestamp 1755519375
transform -1 0 24929 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_252
timestamp 1755519375
transform -1 0 30509 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_253
timestamp 1755519375
transform -1 0 36089 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_254
timestamp 1755519375
transform -1 0 41669 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_255
timestamp 1755519375
transform -1 0 47249 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_256
timestamp 1755519375
transform -1 0 52829 0 1 25296
box -2619 -281 2641 281
use switch  switch_0
timestamp 1753542193
transform 1 0 5896 0 -1 3064
box 1296 -1584 3268 244
use switch  switch_1
timestamp 1753542193
transform 1 0 5896 0 1 -954
box 1296 -1584 3268 244
use switch  switch_2
timestamp 1753542193
transform 1 0 5896 0 -1 -512
box 1296 -1584 3268 244
use switch  switch_5
timestamp 1753542193
transform 1 0 5896 0 -1 6636
box 1296 -1584 3268 244
use switch  switch_6
timestamp 1753542193
transform 1 0 5896 0 -1 17352
box 1296 -1584 3268 244
use switch  switch_7
timestamp 1753542193
transform 1 0 5896 0 -1 13780
box 1296 -1584 3268 244
use switch  switch_8
timestamp 1753542193
transform 1 0 5896 0 -1 24055
box 1296 -1584 3268 244
use switch  switch_9
timestamp 1753542193
transform 1 0 5896 0 -1 20924
box 1296 -1584 3268 244
<< labels >>
flabel metal1 7100 -2538 7146 25639 0 FreeSans 160 90 0 0 VDD
port 9 nsew
flabel space 11128 11 16388 573 0 FreeSans 4800 180 0 0 1
flabel space 11128 1797 16388 4145 0 FreeSans 16000 180 0 0 2
flabel space 11128 5369 16388 11289 0 FreeSans 16000 180 0 0 3
flabel space 11128 12513 16388 25577 0 FreeSans 16000 180 0 0 4
flabel space 16708 -1775 21968 25577 0 FreeSans 16000 180 0 0 5
flabel space 22288 -1775 33128 25577 0 FreeSans 16000 180 0 0 6
flabel space 33448 -1775 55448 25577 0 FreeSans 16000 180 0 0 7
flabel space -39092 -1775 -17092 25577 0 FreeSans 16000 0 0 0 7
flabel space -16772 -1775 -5932 25577 0 FreeSans 16000 0 0 0 6
flabel space -5612 -1775 -352 25577 0 FreeSans 16000 0 0 0 5
flabel space -32 12513 5228 25577 0 FreeSans 16000 0 0 0 4
flabel space -32 5369 5228 11289 0 FreeSans 16000 0 0 0 3
flabel space -32 1797 5228 4145 0 FreeSans 16000 0 0 0 2
flabel space -32 11 5228 573 0 FreeSans 4800 0 0 0 1
flabel space -32 -1775 5228 -1213 0 FreeSans 4800 0 0 0 0
flabel metal1 9210 -2538 9256 25639 0 FreeSans 160 90 0 0 GND
port 8 nsew
flabel metal5 52938 -1894 53258 26024 0 FreeSans 160 90 0 0 OUT
port 10 nsew
flabel metal1 8155 -1686 8815 -1640 0 FreeSans 160 0 0 0 b0
port 12 nsew
flabel metal1 8155 174 8815 220 0 FreeSans 160 0 0 0 b1
port 13 nsew
flabel metal1 8155 3750 8815 3796 0 FreeSans 160 0 0 0 b2
port 14 nsew
flabel metal1 8155 7322 8815 7368 0 FreeSans 160 0 0 0 b3
port 15 nsew
flabel metal1 8155 14466 8815 14512 0 FreeSans 160 0 0 0 b4
port 16 nsew
flabel metal1 8155 18038 8815 18084 0 FreeSans 160 0 0 0 b5
port 17 nsew
flabel metal1 8155 21610 8815 21656 0 FreeSans 160 0 0 0 b6
port 18 nsew
flabel metal1 8155 24741 8815 24787 0 FreeSans 160 0 0 0 b7
port 19 nsew
<< end >>
