** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-11_04-53-17/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.31764705875 8.5u 0.31764705875 8.500001u 0.319411764625 17.0u 0.319411764625 17.000001u 0.3211764705 25.5u
+ 0.3211764705 25.500001u 0.322941176375 34.0u 0.322941176375 34.000001u 0.32470588225 42.5u 0.32470588225 42.500001u 0.326470588125 51.0u
+ 0.326470588125 51.000001u 0.328235294 59.5u 0.328235294 59.500001u 0.33 68.0u 0.33 68.000001u 0.331764705875 76.5u 0.331764705875 76.500001u
+ 0.33352941175 85.0u 0.33352941175 85.000001u 0.335294117625 93.5u 0.335294117625 93.500001u 0.3370588235 102.0u 0.3370588235 102.000001u
+ 0.338823529375 110.5u 0.338823529375 110.500001u 0.34058823525 119.0u 0.34058823525 119.000001u 0.342352941125 127.5u 0.342352941125 127.500001u
+ 0.344117647 136.0u 0.344117647 136.000001u 0.345882352875 144.5u 0.345882352875 144.500001u 0.34764705875 153.0u 0.34764705875 153.000001u
+ 0.349411764625 161.5u 0.349411764625 161.500001u 0.3511764705 170.0u 0.3511764705 170.000001u 0.352941176375 178.5u 0.352941176375)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ff

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 178.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-11_04-53-17/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
