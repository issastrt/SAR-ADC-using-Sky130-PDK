magic
tech sky130A
magscale 1 2
timestamp 1753268444
<< nwell >>
rect 2023 -528 2065 354
rect 3953 -528 3995 354
<< locali >>
rect 2239 394 2551 400
rect 2239 360 2245 394
rect 2545 360 2551 394
rect 2239 242 2551 360
rect 2853 394 3165 400
rect 2853 360 2859 394
rect 3159 360 3165 394
rect 2853 242 3165 360
rect 3467 394 3779 400
rect 3467 360 3473 394
rect 3773 360 3779 394
rect 3467 242 3779 360
rect 2167 -1388 2623 -1300
rect 2167 -1422 2173 -1388
rect 2617 -1422 2623 -1388
rect 2167 -1428 2623 -1422
rect 2781 -1388 3237 -1300
rect 2781 -1422 2787 -1388
rect 3231 -1422 3237 -1388
rect 2781 -1428 3237 -1422
rect 3395 -1388 3851 -1300
rect 3395 -1422 3401 -1388
rect 3845 -1422 3851 -1388
rect 3395 -1428 3851 -1422
<< viali >>
rect 2245 360 2545 394
rect 2859 360 3159 394
rect 3473 360 3773 394
rect 2173 -1422 2617 -1388
rect 2787 -1422 3231 -1388
rect 3401 -1422 3845 -1388
<< metal1 >>
rect 2023 394 3995 400
rect 2023 360 2245 394
rect 2545 360 2859 394
rect 3159 360 3473 394
rect 3773 360 3995 394
rect 2023 354 3995 360
rect 2221 57 2267 354
rect 3293 57 3339 354
rect 2221 11 2317 57
rect 2473 11 2931 57
rect 3087 11 3545 57
rect 2876 -173 2940 -167
rect 2876 -225 2882 -173
rect 2934 -225 2940 -173
rect 2876 -231 2940 -225
rect 3692 -173 3756 -167
rect 3692 -225 3698 -173
rect 3750 -185 3756 -173
rect 3750 -225 3869 -185
rect 3692 -231 3869 -225
rect 2372 -804 2418 -272
rect 2986 -804 3032 -272
rect 3600 -804 3646 -272
rect 3823 -836 3869 -231
rect 3773 -882 3869 -836
rect 2148 -1124 2245 -1078
rect 2545 -1124 2859 -1078
rect 3159 -1124 3473 -1078
rect 2149 -1382 2195 -1124
rect 2023 -1388 3995 -1382
rect 2023 -1422 2173 -1388
rect 2617 -1422 2787 -1388
rect 3231 -1422 3401 -1388
rect 3845 -1422 3995 -1388
rect 2023 -1428 3995 -1422
<< via1 >>
rect 2882 -225 2934 -173
rect 3698 -225 3750 -173
<< metal2 >>
rect 2876 -173 2940 -167
rect 2876 -225 2882 -173
rect 2934 -176 2940 -173
rect 3692 -173 3756 -167
rect 3692 -176 3698 -173
rect 2934 -222 3698 -176
rect 2934 -225 2940 -222
rect 2876 -231 2940 -225
rect 3692 -225 3698 -222
rect 3750 -225 3756 -173
rect 3692 -231 3756 -225
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1 /foss/designs
timestamp 1753266908
transform 1 0 3623 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM2
timestamp 1753266908
transform 1 0 3009 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM3
timestamp 1753266908
transform 1 0 2395 0 1 -87
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4 /foss/designs
timestamp 1753266908
transform 1 0 3623 0 1 -980
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM5
timestamp 1753266908
transform 1 0 3009 0 1 -980
box -372 -402 372 402
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM6
timestamp 1753266908
transform 1 0 2395 0 1 -980
box -372 -402 372 402
<< labels >>
flabel metal1 2023 -1428 3995 -1382 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 2023 354 3995 400 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 2372 -804 2418 -272 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 2986 -804 3032 -272 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal1 3600 -804 3646 -272 0 FreeSans 160 0 0 0 C
port 4 nsew
flabel metal1 3823 -882 3869 -185 0 FreeSans 160 90 0 0 Vout
port 5 nsew
<< end >>
