** sch_path: /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_22-13-40/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.836470588125 8.5u 0.836470588125 8.500001u 0.838235294000 17u 0.838235294000 17.000001u 0.840000000000 25.5u
+ 0.840000000000 25.500001u 0.841764705875 34u 0.841764705875 34.000001u 0.843529411750 42.5u 0.843529411750 42.500001u 0.845294117625 51u
+ 0.845294117625 51.000001u 0.847058823500 59.5u 0.847058823500 59.500001u 0.848823529375 68u 0.848823529375 68.000001u 0.850588235250 76.5u
+ 0.850588235250 76.500001u 0.852352941125 85u 0.852352941125 85.000001u 0.854117647000 93.5u 0.854117647000 93.500001u 0.855882352875 102u
+ 0.855882352875 102.000001u 0.857647058750 110.5u 0.857647058750 110.500001u 0.859411764625 119u 0.859411764625 119.000001u 0.861176470500 127.5u
+ 0.861176470500 127.500001u 0.862941176375 136u 0.862941176375 136.000001u 0.864705882250 144.5u 0.864705882250 144.500001u 0.866470588125 153u
+ 0.866470588125 153.000001u 0.868235294000 161.5u 0.868235294000 161.500001u 0.870000000000 170u 0.870000000000 170.000001u 0.871764705875 178.5u
+ 0.871764705875 178.500001u 0.873529411750 187u 0.873529411750 187.000001u 0.875294117625 195.5u 0.875294117625 195.500001u 0.877058823500 204u
+ 0.877058823500 204.000001u 0.878823529375 212.5u 0.878823529375 212.500001u 0.880588235250 221u 0.880588235250 221.000001u 0.882352941125 229.5u
+ 0.882352941125 229.500001u 0.884117647000 238u 0.884117647000 238.000001u 0.885882352875 246.5u 0.885882352875 246.500001u 0.887647058750 255u
+ 0.887647058750 255.000001u 0.889411764625 263.5u 0.889411764625 263.500001u 0.891176470500 272u 0.891176470500 272.000001u 0.892941176375 280.5u
+ 0.892941176375 280.500001u 0.894705882250 289u 0.894705882250 289.000001u 0.896470588125 297.5u 0.896470588125 297.500001u 0.898235294000 306u
+ 0.898235294000 306.000001u 0.900000000000 314.5u 0.900000000000 314.500001u 0.901764705875 323u 0.901764705875 323.000001u 0.903529411750 331.5u
+ 0.903529411750 331.500001u 0.905294117625 340u 0.905294117625 340.000001u 0.907058823500 348.5u 0.907058823500 348.500001u 0.908823529375 357u
+ 0.908823529375 357.000001u 0.910588235250 365.5u 0.910588235250 365.500001u 0.912352941125 374u 0.912352941125 374.000001u 0.914117647000 382.5u
+ 0.914117647000 382.500001u 0.915882352875 391u 0.915882352875 391.000001u 0.917647058750 399.5u 0.917647058750 399.500001u 0.919411764625 408u
+ 0.919411764625 408.000001u 0.921176470500 416.5u 0.921176470500 416.500001u 0.922941176375 425u 0.922941176375 425.000001u 0.924705882250 433.5u
+ 0.924705882250 433.500001u 0.926470588125 442u 0.926470588125 442.000001u 0.928235294000 450.5u 0.928235294000 450.500001u 0.930000000000 459u
+ 0.930000000000 459.000001u 0.931764705875 467.5u 0.931764705875 467.500001u 0.933529411750 476u 0.933529411750 476.000001u 0.935294117625 484.5u
+ 0.935294117625 484.500001u 0.937058823500 493u 0.937058823500 493.000001u 0.938823529375 501.5u 0.938823529375 501.500001u 0.940588235250 510u
+ 0.940588235250 510.000001u 0.942352941125 518.5u 0.942352941125 518.500001u 0.944117647000 527u 0.944117647000 527.000001u 0.945882352875 535.5u
+ 0.945882352875 535.500001u 0.947647058750 544u 0.947647058750 544.000001u 0.949411764625 552.5u 0.949411764625 552.500001u 0.951176470500 561u
+ 0.951176470500 561.000001u 0.952941176375 569.5u 0.952941176375 569.500001u 0.954705882250 578u 0.954705882250 578.000001u 0.956470588125 586.5u
+ 0.956470588125 586.500001u 0.958235294000 595u 0.958235294000 595.000001u 0.960000000000 603.5u 0.960000000000 603.500001u 0.961764705875 612u
+ 0.961764705875 612.000001u 0.963529411750 620.5u 0.963529411750 620.500001u 0.965294117625 629u 0.965294117625 629.000001u 0.967058823500 637.5u
+ 0.967058823500 637.500001u 0.968823529375 646u 0.968823529375 646.000001u 0.970588235250 654.5u 0.970588235250 654.500001u 0.972352941125 663u
+ 0.972352941125 663.000001u 0.974117647000 671.5u 0.974117647000 671.500001u 0.975882352875 680u 0.975882352875)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/samantha/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 680u uic
  wrdata /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_22-13-40/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
