** sch_path: /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-10_11-35-26/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 1.658823529375 8.5u 1.658823529375 8.500001u 1.66058823525 17.0u 1.66058823525 17.000001u 1.662352941125 25.5u
+ 1.662352941125 25.500001u 1.664117647 34.0u 1.664117647 34.000001u 1.665882352875 42.5u 1.665882352875 42.500001u 1.66764705875 51.0u
+ 1.66764705875 51.000001u 1.669411764625 59.5u 1.669411764625 59.500001u 1.6711764705 68.0u 1.6711764705 68.000001u 1.672941176375 76.5u
+ 1.672941176375 76.500001u 1.67470588225 85.0u 1.67470588225 85.000001u 1.676470588125 93.5u 1.676470588125 93.500001u 1.678235294 102.0u
+ 1.678235294 102.000001u 1.68 110.5u 1.68 110.500001u 1.681764705875 119.0u 1.681764705875 119.000001u 1.68352941175 127.5u 1.68352941175
+ 127.500001u 1.685294117625 136.0u 1.685294117625 136.000001u 1.6870588235 144.5u 1.6870588235 144.500001u 1.688823529375 153.0u
+ 1.688823529375 153.000001u 1.69058823525 161.5u 1.69058823525 161.500001u 1.692352941125 170.0u 1.692352941125 170.000001u 1.694117647 178.5u
+ 1.694117647)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/madra/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 178.5u uic
  wrdata /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-10_11-35-26/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
