** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_04-35-14/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.0352941175 8.5u 0.0352941175 8.500001u 0.037058823375 17u 0.037058823375 17.000001u 0.03882352925 25.5u
+ 0.03882352925 25.500001u 0.040588235125 34u 0.040588235125 34.000001u 0.08470588225 42.5u 0.08470588225 42.500001u 0.086470588125 51u
+ 0.086470588125 51.000001u 0.088235294 59.5u 0.088235294 59.500001u 0.09 68u 0.09 68.000001u 0.148235294 76.5u 0.148235294 76.500001u 0.15 85u
+ 0.15 85.000001u 0.151764705875 93.5u 0.151764705875 93.500001u 0.15352941175 102u 0.15352941175 102.000001u 0.20470588225 110.5u
+ 0.20470588225 110.500001u 0.206470588125 119u 0.206470588125 119.000001u 0.208235294 127.5u 0.208235294 127.500001u 0.21 136u 0.21 136.000001u
+ 0.211764705875 144.5u 0.211764705875 144.500001u 0.2611764705 153u 0.2611764705 153.000001u 0.262941176375 161.5u 0.262941176375 161.500001u
+ 0.26470588225 170u 0.26470588225 170.000001u 0.266470588125 178.5u 0.266470588125 178.500001u 0.31764705875 187u 0.31764705875 187.000001u
+ 0.319411764625 195.5u 0.319411764625 195.500001u 0.3211764705 204u 0.3211764705 204.000001u 0.322941176375 212.5u 0.322941176375 212.500001u
+ 0.374117647 221u 0.374117647 221.000001u 0.375882352875 229.5u 0.375882352875 229.500001u 0.37764705875 238u 0.37764705875 238.000001u
+ 0.379411764625 246.5u 0.379411764625 246.500001u 0.43058823525 255u 0.43058823525 255.000001u 0.432352941125 263.5u 0.432352941125 263.500001u
+ 0.434117647 272u 0.434117647 272.000001u 0.435882352875 280.5u 0.435882352875)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=125
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 280.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_04-35-14/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
