magic
tech sky130A
magscale 1 2
timestamp 1757103913
<< nwell >>
rect -2163 -5014 -2089 -5000
rect 1781 -5014 1855 -5000
rect 5725 -5014 5799 -5000
rect 9669 -5014 9743 -5000
rect 13613 -5014 13687 -5000
rect 17557 -5014 17631 -5000
rect 21501 -5014 21575 -5000
<< pwell >>
rect -1873 -6736 -1799 -6722
rect 2071 -6736 2145 -6722
rect 6015 -6736 6089 -6722
rect 9959 -6736 10033 -6722
rect 13903 -6736 13977 -6722
rect 17847 -6736 17921 -6722
rect 21791 -6736 21865 -6722
<< metal1 >>
rect -6102 -4951 -6038 -4945
rect -6102 -4954 -6096 -4951
rect -6604 -5000 -6096 -4954
rect -6102 -5003 -6096 -5000
rect -6044 -4954 -6038 -4951
rect -2158 -4951 -2094 -4945
rect -2158 -4954 -2152 -4951
rect -6044 -5000 -2152 -4954
rect -6044 -5003 -6038 -5000
rect -6102 -5009 -6038 -5003
rect -2158 -5003 -2152 -5000
rect -2100 -4954 -2094 -4951
rect 1786 -4951 1850 -4945
rect 1786 -4954 1792 -4951
rect -2100 -5000 1792 -4954
rect -2100 -5003 -2094 -5000
rect -2158 -5009 -2094 -5003
rect 1786 -5003 1792 -5000
rect 1844 -4954 1850 -4951
rect 5730 -4951 5794 -4945
rect 5730 -4954 5736 -4951
rect 1844 -5000 5736 -4954
rect 1844 -5003 1850 -5000
rect 1786 -5009 1850 -5003
rect 5730 -5003 5736 -5000
rect 5788 -4954 5794 -4951
rect 9674 -4951 9738 -4945
rect 9674 -4954 9680 -4951
rect 5788 -5000 9680 -4954
rect 5788 -5003 5794 -5000
rect 5730 -5009 5794 -5003
rect 9674 -5003 9680 -5000
rect 9732 -4954 9738 -4951
rect 13618 -4951 13682 -4945
rect 13618 -4954 13624 -4951
rect 9732 -5000 13624 -4954
rect 9732 -5003 9738 -5000
rect 9674 -5009 9738 -5003
rect 13618 -5003 13624 -5000
rect 13676 -4954 13682 -4951
rect 17562 -4951 17626 -4945
rect 17562 -4954 17568 -4951
rect 13676 -5000 17568 -4954
rect 13676 -5003 13682 -5000
rect 13618 -5009 13682 -5003
rect 17562 -5003 17568 -5000
rect 17620 -4954 17626 -4951
rect 21506 -4951 21570 -4945
rect 21506 -4954 21512 -4951
rect 17620 -5000 21512 -4954
rect 17620 -5003 17626 -5000
rect 17562 -5009 17626 -5003
rect 21506 -5003 21512 -5000
rect 21564 -4954 21570 -4951
rect 21564 -5000 22976 -4954
rect 21564 -5003 21570 -5000
rect 21506 -5009 21570 -5003
rect 21445 -5392 21509 -5386
rect 2137 -5416 2201 -5410
rect 2137 -5468 2143 -5416
rect 2195 -5468 2201 -5416
rect 21445 -5444 21451 -5392
rect 21503 -5444 21509 -5392
rect 21445 -5450 21509 -5444
rect 2137 -5474 2201 -5468
rect 5875 -5536 5939 -5530
rect 5875 -5588 5881 -5536
rect 5933 -5588 5939 -5536
rect 5875 -5594 5939 -5588
rect 9819 -5536 9883 -5530
rect 9819 -5588 9825 -5536
rect 9877 -5588 9883 -5536
rect 9819 -5594 9883 -5588
rect 17707 -5678 17771 -5672
rect 17707 -5730 17713 -5678
rect 17765 -5730 17771 -5678
rect 17707 -5736 17771 -5730
rect -5641 -5930 -4981 -5884
rect -1697 -5930 -1037 -5884
rect 2247 -5930 2907 -5884
rect 6191 -5930 6851 -5884
rect 10135 -5930 10795 -5884
rect 14079 -5930 14739 -5884
rect 18023 -5930 18683 -5884
rect 21967 -5930 22627 -5884
rect -2013 -6012 -1949 -6006
rect -2013 -6064 -2007 -6012
rect -1955 -6064 -1949 -6012
rect -2013 -6070 -1949 -6064
rect -5823 -6317 -5759 -6311
rect -5823 -6369 -5817 -6317
rect -5765 -6369 -5759 -6317
rect -5823 -6375 -5759 -6369
rect 13629 -6318 13693 -6312
rect 13629 -6370 13635 -6318
rect 13687 -6370 13693 -6318
rect 13629 -6376 13693 -6370
rect -5812 -6733 -5748 -6727
rect -5812 -6736 -5806 -6733
rect -6604 -6782 -5806 -6736
rect -5812 -6785 -5806 -6782
rect -5754 -6736 -5748 -6733
rect -1868 -6733 -1804 -6727
rect -1868 -6736 -1862 -6733
rect -5754 -6782 -1862 -6736
rect -5754 -6785 -5748 -6782
rect -5812 -6791 -5748 -6785
rect -1868 -6785 -1862 -6782
rect -1810 -6736 -1804 -6733
rect 2076 -6733 2140 -6727
rect 2076 -6736 2082 -6733
rect -1810 -6782 2082 -6736
rect -1810 -6785 -1804 -6782
rect -1868 -6791 -1804 -6785
rect 2076 -6785 2082 -6782
rect 2134 -6736 2140 -6733
rect 6020 -6733 6084 -6727
rect 6020 -6736 6026 -6733
rect 2134 -6782 6026 -6736
rect 2134 -6785 2140 -6782
rect 2076 -6791 2140 -6785
rect 6020 -6785 6026 -6782
rect 6078 -6736 6084 -6733
rect 9964 -6733 10028 -6727
rect 9964 -6736 9970 -6733
rect 6078 -6782 9970 -6736
rect 6078 -6785 6084 -6782
rect 6020 -6791 6084 -6785
rect 9964 -6785 9970 -6782
rect 10022 -6736 10028 -6733
rect 13908 -6733 13972 -6727
rect 13908 -6736 13914 -6733
rect 10022 -6782 13914 -6736
rect 10022 -6785 10028 -6782
rect 9964 -6791 10028 -6785
rect 13908 -6785 13914 -6782
rect 13966 -6736 13972 -6733
rect 17852 -6733 17916 -6727
rect 17852 -6736 17858 -6733
rect 13966 -6782 17858 -6736
rect 13966 -6785 13972 -6782
rect 13908 -6791 13972 -6785
rect 17852 -6785 17858 -6782
rect 17910 -6736 17916 -6733
rect 21796 -6733 21860 -6727
rect 21796 -6736 21802 -6733
rect 17910 -6782 21802 -6736
rect 17910 -6785 17916 -6782
rect 17852 -6791 17916 -6785
rect 21796 -6785 21802 -6782
rect 21854 -6736 21860 -6733
rect 21854 -6782 22976 -6736
rect 21854 -6785 21860 -6782
rect 21796 -6791 21860 -6785
<< via1 >>
rect -6096 -5003 -6044 -4951
rect -2152 -5003 -2100 -4951
rect 1792 -5003 1844 -4951
rect 5736 -5003 5788 -4951
rect 9680 -5003 9732 -4951
rect 13624 -5003 13676 -4951
rect 17568 -5003 17620 -4951
rect 21512 -5003 21564 -4951
rect 2143 -5468 2195 -5416
rect 21451 -5444 21503 -5392
rect 5881 -5588 5933 -5536
rect 9825 -5588 9877 -5536
rect 17713 -5730 17765 -5678
rect -2007 -6064 -1955 -6012
rect -5817 -6369 -5765 -6317
rect 13635 -6370 13687 -6318
rect -5806 -6785 -5754 -6733
rect -1862 -6785 -1810 -6733
rect 2082 -6785 2134 -6733
rect 6026 -6785 6078 -6733
rect 9970 -6785 10022 -6733
rect 13914 -6785 13966 -6733
rect 17858 -6785 17910 -6733
rect 21802 -6785 21854 -6733
<< metal2 >>
rect -6107 -4949 -6033 -4940
rect -6107 -5005 -6098 -4949
rect -6042 -5005 -6033 -4949
rect -6107 -5014 -6033 -5005
rect -2163 -4949 -2089 -4940
rect -2163 -5005 -2154 -4949
rect -2098 -5005 -2089 -4949
rect -2163 -5014 -2089 -5005
rect 1781 -4949 1855 -4940
rect 1781 -5005 1790 -4949
rect 1846 -5005 1855 -4949
rect 1781 -5014 1855 -5005
rect 5725 -4949 5799 -4940
rect 5725 -5005 5734 -4949
rect 5790 -5005 5799 -4949
rect 5725 -5014 5799 -5005
rect 9669 -4949 9743 -4940
rect 9669 -5005 9678 -4949
rect 9734 -5005 9743 -4949
rect 9669 -5014 9743 -5005
rect 13613 -4949 13687 -4940
rect 13613 -5005 13622 -4949
rect 13678 -5005 13687 -4949
rect 13613 -5014 13687 -5005
rect 17557 -4949 17631 -4940
rect 17557 -5005 17566 -4949
rect 17622 -5005 17631 -4949
rect 17557 -5014 17631 -5005
rect 21501 -4949 21575 -4940
rect 21501 -5005 21510 -4949
rect 21566 -5005 21575 -4949
rect 21501 -5014 21575 -5005
rect 10912 -5390 10986 -5381
rect 2137 -5416 2201 -5410
rect 2137 -5468 2143 -5416
rect 2195 -5419 2201 -5416
rect 5563 -5414 5637 -5405
rect 5563 -5419 5572 -5414
rect 2195 -5465 5572 -5419
rect 2195 -5468 2201 -5465
rect 2137 -5474 2201 -5468
rect 5563 -5470 5572 -5465
rect 5628 -5470 5637 -5414
rect 10912 -5446 10921 -5390
rect 10977 -5395 10986 -5390
rect 21445 -5392 21509 -5386
rect 21445 -5395 21451 -5392
rect 10977 -5441 21451 -5395
rect 10977 -5446 10986 -5441
rect 10912 -5455 10986 -5446
rect 21445 -5444 21451 -5441
rect 21503 -5444 21509 -5392
rect 21445 -5450 21509 -5444
rect 5563 -5479 5637 -5470
rect 5870 -5534 5944 -5525
rect 5870 -5590 5879 -5534
rect 5935 -5590 5944 -5534
rect 5870 -5599 5944 -5590
rect 9814 -5534 9888 -5525
rect 9814 -5590 9823 -5534
rect 9879 -5590 9888 -5534
rect 9814 -5599 9888 -5590
rect 10625 -5676 10699 -5667
rect 10625 -5732 10634 -5676
rect 10690 -5681 10699 -5676
rect 17707 -5678 17771 -5672
rect 17707 -5681 17713 -5678
rect 10690 -5727 17713 -5681
rect 10690 -5732 10699 -5727
rect 10625 -5741 10699 -5732
rect 17707 -5730 17713 -5727
rect 17765 -5730 17771 -5678
rect 17707 -5736 17771 -5730
rect -2013 -6012 -1949 -6006
rect -2013 -6064 -2007 -6012
rect -1955 -6015 -1949 -6012
rect 5341 -6010 5415 -6001
rect 5341 -6015 5350 -6010
rect -1955 -6061 5350 -6015
rect -1955 -6064 -1949 -6061
rect -2013 -6070 -1949 -6064
rect 5341 -6066 5350 -6061
rect 5406 -6066 5415 -6010
rect 5341 -6075 5415 -6066
rect -5823 -6317 -5759 -6311
rect -5823 -6369 -5817 -6317
rect -5765 -6320 -5759 -6317
rect 5033 -6315 5107 -6306
rect 5033 -6320 5042 -6315
rect -5765 -6366 5042 -6320
rect -5765 -6369 -5759 -6366
rect -5823 -6375 -5759 -6369
rect 5033 -6371 5042 -6366
rect 5098 -6371 5107 -6315
rect 5033 -6380 5107 -6371
rect 10121 -6316 10195 -6307
rect 10121 -6372 10130 -6316
rect 10186 -6321 10195 -6316
rect 13629 -6318 13693 -6312
rect 13629 -6321 13635 -6318
rect 10186 -6367 13635 -6321
rect 10186 -6372 10195 -6367
rect 10121 -6381 10195 -6372
rect 13629 -6370 13635 -6367
rect 13687 -6370 13693 -6318
rect 13629 -6376 13693 -6370
rect -5817 -6731 -5743 -6722
rect -5817 -6787 -5808 -6731
rect -5752 -6787 -5743 -6731
rect -5817 -6796 -5743 -6787
rect -1873 -6731 -1799 -6722
rect -1873 -6787 -1864 -6731
rect -1808 -6787 -1799 -6731
rect -1873 -6796 -1799 -6787
rect 2071 -6731 2145 -6722
rect 2071 -6787 2080 -6731
rect 2136 -6787 2145 -6731
rect 2071 -6796 2145 -6787
rect 6015 -6731 6089 -6722
rect 6015 -6787 6024 -6731
rect 6080 -6787 6089 -6731
rect 6015 -6796 6089 -6787
rect 9959 -6731 10033 -6722
rect 9959 -6787 9968 -6731
rect 10024 -6787 10033 -6731
rect 9959 -6796 10033 -6787
rect 13903 -6731 13977 -6722
rect 13903 -6787 13912 -6731
rect 13968 -6787 13977 -6731
rect 13903 -6796 13977 -6787
rect 17847 -6731 17921 -6722
rect 17847 -6787 17856 -6731
rect 17912 -6787 17921 -6731
rect 17847 -6796 17921 -6787
rect 21791 -6731 21865 -6722
rect 21791 -6787 21800 -6731
rect 21856 -6787 21865 -6731
rect 21791 -6796 21865 -6787
<< via2 >>
rect -6098 -4951 -6042 -4949
rect -6098 -5003 -6096 -4951
rect -6096 -5003 -6044 -4951
rect -6044 -5003 -6042 -4951
rect -6098 -5005 -6042 -5003
rect -2154 -4951 -2098 -4949
rect -2154 -5003 -2152 -4951
rect -2152 -5003 -2100 -4951
rect -2100 -5003 -2098 -4951
rect -2154 -5005 -2098 -5003
rect 1790 -4951 1846 -4949
rect 1790 -5003 1792 -4951
rect 1792 -5003 1844 -4951
rect 1844 -5003 1846 -4951
rect 1790 -5005 1846 -5003
rect 5734 -4951 5790 -4949
rect 5734 -5003 5736 -4951
rect 5736 -5003 5788 -4951
rect 5788 -5003 5790 -4951
rect 5734 -5005 5790 -5003
rect 9678 -4951 9734 -4949
rect 9678 -5003 9680 -4951
rect 9680 -5003 9732 -4951
rect 9732 -5003 9734 -4951
rect 9678 -5005 9734 -5003
rect 13622 -4951 13678 -4949
rect 13622 -5003 13624 -4951
rect 13624 -5003 13676 -4951
rect 13676 -5003 13678 -4951
rect 13622 -5005 13678 -5003
rect 17566 -4951 17622 -4949
rect 17566 -5003 17568 -4951
rect 17568 -5003 17620 -4951
rect 17620 -5003 17622 -4951
rect 17566 -5005 17622 -5003
rect 21510 -4951 21566 -4949
rect 21510 -5003 21512 -4951
rect 21512 -5003 21564 -4951
rect 21564 -5003 21566 -4951
rect 21510 -5005 21566 -5003
rect 5572 -5470 5628 -5414
rect 10921 -5446 10977 -5390
rect 5879 -5536 5935 -5534
rect 5879 -5588 5881 -5536
rect 5881 -5588 5933 -5536
rect 5933 -5588 5935 -5536
rect 5879 -5590 5935 -5588
rect 9823 -5536 9879 -5534
rect 9823 -5588 9825 -5536
rect 9825 -5588 9877 -5536
rect 9877 -5588 9879 -5536
rect 9823 -5590 9879 -5588
rect 10634 -5732 10690 -5676
rect 5350 -6066 5406 -6010
rect 5042 -6371 5098 -6315
rect 10130 -6372 10186 -6316
rect -5808 -6733 -5752 -6731
rect -5808 -6785 -5806 -6733
rect -5806 -6785 -5754 -6733
rect -5754 -6785 -5752 -6733
rect -5808 -6787 -5752 -6785
rect -1864 -6733 -1808 -6731
rect -1864 -6785 -1862 -6733
rect -1862 -6785 -1810 -6733
rect -1810 -6785 -1808 -6733
rect -1864 -6787 -1808 -6785
rect 2080 -6733 2136 -6731
rect 2080 -6785 2082 -6733
rect 2082 -6785 2134 -6733
rect 2134 -6785 2136 -6733
rect 2080 -6787 2136 -6785
rect 6024 -6733 6080 -6731
rect 6024 -6785 6026 -6733
rect 6026 -6785 6078 -6733
rect 6078 -6785 6080 -6733
rect 6024 -6787 6080 -6785
rect 9968 -6733 10024 -6731
rect 9968 -6785 9970 -6733
rect 9970 -6785 10022 -6733
rect 10022 -6785 10024 -6733
rect 9968 -6787 10024 -6785
rect 13912 -6733 13968 -6731
rect 13912 -6785 13914 -6733
rect 13914 -6785 13966 -6733
rect 13966 -6785 13968 -6733
rect 13912 -6787 13968 -6785
rect 17856 -6733 17912 -6731
rect 17856 -6785 17858 -6733
rect 17858 -6785 17910 -6733
rect 17910 -6785 17912 -6733
rect 17856 -6787 17912 -6785
rect 21800 -6733 21856 -6731
rect 21800 -6785 21802 -6733
rect 21802 -6785 21854 -6733
rect 21854 -6785 21856 -6733
rect 21800 -6787 21856 -6785
<< metal3 >>
rect 9813 14023 9889 14029
rect 9813 13959 9819 14023
rect 9883 13959 9889 14023
rect 9813 13953 9889 13959
rect 5869 10523 5945 10529
rect 5869 10459 5875 10523
rect 5939 10459 5945 10523
rect 5869 10453 5945 10459
rect 5562 3312 5638 3318
rect 5562 3248 5568 3312
rect 5632 3248 5638 3312
rect 5562 3242 5638 3248
rect 5340 -252 5416 -246
rect 5340 -316 5346 -252
rect 5410 -316 5416 -252
rect 5340 -322 5416 -316
rect 5032 -1975 5108 -1969
rect 5032 -2039 5038 -1975
rect 5102 -2039 5108 -1975
rect 5032 -2045 5108 -2039
rect -6103 -4949 -6037 -4944
rect -6103 -5005 -6098 -4949
rect -6042 -5005 -6037 -4949
rect -6103 -5010 -6037 -5005
rect -2159 -4949 -2093 -4944
rect -2159 -5005 -2154 -4949
rect -2098 -5005 -2093 -4949
rect -2159 -5010 -2093 -5005
rect 1785 -4949 1851 -4944
rect 1785 -5005 1790 -4949
rect 1846 -5005 1851 -4949
rect 1785 -5010 1851 -5005
rect -6100 -5581 -6040 -5010
rect -2156 -5581 -2096 -5010
rect 1788 -5581 1848 -5010
rect -5810 -6726 -5750 -6190
rect -1866 -6726 -1806 -6190
rect 2078 -6726 2138 -6190
rect 5040 -6310 5100 -2045
rect 5348 -6005 5408 -322
rect 5570 -5409 5630 3242
rect 5729 -4949 5795 -4944
rect 5729 -5005 5734 -4949
rect 5790 -5005 5795 -4949
rect 5729 -5010 5795 -5005
rect 5567 -5414 5633 -5409
rect 5567 -5470 5572 -5414
rect 5628 -5470 5633 -5414
rect 5567 -5475 5633 -5470
rect 5732 -5581 5792 -5010
rect 5877 -5529 5937 10453
rect 9673 -4949 9739 -4944
rect 9673 -5005 9678 -4949
rect 9734 -5005 9739 -4949
rect 9673 -5010 9739 -5005
rect 5874 -5534 5940 -5529
rect 5874 -5590 5879 -5534
rect 5935 -5590 5940 -5534
rect 9676 -5581 9736 -5010
rect 9821 -5529 9881 13953
rect 10911 12235 10987 12241
rect 10911 12171 10917 12235
rect 10981 12171 10987 12235
rect 10911 12165 10987 12171
rect 10624 8662 10700 8668
rect 10624 8598 10630 8662
rect 10694 8598 10700 8662
rect 10624 8592 10700 8598
rect 10120 5096 10196 5102
rect 10120 5032 10126 5096
rect 10190 5032 10196 5096
rect 10120 5026 10196 5032
rect 9818 -5534 9884 -5529
rect 5874 -5595 5940 -5590
rect 9818 -5590 9823 -5534
rect 9879 -5590 9884 -5534
rect 9818 -5595 9884 -5590
rect 5345 -6010 5411 -6005
rect 5345 -6066 5350 -6010
rect 5406 -6066 5411 -6010
rect 5345 -6071 5411 -6066
rect 5037 -6315 5103 -6310
rect 5037 -6371 5042 -6315
rect 5098 -6371 5103 -6315
rect 5037 -6376 5103 -6371
rect 6022 -6726 6082 -6190
rect 9966 -6726 10026 -6190
rect 10128 -6311 10188 5026
rect 10632 -5671 10692 8592
rect 10919 -5385 10979 12165
rect 13617 -4949 13683 -4944
rect 13617 -5005 13622 -4949
rect 13678 -5005 13683 -4949
rect 13617 -5010 13683 -5005
rect 17561 -4949 17627 -4944
rect 17561 -5005 17566 -4949
rect 17622 -5005 17627 -4949
rect 17561 -5010 17627 -5005
rect 21505 -4949 21571 -4944
rect 21505 -5005 21510 -4949
rect 21566 -5005 21571 -4949
rect 21505 -5010 21571 -5005
rect 10916 -5390 10982 -5385
rect 10916 -5446 10921 -5390
rect 10977 -5446 10982 -5390
rect 10916 -5451 10982 -5446
rect 13620 -5581 13680 -5010
rect 17564 -5581 17624 -5010
rect 21508 -5581 21568 -5010
rect 10629 -5676 10695 -5671
rect 10629 -5732 10634 -5676
rect 10690 -5732 10695 -5676
rect 10629 -5737 10695 -5732
rect 10125 -6316 10191 -6311
rect 10125 -6372 10130 -6316
rect 10186 -6372 10191 -6316
rect 10125 -6377 10191 -6372
rect 13910 -6726 13970 -6190
rect 17854 -6726 17914 -6190
rect 21798 -6726 21858 -6190
rect -5813 -6731 -5747 -6726
rect -5813 -6787 -5808 -6731
rect -5752 -6787 -5747 -6731
rect -5813 -6792 -5747 -6787
rect -1869 -6731 -1803 -6726
rect -1869 -6787 -1864 -6731
rect -1808 -6787 -1803 -6731
rect -1869 -6792 -1803 -6787
rect 2075 -6731 2141 -6726
rect 2075 -6787 2080 -6731
rect 2136 -6787 2141 -6731
rect 2075 -6792 2141 -6787
rect 6019 -6731 6085 -6726
rect 6019 -6787 6024 -6731
rect 6080 -6787 6085 -6731
rect 6019 -6792 6085 -6787
rect 9963 -6731 10029 -6726
rect 9963 -6787 9968 -6731
rect 10024 -6787 10029 -6731
rect 9963 -6792 10029 -6787
rect 13907 -6731 13973 -6726
rect 13907 -6787 13912 -6731
rect 13968 -6787 13973 -6731
rect 13907 -6792 13973 -6787
rect 17851 -6731 17917 -6726
rect 17851 -6787 17856 -6731
rect 17912 -6787 17917 -6731
rect 17851 -6792 17917 -6787
rect 21795 -6731 21861 -6726
rect 21795 -6787 21800 -6731
rect 21856 -6787 21861 -6731
rect 21795 -6792 21861 -6787
<< via3 >>
rect 9819 13959 9883 14023
rect 5875 10459 5939 10523
rect 5568 3248 5632 3312
rect 5346 -316 5410 -252
rect 5038 -2039 5102 -1975
rect 10917 12171 10981 12235
rect 10630 8598 10694 8662
rect 10126 5032 10190 5096
<< metal4 >>
rect -36624 25764 -31280 26000
rect -31044 25764 -25700 26000
rect -25464 25764 -20120 26000
rect -19884 25764 -14540 26000
rect -14304 25764 -8960 26000
rect -8724 25764 -3380 26000
rect -3144 25764 2200 26000
rect 2436 25764 13920 26000
rect 14156 25764 19500 26000
rect 19736 25764 25080 26000
rect 25316 25764 30660 26000
rect 30896 25764 36240 26000
rect 36476 25764 41820 26000
rect 42056 25764 47400 26000
rect 47636 25764 52980 26000
rect -36624 23978 -31280 24214
rect -31044 23978 -25700 24214
rect -25464 23978 -20120 24214
rect -19884 23978 -14540 24214
rect -14304 23978 -8960 24214
rect -8724 23978 -3380 24214
rect -3144 23978 2200 24214
rect 2436 23978 13920 24214
rect 14156 23978 19500 24214
rect 19736 23978 25080 24214
rect 25316 23978 30660 24214
rect 30896 23978 36240 24214
rect 36476 23978 41820 24214
rect 42056 23978 47400 24214
rect 47636 23978 52980 24214
rect -11554 22805 -6210 23041
rect -5974 22805 22330 23041
rect 22566 22805 27910 23041
rect -36624 22192 -31280 22428
rect -31044 22192 -25700 22428
rect -25464 22192 -20120 22428
rect -19884 22192 -14540 22428
rect -14304 22192 -8960 22428
rect -8724 22192 -3380 22428
rect -3144 22192 2200 22428
rect 2436 22192 13920 22428
rect 14156 22192 19500 22428
rect 19736 22192 25080 22428
rect 25316 22192 30660 22428
rect 30896 22192 36240 22428
rect 36476 22192 41820 22428
rect 42056 22192 47400 22428
rect 47636 22192 52980 22428
rect 5186 21019 11170 21255
rect -36624 20406 -31280 20642
rect -31044 20406 -25700 20642
rect -25464 20406 -20120 20642
rect -19884 20406 -14540 20642
rect -14304 20406 -8960 20642
rect -8724 20406 -3380 20642
rect -3144 20406 2200 20642
rect 2436 20406 13920 20642
rect 14156 20406 19500 20642
rect 19736 20406 25080 20642
rect 25316 20406 30660 20642
rect 30896 20406 36240 20642
rect 36476 20406 41820 20642
rect 42056 20406 47400 20642
rect 47636 20406 52980 20642
rect -394 19233 16750 19469
rect -36624 18620 -31280 18856
rect -31044 18620 -25700 18856
rect -25464 18620 -20120 18856
rect -19884 18620 -14540 18856
rect -14304 18620 -8960 18856
rect -8724 18620 -3380 18856
rect -3144 18620 2200 18856
rect 2436 18620 13920 18856
rect 14156 18620 19500 18856
rect 19736 18620 25080 18856
rect 25316 18620 30660 18856
rect 30896 18620 36240 18856
rect 36476 18620 41820 18856
rect 42056 18620 47400 18856
rect 47636 18620 52980 18856
rect -36624 16834 -31280 17070
rect -31044 16834 -25700 17070
rect -25464 16834 -20120 17070
rect -19884 16834 -14540 17070
rect -14304 16834 -8960 17070
rect -8724 16834 -3380 17070
rect -3144 16834 2200 17070
rect 2436 16834 13920 17070
rect 14156 16834 19500 17070
rect 19736 16834 25080 17070
rect 25316 16834 30660 17070
rect 30896 16834 36240 17070
rect 36476 16834 41820 17070
rect 42056 16834 47400 17070
rect 47636 16834 52980 17070
rect -36624 15048 -31280 15284
rect -31044 15048 -25700 15284
rect -25464 15048 -20120 15284
rect -19884 15048 -14540 15284
rect -14304 15048 -8960 15284
rect -8724 15048 -3380 15284
rect -3144 15048 2200 15284
rect 2436 15048 13920 15284
rect 14156 15048 19500 15284
rect 19736 15048 25080 15284
rect 25316 15048 30660 15284
rect 30896 15048 36240 15284
rect 36476 15048 41820 15284
rect 42056 15048 47400 15284
rect 47636 15048 52980 15284
rect 5186 14023 11170 14111
rect 5186 13959 9819 14023
rect 9883 13959 11170 14023
rect 5186 13875 11170 13959
rect -36624 13262 -31280 13498
rect -31044 13262 -25700 13498
rect -25464 13262 -20120 13498
rect -19884 13262 -14540 13498
rect -14304 13262 -8960 13498
rect -8724 13262 -3380 13498
rect -3144 13262 2200 13498
rect 2436 13262 13920 13498
rect 14156 13262 19500 13498
rect 19736 13262 25080 13498
rect 25316 13262 30660 13498
rect 30896 13262 36240 13498
rect 36476 13262 41820 13498
rect 42056 13262 47400 13498
rect 47636 13262 52980 13498
rect -33874 12089 -28530 12325
rect -28294 12089 -22950 12325
rect -22714 12089 -17370 12325
rect -17134 12235 33490 12325
rect -17134 12171 10917 12235
rect 10981 12171 33490 12235
rect -17134 12089 33490 12171
rect 33726 12089 39070 12325
rect 39306 12089 44650 12325
rect 44886 12089 50230 12325
rect -36624 11476 -31280 11712
rect -31044 11476 -25700 11712
rect -25464 11476 -20120 11712
rect -19884 11476 -14540 11712
rect -14304 11476 -8960 11712
rect -8724 11476 -3380 11712
rect -3144 11476 2200 11712
rect 2436 11476 13920 11712
rect 14156 11476 19500 11712
rect 19736 11476 25080 11712
rect 25316 11476 30660 11712
rect 30896 11476 36240 11712
rect 36476 11476 41820 11712
rect 42056 11476 47400 11712
rect 47636 11476 52980 11712
rect 5186 10523 11170 10608
rect 5186 10459 5875 10523
rect 5939 10459 11170 10523
rect 5186 10372 11170 10459
rect -36624 9690 -31280 9926
rect -31044 9690 -25700 9926
rect -25464 9690 -20120 9926
rect -19884 9690 -14540 9926
rect -14304 9690 -8960 9926
rect -8724 9690 -3380 9926
rect -3144 9690 2200 9926
rect 2436 9690 13920 9926
rect 14156 9690 19500 9926
rect 19736 9690 25080 9926
rect 25316 9690 30660 9926
rect 30896 9690 36240 9926
rect 36476 9690 41820 9926
rect 42056 9690 47400 9926
rect 47636 9690 52980 9926
rect -11554 8517 -6210 8753
rect -5974 8662 22330 8753
rect -5974 8598 10630 8662
rect 10694 8598 22330 8662
rect -5974 8517 22330 8598
rect 22566 8517 27910 8753
rect -36624 7904 -31280 8140
rect -31044 7904 -25700 8140
rect -25464 7904 -20120 8140
rect -19884 7904 -14540 8140
rect -14304 7904 -8960 8140
rect -8724 7904 -3380 8140
rect -3144 7904 2200 8140
rect 2436 7904 13920 8140
rect 14156 7904 19500 8140
rect 19736 7904 25080 8140
rect 25316 7904 30660 8140
rect 30896 7904 36240 8140
rect 36476 7904 41820 8140
rect 42056 7904 47400 8140
rect 47636 7904 52980 8140
rect 5186 6800 11170 7036
rect -36624 6118 -31280 6354
rect -31044 6118 -25700 6354
rect -25464 6118 -20120 6354
rect -19884 6118 -14540 6354
rect -14304 6118 -8960 6354
rect -8724 6118 -3380 6354
rect -3144 6118 2200 6354
rect 2436 6118 13920 6354
rect 14156 6118 19500 6354
rect 19736 6118 25080 6354
rect 25316 6118 30660 6354
rect 30896 6118 36240 6354
rect 36476 6118 41820 6354
rect 42056 6118 47400 6354
rect 47636 6118 52980 6354
rect -394 5096 16750 5181
rect -394 5032 10126 5096
rect 10190 5032 16750 5096
rect -394 4945 16750 5032
rect -36624 4332 -31280 4568
rect -31044 4332 -25700 4568
rect -25464 4332 -20120 4568
rect -19884 4332 -14540 4568
rect -14304 4332 -8960 4568
rect -8724 4332 -3380 4568
rect -3144 4332 2200 4568
rect 2436 4332 13920 4568
rect 14156 4332 19500 4568
rect 19736 4332 25080 4568
rect 25316 4332 30660 4568
rect 30896 4332 36240 4568
rect 36476 4332 41820 4568
rect 42056 4332 47400 4568
rect 47636 4332 52980 4568
rect 5186 3312 11170 3395
rect 5186 3248 5568 3312
rect 5632 3248 11170 3312
rect 5186 3159 11170 3248
rect -36624 2546 -31280 2782
rect -31044 2546 -25700 2782
rect -25464 2546 -20120 2782
rect -19884 2546 -14540 2782
rect -14304 2546 -8960 2782
rect -8724 2546 -3380 2782
rect -3144 2546 2200 2782
rect 2436 2546 13920 2782
rect 14156 2546 19500 2782
rect 19736 2546 25080 2782
rect 25316 2546 30660 2782
rect 30896 2546 36240 2782
rect 36476 2546 41820 2782
rect 42056 2546 47400 2782
rect 47636 2546 52980 2782
rect 5186 1373 11170 1609
rect -36624 760 -31280 996
rect -31044 760 -25700 996
rect -25464 760 -20120 996
rect -19884 760 -14540 996
rect -14304 760 -8960 996
rect -8724 760 -3380 996
rect -3144 760 2200 996
rect 2436 760 13920 996
rect 14156 760 19500 996
rect 19736 760 25080 996
rect 25316 760 30660 996
rect 30896 760 36240 996
rect 36476 760 41820 996
rect 42056 760 47400 996
rect 47636 760 52980 996
rect 5186 -252 11170 -177
rect 5186 -316 5346 -252
rect 5410 -316 11170 -252
rect 5186 -413 11170 -316
rect -36624 -1026 -31280 -790
rect -31044 -1026 -25700 -790
rect -25464 -1026 -20120 -790
rect -19884 -1026 -14540 -790
rect -14304 -1026 -8960 -790
rect -8724 -1026 -3380 -790
rect -3144 -1026 2200 -790
rect 2436 -1026 19500 -790
rect 19736 -1026 25080 -790
rect 25316 -1026 30660 -790
rect 30896 -1026 36240 -790
rect 36476 -1026 41820 -790
rect 42056 -1026 47400 -790
rect 47636 -1026 52980 -790
<< via4 >>
rect -36860 25764 -36624 26000
rect -31280 25764 -31044 26000
rect -25700 25764 -25464 26000
rect -20120 25764 -19884 26000
rect -14540 25764 -14304 26000
rect -8960 25764 -8724 26000
rect -3380 25764 -3144 26000
rect 2200 25764 2436 26000
rect 13920 25764 14156 26000
rect 19500 25764 19736 26000
rect 25080 25764 25316 26000
rect 30660 25764 30896 26000
rect 36240 25764 36476 26000
rect 41820 25764 42056 26000
rect 47400 25764 47636 26000
rect 52980 25764 53216 26000
rect -36860 23978 -36624 24214
rect -31280 23978 -31044 24214
rect -25700 23978 -25464 24214
rect -20120 23978 -19884 24214
rect -14540 23978 -14304 24214
rect -8960 23978 -8724 24214
rect -3380 23978 -3144 24214
rect 2200 23978 2436 24214
rect 13920 23978 14156 24214
rect 19500 23978 19736 24214
rect 25080 23978 25316 24214
rect 30660 23978 30896 24214
rect 36240 23978 36476 24214
rect 41820 23978 42056 24214
rect 47400 23978 47636 24214
rect 52980 23978 53216 24214
rect -11790 22805 -11554 23041
rect -6210 22805 -5974 23041
rect 22330 22805 22566 23041
rect 27910 22805 28146 23041
rect -36860 22192 -36624 22428
rect -31280 22192 -31044 22428
rect -25700 22192 -25464 22428
rect -20120 22192 -19884 22428
rect -14540 22192 -14304 22428
rect -8960 22192 -8724 22428
rect -3380 22192 -3144 22428
rect 2200 22192 2436 22428
rect 13920 22192 14156 22428
rect 19500 22192 19736 22428
rect 25080 22192 25316 22428
rect 30660 22192 30896 22428
rect 36240 22192 36476 22428
rect 41820 22192 42056 22428
rect 47400 22192 47636 22428
rect 52980 22192 53216 22428
rect 4950 21019 5186 21255
rect 11170 21019 11406 21255
rect -36860 20406 -36624 20642
rect -31280 20406 -31044 20642
rect -25700 20406 -25464 20642
rect -20120 20406 -19884 20642
rect -14540 20406 -14304 20642
rect -8960 20406 -8724 20642
rect -3380 20406 -3144 20642
rect 2200 20406 2436 20642
rect 13920 20406 14156 20642
rect 19500 20406 19736 20642
rect 25080 20406 25316 20642
rect 30660 20406 30896 20642
rect 36240 20406 36476 20642
rect 41820 20406 42056 20642
rect 47400 20406 47636 20642
rect 52980 20406 53216 20642
rect -630 19233 -394 19469
rect 16750 19233 16986 19469
rect -36860 18620 -36624 18856
rect -31280 18620 -31044 18856
rect -25700 18620 -25464 18856
rect -20120 18620 -19884 18856
rect -14540 18620 -14304 18856
rect -8960 18620 -8724 18856
rect -3380 18620 -3144 18856
rect 2200 18620 2436 18856
rect 13920 18620 14156 18856
rect 19500 18620 19736 18856
rect 25080 18620 25316 18856
rect 30660 18620 30896 18856
rect 36240 18620 36476 18856
rect 41820 18620 42056 18856
rect 47400 18620 47636 18856
rect 52980 18620 53216 18856
rect -36860 16834 -36624 17070
rect -31280 16834 -31044 17070
rect -25700 16834 -25464 17070
rect -20120 16834 -19884 17070
rect -14540 16834 -14304 17070
rect -8960 16834 -8724 17070
rect -3380 16834 -3144 17070
rect 2200 16834 2436 17070
rect 13920 16834 14156 17070
rect 19500 16834 19736 17070
rect 25080 16834 25316 17070
rect 30660 16834 30896 17070
rect 36240 16834 36476 17070
rect 41820 16834 42056 17070
rect 47400 16834 47636 17070
rect 52980 16834 53216 17070
rect -36860 15048 -36624 15284
rect -31280 15048 -31044 15284
rect -25700 15048 -25464 15284
rect -20120 15048 -19884 15284
rect -14540 15048 -14304 15284
rect -8960 15048 -8724 15284
rect -3380 15048 -3144 15284
rect 2200 15048 2436 15284
rect 13920 15048 14156 15284
rect 19500 15048 19736 15284
rect 25080 15048 25316 15284
rect 30660 15048 30896 15284
rect 36240 15048 36476 15284
rect 41820 15048 42056 15284
rect 47400 15048 47636 15284
rect 52980 15048 53216 15284
rect 4950 13875 5186 14111
rect 11170 13875 11406 14111
rect -36860 13262 -36624 13498
rect -31280 13262 -31044 13498
rect -25700 13262 -25464 13498
rect -20120 13262 -19884 13498
rect -14540 13262 -14304 13498
rect -8960 13262 -8724 13498
rect -3380 13262 -3144 13498
rect 2200 13262 2436 13498
rect 13920 13262 14156 13498
rect 19500 13262 19736 13498
rect 25080 13262 25316 13498
rect 30660 13262 30896 13498
rect 36240 13262 36476 13498
rect 41820 13262 42056 13498
rect 47400 13262 47636 13498
rect 52980 13262 53216 13498
rect -34110 12089 -33874 12325
rect -28530 12089 -28294 12325
rect -22950 12089 -22714 12325
rect -17370 12089 -17134 12325
rect 33490 12089 33726 12325
rect 39070 12089 39306 12325
rect 44650 12089 44886 12325
rect 50230 12089 50466 12325
rect -36860 11476 -36624 11712
rect -31280 11476 -31044 11712
rect -25700 11476 -25464 11712
rect -20120 11476 -19884 11712
rect -14540 11476 -14304 11712
rect -8960 11476 -8724 11712
rect -3380 11476 -3144 11712
rect 2200 11476 2436 11712
rect 13920 11476 14156 11712
rect 19500 11476 19736 11712
rect 25080 11476 25316 11712
rect 30660 11476 30896 11712
rect 36240 11476 36476 11712
rect 41820 11476 42056 11712
rect 47400 11476 47636 11712
rect 52980 11476 53216 11712
rect 4950 10372 5186 10608
rect 11170 10372 11406 10608
rect -36860 9690 -36624 9926
rect -31280 9690 -31044 9926
rect -25700 9690 -25464 9926
rect -20120 9690 -19884 9926
rect -14540 9690 -14304 9926
rect -8960 9690 -8724 9926
rect -3380 9690 -3144 9926
rect 2200 9690 2436 9926
rect 13920 9690 14156 9926
rect 19500 9690 19736 9926
rect 25080 9690 25316 9926
rect 30660 9690 30896 9926
rect 36240 9690 36476 9926
rect 41820 9690 42056 9926
rect 47400 9690 47636 9926
rect 52980 9690 53216 9926
rect -11790 8517 -11554 8753
rect -6210 8517 -5974 8753
rect 22330 8517 22566 8753
rect 27910 8517 28146 8753
rect -36860 7904 -36624 8140
rect -31280 7904 -31044 8140
rect -25700 7904 -25464 8140
rect -20120 7904 -19884 8140
rect -14540 7904 -14304 8140
rect -8960 7904 -8724 8140
rect -3380 7904 -3144 8140
rect 2200 7904 2436 8140
rect 13920 7904 14156 8140
rect 19500 7904 19736 8140
rect 25080 7904 25316 8140
rect 30660 7904 30896 8140
rect 36240 7904 36476 8140
rect 41820 7904 42056 8140
rect 47400 7904 47636 8140
rect 52980 7904 53216 8140
rect 4950 6800 5186 7036
rect 11170 6800 11406 7036
rect -36860 6118 -36624 6354
rect -31280 6118 -31044 6354
rect -25700 6118 -25464 6354
rect -20120 6118 -19884 6354
rect -14540 6118 -14304 6354
rect -8960 6118 -8724 6354
rect -3380 6118 -3144 6354
rect 2200 6118 2436 6354
rect 13920 6118 14156 6354
rect 19500 6118 19736 6354
rect 25080 6118 25316 6354
rect 30660 6118 30896 6354
rect 36240 6118 36476 6354
rect 41820 6118 42056 6354
rect 47400 6118 47636 6354
rect 52980 6118 53216 6354
rect -630 4945 -394 5181
rect 16750 4945 16986 5181
rect -36860 4332 -36624 4568
rect -31280 4332 -31044 4568
rect -25700 4332 -25464 4568
rect -20120 4332 -19884 4568
rect -14540 4332 -14304 4568
rect -8960 4332 -8724 4568
rect -3380 4332 -3144 4568
rect 2200 4332 2436 4568
rect 13920 4332 14156 4568
rect 19500 4332 19736 4568
rect 25080 4332 25316 4568
rect 30660 4332 30896 4568
rect 36240 4332 36476 4568
rect 41820 4332 42056 4568
rect 47400 4332 47636 4568
rect 52980 4332 53216 4568
rect 4950 3159 5186 3395
rect 11170 3159 11406 3395
rect -36860 2546 -36624 2782
rect -31280 2546 -31044 2782
rect -25700 2546 -25464 2782
rect -20120 2546 -19884 2782
rect -14540 2546 -14304 2782
rect -8960 2546 -8724 2782
rect -3380 2546 -3144 2782
rect 2200 2546 2436 2782
rect 13920 2546 14156 2782
rect 19500 2546 19736 2782
rect 25080 2546 25316 2782
rect 30660 2546 30896 2782
rect 36240 2546 36476 2782
rect 41820 2546 42056 2782
rect 47400 2546 47636 2782
rect 52980 2546 53216 2782
rect 4950 1373 5186 1609
rect 11170 1373 11406 1609
rect -36860 760 -36624 996
rect -31280 760 -31044 996
rect -25700 760 -25464 996
rect -20120 760 -19884 996
rect -14540 760 -14304 996
rect -8960 760 -8724 996
rect -3380 760 -3144 996
rect 2200 760 2436 996
rect 13920 760 14156 996
rect 19500 760 19736 996
rect 25080 760 25316 996
rect 30660 760 30896 996
rect 36240 760 36476 996
rect 41820 760 42056 996
rect 47400 760 47636 996
rect 52980 760 53216 996
rect 4950 -413 5186 -177
rect 11170 -413 11406 -177
rect -36860 -1026 -36624 -790
rect -31280 -1026 -31044 -790
rect -25700 -1026 -25464 -790
rect -20120 -1026 -19884 -790
rect -14540 -1026 -14304 -790
rect -8960 -1026 -8724 -790
rect -3380 -1026 -3144 -790
rect 2200 -1026 2436 -790
rect 19500 -1026 19736 -790
rect 25080 -1026 25316 -790
rect 30660 -1026 30896 -790
rect 36240 -1026 36476 -790
rect 41820 -1026 42056 -790
rect 47400 -1026 47636 -790
rect 52980 -1026 53216 -790
rect -34110 -2130 -33874 -1894
rect -28530 -2130 -28294 -1894
rect -22950 -2130 -22714 -1894
rect -17370 -2130 -17134 -1894
rect -11790 -2130 -11554 -1894
rect -6210 -2130 -5974 -1894
rect -630 -2130 -394 -1894
rect 4950 -1975 5186 -1894
rect 4950 -2039 5038 -1975
rect 5038 -2039 5102 -1975
rect 5102 -2039 5186 -1975
rect 4950 -2130 5186 -2039
rect 16750 -2130 16986 -1894
rect 22330 -2130 22566 -1894
rect 27910 -2130 28146 -1894
rect 33490 -2130 33726 -1894
rect 39070 -2130 39306 -1894
rect 44650 -2130 44886 -1894
rect 50230 -2130 50466 -1894
<< metal5 >>
rect -36902 26000 -36582 26024
rect -36902 25764 -36860 26000
rect -36624 25764 -36582 26000
rect -36902 24214 -36582 25764
rect -31322 26000 -31002 26024
rect -31322 25764 -31280 26000
rect -31044 25764 -31002 26000
rect -36902 23978 -36860 24214
rect -36624 23978 -36582 24214
rect -36902 22428 -36582 23978
rect -36902 22192 -36860 22428
rect -36624 22192 -36582 22428
rect -36902 20642 -36582 22192
rect -36902 20406 -36860 20642
rect -36624 20406 -36582 20642
rect -36902 18856 -36582 20406
rect -36902 18620 -36860 18856
rect -36624 18620 -36582 18856
rect -36902 17070 -36582 18620
rect -36902 16834 -36860 17070
rect -36624 16834 -36582 17070
rect -36902 15284 -36582 16834
rect -36902 15048 -36860 15284
rect -36624 15048 -36582 15284
rect -36902 13498 -36582 15048
rect -36902 13262 -36860 13498
rect -36624 13262 -36582 13498
rect -36902 11712 -36582 13262
rect -36902 11476 -36860 11712
rect -36624 11476 -36582 11712
rect -36902 9926 -36582 11476
rect -36902 9690 -36860 9926
rect -36624 9690 -36582 9926
rect -36902 8140 -36582 9690
rect -36902 7904 -36860 8140
rect -36624 7904 -36582 8140
rect -36902 6354 -36582 7904
rect -36902 6118 -36860 6354
rect -36624 6118 -36582 6354
rect -36902 4568 -36582 6118
rect -36902 4332 -36860 4568
rect -36624 4332 -36582 4568
rect -36902 2782 -36582 4332
rect -36902 2546 -36860 2782
rect -36624 2546 -36582 2782
rect -36902 996 -36582 2546
rect -36902 760 -36860 996
rect -36624 760 -36582 996
rect -36902 -790 -36582 760
rect -36902 -1026 -36860 -790
rect -36624 -1026 -36582 -790
rect -36902 -1894 -36582 -1026
rect -34152 12325 -33832 25696
rect -34152 12089 -34110 12325
rect -33874 12089 -33832 12325
rect -34152 -1894 -33832 12089
rect -31322 24214 -31002 25764
rect -25742 26000 -25422 26024
rect -25742 25764 -25700 26000
rect -25464 25764 -25422 26000
rect -31322 23978 -31280 24214
rect -31044 23978 -31002 24214
rect -31322 22428 -31002 23978
rect -31322 22192 -31280 22428
rect -31044 22192 -31002 22428
rect -31322 20642 -31002 22192
rect -31322 20406 -31280 20642
rect -31044 20406 -31002 20642
rect -31322 18856 -31002 20406
rect -31322 18620 -31280 18856
rect -31044 18620 -31002 18856
rect -31322 17070 -31002 18620
rect -31322 16834 -31280 17070
rect -31044 16834 -31002 17070
rect -31322 15284 -31002 16834
rect -31322 15048 -31280 15284
rect -31044 15048 -31002 15284
rect -31322 13498 -31002 15048
rect -31322 13262 -31280 13498
rect -31044 13262 -31002 13498
rect -31322 11712 -31002 13262
rect -31322 11476 -31280 11712
rect -31044 11476 -31002 11712
rect -31322 9926 -31002 11476
rect -31322 9690 -31280 9926
rect -31044 9690 -31002 9926
rect -31322 8140 -31002 9690
rect -31322 7904 -31280 8140
rect -31044 7904 -31002 8140
rect -31322 6354 -31002 7904
rect -31322 6118 -31280 6354
rect -31044 6118 -31002 6354
rect -31322 4568 -31002 6118
rect -31322 4332 -31280 4568
rect -31044 4332 -31002 4568
rect -31322 2782 -31002 4332
rect -31322 2546 -31280 2782
rect -31044 2546 -31002 2782
rect -31322 996 -31002 2546
rect -31322 760 -31280 996
rect -31044 760 -31002 996
rect -31322 -790 -31002 760
rect -31322 -1026 -31280 -790
rect -31044 -1026 -31002 -790
rect -31322 -1894 -31002 -1026
rect -28572 12325 -28252 25696
rect -28572 12089 -28530 12325
rect -28294 12089 -28252 12325
rect -28572 -1894 -28252 12089
rect -25742 24214 -25422 25764
rect -20162 26000 -19842 26024
rect -20162 25764 -20120 26000
rect -19884 25764 -19842 26000
rect -25742 23978 -25700 24214
rect -25464 23978 -25422 24214
rect -25742 22428 -25422 23978
rect -25742 22192 -25700 22428
rect -25464 22192 -25422 22428
rect -25742 20642 -25422 22192
rect -25742 20406 -25700 20642
rect -25464 20406 -25422 20642
rect -25742 18856 -25422 20406
rect -25742 18620 -25700 18856
rect -25464 18620 -25422 18856
rect -25742 17070 -25422 18620
rect -25742 16834 -25700 17070
rect -25464 16834 -25422 17070
rect -25742 15284 -25422 16834
rect -25742 15048 -25700 15284
rect -25464 15048 -25422 15284
rect -25742 13498 -25422 15048
rect -25742 13262 -25700 13498
rect -25464 13262 -25422 13498
rect -25742 11712 -25422 13262
rect -25742 11476 -25700 11712
rect -25464 11476 -25422 11712
rect -25742 9926 -25422 11476
rect -25742 9690 -25700 9926
rect -25464 9690 -25422 9926
rect -25742 8140 -25422 9690
rect -25742 7904 -25700 8140
rect -25464 7904 -25422 8140
rect -25742 6354 -25422 7904
rect -25742 6118 -25700 6354
rect -25464 6118 -25422 6354
rect -25742 4568 -25422 6118
rect -25742 4332 -25700 4568
rect -25464 4332 -25422 4568
rect -25742 2782 -25422 4332
rect -25742 2546 -25700 2782
rect -25464 2546 -25422 2782
rect -25742 996 -25422 2546
rect -25742 760 -25700 996
rect -25464 760 -25422 996
rect -25742 -790 -25422 760
rect -25742 -1026 -25700 -790
rect -25464 -1026 -25422 -790
rect -25742 -1894 -25422 -1026
rect -22992 12325 -22672 25696
rect -22992 12089 -22950 12325
rect -22714 12089 -22672 12325
rect -22992 -1894 -22672 12089
rect -20162 24214 -19842 25764
rect -14582 26000 -14262 26024
rect -14582 25764 -14540 26000
rect -14304 25764 -14262 26000
rect -20162 23978 -20120 24214
rect -19884 23978 -19842 24214
rect -20162 22428 -19842 23978
rect -20162 22192 -20120 22428
rect -19884 22192 -19842 22428
rect -20162 20642 -19842 22192
rect -20162 20406 -20120 20642
rect -19884 20406 -19842 20642
rect -20162 18856 -19842 20406
rect -20162 18620 -20120 18856
rect -19884 18620 -19842 18856
rect -20162 17070 -19842 18620
rect -20162 16834 -20120 17070
rect -19884 16834 -19842 17070
rect -20162 15284 -19842 16834
rect -20162 15048 -20120 15284
rect -19884 15048 -19842 15284
rect -20162 13498 -19842 15048
rect -20162 13262 -20120 13498
rect -19884 13262 -19842 13498
rect -20162 11712 -19842 13262
rect -20162 11476 -20120 11712
rect -19884 11476 -19842 11712
rect -20162 9926 -19842 11476
rect -20162 9690 -20120 9926
rect -19884 9690 -19842 9926
rect -20162 8140 -19842 9690
rect -20162 7904 -20120 8140
rect -19884 7904 -19842 8140
rect -20162 6354 -19842 7904
rect -20162 6118 -20120 6354
rect -19884 6118 -19842 6354
rect -20162 4568 -19842 6118
rect -20162 4332 -20120 4568
rect -19884 4332 -19842 4568
rect -20162 2782 -19842 4332
rect -20162 2546 -20120 2782
rect -19884 2546 -19842 2782
rect -20162 996 -19842 2546
rect -20162 760 -20120 996
rect -19884 760 -19842 996
rect -20162 -790 -19842 760
rect -20162 -1026 -20120 -790
rect -19884 -1026 -19842 -790
rect -20162 -1894 -19842 -1026
rect -17412 12325 -17092 25696
rect -17412 12089 -17370 12325
rect -17134 12089 -17092 12325
rect -17412 -1894 -17092 12089
rect -14582 24214 -14262 25764
rect -9002 26000 -8682 26024
rect -9002 25764 -8960 26000
rect -8724 25764 -8682 26000
rect -14582 23978 -14540 24214
rect -14304 23978 -14262 24214
rect -14582 22428 -14262 23978
rect -14582 22192 -14540 22428
rect -14304 22192 -14262 22428
rect -14582 20642 -14262 22192
rect -14582 20406 -14540 20642
rect -14304 20406 -14262 20642
rect -14582 18856 -14262 20406
rect -14582 18620 -14540 18856
rect -14304 18620 -14262 18856
rect -14582 17070 -14262 18620
rect -14582 16834 -14540 17070
rect -14304 16834 -14262 17070
rect -14582 15284 -14262 16834
rect -14582 15048 -14540 15284
rect -14304 15048 -14262 15284
rect -14582 13498 -14262 15048
rect -14582 13262 -14540 13498
rect -14304 13262 -14262 13498
rect -14582 11712 -14262 13262
rect -14582 11476 -14540 11712
rect -14304 11476 -14262 11712
rect -14582 9926 -14262 11476
rect -14582 9690 -14540 9926
rect -14304 9690 -14262 9926
rect -14582 8140 -14262 9690
rect -14582 7904 -14540 8140
rect -14304 7904 -14262 8140
rect -14582 6354 -14262 7904
rect -14582 6118 -14540 6354
rect -14304 6118 -14262 6354
rect -14582 4568 -14262 6118
rect -14582 4332 -14540 4568
rect -14304 4332 -14262 4568
rect -14582 2782 -14262 4332
rect -14582 2546 -14540 2782
rect -14304 2546 -14262 2782
rect -14582 996 -14262 2546
rect -14582 760 -14540 996
rect -14304 760 -14262 996
rect -14582 -790 -14262 760
rect -14582 -1026 -14540 -790
rect -14304 -1026 -14262 -790
rect -14582 -1894 -14262 -1026
rect -11832 23041 -11512 25696
rect -11832 22805 -11790 23041
rect -11554 22805 -11512 23041
rect -11832 8753 -11512 22805
rect -11832 8517 -11790 8753
rect -11554 8517 -11512 8753
rect -11832 -1894 -11512 8517
rect -9002 24214 -8682 25764
rect -3422 26000 -3102 26024
rect -3422 25764 -3380 26000
rect -3144 25764 -3102 26000
rect -9002 23978 -8960 24214
rect -8724 23978 -8682 24214
rect -9002 22428 -8682 23978
rect -9002 22192 -8960 22428
rect -8724 22192 -8682 22428
rect -9002 20642 -8682 22192
rect -9002 20406 -8960 20642
rect -8724 20406 -8682 20642
rect -9002 18856 -8682 20406
rect -9002 18620 -8960 18856
rect -8724 18620 -8682 18856
rect -9002 17070 -8682 18620
rect -9002 16834 -8960 17070
rect -8724 16834 -8682 17070
rect -9002 15284 -8682 16834
rect -9002 15048 -8960 15284
rect -8724 15048 -8682 15284
rect -9002 13498 -8682 15048
rect -9002 13262 -8960 13498
rect -8724 13262 -8682 13498
rect -9002 11712 -8682 13262
rect -9002 11476 -8960 11712
rect -8724 11476 -8682 11712
rect -9002 9926 -8682 11476
rect -9002 9690 -8960 9926
rect -8724 9690 -8682 9926
rect -9002 8140 -8682 9690
rect -9002 7904 -8960 8140
rect -8724 7904 -8682 8140
rect -9002 6354 -8682 7904
rect -9002 6118 -8960 6354
rect -8724 6118 -8682 6354
rect -9002 4568 -8682 6118
rect -9002 4332 -8960 4568
rect -8724 4332 -8682 4568
rect -9002 2782 -8682 4332
rect -9002 2546 -8960 2782
rect -8724 2546 -8682 2782
rect -9002 996 -8682 2546
rect -9002 760 -8960 996
rect -8724 760 -8682 996
rect -9002 -790 -8682 760
rect -9002 -1026 -8960 -790
rect -8724 -1026 -8682 -790
rect -9002 -1894 -8682 -1026
rect -6252 23041 -5932 25696
rect -6252 22805 -6210 23041
rect -5974 22805 -5932 23041
rect -6252 8753 -5932 22805
rect -6252 8517 -6210 8753
rect -5974 8517 -5932 8753
rect -6252 -1894 -5932 8517
rect -3422 24214 -3102 25764
rect 2158 26000 2478 26024
rect 2158 25764 2200 26000
rect 2436 25764 2478 26000
rect -3422 23978 -3380 24214
rect -3144 23978 -3102 24214
rect -3422 22428 -3102 23978
rect -3422 22192 -3380 22428
rect -3144 22192 -3102 22428
rect -3422 20642 -3102 22192
rect -3422 20406 -3380 20642
rect -3144 20406 -3102 20642
rect -3422 18856 -3102 20406
rect -3422 18620 -3380 18856
rect -3144 18620 -3102 18856
rect -3422 17070 -3102 18620
rect -3422 16834 -3380 17070
rect -3144 16834 -3102 17070
rect -3422 15284 -3102 16834
rect -3422 15048 -3380 15284
rect -3144 15048 -3102 15284
rect -3422 13498 -3102 15048
rect -3422 13262 -3380 13498
rect -3144 13262 -3102 13498
rect -3422 11712 -3102 13262
rect -3422 11476 -3380 11712
rect -3144 11476 -3102 11712
rect -3422 9926 -3102 11476
rect -3422 9690 -3380 9926
rect -3144 9690 -3102 9926
rect -3422 8140 -3102 9690
rect -3422 7904 -3380 8140
rect -3144 7904 -3102 8140
rect -3422 6354 -3102 7904
rect -3422 6118 -3380 6354
rect -3144 6118 -3102 6354
rect -3422 4568 -3102 6118
rect -3422 4332 -3380 4568
rect -3144 4332 -3102 4568
rect -3422 2782 -3102 4332
rect -3422 2546 -3380 2782
rect -3144 2546 -3102 2782
rect -3422 996 -3102 2546
rect -3422 760 -3380 996
rect -3144 760 -3102 996
rect -3422 -790 -3102 760
rect -3422 -1026 -3380 -790
rect -3144 -1026 -3102 -790
rect -3422 -1894 -3102 -1026
rect -672 19469 -352 25696
rect -672 19233 -630 19469
rect -394 19233 -352 19469
rect -672 5181 -352 19233
rect -672 4945 -630 5181
rect -394 4945 -352 5181
rect -672 -1894 -352 4945
rect 2158 24214 2478 25764
rect 13878 26000 14198 26024
rect 13878 25764 13920 26000
rect 14156 25764 14198 26000
rect 2158 23978 2200 24214
rect 2436 23978 2478 24214
rect 2158 22428 2478 23978
rect 2158 22192 2200 22428
rect 2436 22192 2478 22428
rect 2158 20642 2478 22192
rect 2158 20406 2200 20642
rect 2436 20406 2478 20642
rect 2158 18856 2478 20406
rect 2158 18620 2200 18856
rect 2436 18620 2478 18856
rect 2158 17070 2478 18620
rect 2158 16834 2200 17070
rect 2436 16834 2478 17070
rect 2158 15284 2478 16834
rect 2158 15048 2200 15284
rect 2436 15048 2478 15284
rect 2158 13498 2478 15048
rect 2158 13262 2200 13498
rect 2436 13262 2478 13498
rect 2158 11712 2478 13262
rect 4908 21255 5228 25696
rect 4908 21019 4950 21255
rect 5186 21019 5228 21255
rect 4908 14111 5228 21019
rect 4908 13875 4950 14111
rect 5186 13875 5228 14111
rect 4908 12134 5228 13875
rect 11128 21255 11448 25696
rect 11128 21019 11170 21255
rect 11406 21019 11448 21255
rect 11128 14111 11448 21019
rect 11128 13875 11170 14111
rect 11406 13875 11448 14111
rect 11128 12134 11448 13875
rect 13878 24214 14198 25764
rect 19458 26000 19778 26024
rect 19458 25764 19500 26000
rect 19736 25764 19778 26000
rect 13878 23978 13920 24214
rect 14156 23978 14198 24214
rect 13878 22428 14198 23978
rect 13878 22192 13920 22428
rect 14156 22192 14198 22428
rect 13878 20642 14198 22192
rect 13878 20406 13920 20642
rect 14156 20406 14198 20642
rect 13878 18856 14198 20406
rect 13878 18620 13920 18856
rect 14156 18620 14198 18856
rect 13878 17070 14198 18620
rect 13878 16834 13920 17070
rect 14156 16834 14198 17070
rect 13878 15284 14198 16834
rect 13878 15048 13920 15284
rect 14156 15048 14198 15284
rect 13878 13498 14198 15048
rect 13878 13262 13920 13498
rect 14156 13262 14198 13498
rect 2158 11476 2200 11712
rect 2436 11476 2478 11712
rect 2158 9926 2478 11476
rect 13878 11712 14198 13262
rect 13878 11476 13920 11712
rect 14156 11476 14198 11712
rect 2158 9690 2200 9926
rect 2436 9690 2478 9926
rect 2158 8140 2478 9690
rect 2158 7904 2200 8140
rect 2436 7904 2478 8140
rect 2158 6354 2478 7904
rect 2158 6118 2200 6354
rect 2436 6118 2478 6354
rect 2158 4568 2478 6118
rect 4908 10608 5228 11408
rect 4908 10372 4950 10608
rect 5186 10372 5228 10608
rect 4908 7036 5228 10372
rect 4908 6800 4950 7036
rect 5186 6800 5228 7036
rect 4908 5250 5228 6800
rect 11128 10608 11448 11408
rect 11128 10372 11170 10608
rect 11406 10372 11448 10608
rect 11128 7036 11448 10372
rect 11128 6800 11170 7036
rect 11406 6800 11448 7036
rect 11128 5250 11448 6800
rect 13878 9926 14198 11476
rect 13878 9690 13920 9926
rect 14156 9690 14198 9926
rect 13878 8140 14198 9690
rect 13878 7904 13920 8140
rect 14156 7904 14198 8140
rect 13878 6354 14198 7904
rect 13878 6118 13920 6354
rect 14156 6118 14198 6354
rect 2158 4332 2200 4568
rect 2436 4332 2478 4568
rect 2158 2782 2478 4332
rect 13878 4568 14198 6118
rect 13878 4332 13920 4568
rect 14156 4332 14198 4568
rect 2158 2546 2200 2782
rect 2436 2546 2478 2782
rect 2158 996 2478 2546
rect 4908 3395 5228 4264
rect 4908 3159 4950 3395
rect 5186 3159 5228 3395
rect 4908 1609 5228 3159
rect 4908 1373 4950 1609
rect 5186 1373 5228 1609
rect 4908 1349 5228 1373
rect 11128 3395 11448 4264
rect 11128 3159 11170 3395
rect 11406 3159 11448 3395
rect 11128 1609 11448 3159
rect 11128 1373 11170 1609
rect 11406 1373 11448 1609
rect 11128 1349 11448 1373
rect 13878 2782 14198 4332
rect 13878 2546 13920 2782
rect 14156 2546 14198 2782
rect 2158 760 2200 996
rect 2436 760 2478 996
rect 2158 -790 2478 760
rect 13878 996 14198 2546
rect 13878 760 13920 996
rect 14156 760 14198 996
rect 4908 -177 5228 692
rect 4908 -413 4950 -177
rect 5186 -413 5228 -177
rect 4908 -437 5228 -413
rect 11128 -177 11448 692
rect 13878 -108 14198 760
rect 16708 19469 17028 25696
rect 16708 19233 16750 19469
rect 16986 19233 17028 19469
rect 16708 5181 17028 19233
rect 16708 4945 16750 5181
rect 16986 4945 17028 5181
rect 11128 -413 11170 -177
rect 11406 -413 11448 -177
rect 11128 -437 11448 -413
rect 2158 -1026 2200 -790
rect 2436 -1026 2478 -790
rect 2158 -1894 2478 -1026
rect 4908 -1894 5228 -1094
rect -34152 -2130 -34110 -1894
rect -33874 -2130 -33832 -1894
rect -34152 -2154 -33832 -2130
rect -28572 -2130 -28530 -1894
rect -28294 -2130 -28252 -1894
rect -28572 -2154 -28252 -2130
rect -22992 -2130 -22950 -1894
rect -22714 -2130 -22672 -1894
rect -22992 -2154 -22672 -2130
rect -17412 -2130 -17370 -1894
rect -17134 -2130 -17092 -1894
rect -17412 -2154 -17092 -2130
rect -11832 -2130 -11790 -1894
rect -11554 -2130 -11512 -1894
rect -11832 -2154 -11512 -2130
rect -6252 -2130 -6210 -1894
rect -5974 -2130 -5932 -1894
rect -6252 -2154 -5932 -2130
rect -672 -2130 -630 -1894
rect -394 -2130 -352 -1894
rect -672 -2154 -352 -2130
rect 4908 -2130 4950 -1894
rect 5186 -2130 5228 -1894
rect 4908 -2154 5228 -2130
rect 16708 -1894 17028 4945
rect 19458 24214 19778 25764
rect 25038 26000 25358 26024
rect 25038 25764 25080 26000
rect 25316 25764 25358 26000
rect 19458 23978 19500 24214
rect 19736 23978 19778 24214
rect 19458 22428 19778 23978
rect 19458 22192 19500 22428
rect 19736 22192 19778 22428
rect 19458 20642 19778 22192
rect 19458 20406 19500 20642
rect 19736 20406 19778 20642
rect 19458 18856 19778 20406
rect 19458 18620 19500 18856
rect 19736 18620 19778 18856
rect 19458 17070 19778 18620
rect 19458 16834 19500 17070
rect 19736 16834 19778 17070
rect 19458 15284 19778 16834
rect 19458 15048 19500 15284
rect 19736 15048 19778 15284
rect 19458 13498 19778 15048
rect 19458 13262 19500 13498
rect 19736 13262 19778 13498
rect 19458 11712 19778 13262
rect 19458 11476 19500 11712
rect 19736 11476 19778 11712
rect 19458 9926 19778 11476
rect 19458 9690 19500 9926
rect 19736 9690 19778 9926
rect 19458 8140 19778 9690
rect 19458 7904 19500 8140
rect 19736 7904 19778 8140
rect 19458 6354 19778 7904
rect 19458 6118 19500 6354
rect 19736 6118 19778 6354
rect 19458 4568 19778 6118
rect 19458 4332 19500 4568
rect 19736 4332 19778 4568
rect 19458 2782 19778 4332
rect 19458 2546 19500 2782
rect 19736 2546 19778 2782
rect 19458 996 19778 2546
rect 19458 760 19500 996
rect 19736 760 19778 996
rect 19458 -790 19778 760
rect 19458 -1026 19500 -790
rect 19736 -1026 19778 -790
rect 19458 -1894 19778 -1026
rect 22288 23041 22608 25696
rect 22288 22805 22330 23041
rect 22566 22805 22608 23041
rect 22288 8753 22608 22805
rect 22288 8517 22330 8753
rect 22566 8517 22608 8753
rect 22288 -1894 22608 8517
rect 25038 24214 25358 25764
rect 30618 26000 30938 26024
rect 30618 25764 30660 26000
rect 30896 25764 30938 26000
rect 25038 23978 25080 24214
rect 25316 23978 25358 24214
rect 25038 22428 25358 23978
rect 25038 22192 25080 22428
rect 25316 22192 25358 22428
rect 25038 20642 25358 22192
rect 25038 20406 25080 20642
rect 25316 20406 25358 20642
rect 25038 18856 25358 20406
rect 25038 18620 25080 18856
rect 25316 18620 25358 18856
rect 25038 17070 25358 18620
rect 25038 16834 25080 17070
rect 25316 16834 25358 17070
rect 25038 15284 25358 16834
rect 25038 15048 25080 15284
rect 25316 15048 25358 15284
rect 25038 13498 25358 15048
rect 25038 13262 25080 13498
rect 25316 13262 25358 13498
rect 25038 11712 25358 13262
rect 25038 11476 25080 11712
rect 25316 11476 25358 11712
rect 25038 9926 25358 11476
rect 25038 9690 25080 9926
rect 25316 9690 25358 9926
rect 25038 8140 25358 9690
rect 25038 7904 25080 8140
rect 25316 7904 25358 8140
rect 25038 6354 25358 7904
rect 25038 6118 25080 6354
rect 25316 6118 25358 6354
rect 25038 4568 25358 6118
rect 25038 4332 25080 4568
rect 25316 4332 25358 4568
rect 25038 2782 25358 4332
rect 25038 2546 25080 2782
rect 25316 2546 25358 2782
rect 25038 996 25358 2546
rect 25038 760 25080 996
rect 25316 760 25358 996
rect 25038 -790 25358 760
rect 25038 -1026 25080 -790
rect 25316 -1026 25358 -790
rect 25038 -1894 25358 -1026
rect 27868 23041 28188 25696
rect 27868 22805 27910 23041
rect 28146 22805 28188 23041
rect 27868 8753 28188 22805
rect 27868 8517 27910 8753
rect 28146 8517 28188 8753
rect 27868 -1894 28188 8517
rect 30618 24214 30938 25764
rect 36198 26000 36518 26024
rect 36198 25764 36240 26000
rect 36476 25764 36518 26000
rect 30618 23978 30660 24214
rect 30896 23978 30938 24214
rect 30618 22428 30938 23978
rect 30618 22192 30660 22428
rect 30896 22192 30938 22428
rect 30618 20642 30938 22192
rect 30618 20406 30660 20642
rect 30896 20406 30938 20642
rect 30618 18856 30938 20406
rect 30618 18620 30660 18856
rect 30896 18620 30938 18856
rect 30618 17070 30938 18620
rect 30618 16834 30660 17070
rect 30896 16834 30938 17070
rect 30618 15284 30938 16834
rect 30618 15048 30660 15284
rect 30896 15048 30938 15284
rect 30618 13498 30938 15048
rect 30618 13262 30660 13498
rect 30896 13262 30938 13498
rect 30618 11712 30938 13262
rect 30618 11476 30660 11712
rect 30896 11476 30938 11712
rect 30618 9926 30938 11476
rect 30618 9690 30660 9926
rect 30896 9690 30938 9926
rect 30618 8140 30938 9690
rect 30618 7904 30660 8140
rect 30896 7904 30938 8140
rect 30618 6354 30938 7904
rect 30618 6118 30660 6354
rect 30896 6118 30938 6354
rect 30618 4568 30938 6118
rect 30618 4332 30660 4568
rect 30896 4332 30938 4568
rect 30618 2782 30938 4332
rect 30618 2546 30660 2782
rect 30896 2546 30938 2782
rect 30618 996 30938 2546
rect 30618 760 30660 996
rect 30896 760 30938 996
rect 30618 -790 30938 760
rect 30618 -1026 30660 -790
rect 30896 -1026 30938 -790
rect 30618 -1894 30938 -1026
rect 33448 12325 33768 25696
rect 33448 12089 33490 12325
rect 33726 12089 33768 12325
rect 33448 -1894 33768 12089
rect 36198 24214 36518 25764
rect 41778 26000 42098 26024
rect 41778 25764 41820 26000
rect 42056 25764 42098 26000
rect 36198 23978 36240 24214
rect 36476 23978 36518 24214
rect 36198 22428 36518 23978
rect 36198 22192 36240 22428
rect 36476 22192 36518 22428
rect 36198 20642 36518 22192
rect 36198 20406 36240 20642
rect 36476 20406 36518 20642
rect 36198 18856 36518 20406
rect 36198 18620 36240 18856
rect 36476 18620 36518 18856
rect 36198 17070 36518 18620
rect 36198 16834 36240 17070
rect 36476 16834 36518 17070
rect 36198 15284 36518 16834
rect 36198 15048 36240 15284
rect 36476 15048 36518 15284
rect 36198 13498 36518 15048
rect 36198 13262 36240 13498
rect 36476 13262 36518 13498
rect 36198 11712 36518 13262
rect 36198 11476 36240 11712
rect 36476 11476 36518 11712
rect 36198 9926 36518 11476
rect 36198 9690 36240 9926
rect 36476 9690 36518 9926
rect 36198 8140 36518 9690
rect 36198 7904 36240 8140
rect 36476 7904 36518 8140
rect 36198 6354 36518 7904
rect 36198 6118 36240 6354
rect 36476 6118 36518 6354
rect 36198 4568 36518 6118
rect 36198 4332 36240 4568
rect 36476 4332 36518 4568
rect 36198 2782 36518 4332
rect 36198 2546 36240 2782
rect 36476 2546 36518 2782
rect 36198 996 36518 2546
rect 36198 760 36240 996
rect 36476 760 36518 996
rect 36198 -790 36518 760
rect 36198 -1026 36240 -790
rect 36476 -1026 36518 -790
rect 36198 -1894 36518 -1026
rect 39028 12325 39348 25696
rect 39028 12089 39070 12325
rect 39306 12089 39348 12325
rect 39028 -1894 39348 12089
rect 41778 24214 42098 25764
rect 47358 26000 47678 26024
rect 47358 25764 47400 26000
rect 47636 25764 47678 26000
rect 41778 23978 41820 24214
rect 42056 23978 42098 24214
rect 41778 22428 42098 23978
rect 41778 22192 41820 22428
rect 42056 22192 42098 22428
rect 41778 20642 42098 22192
rect 41778 20406 41820 20642
rect 42056 20406 42098 20642
rect 41778 18856 42098 20406
rect 41778 18620 41820 18856
rect 42056 18620 42098 18856
rect 41778 17070 42098 18620
rect 41778 16834 41820 17070
rect 42056 16834 42098 17070
rect 41778 15284 42098 16834
rect 41778 15048 41820 15284
rect 42056 15048 42098 15284
rect 41778 13498 42098 15048
rect 41778 13262 41820 13498
rect 42056 13262 42098 13498
rect 41778 11712 42098 13262
rect 41778 11476 41820 11712
rect 42056 11476 42098 11712
rect 41778 9926 42098 11476
rect 41778 9690 41820 9926
rect 42056 9690 42098 9926
rect 41778 8140 42098 9690
rect 41778 7904 41820 8140
rect 42056 7904 42098 8140
rect 41778 6354 42098 7904
rect 41778 6118 41820 6354
rect 42056 6118 42098 6354
rect 41778 4568 42098 6118
rect 41778 4332 41820 4568
rect 42056 4332 42098 4568
rect 41778 2782 42098 4332
rect 41778 2546 41820 2782
rect 42056 2546 42098 2782
rect 41778 996 42098 2546
rect 41778 760 41820 996
rect 42056 760 42098 996
rect 41778 -790 42098 760
rect 41778 -1026 41820 -790
rect 42056 -1026 42098 -790
rect 41778 -1894 42098 -1026
rect 44608 12325 44928 25696
rect 44608 12089 44650 12325
rect 44886 12089 44928 12325
rect 44608 -1894 44928 12089
rect 47358 24214 47678 25764
rect 52938 26000 53258 26024
rect 52938 25764 52980 26000
rect 53216 25764 53258 26000
rect 47358 23978 47400 24214
rect 47636 23978 47678 24214
rect 47358 22428 47678 23978
rect 47358 22192 47400 22428
rect 47636 22192 47678 22428
rect 47358 20642 47678 22192
rect 47358 20406 47400 20642
rect 47636 20406 47678 20642
rect 47358 18856 47678 20406
rect 47358 18620 47400 18856
rect 47636 18620 47678 18856
rect 47358 17070 47678 18620
rect 47358 16834 47400 17070
rect 47636 16834 47678 17070
rect 47358 15284 47678 16834
rect 47358 15048 47400 15284
rect 47636 15048 47678 15284
rect 47358 13498 47678 15048
rect 47358 13262 47400 13498
rect 47636 13262 47678 13498
rect 47358 11712 47678 13262
rect 47358 11476 47400 11712
rect 47636 11476 47678 11712
rect 47358 9926 47678 11476
rect 47358 9690 47400 9926
rect 47636 9690 47678 9926
rect 47358 8140 47678 9690
rect 47358 7904 47400 8140
rect 47636 7904 47678 8140
rect 47358 6354 47678 7904
rect 47358 6118 47400 6354
rect 47636 6118 47678 6354
rect 47358 4568 47678 6118
rect 47358 4332 47400 4568
rect 47636 4332 47678 4568
rect 47358 2782 47678 4332
rect 47358 2546 47400 2782
rect 47636 2546 47678 2782
rect 47358 996 47678 2546
rect 47358 760 47400 996
rect 47636 760 47678 996
rect 47358 -790 47678 760
rect 47358 -1026 47400 -790
rect 47636 -1026 47678 -790
rect 47358 -1894 47678 -1026
rect 50188 12325 50508 25696
rect 50188 12089 50230 12325
rect 50466 12089 50508 12325
rect 50188 -1894 50508 12089
rect 52938 24214 53258 25764
rect 52938 23978 52980 24214
rect 53216 23978 53258 24214
rect 52938 22428 53258 23978
rect 52938 22192 52980 22428
rect 53216 22192 53258 22428
rect 52938 20642 53258 22192
rect 52938 20406 52980 20642
rect 53216 20406 53258 20642
rect 52938 18856 53258 20406
rect 52938 18620 52980 18856
rect 53216 18620 53258 18856
rect 52938 17070 53258 18620
rect 52938 16834 52980 17070
rect 53216 16834 53258 17070
rect 52938 15284 53258 16834
rect 52938 15048 52980 15284
rect 53216 15048 53258 15284
rect 52938 13498 53258 15048
rect 52938 13262 52980 13498
rect 53216 13262 53258 13498
rect 52938 11712 53258 13262
rect 52938 11476 52980 11712
rect 53216 11476 53258 11712
rect 52938 9926 53258 11476
rect 52938 9690 52980 9926
rect 53216 9690 53258 9926
rect 52938 8140 53258 9690
rect 52938 7904 52980 8140
rect 53216 7904 53258 8140
rect 52938 6354 53258 7904
rect 52938 6118 52980 6354
rect 53216 6118 53258 6354
rect 52938 4568 53258 6118
rect 52938 4332 52980 4568
rect 53216 4332 53258 4568
rect 52938 2782 53258 4332
rect 52938 2546 52980 2782
rect 53216 2546 53258 2782
rect 52938 996 53258 2546
rect 52938 760 52980 996
rect 53216 760 53258 996
rect 52938 -790 53258 760
rect 52938 -1026 52980 -790
rect 53216 -1026 53258 -790
rect 52938 -1894 53258 -1026
rect 16708 -2130 16750 -1894
rect 16986 -2130 17028 -1894
rect 16708 -2154 17028 -2130
rect 22288 -2130 22330 -1894
rect 22566 -2130 22608 -1894
rect 22288 -2154 22608 -2130
rect 27868 -2130 27910 -1894
rect 28146 -2130 28188 -1894
rect 27868 -2154 28188 -2130
rect 33448 -2130 33490 -1894
rect 33726 -2130 33768 -1894
rect 33448 -2154 33768 -2130
rect 39028 -2130 39070 -1894
rect 39306 -2130 39348 -1894
rect 39028 -2154 39348 -2130
rect 44608 -2130 44650 -1894
rect 44886 -2130 44928 -1894
rect 44608 -2154 44928 -2130
rect 50188 -2130 50230 -1894
rect 50466 -2130 50508 -1894
rect 50188 -2154 50508 -2130
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_0
timestamp 1757093863
transform 1 0 -8573 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_1
timestamp 1757093863
transform 1 0 -8573 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_2
timestamp 1757093863
transform 1 0 -8573 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_3
timestamp 1757093863
transform 1 0 -8573 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_4
timestamp 1757093863
transform 1 0 -8573 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_5
timestamp 1757093863
transform 1 0 -8573 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_6
timestamp 1757093863
transform 1 0 -8573 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_7
timestamp 1757093863
transform 1 0 -8573 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_8
timestamp 1757093863
transform 1 0 -8573 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_9
timestamp 1757093863
transform 1 0 -8573 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_10
timestamp 1757093863
transform 1 0 -8573 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_11
timestamp 1757093863
transform 1 0 -8573 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_12
timestamp 1757093863
transform 1 0 -8573 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_13
timestamp 1757093863
transform 1 0 -8573 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_14
timestamp 1757093863
transform 1 0 -8573 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_15
timestamp 1757093863
transform 1 0 -30893 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_16
timestamp 1757093863
transform -1 0 19349 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_17
timestamp 1757093863
transform 1 0 2587 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_18
timestamp 1757093863
transform 1 0 2587 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_19
timestamp 1757093863
transform 1 0 2587 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_20
timestamp 1757093863
transform 1 0 2587 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_21
timestamp 1757093863
transform 1 0 2587 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_22
timestamp 1757093863
transform 1 0 2587 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_23
timestamp 1757093863
transform 1 0 2587 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_24
timestamp 1757093863
transform 1 0 2587 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_25
timestamp 1757093863
transform 1 0 2587 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_26
timestamp 1757093863
transform 1 0 2587 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_27
timestamp 1757093863
transform 1 0 2587 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_28
timestamp 1757093863
transform 1 0 2587 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_29
timestamp 1757093863
transform 1 0 2587 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_30
timestamp 1757093863
transform 1 0 2587 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_31
timestamp 1757093863
transform 1 0 2587 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_32
timestamp 1757093863
transform 1 0 -30893 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_33
timestamp 1757093863
transform 1 0 -2993 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_34
timestamp 1757093863
transform 1 0 -2993 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_35
timestamp 1757093863
transform 1 0 -2993 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_36
timestamp 1757093863
transform 1 0 -2993 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_37
timestamp 1757093863
transform 1 0 -2993 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_38
timestamp 1757093863
transform 1 0 -2993 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_39
timestamp 1757093863
transform 1 0 -2993 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_40
timestamp 1757093863
transform 1 0 -2993 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_41
timestamp 1757093863
transform 1 0 -2993 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_42
timestamp 1757093863
transform 1 0 -2993 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_43
timestamp 1757093863
transform 1 0 -2993 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_44
timestamp 1757093863
transform 1 0 -2993 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_45
timestamp 1757093863
transform 1 0 -2993 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_46
timestamp 1757093863
transform 1 0 -2993 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_47
timestamp 1757093863
transform 1 0 -2993 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_48
timestamp 1757093863
transform 1 0 -36473 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_49
timestamp 1757093863
transform 1 0 -14153 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_50
timestamp 1757093863
transform 1 0 -14153 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_51
timestamp 1757093863
transform 1 0 -36473 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_52
timestamp 1757093863
transform 1 0 -14153 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_53
timestamp 1757093863
transform 1 0 -14153 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_54
timestamp 1757093863
transform 1 0 -14153 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_55
timestamp 1757093863
transform 1 0 -14153 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_56
timestamp 1757093863
transform 1 0 -14153 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_57
timestamp 1757093863
transform 1 0 -14153 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_58
timestamp 1757093863
transform 1 0 -14153 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_59
timestamp 1757093863
transform 1 0 -14153 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_60
timestamp 1757093863
transform 1 0 -14153 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_61
timestamp 1757093863
transform 1 0 -14153 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_62
timestamp 1757093863
transform 1 0 -14153 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_63
timestamp 1757093863
transform 1 0 -14153 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_64
timestamp 1757093863
transform 1 0 -14153 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_65
timestamp 1757093863
transform 1 0 2587 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_66
timestamp 1757093863
transform 1 0 -2993 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_67
timestamp 1757093863
transform 1 0 -8573 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_68
timestamp 1757093863
transform 1 0 -14153 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_69
timestamp 1757093863
transform 1 0 -30893 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_70
timestamp 1757093863
transform 1 0 -30893 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_71
timestamp 1757093863
transform 1 0 -36473 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_72
timestamp 1757093863
transform 1 0 -36473 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_73
timestamp 1757093863
transform 1 0 -30893 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_74
timestamp 1757093863
transform 1 0 -30893 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_75
timestamp 1757093863
transform 1 0 -36473 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_76
timestamp 1757093863
transform 1 0 -36473 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_77
timestamp 1757093863
transform 1 0 -30893 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_78
timestamp 1757093863
transform 1 0 -30893 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_79
timestamp 1757093863
transform 1 0 -36473 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_80
timestamp 1757093863
transform 1 0 -36473 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_81
timestamp 1757093863
transform 1 0 -30893 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_82
timestamp 1757093863
transform 1 0 -30893 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_83
timestamp 1757093863
transform 1 0 -36473 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_84
timestamp 1757093863
transform 1 0 -36473 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_85
timestamp 1757093863
transform 1 0 -30893 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_86
timestamp 1757093863
transform 1 0 -30893 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_87
timestamp 1757093863
transform 1 0 -36473 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_88
timestamp 1757093863
transform 1 0 -36473 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_89
timestamp 1757093863
transform 1 0 -30893 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_90
timestamp 1757093863
transform 1 0 -30893 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_91
timestamp 1757093863
transform 1 0 -36473 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_92
timestamp 1757093863
transform 1 0 -36473 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_93
timestamp 1757093863
transform 1 0 -30893 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_94
timestamp 1757093863
transform 1 0 -30893 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_95
timestamp 1757093863
transform 1 0 -36473 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_96
timestamp 1757093863
transform 1 0 -36473 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_97
timestamp 1757093863
transform 1 0 -25313 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_98
timestamp 1757093863
transform 1 0 -25313 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_99
timestamp 1757093863
transform 1 0 -25313 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_100
timestamp 1757093863
transform 1 0 -25313 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_101
timestamp 1757093863
transform 1 0 -19733 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_102
timestamp 1757093863
transform 1 0 -19733 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_103
timestamp 1757093863
transform 1 0 -19733 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_104
timestamp 1757093863
transform 1 0 -19733 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_105
timestamp 1757093863
transform 1 0 -25313 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_106
timestamp 1757093863
transform 1 0 -25313 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_107
timestamp 1757093863
transform 1 0 -25313 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_108
timestamp 1757093863
transform 1 0 -25313 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_109
timestamp 1757093863
transform 1 0 -19733 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_110
timestamp 1757093863
transform 1 0 -19733 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_111
timestamp 1757093863
transform 1 0 -19733 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_112
timestamp 1757093863
transform 1 0 -19733 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_113
timestamp 1757093863
transform 1 0 -25313 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_114
timestamp 1757093863
transform 1 0 -25313 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_115
timestamp 1757093863
transform 1 0 -25313 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_116
timestamp 1757093863
transform 1 0 -19733 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_117
timestamp 1757093863
transform 1 0 -19733 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_118
timestamp 1757093863
transform 1 0 -19733 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_119
timestamp 1757093863
transform 1 0 -25313 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_120
timestamp 1757093863
transform 1 0 -25313 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_121
timestamp 1757093863
transform 1 0 -25313 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_122
timestamp 1757093863
transform 1 0 -25313 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_123
timestamp 1757093863
transform 1 0 -19733 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_124
timestamp 1757093863
transform 1 0 -19733 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_125
timestamp 1757093863
transform 1 0 -19733 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_126
timestamp 1757093863
transform 1 0 -19733 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_127
timestamp 1757093863
transform 1 0 -25313 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_128
timestamp 1757093863
transform 1 0 -19733 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_129
timestamp 1757093863
transform -1 0 52829 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_130
timestamp 1757093863
transform -1 0 47249 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_131
timestamp 1757093863
transform -1 0 41669 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_132
timestamp 1757093863
transform -1 0 36089 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_133
timestamp 1757093863
transform -1 0 30509 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_134
timestamp 1757093863
transform -1 0 24929 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_135
timestamp 1757093863
transform -1 0 19349 0 1 -1494
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_137
timestamp 1757093863
transform -1 0 52829 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_138
timestamp 1757093863
transform -1 0 47249 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_139
timestamp 1757093863
transform -1 0 41669 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_140
timestamp 1757093863
transform -1 0 36089 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_141
timestamp 1757093863
transform -1 0 30509 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_142
timestamp 1757093863
transform -1 0 24929 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_143
timestamp 1757093863
transform -1 0 19349 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_144
timestamp 1757093863
transform -1 0 13769 0 1 292
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_145
timestamp 1757093863
transform -1 0 52829 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_146
timestamp 1757093863
transform -1 0 47249 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_147
timestamp 1757093863
transform -1 0 41669 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_148
timestamp 1757093863
transform -1 0 36089 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_149
timestamp 1757093863
transform -1 0 30509 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_150
timestamp 1757093863
transform -1 0 24929 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_152
timestamp 1757093863
transform -1 0 13769 0 1 2078
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_153
timestamp 1757093863
transform -1 0 52829 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_154
timestamp 1757093863
transform -1 0 47249 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_155
timestamp 1757093863
transform -1 0 41669 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_156
timestamp 1757093863
transform -1 0 36089 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_157
timestamp 1757093863
transform -1 0 30509 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_158
timestamp 1757093863
transform -1 0 24929 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_159
timestamp 1757093863
transform -1 0 19349 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_160
timestamp 1757093863
transform -1 0 13769 0 1 3864
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_161
timestamp 1757093863
transform -1 0 52829 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_162
timestamp 1757093863
transform -1 0 47249 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_163
timestamp 1757093863
transform -1 0 41669 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_164
timestamp 1757093863
transform -1 0 36089 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_165
timestamp 1757093863
transform -1 0 30509 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_166
timestamp 1757093863
transform -1 0 24929 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_167
timestamp 1757093863
transform -1 0 19349 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_168
timestamp 1757093863
transform -1 0 13769 0 1 5650
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_169
timestamp 1757093863
transform -1 0 52829 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_170
timestamp 1757093863
transform -1 0 47249 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_171
timestamp 1757093863
transform -1 0 41669 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_172
timestamp 1757093863
transform -1 0 36089 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_173
timestamp 1757093863
transform -1 0 30509 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_174
timestamp 1757093863
transform -1 0 24929 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_175
timestamp 1757093863
transform -1 0 19349 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_176
timestamp 1757093863
transform -1 0 13769 0 1 7436
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_177
timestamp 1757093863
transform -1 0 52829 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_178
timestamp 1757093863
transform -1 0 47249 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_179
timestamp 1757093863
transform -1 0 41669 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_180
timestamp 1757093863
transform -1 0 36089 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_181
timestamp 1757093863
transform -1 0 30509 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_182
timestamp 1757093863
transform -1 0 24929 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_183
timestamp 1757093863
transform -1 0 19349 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_184
timestamp 1757093863
transform -1 0 13769 0 1 9222
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_185
timestamp 1757093863
transform -1 0 52829 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_186
timestamp 1757093863
transform -1 0 47249 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_187
timestamp 1757093863
transform -1 0 41669 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_188
timestamp 1757093863
transform -1 0 36089 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_189
timestamp 1757093863
transform -1 0 30509 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_190
timestamp 1757093863
transform -1 0 24929 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_191
timestamp 1757093863
transform -1 0 19349 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_192
timestamp 1757093863
transform -1 0 13769 0 1 11008
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_193
timestamp 1757093863
transform -1 0 52829 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_194
timestamp 1757093863
transform -1 0 47249 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_195
timestamp 1757093863
transform -1 0 41669 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_196
timestamp 1757093863
transform -1 0 36089 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_197
timestamp 1757093863
transform -1 0 30509 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_198
timestamp 1757093863
transform -1 0 24929 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_199
timestamp 1757093863
transform -1 0 19349 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_200
timestamp 1757093863
transform -1 0 13769 0 1 12794
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_201
timestamp 1757093863
transform -1 0 52829 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_202
timestamp 1757093863
transform -1 0 47249 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_203
timestamp 1757093863
transform -1 0 41669 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_204
timestamp 1757093863
transform -1 0 36089 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_205
timestamp 1757093863
transform -1 0 30509 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_206
timestamp 1757093863
transform -1 0 24929 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_207
timestamp 1757093863
transform -1 0 19349 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_208
timestamp 1757093863
transform -1 0 13769 0 1 14580
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_209
timestamp 1757093863
transform -1 0 52829 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_210
timestamp 1757093863
transform -1 0 47249 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_211
timestamp 1757093863
transform -1 0 41669 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_212
timestamp 1757093863
transform -1 0 36089 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_213
timestamp 1757093863
transform -1 0 30509 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_214
timestamp 1757093863
transform -1 0 24929 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_215
timestamp 1757093863
transform -1 0 19349 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_216
timestamp 1757093863
transform -1 0 13769 0 1 16366
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_217
timestamp 1757093863
transform -1 0 52829 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_218
timestamp 1757093863
transform -1 0 47249 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_219
timestamp 1757093863
transform -1 0 41669 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_220
timestamp 1757093863
transform -1 0 36089 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_221
timestamp 1757093863
transform -1 0 30509 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_222
timestamp 1757093863
transform -1 0 24929 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_223
timestamp 1757093863
transform -1 0 19349 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_224
timestamp 1757093863
transform -1 0 13769 0 1 18152
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_225
timestamp 1757093863
transform -1 0 52829 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_226
timestamp 1757093863
transform -1 0 47249 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_227
timestamp 1757093863
transform -1 0 41669 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_228
timestamp 1757093863
transform -1 0 36089 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_229
timestamp 1757093863
transform -1 0 30509 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_230
timestamp 1757093863
transform -1 0 24929 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_231
timestamp 1757093863
transform -1 0 19349 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_232
timestamp 1757093863
transform -1 0 13769 0 1 19938
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_233
timestamp 1757093863
transform -1 0 52829 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_234
timestamp 1757093863
transform -1 0 47249 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_235
timestamp 1757093863
transform -1 0 41669 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_236
timestamp 1757093863
transform -1 0 36089 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_237
timestamp 1757093863
transform -1 0 30509 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_238
timestamp 1757093863
transform -1 0 24929 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_239
timestamp 1757093863
transform -1 0 19349 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_240
timestamp 1757093863
transform -1 0 13769 0 1 21724
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_241
timestamp 1757093863
transform -1 0 52829 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_242
timestamp 1757093863
transform -1 0 47249 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_243
timestamp 1757093863
transform -1 0 41669 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_244
timestamp 1757093863
transform -1 0 36089 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_245
timestamp 1757093863
transform -1 0 30509 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_246
timestamp 1757093863
transform -1 0 24929 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_247
timestamp 1757093863
transform -1 0 19349 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_248
timestamp 1757093863
transform -1 0 13769 0 1 23510
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_249
timestamp 1757093863
transform -1 0 13769 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_250
timestamp 1757093863
transform -1 0 19349 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_251
timestamp 1757093863
transform -1 0 24929 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_252
timestamp 1757093863
transform -1 0 30509 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_253
timestamp 1757093863
transform -1 0 36089 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_254
timestamp 1757093863
transform -1 0 41669 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_255
timestamp 1757093863
transform -1 0 47249 0 1 25296
box -2619 -281 2641 281
use sky130_fd_pr__cap_mim_m3_2_XAJUMH  sky130_fd_pr__cap_mim_m3_2_XAJUMH_256
timestamp 1757093863
transform -1 0 52829 0 1 25296
box -2619 -281 2641 281
use switch  switch_0
timestamp 1757093863
transform 1 0 7876 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_1
timestamp 1757093863
transform 1 0 19708 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_2
timestamp 1757093863
transform 1 0 11820 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_3
timestamp 1757093863
transform 1 0 -7900 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_4
timestamp 1757093863
transform 1 0 3932 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_5
timestamp 1757093863
transform 1 0 -12 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_6
timestamp 1757093863
transform 1 0 -3956 0 1 -5198
box 1296 -1584 3268 244
use switch  switch_7
timestamp 1757093863
transform 1 0 15764 0 1 -5198
box 1296 -1584 3268 244
<< labels >>
flabel metal5 52938 -1894 53258 26024 0 FreeSans 160 90 0 0 OUT
port 9 nsew
flabel metal1 -6604 -5000 22976 -4954 0 FreeSans 160 0 0 0 VDD
port 10 nsew
flabel metal1 -6604 -6782 22976 -6736 0 FreeSans 160 0 0 0 GND
port 8 nsew
flabel metal1 -5641 -5930 -4981 -5884 0 FreeSans 160 0 0 0 b0
port 0 nsew
flabel metal1 -1697 -5930 -1037 -5884 0 FreeSans 160 0 0 0 b1
port 1 nsew
flabel metal1 2247 -5930 2907 -5884 0 FreeSans 160 0 0 0 b2
port 2 nsew
flabel metal1 6191 -5930 6851 -5884 0 FreeSans 160 0 0 0 b3
port 3 nsew
flabel metal1 10135 -5930 10795 -5884 0 FreeSans 160 0 0 0 b4
port 4 nsew
flabel metal1 14079 -5930 14739 -5884 0 FreeSans 160 0 0 0 b5
port 5 nsew
flabel metal1 18023 -5930 18683 -5884 0 FreeSans 160 0 0 0 b6
port 6 nsew
flabel metal1 21967 -5930 22627 -5884 0 FreeSans 160 0 0 0 b7
port 7 nsew
<< end >>
