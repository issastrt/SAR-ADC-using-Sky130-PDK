magic
tech sky130A
magscale 1 2
timestamp 1756382177
<< nwell >>
rect 29235 16606 29951 18606
<< pwell >>
rect 27899 -2020 27965 -1964
rect 28952 -2020 29018 -1964
<< locali >>
rect 27657 29240 28743 29246
rect 27657 29206 27663 29240
rect 28737 29206 28743 29240
rect 27657 29088 28743 29206
rect 29313 29240 29873 29246
rect 29313 29206 29319 29240
rect 29867 29206 29873 29240
rect 29313 29088 29873 29206
rect 25211 -1970 26617 -1894
rect 25211 -2004 25217 -1970
rect 26611 -2004 26617 -1970
rect 25211 -2010 26617 -2004
rect 27523 -1970 28609 -1882
rect 27523 -2004 27529 -1970
rect 28603 -2004 28609 -1970
rect 27523 -2010 28609 -2004
rect 29361 -1970 29921 -1882
rect 29361 -2004 29367 -1970
rect 29915 -2004 29921 -1970
rect 29361 -2010 29921 -2004
<< viali >>
rect 27663 29206 28737 29240
rect 29319 29206 29867 29240
rect 25217 -2004 26611 -1970
rect 27529 -2004 28603 -1970
rect 29367 -2004 29915 -1970
<< metal1 >>
rect 25175 29240 29951 29246
rect 25175 29206 27663 29240
rect 28737 29206 29319 29240
rect 29867 29206 29951 29240
rect 25175 29200 29951 29206
rect 25341 28832 26487 29200
rect 28177 28903 28223 29200
rect 29391 28903 29437 29200
rect 28089 28857 28311 28903
rect 29391 28857 29441 28903
rect 26057 28818 26103 28832
rect 27776 18957 27840 18963
rect 27776 18905 27782 18957
rect 27834 18905 27840 18957
rect 27776 18899 27840 18905
rect 28560 18957 28624 18963
rect 28560 18905 28566 18957
rect 28618 18905 28624 18957
rect 28560 18899 28624 18905
rect 27905 18865 27969 18871
rect 27905 18813 27911 18865
rect 27963 18813 27969 18865
rect 27905 18807 27969 18813
rect 28431 18865 28495 18871
rect 28431 18813 28437 18865
rect 28489 18813 28495 18865
rect 28431 18807 28495 18813
rect 29690 16957 29754 16963
rect 29690 16905 29696 16957
rect 29748 16905 29754 16957
rect 29690 16899 29754 16905
rect 29561 16865 29625 16871
rect 29561 16813 29567 16865
rect 29619 16813 29625 16865
rect 29561 16807 29625 16813
rect 27905 12160 27969 12166
rect 27905 12108 27911 12160
rect 27963 12108 27969 12160
rect 27905 12102 27969 12108
rect 27776 12077 27840 12083
rect 27776 12025 27782 12077
rect 27834 12025 27840 12077
rect 27776 12019 27840 12025
rect 28560 12077 28624 12083
rect 28560 12025 28566 12077
rect 28618 12025 28624 12077
rect 28560 12019 28624 12025
rect 28034 9133 28098 9139
rect 28034 9081 28040 9133
rect 28092 9081 28098 9133
rect 28034 9075 28098 9081
rect 28302 9133 28366 9139
rect 28302 9081 28308 9133
rect 28360 9081 28366 9133
rect 28302 9075 28366 9081
rect 28431 9050 28495 9056
rect 28431 8998 28437 9050
rect 28489 8998 28495 9050
rect 28431 8992 28495 8998
rect 28167 2292 28231 2298
rect 28167 2240 28173 2292
rect 28225 2240 28231 2292
rect 28167 2234 28231 2240
rect 29738 292 29802 298
rect 29738 240 29744 292
rect 29796 240 29802 292
rect 29738 234 29802 240
rect 26378 -1652 26442 -1646
rect 26378 -1704 26384 -1652
rect 26436 -1704 26442 -1652
rect 26378 -1710 26442 -1704
rect 27642 -1652 27706 -1646
rect 27642 -1704 27648 -1652
rect 27700 -1704 27706 -1652
rect 27642 -1710 27706 -1704
rect 27900 -1652 27964 -1646
rect 27900 -1704 27906 -1652
rect 27958 -1704 27964 -1652
rect 27900 -1710 27964 -1704
rect 28426 -1652 28490 -1646
rect 28426 -1704 28432 -1652
rect 28484 -1704 28490 -1652
rect 28426 -1710 28490 -1704
rect 29480 -1652 29544 -1646
rect 29480 -1704 29486 -1652
rect 29538 -1704 29544 -1652
rect 29480 -1710 29544 -1704
rect 27651 -1738 27697 -1710
rect 27651 -1784 29737 -1738
rect 27900 -1961 27964 -1955
rect 27900 -1964 27906 -1961
rect 25175 -1970 27906 -1964
rect 27958 -1964 27964 -1961
rect 28953 -1961 29017 -1955
rect 28953 -1964 28959 -1961
rect 27958 -1970 28959 -1964
rect 25175 -2004 25217 -1970
rect 26611 -2004 27529 -1970
rect 28603 -2004 28959 -1970
rect 25175 -2010 27906 -2004
rect 27900 -2013 27906 -2010
rect 27958 -2010 28959 -2004
rect 27958 -2013 27964 -2010
rect 27900 -2019 27964 -2013
rect 28953 -2013 28959 -2010
rect 29011 -1964 29017 -1961
rect 29011 -1970 29969 -1964
rect 29011 -2004 29367 -1970
rect 29915 -2004 29969 -1970
rect 29011 -2010 29969 -2004
rect 29011 -2013 29017 -2010
rect 28953 -2019 29017 -2013
<< via1 >>
rect 27782 18905 27834 18957
rect 28566 18905 28618 18957
rect 27911 18813 27963 18865
rect 28437 18813 28489 18865
rect 29696 16905 29748 16957
rect 29567 16813 29619 16865
rect 27911 12108 27963 12160
rect 27782 12025 27834 12077
rect 28566 12025 28618 12077
rect 28040 9081 28092 9133
rect 28308 9081 28360 9133
rect 28437 8998 28489 9050
rect 28173 2240 28225 2292
rect 29744 240 29796 292
rect 26384 -1704 26436 -1652
rect 27648 -1704 27700 -1652
rect 27906 -1704 27958 -1652
rect 28432 -1704 28484 -1652
rect 29486 -1704 29538 -1652
rect 27906 -1970 27958 -1961
rect 27906 -2004 27958 -1970
rect 27906 -2013 27958 -2004
rect 28959 -2013 29011 -1961
<< metal2 >>
rect 27771 18959 27845 18968
rect 27771 18903 27780 18959
rect 27836 18903 27845 18959
rect 27771 18867 27845 18903
rect 28555 18959 28629 18968
rect 28555 18903 28564 18959
rect 28620 18903 28629 18959
rect 28555 18894 28629 18903
rect 27771 18811 27780 18867
rect 27836 18862 27845 18867
rect 27905 18865 27969 18871
rect 27905 18862 27911 18865
rect 27836 18816 27911 18862
rect 27836 18811 27845 18816
rect 27771 18802 27845 18811
rect 27905 18813 27911 18816
rect 27963 18862 27969 18865
rect 28431 18865 28495 18871
rect 28431 18862 28437 18865
rect 27963 18816 28437 18862
rect 27963 18813 27969 18816
rect 27905 18807 27969 18813
rect 28431 18813 28437 18816
rect 28489 18813 28495 18865
rect 28431 18807 28495 18813
rect 29690 16957 29754 16963
rect 29690 16905 29696 16957
rect 29748 16954 29754 16957
rect 30164 16959 30238 16968
rect 30164 16954 30173 16959
rect 29748 16908 30173 16954
rect 29748 16905 29754 16908
rect 29690 16899 29754 16905
rect 30164 16903 30173 16908
rect 30229 16903 30238 16959
rect 30164 16894 30238 16903
rect 28555 16867 28629 16876
rect 28555 16811 28564 16867
rect 28620 16862 28629 16867
rect 29556 16867 29630 16876
rect 29556 16862 29565 16867
rect 28620 16816 29565 16862
rect 28620 16811 28629 16816
rect 28555 16802 28629 16811
rect 29556 16811 29565 16816
rect 29621 16811 29630 16867
rect 29556 16802 29630 16811
rect 27900 12162 27974 12171
rect 27900 12106 27909 12162
rect 27965 12106 27974 12162
rect 27900 12097 27974 12106
rect 27771 12079 27845 12088
rect 27771 12023 27780 12079
rect 27836 12023 27845 12079
rect 27771 12014 27845 12023
rect 28555 12079 28629 12088
rect 28555 12023 28564 12079
rect 28620 12023 28629 12079
rect 28555 12014 28629 12023
rect 28034 9133 28098 9139
rect 28034 9081 28040 9133
rect 28092 9130 28098 9133
rect 28163 9135 28237 9144
rect 28163 9130 28172 9135
rect 28092 9084 28172 9130
rect 28092 9081 28098 9084
rect 28034 9075 28098 9081
rect 28163 9079 28172 9084
rect 28228 9130 28237 9135
rect 28302 9133 28366 9139
rect 28302 9130 28308 9133
rect 28228 9084 28308 9130
rect 28228 9079 28237 9084
rect 28163 9070 28237 9079
rect 28302 9081 28308 9084
rect 28360 9081 28366 9133
rect 28302 9075 28366 9081
rect 28426 9052 28500 9061
rect 28426 8996 28435 9052
rect 28491 8996 28500 9052
rect 28426 8987 28500 8996
rect 28162 2294 28236 2303
rect 28162 2238 28171 2294
rect 28227 2238 28236 2294
rect 28162 2229 28236 2238
rect 29738 292 29802 298
rect 29738 240 29744 292
rect 29796 289 29802 292
rect 30164 294 30238 303
rect 30164 289 30173 294
rect 29796 243 30173 289
rect 29796 240 29802 243
rect 29738 234 29802 240
rect 30164 238 30173 243
rect 30229 238 30238 294
rect 30164 229 30238 238
rect 26378 -1652 26442 -1646
rect 26378 -1704 26384 -1652
rect 26436 -1655 26442 -1652
rect 27642 -1652 27706 -1646
rect 27642 -1655 27648 -1652
rect 26436 -1701 27648 -1655
rect 26436 -1704 26442 -1701
rect 26378 -1710 26442 -1704
rect 27642 -1704 27648 -1701
rect 27700 -1704 27706 -1652
rect 27642 -1710 27706 -1704
rect 27895 -1650 27969 -1641
rect 27895 -1706 27904 -1650
rect 27960 -1655 27969 -1650
rect 28426 -1652 28490 -1646
rect 28426 -1655 28432 -1652
rect 27960 -1701 28432 -1655
rect 27960 -1706 27969 -1701
rect 27895 -1715 27969 -1706
rect 28426 -1704 28432 -1701
rect 28484 -1655 28490 -1652
rect 28948 -1650 29022 -1641
rect 28948 -1655 28957 -1650
rect 28484 -1701 28957 -1655
rect 28484 -1704 28490 -1701
rect 28426 -1710 28490 -1704
rect 28948 -1706 28957 -1701
rect 29013 -1655 29022 -1650
rect 29480 -1652 29544 -1646
rect 29480 -1655 29486 -1652
rect 29013 -1701 29486 -1655
rect 29013 -1706 29022 -1701
rect 28948 -1715 29022 -1706
rect 29480 -1704 29486 -1701
rect 29538 -1704 29544 -1652
rect 29480 -1710 29544 -1704
rect 27895 -1959 27969 -1950
rect 27895 -2015 27904 -1959
rect 27960 -2015 27969 -1959
rect 27895 -2024 27969 -2015
rect 28948 -1959 29022 -1950
rect 28948 -2015 28957 -1959
rect 29013 -2015 29022 -1959
rect 28948 -2024 29022 -2015
<< via2 >>
rect 27780 18957 27836 18959
rect 27780 18905 27782 18957
rect 27782 18905 27834 18957
rect 27834 18905 27836 18957
rect 27780 18903 27836 18905
rect 28564 18957 28620 18959
rect 28564 18905 28566 18957
rect 28566 18905 28618 18957
rect 28618 18905 28620 18957
rect 28564 18903 28620 18905
rect 27780 18811 27836 18867
rect 30173 16903 30229 16959
rect 28564 16811 28620 16867
rect 29565 16865 29621 16867
rect 29565 16813 29567 16865
rect 29567 16813 29619 16865
rect 29619 16813 29621 16865
rect 29565 16811 29621 16813
rect 27909 12160 27965 12162
rect 27909 12108 27911 12160
rect 27911 12108 27963 12160
rect 27963 12108 27965 12160
rect 27909 12106 27965 12108
rect 27780 12077 27836 12079
rect 27780 12025 27782 12077
rect 27782 12025 27834 12077
rect 27834 12025 27836 12077
rect 27780 12023 27836 12025
rect 28564 12077 28620 12079
rect 28564 12025 28566 12077
rect 28566 12025 28618 12077
rect 28618 12025 28620 12077
rect 28564 12023 28620 12025
rect 28172 9079 28228 9135
rect 28435 9050 28491 9052
rect 28435 8998 28437 9050
rect 28437 8998 28489 9050
rect 28489 8998 28491 9050
rect 28435 8996 28491 8998
rect 28171 2292 28227 2294
rect 28171 2240 28173 2292
rect 28173 2240 28225 2292
rect 28225 2240 28227 2292
rect 28171 2238 28227 2240
rect 30173 238 30229 294
rect 27904 -1652 27960 -1650
rect 27904 -1704 27906 -1652
rect 27906 -1704 27958 -1652
rect 27958 -1704 27960 -1652
rect 27904 -1706 27960 -1704
rect 28957 -1706 29013 -1650
rect 27904 -1961 27960 -1959
rect 27904 -2013 27906 -1961
rect 27906 -2013 27958 -1961
rect 27958 -2013 27960 -1961
rect 27904 -2015 27960 -2013
rect 28957 -1961 29013 -1959
rect 28957 -2013 28959 -1961
rect 28959 -2013 29011 -1961
rect 29011 -2013 29013 -1961
rect 28957 -2015 29013 -2013
<< metal3 >>
rect 27775 18959 27841 18964
rect 27775 18903 27780 18959
rect 27836 18903 27841 18959
rect 27775 18867 27841 18903
rect 28559 18959 28625 18964
rect 28559 18903 28564 18959
rect 28620 18903 28625 18959
rect 28559 18898 28625 18903
rect 27775 18811 27780 18867
rect 27836 18811 27841 18867
rect 27775 18806 27841 18811
rect 27778 12084 27838 18806
rect 28562 16872 28622 18898
rect 30168 16959 30234 16964
rect 30168 16903 30173 16959
rect 30229 16903 30234 16959
rect 30168 16898 30234 16903
rect 28559 16867 28625 16872
rect 28559 16811 28564 16867
rect 28620 16811 28625 16867
rect 28559 16806 28625 16811
rect 29560 16867 29626 16872
rect 29560 16811 29565 16867
rect 29621 16811 29626 16867
rect 29560 16806 29626 16811
rect 27899 12475 27975 12481
rect 27899 12411 27905 12475
rect 27969 12411 27975 12475
rect 27899 12405 27975 12411
rect 27907 12167 27967 12405
rect 27904 12162 27970 12167
rect 27904 12106 27909 12162
rect 27965 12106 27970 12162
rect 27904 12101 27970 12106
rect 28562 12084 28622 16806
rect 29563 13429 29623 16806
rect 29555 13423 29631 13429
rect 29555 13359 29561 13423
rect 29625 13359 29631 13423
rect 29555 13353 29631 13359
rect 27775 12079 27841 12084
rect 27775 12023 27780 12079
rect 27836 12023 27841 12079
rect 27775 12018 27841 12023
rect 28559 12079 28625 12084
rect 28559 12023 28564 12079
rect 28620 12023 28625 12079
rect 28559 12018 28625 12023
rect 30171 11311 30231 16898
rect 30163 11305 30239 11311
rect 30163 11241 30169 11305
rect 30233 11241 30239 11305
rect 30163 11235 30239 11241
rect 28167 9135 28233 9140
rect 28167 9079 28172 9135
rect 28228 9079 28233 9135
rect 28167 9074 28233 9079
rect 28170 2299 28230 9074
rect 28430 9052 28496 9057
rect 28430 8996 28435 9052
rect 28491 8996 28496 9052
rect 28430 8991 28496 8996
rect 28433 8753 28493 8991
rect 28425 8747 28501 8753
rect 28425 8683 28431 8747
rect 28495 8683 28501 8747
rect 28425 8677 28501 8683
rect 28947 5357 29023 5363
rect 28947 5293 28953 5357
rect 29017 5293 29023 5357
rect 28947 5287 29023 5293
rect 28166 2294 28232 2299
rect 28166 2238 28171 2294
rect 28227 2238 28232 2294
rect 28166 2233 28232 2238
rect 28955 -1645 29015 5287
rect 30171 299 30231 11235
rect 30168 294 30234 299
rect 30168 238 30173 294
rect 30229 238 30234 294
rect 30168 233 30234 238
rect 27899 -1650 27965 -1645
rect 27899 -1706 27904 -1650
rect 27960 -1706 27965 -1650
rect 27899 -1711 27965 -1706
rect 28952 -1650 29018 -1645
rect 28952 -1706 28957 -1650
rect 29013 -1706 29018 -1650
rect 28952 -1711 29018 -1706
rect 27902 -1954 27962 -1711
rect 28955 -1954 29015 -1711
rect 27899 -1959 27965 -1954
rect 27899 -2015 27904 -1959
rect 27960 -2015 27965 -1959
rect 27899 -2020 27965 -2015
rect 28952 -1959 29018 -1954
rect 28952 -2015 28957 -1959
rect 29013 -2015 29018 -1959
rect 28952 -2020 29018 -2015
<< via3 >>
rect 27905 12411 27969 12475
rect 29561 13359 29625 13423
rect 30169 11241 30233 11305
rect 28431 8683 28495 8747
rect 28953 5293 29017 5357
<< via4 >>
rect 29475 13423 29711 13509
rect 29475 13359 29561 13423
rect 29561 13359 29625 13423
rect 29625 13359 29711 13423
rect 29475 13273 29711 13359
rect 27819 12475 28055 12561
rect 27819 12411 27905 12475
rect 27905 12411 27969 12475
rect 27969 12411 28055 12475
rect 27819 12325 28055 12411
rect 30083 11305 30319 11391
rect 30083 11241 30169 11305
rect 30169 11241 30233 11305
rect 30233 11241 30319 11305
rect 30083 11155 30319 11241
rect 28345 8747 28581 8833
rect 28345 8683 28431 8747
rect 28431 8683 28495 8747
rect 28495 8683 28581 8747
rect 28345 8597 28581 8683
rect 28867 5357 29103 5443
rect 28867 5293 28953 5357
rect 28953 5293 29017 5357
rect 29017 5293 29103 5357
rect 28867 5207 29103 5293
<< metal5 >>
rect 29433 13509 29753 13533
rect 29433 13273 29475 13509
rect 29711 13273 29753 13509
rect 27777 12561 28097 12881
rect 27777 12325 27819 12561
rect 28055 12325 28097 12561
rect 27777 12301 28097 12325
rect 29433 12128 29753 13273
rect 29103 11391 30343 11433
rect 29103 11155 30083 11391
rect 30319 11155 30343 11391
rect 29103 11113 30343 11155
rect 28303 8833 28623 8857
rect 28303 8597 28345 8833
rect 28581 8597 28623 8833
rect 28303 8277 28623 8597
rect 29433 6180 29753 11113
rect 28835 5443 30165 5485
rect 28835 5207 28867 5443
rect 29103 5207 30165 5443
rect 28835 5165 30165 5207
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_0
timestamp 1755260286
transform 0 1 29593 -1 0 6071
box -884 -281 906 281
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_1
timestamp 1755260286
transform 0 1 29593 -1 0 12019
box -884 -281 906 281
use sky130_fd_pr__res_xhigh_po_5p73_2WP2GG  sky130_fd_pr__res_xhigh_po_5p73_2WP2GG_0
timestamp 1756382177
transform 1 0 25914 0 1 13618
box -739 -15582 739 15582
use sky130_fd_pr__nfet_g5v0d10v5_Q3MXVW  XM1
timestamp 1755260286
transform 1 0 27937 0 1 10579
box -328 -1758 328 1758
use sky130_fd_pr__nfet_g5v0d10v5_Q3MXVW  XM2
timestamp 1755260286
transform 1 0 28463 0 1 10579
box -328 -1758 328 1758
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM3
timestamp 1755260286
transform 1 0 27937 0 1 23903
box -358 -5297 358 5297
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM4
timestamp 1755260286
transform 1 0 28463 0 1 23903
box -358 -5297 358 5297
use sky130_fd_pr__nfet_g5v0d10v5_53M7DK  XM5
timestamp 1755260286
transform 1 0 28329 0 1 294
box -328 -2258 328 2258
use sky130_fd_pr__nfet_g5v0d10v5_Q3M7H8  XM6
timestamp 1755260286
transform 1 0 29641 0 1 -706
box -328 -1258 328 1258
use sky130_fd_pr__nfet_g5v0d10v5_53M7DK  XM7
timestamp 1755260286
transform 1 0 27803 0 1 294
box -328 -2258 328 2258
use sky130_fd_pr__pfet_g5v0d10v5_UX3D7Q  XM9
timestamp 1755260286
transform 1 0 29593 0 1 22903
box -358 -6297 358 6297
<< labels >>
flabel metal5 27777 12561 28097 12881 0 FreeSans 800 0 0 0 Vinm
port 3 nsew
flabel metal5 28303 8277 28623 8597 0 FreeSans 800 0 0 0 Vinp
port 4 nsew
flabel metal5 29433 6180 29753 10857 0 FreeSans 800 0 0 0 Vout
port 5 nsew
flabel metal1 25341 29200 29951 29246 0 FreeSans 160 0 0 0 VDD
port 2 nsew
flabel metal1 25175 -2010 27906 -1964 0 FreeSans 160 0 0 0 VSS
port 6 nsew
<< end >>
