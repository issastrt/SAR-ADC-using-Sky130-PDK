magic
tech sky130A
magscale 1 2
timestamp 1757226903
<< metal1 >>
rect 1861 -9936 1925 -9930
rect 1861 -9988 1867 -9936
rect 1919 -9988 1925 -9936
rect 1861 -9994 1925 -9988
rect 2304 -11944 2368 -11938
rect 2304 -11996 2310 -11944
rect 2362 -11996 2368 -11944
rect 2304 -12002 2368 -11996
rect 2010 -13500 2074 -13494
rect 2010 -13503 2016 -13500
rect 2005 -13549 2016 -13503
rect 2010 -13552 2016 -13549
rect 2068 -13503 2074 -13500
rect 2068 -13549 2079 -13503
rect 2068 -13552 2074 -13549
rect 2010 -13558 2074 -13552
rect 2304 -15508 2368 -15502
rect 2304 -15560 2310 -15508
rect 2362 -15560 2368 -15508
rect 2304 -15566 2368 -15560
rect 2010 -17064 2074 -17058
rect 2010 -17067 2016 -17064
rect 2005 -17113 2016 -17067
rect 2010 -17116 2016 -17113
rect 2068 -17067 2074 -17064
rect 2068 -17113 2079 -17067
rect 2068 -17116 2074 -17113
rect 2010 -17122 2074 -17116
rect 2304 -19072 2368 -19066
rect 2304 -19124 2310 -19072
rect 2362 -19124 2368 -19072
rect 2304 -19130 2368 -19124
rect 2010 -20628 2074 -20622
rect 2010 -20631 2016 -20628
rect 2005 -20677 2016 -20631
rect 2010 -20680 2016 -20677
rect 2068 -20631 2074 -20628
rect 2068 -20677 2079 -20631
rect 2068 -20680 2074 -20677
rect 2010 -20686 2074 -20680
rect 2304 -22636 2368 -22630
rect 2304 -22688 2310 -22636
rect 2362 -22688 2368 -22636
rect 2304 -22694 2368 -22688
rect 2010 -24192 2074 -24186
rect 2010 -24195 2016 -24192
rect 2005 -24241 2016 -24195
rect 2010 -24244 2016 -24241
rect 2068 -24195 2074 -24192
rect 2068 -24241 2079 -24195
rect 2068 -24244 2074 -24241
rect 2010 -24250 2074 -24244
rect 2304 -26200 2368 -26194
rect 2304 -26252 2310 -26200
rect 2362 -26252 2368 -26200
rect 2304 -26258 2368 -26252
rect 2010 -27756 2074 -27750
rect 2010 -27759 2016 -27756
rect 2005 -27805 2016 -27759
rect 2010 -27808 2016 -27805
rect 2068 -27759 2074 -27756
rect 2068 -27805 2079 -27759
rect 2068 -27808 2074 -27805
rect 2010 -27814 2074 -27808
rect 2304 -29764 2368 -29758
rect 2304 -29816 2310 -29764
rect 2362 -29816 2368 -29764
rect 2304 -29822 2368 -29816
rect 2010 -31320 2074 -31314
rect 2010 -31323 2016 -31320
rect 2005 -31369 2016 -31323
rect 2010 -31372 2016 -31369
rect 2068 -31323 2074 -31320
rect 2068 -31369 2079 -31323
rect 2068 -31372 2074 -31369
rect 2010 -31378 2074 -31372
rect 2304 -33328 2368 -33322
rect 2304 -33380 2310 -33328
rect 2362 -33380 2368 -33328
rect 2304 -33386 2368 -33380
rect 2010 -34884 2074 -34878
rect 2010 -34887 2016 -34884
rect 2005 -34933 2016 -34887
rect 2010 -34936 2016 -34933
rect 2068 -34887 2074 -34884
rect 2068 -34933 2079 -34887
rect 2068 -34936 2074 -34933
rect 2010 -34942 2074 -34936
rect 2304 -36892 2368 -36886
rect 2304 -36944 2310 -36892
rect 2362 -36944 2368 -36892
rect 2304 -36950 2368 -36944
rect 2010 -38448 2074 -38442
rect 2010 -38451 2016 -38448
rect 2005 -38497 2016 -38451
rect 2010 -38500 2016 -38497
rect 2068 -38451 2074 -38448
rect 2068 -38497 2079 -38451
rect 2068 -38500 2074 -38497
rect 2010 -38506 2074 -38500
rect 2304 -40456 2368 -40450
rect 2304 -40508 2310 -40456
rect 2362 -40508 2368 -40456
rect 2304 -40514 2368 -40508
rect 2010 -42012 2074 -42006
rect 2010 -42015 2016 -42012
rect 2005 -42061 2016 -42015
rect 2010 -42064 2016 -42061
rect 2068 -42015 2074 -42012
rect 2068 -42061 2079 -42015
rect 2068 -42064 2074 -42061
rect 2010 -42070 2074 -42064
rect 2304 -44020 2368 -44014
rect 2304 -44072 2310 -44020
rect 2362 -44072 2368 -44020
rect 2304 -44078 2368 -44072
rect 2010 -45576 2074 -45570
rect 2010 -45579 2016 -45576
rect 2005 -45625 2016 -45579
rect 2010 -45628 2016 -45625
rect 2068 -45579 2074 -45576
rect 2068 -45625 2079 -45579
rect 2068 -45628 2074 -45625
rect 2010 -45634 2074 -45628
rect 2304 -47584 2368 -47578
rect 2304 -47636 2310 -47584
rect 2362 -47636 2368 -47584
rect 2304 -47642 2368 -47636
rect 2010 -49140 2074 -49134
rect 2010 -49143 2016 -49140
rect 2005 -49189 2016 -49143
rect 2010 -49192 2016 -49189
rect 2068 -49143 2074 -49140
rect 2068 -49189 2079 -49143
rect 2068 -49192 2074 -49189
rect 2010 -49198 2074 -49192
rect 2304 -51148 2368 -51142
rect 2304 -51200 2310 -51148
rect 2362 -51200 2368 -51148
rect 2304 -51206 2368 -51200
rect 2010 -52704 2074 -52698
rect 2010 -52707 2016 -52704
rect 2005 -52753 2016 -52707
rect 2010 -52756 2016 -52753
rect 2068 -52707 2074 -52704
rect 2068 -52753 2079 -52707
rect 2068 -52756 2074 -52753
rect 2010 -52762 2074 -52756
rect 2304 -54712 2368 -54706
rect 2304 -54764 2310 -54712
rect 2362 -54764 2368 -54712
rect 2304 -54770 2368 -54764
rect 2010 -56268 2074 -56262
rect 2010 -56271 2016 -56268
rect 2005 -56317 2016 -56271
rect 2010 -56320 2016 -56317
rect 2068 -56271 2074 -56268
rect 2068 -56317 2079 -56271
rect 2068 -56320 2074 -56317
rect 2010 -56326 2074 -56320
rect 2304 -58276 2368 -58270
rect 2304 -58328 2310 -58276
rect 2362 -58328 2368 -58276
rect 2304 -58334 2368 -58328
rect 2010 -59832 2074 -59826
rect 2010 -59835 2016 -59832
rect 2005 -59881 2016 -59835
rect 2010 -59884 2016 -59881
rect 2068 -59835 2074 -59832
rect 2068 -59881 2079 -59835
rect 2068 -59884 2074 -59881
rect 2010 -59890 2074 -59884
rect 2304 -61840 2368 -61834
rect 2304 -61892 2310 -61840
rect 2362 -61892 2368 -61840
rect 2304 -61898 2368 -61892
rect 2010 -63396 2074 -63390
rect 2010 -63399 2016 -63396
rect 2005 -63445 2016 -63399
rect 2010 -63448 2016 -63445
rect 2068 -63399 2074 -63396
rect 2068 -63445 2079 -63399
rect 2068 -63448 2074 -63445
rect 2010 -63454 2074 -63448
rect 2304 -65404 2368 -65398
rect 2304 -65456 2310 -65404
rect 2362 -65456 2368 -65404
rect 2304 -65462 2368 -65456
rect 2010 -66960 2074 -66954
rect 2010 -67012 2016 -66960
rect 2068 -67012 2074 -66960
rect 2010 -67018 2074 -67012
<< via1 >>
rect 1867 -9988 1919 -9936
rect 2310 -11996 2362 -11944
rect 2016 -13552 2068 -13500
rect 2310 -15560 2362 -15508
rect 2016 -17116 2068 -17064
rect 2310 -19124 2362 -19072
rect 2016 -20680 2068 -20628
rect 2310 -22688 2362 -22636
rect 2016 -24244 2068 -24192
rect 2310 -26252 2362 -26200
rect 2016 -27808 2068 -27756
rect 2310 -29816 2362 -29764
rect 2016 -31372 2068 -31320
rect 2310 -33380 2362 -33328
rect 2016 -34936 2068 -34884
rect 2310 -36944 2362 -36892
rect 2016 -38500 2068 -38448
rect 2310 -40508 2362 -40456
rect 2016 -42064 2068 -42012
rect 2310 -44072 2362 -44020
rect 2016 -45628 2068 -45576
rect 2310 -47636 2362 -47584
rect 2016 -49192 2068 -49140
rect 2310 -51200 2362 -51148
rect 2016 -52756 2068 -52704
rect 2310 -54764 2362 -54712
rect 2016 -56320 2068 -56268
rect 2310 -58328 2362 -58276
rect 2016 -59884 2068 -59832
rect 2310 -61892 2362 -61840
rect 2016 -63448 2068 -63396
rect 2310 -65456 2362 -65404
rect 2016 -67012 2068 -66960
<< metal2 >>
rect 2299 -9004 2373 -8995
rect 2299 -9060 2308 -9004
rect 2364 -9060 2373 -9004
rect 2299 -9069 2373 -9060
rect 1856 -9934 1930 -9925
rect 1856 -9990 1865 -9934
rect 1921 -9990 1930 -9934
rect 1856 -9999 1930 -9990
rect 1721 -10190 1795 -10181
rect 1721 -10246 1730 -10190
rect 1786 -10246 1795 -10190
rect 1721 -10255 1795 -10246
rect 2304 -11944 2368 -11938
rect 2304 -11996 2310 -11944
rect 2362 -11947 2368 -11944
rect 9060 -11942 9134 -11933
rect 9060 -11947 9069 -11942
rect 2362 -11993 9069 -11947
rect 2362 -11996 2368 -11993
rect 2304 -12002 2368 -11996
rect 9060 -11998 9069 -11993
rect 9125 -11998 9134 -11942
rect 9060 -12007 9134 -11998
rect 2005 -12688 2079 -12679
rect 2005 -12744 2014 -12688
rect 2070 -12744 2079 -12688
rect 2005 -12753 2079 -12744
rect 1721 -13242 1795 -13233
rect 1721 -13298 1730 -13242
rect 1786 -13298 1795 -13242
rect 1721 -13307 1795 -13298
rect 2005 -13498 2079 -13489
rect 2005 -13554 2014 -13498
rect 2070 -13554 2079 -13498
rect 2005 -13563 2079 -13554
rect 2304 -15508 2368 -15502
rect 2304 -15560 2310 -15508
rect 2362 -15511 2368 -15508
rect 9060 -15506 9134 -15497
rect 9060 -15511 9069 -15506
rect 2362 -15557 9069 -15511
rect 2362 -15560 2368 -15557
rect 2304 -15566 2368 -15560
rect 9060 -15562 9069 -15557
rect 9125 -15562 9134 -15506
rect 9060 -15571 9134 -15562
rect 2005 -17062 2079 -17053
rect 2005 -17118 2014 -17062
rect 2070 -17118 2079 -17062
rect 2005 -17127 2079 -17118
rect 2304 -19072 2368 -19066
rect 2304 -19124 2310 -19072
rect 2362 -19075 2368 -19072
rect 9060 -19070 9134 -19061
rect 9060 -19075 9069 -19070
rect 2362 -19121 9069 -19075
rect 2362 -19124 2368 -19121
rect 2304 -19130 2368 -19124
rect 9060 -19126 9069 -19121
rect 9125 -19126 9134 -19070
rect 9060 -19135 9134 -19126
rect 2005 -20626 2079 -20617
rect 2005 -20682 2014 -20626
rect 2070 -20682 2079 -20626
rect 2005 -20691 2079 -20682
rect 2304 -22636 2368 -22630
rect 2304 -22688 2310 -22636
rect 2362 -22639 2368 -22636
rect 9060 -22634 9134 -22625
rect 9060 -22639 9069 -22634
rect 2362 -22685 9069 -22639
rect 2362 -22688 2368 -22685
rect 2304 -22694 2368 -22688
rect 9060 -22690 9069 -22685
rect 9125 -22690 9134 -22634
rect 9060 -22699 9134 -22690
rect 2005 -24190 2079 -24181
rect 2005 -24246 2014 -24190
rect 2070 -24246 2079 -24190
rect 2005 -24255 2079 -24246
rect 2304 -26200 2368 -26194
rect 2304 -26252 2310 -26200
rect 2362 -26203 2368 -26200
rect 9060 -26198 9134 -26189
rect 9060 -26203 9069 -26198
rect 2362 -26249 9069 -26203
rect 2362 -26252 2368 -26249
rect 2304 -26258 2368 -26252
rect 9060 -26254 9069 -26249
rect 9125 -26254 9134 -26198
rect 9060 -26263 9134 -26254
rect 2005 -27754 2079 -27745
rect 2005 -27810 2014 -27754
rect 2070 -27810 2079 -27754
rect 2005 -27819 2079 -27810
rect 2304 -29764 2368 -29758
rect 2304 -29816 2310 -29764
rect 2362 -29767 2368 -29764
rect 9060 -29762 9134 -29753
rect 9060 -29767 9069 -29762
rect 2362 -29813 9069 -29767
rect 2362 -29816 2368 -29813
rect 2304 -29822 2368 -29816
rect 9060 -29818 9069 -29813
rect 9125 -29818 9134 -29762
rect 9060 -29827 9134 -29818
rect 2005 -31318 2079 -31309
rect 2005 -31374 2014 -31318
rect 2070 -31374 2079 -31318
rect 2005 -31383 2079 -31374
rect 2304 -33328 2368 -33322
rect 2304 -33380 2310 -33328
rect 2362 -33331 2368 -33328
rect 9060 -33326 9134 -33317
rect 9060 -33331 9069 -33326
rect 2362 -33377 9069 -33331
rect 2362 -33380 2368 -33377
rect 2304 -33386 2368 -33380
rect 9060 -33382 9069 -33377
rect 9125 -33382 9134 -33326
rect 9060 -33391 9134 -33382
rect 2005 -34882 2079 -34873
rect 2005 -34938 2014 -34882
rect 2070 -34938 2079 -34882
rect 2005 -34947 2079 -34938
rect 2304 -36892 2368 -36886
rect 2304 -36944 2310 -36892
rect 2362 -36895 2368 -36892
rect 9060 -36890 9134 -36881
rect 9060 -36895 9069 -36890
rect 2362 -36941 9069 -36895
rect 2362 -36944 2368 -36941
rect 2304 -36950 2368 -36944
rect 9060 -36946 9069 -36941
rect 9125 -36946 9134 -36890
rect 9060 -36955 9134 -36946
rect 2005 -38446 2079 -38437
rect 2005 -38502 2014 -38446
rect 2070 -38502 2079 -38446
rect 2005 -38511 2079 -38502
rect 2304 -40456 2368 -40450
rect 2304 -40508 2310 -40456
rect 2362 -40459 2368 -40456
rect 9060 -40454 9134 -40445
rect 9060 -40459 9069 -40454
rect 2362 -40505 9069 -40459
rect 2362 -40508 2368 -40505
rect 2304 -40514 2368 -40508
rect 9060 -40510 9069 -40505
rect 9125 -40510 9134 -40454
rect 9060 -40519 9134 -40510
rect 2005 -42010 2079 -42001
rect 2005 -42066 2014 -42010
rect 2070 -42066 2079 -42010
rect 2005 -42075 2079 -42066
rect 2304 -44020 2368 -44014
rect 2304 -44072 2310 -44020
rect 2362 -44023 2368 -44020
rect 9060 -44018 9134 -44009
rect 9060 -44023 9069 -44018
rect 2362 -44069 9069 -44023
rect 2362 -44072 2368 -44069
rect 2304 -44078 2368 -44072
rect 9060 -44074 9069 -44069
rect 9125 -44074 9134 -44018
rect 9060 -44083 9134 -44074
rect 2005 -45574 2079 -45565
rect 2005 -45630 2014 -45574
rect 2070 -45630 2079 -45574
rect 2005 -45639 2079 -45630
rect 2304 -47584 2368 -47578
rect 2304 -47636 2310 -47584
rect 2362 -47587 2368 -47584
rect 9060 -47582 9134 -47573
rect 9060 -47587 9069 -47582
rect 2362 -47633 9069 -47587
rect 2362 -47636 2368 -47633
rect 2304 -47642 2368 -47636
rect 9060 -47638 9069 -47633
rect 9125 -47638 9134 -47582
rect 9060 -47647 9134 -47638
rect 2005 -49138 2079 -49129
rect 2005 -49194 2014 -49138
rect 2070 -49194 2079 -49138
rect 2005 -49203 2079 -49194
rect 2304 -51148 2368 -51142
rect 2304 -51200 2310 -51148
rect 2362 -51151 2368 -51148
rect 9060 -51146 9134 -51137
rect 9060 -51151 9069 -51146
rect 2362 -51197 9069 -51151
rect 2362 -51200 2368 -51197
rect 2304 -51206 2368 -51200
rect 9060 -51202 9069 -51197
rect 9125 -51202 9134 -51146
rect 9060 -51211 9134 -51202
rect 2005 -52702 2079 -52693
rect 2005 -52758 2014 -52702
rect 2070 -52758 2079 -52702
rect 2005 -52767 2079 -52758
rect 2304 -54712 2368 -54706
rect 2304 -54764 2310 -54712
rect 2362 -54715 2368 -54712
rect 9060 -54710 9134 -54701
rect 9060 -54715 9069 -54710
rect 2362 -54761 9069 -54715
rect 2362 -54764 2368 -54761
rect 2304 -54770 2368 -54764
rect 9060 -54766 9069 -54761
rect 9125 -54766 9134 -54710
rect 9060 -54775 9134 -54766
rect 2005 -56266 2079 -56257
rect 2005 -56322 2014 -56266
rect 2070 -56322 2079 -56266
rect 2005 -56331 2079 -56322
rect 2304 -58276 2368 -58270
rect 2304 -58328 2310 -58276
rect 2362 -58279 2368 -58276
rect 9060 -58274 9134 -58265
rect 9060 -58279 9069 -58274
rect 2362 -58325 9069 -58279
rect 2362 -58328 2368 -58325
rect 2304 -58334 2368 -58328
rect 9060 -58330 9069 -58325
rect 9125 -58330 9134 -58274
rect 9060 -58339 9134 -58330
rect 2005 -59830 2079 -59821
rect 2005 -59886 2014 -59830
rect 2070 -59886 2079 -59830
rect 2005 -59895 2079 -59886
rect 2304 -61840 2368 -61834
rect 2304 -61892 2310 -61840
rect 2362 -61843 2368 -61840
rect 9060 -61838 9134 -61829
rect 9060 -61843 9069 -61838
rect 2362 -61889 9069 -61843
rect 2362 -61892 2368 -61889
rect 2304 -61898 2368 -61892
rect 9060 -61894 9069 -61889
rect 9125 -61894 9134 -61838
rect 9060 -61903 9134 -61894
rect 2005 -63394 2079 -63385
rect 2005 -63450 2014 -63394
rect 2070 -63450 2079 -63394
rect 2005 -63459 2079 -63450
rect 2304 -65404 2368 -65398
rect 2304 -65456 2310 -65404
rect 2362 -65407 2368 -65404
rect 9060 -65402 9134 -65393
rect 9060 -65407 9069 -65402
rect 2362 -65453 9069 -65407
rect 2362 -65456 2368 -65453
rect 2304 -65462 2368 -65456
rect 9060 -65458 9069 -65453
rect 9125 -65458 9134 -65402
rect 9060 -65467 9134 -65458
rect 2005 -66958 2079 -66949
rect 2005 -67014 2014 -66958
rect 2070 -67014 2079 -66958
rect 2005 -67023 2079 -67014
rect 2299 -66958 2373 -66949
rect 2299 -67014 2308 -66958
rect 2364 -66963 2373 -66958
rect 9060 -66958 9134 -66949
rect 9060 -66963 9069 -66958
rect 2364 -67009 9069 -66963
rect 2364 -67014 2373 -67009
rect 2299 -67023 2373 -67014
rect 9060 -67014 9069 -67009
rect 9125 -67014 9134 -66958
rect 9060 -67023 9134 -67014
<< via2 >>
rect 2308 -9060 2364 -9004
rect 1865 -9936 1921 -9934
rect 1865 -9988 1867 -9936
rect 1867 -9988 1919 -9936
rect 1919 -9988 1921 -9936
rect 1865 -9990 1921 -9988
rect 1730 -10246 1786 -10190
rect 9069 -11998 9125 -11942
rect 2014 -12744 2070 -12688
rect 1730 -13298 1786 -13242
rect 2014 -13500 2070 -13498
rect 2014 -13552 2016 -13500
rect 2016 -13552 2068 -13500
rect 2068 -13552 2070 -13500
rect 2014 -13554 2070 -13552
rect 9069 -15562 9125 -15506
rect 2014 -17064 2070 -17062
rect 2014 -17116 2016 -17064
rect 2016 -17116 2068 -17064
rect 2068 -17116 2070 -17064
rect 2014 -17118 2070 -17116
rect 9069 -19126 9125 -19070
rect 2014 -20628 2070 -20626
rect 2014 -20680 2016 -20628
rect 2016 -20680 2068 -20628
rect 2068 -20680 2070 -20628
rect 2014 -20682 2070 -20680
rect 9069 -22690 9125 -22634
rect 2014 -24192 2070 -24190
rect 2014 -24244 2016 -24192
rect 2016 -24244 2068 -24192
rect 2068 -24244 2070 -24192
rect 2014 -24246 2070 -24244
rect 9069 -26254 9125 -26198
rect 2014 -27756 2070 -27754
rect 2014 -27808 2016 -27756
rect 2016 -27808 2068 -27756
rect 2068 -27808 2070 -27756
rect 2014 -27810 2070 -27808
rect 9069 -29818 9125 -29762
rect 2014 -31320 2070 -31318
rect 2014 -31372 2016 -31320
rect 2016 -31372 2068 -31320
rect 2068 -31372 2070 -31320
rect 2014 -31374 2070 -31372
rect 9069 -33382 9125 -33326
rect 2014 -34884 2070 -34882
rect 2014 -34936 2016 -34884
rect 2016 -34936 2068 -34884
rect 2068 -34936 2070 -34884
rect 2014 -34938 2070 -34936
rect 9069 -36946 9125 -36890
rect 2014 -38448 2070 -38446
rect 2014 -38500 2016 -38448
rect 2016 -38500 2068 -38448
rect 2068 -38500 2070 -38448
rect 2014 -38502 2070 -38500
rect 9069 -40510 9125 -40454
rect 2014 -42012 2070 -42010
rect 2014 -42064 2016 -42012
rect 2016 -42064 2068 -42012
rect 2068 -42064 2070 -42012
rect 2014 -42066 2070 -42064
rect 9069 -44074 9125 -44018
rect 2014 -45576 2070 -45574
rect 2014 -45628 2016 -45576
rect 2016 -45628 2068 -45576
rect 2068 -45628 2070 -45576
rect 2014 -45630 2070 -45628
rect 9069 -47638 9125 -47582
rect 2014 -49140 2070 -49138
rect 2014 -49192 2016 -49140
rect 2016 -49192 2068 -49140
rect 2068 -49192 2070 -49140
rect 2014 -49194 2070 -49192
rect 9069 -51202 9125 -51146
rect 2014 -52704 2070 -52702
rect 2014 -52756 2016 -52704
rect 2016 -52756 2068 -52704
rect 2068 -52756 2070 -52704
rect 2014 -52758 2070 -52756
rect 9069 -54766 9125 -54710
rect 2014 -56268 2070 -56266
rect 2014 -56320 2016 -56268
rect 2016 -56320 2068 -56268
rect 2068 -56320 2070 -56268
rect 2014 -56322 2070 -56320
rect 9069 -58330 9125 -58274
rect 2014 -59832 2070 -59830
rect 2014 -59884 2016 -59832
rect 2016 -59884 2068 -59832
rect 2068 -59884 2070 -59832
rect 2014 -59886 2070 -59884
rect 9069 -61894 9125 -61838
rect 2014 -63396 2070 -63394
rect 2014 -63448 2016 -63396
rect 2016 -63448 2068 -63396
rect 2068 -63448 2070 -63396
rect 2014 -63450 2070 -63448
rect 9069 -65458 9125 -65402
rect 2014 -66960 2070 -66958
rect 2014 -67012 2016 -66960
rect 2016 -67012 2068 -66960
rect 2068 -67012 2070 -66960
rect 2014 -67014 2070 -67012
rect 2308 -67014 2364 -66958
rect 9069 -67014 9125 -66958
<< metal3 >>
rect 635 -68740 695 -8212
rect 2303 -9004 2369 -8999
rect 2303 -9060 2308 -9004
rect 2364 -9060 2369 -9004
rect 2303 -9065 2369 -9060
rect 1860 -9934 1926 -9929
rect 1860 -9990 1865 -9934
rect 1921 -9990 1926 -9934
rect 1860 -9995 1926 -9990
rect 1725 -10190 1791 -10185
rect 1725 -10246 1730 -10190
rect 1786 -10246 1791 -10190
rect 1725 -10251 1791 -10246
rect 1728 -13237 1788 -10251
rect 2012 -12683 2072 -10742
rect 1725 -13242 1791 -13237
rect 1725 -13298 1730 -13242
rect 1786 -13298 1791 -13242
rect 1725 -13303 1791 -13298
rect 1863 -67272 1923 -12686
rect 2009 -12688 2075 -12683
rect 2009 -12744 2014 -12688
rect 2070 -12744 2075 -12688
rect 2009 -12749 2075 -12744
rect 2012 -13493 2072 -13340
rect 2009 -13498 2075 -13493
rect 2009 -13554 2014 -13498
rect 2070 -13554 2075 -13498
rect 2009 -13559 2075 -13554
rect 2012 -17057 2072 -13559
rect 2009 -17062 2075 -17057
rect 2009 -17118 2014 -17062
rect 2070 -17118 2075 -17062
rect 2009 -17123 2075 -17118
rect 2012 -20621 2072 -17123
rect 2009 -20626 2075 -20621
rect 2009 -20682 2014 -20626
rect 2070 -20682 2075 -20626
rect 2009 -20687 2075 -20682
rect 2012 -24185 2072 -20687
rect 2009 -24190 2075 -24185
rect 2009 -24246 2014 -24190
rect 2070 -24246 2075 -24190
rect 2009 -24251 2075 -24246
rect 2012 -27749 2072 -24251
rect 2009 -27754 2075 -27749
rect 2009 -27810 2014 -27754
rect 2070 -27810 2075 -27754
rect 2009 -27815 2075 -27810
rect 2012 -31313 2072 -27815
rect 2009 -31318 2075 -31313
rect 2009 -31374 2014 -31318
rect 2070 -31374 2075 -31318
rect 2009 -31379 2075 -31374
rect 2012 -34877 2072 -31379
rect 2009 -34882 2075 -34877
rect 2009 -34938 2014 -34882
rect 2070 -34938 2075 -34882
rect 2009 -34943 2075 -34938
rect 2012 -38441 2072 -34943
rect 2009 -38446 2075 -38441
rect 2009 -38502 2014 -38446
rect 2070 -38502 2075 -38446
rect 2009 -38507 2075 -38502
rect 2012 -42005 2072 -38507
rect 2009 -42010 2075 -42005
rect 2009 -42066 2014 -42010
rect 2070 -42066 2075 -42010
rect 2009 -42071 2075 -42066
rect 2012 -45569 2072 -42071
rect 2009 -45574 2075 -45569
rect 2009 -45630 2014 -45574
rect 2070 -45630 2075 -45574
rect 2009 -45635 2075 -45630
rect 2012 -49133 2072 -45635
rect 2009 -49138 2075 -49133
rect 2009 -49194 2014 -49138
rect 2070 -49194 2075 -49138
rect 2009 -49199 2075 -49194
rect 2012 -52697 2072 -49199
rect 2009 -52702 2075 -52697
rect 2009 -52758 2014 -52702
rect 2070 -52758 2075 -52702
rect 2009 -52763 2075 -52758
rect 2012 -56261 2072 -52763
rect 2009 -56266 2075 -56261
rect 2009 -56322 2014 -56266
rect 2070 -56322 2075 -56266
rect 2009 -56327 2075 -56322
rect 2012 -59825 2072 -56327
rect 2009 -59830 2075 -59825
rect 2009 -59886 2014 -59830
rect 2070 -59886 2075 -59830
rect 2009 -59891 2075 -59886
rect 2012 -63389 2072 -59891
rect 2009 -63394 2075 -63389
rect 2009 -63450 2014 -63394
rect 2070 -63450 2075 -63394
rect 2009 -63455 2075 -63450
rect 2012 -66953 2072 -63455
rect 2306 -66953 2366 -9065
rect 2009 -66958 2075 -66953
rect 2009 -67014 2014 -66958
rect 2070 -67014 2075 -66958
rect 2009 -67019 2075 -67014
rect 2303 -66958 2369 -66953
rect 2303 -67014 2308 -66958
rect 2364 -67014 2369 -66958
rect 2303 -67019 2369 -67014
rect 2012 -67826 2072 -67019
rect 2920 -67272 2980 -9676
rect 9067 -11937 9127 -9580
rect 9064 -11942 9130 -11937
rect 9064 -11998 9069 -11942
rect 9125 -11998 9130 -11942
rect 9064 -12003 9130 -11998
rect 9067 -15501 9127 -13144
rect 9064 -15506 9130 -15501
rect 9064 -15562 9069 -15506
rect 9125 -15562 9130 -15506
rect 9064 -15567 9130 -15562
rect 9067 -19065 9127 -16708
rect 9064 -19070 9130 -19065
rect 9064 -19126 9069 -19070
rect 9125 -19126 9130 -19070
rect 9064 -19131 9130 -19126
rect 9067 -22629 9127 -20272
rect 9064 -22634 9130 -22629
rect 9064 -22690 9069 -22634
rect 9125 -22690 9130 -22634
rect 9064 -22695 9130 -22690
rect 9067 -26193 9127 -23836
rect 9064 -26198 9130 -26193
rect 9064 -26254 9069 -26198
rect 9125 -26254 9130 -26198
rect 9064 -26259 9130 -26254
rect 9067 -29757 9127 -27400
rect 9064 -29762 9130 -29757
rect 9064 -29818 9069 -29762
rect 9125 -29818 9130 -29762
rect 9064 -29823 9130 -29818
rect 9067 -33321 9127 -30964
rect 9064 -33326 9130 -33321
rect 9064 -33382 9069 -33326
rect 9125 -33382 9130 -33326
rect 9064 -33387 9130 -33382
rect 9067 -36885 9127 -34528
rect 9064 -36890 9130 -36885
rect 9064 -36946 9069 -36890
rect 9125 -36946 9130 -36890
rect 9064 -36951 9130 -36946
rect 9067 -40449 9127 -38092
rect 9064 -40454 9130 -40449
rect 9064 -40510 9069 -40454
rect 9125 -40510 9130 -40454
rect 9064 -40515 9130 -40510
rect 9067 -44013 9127 -41656
rect 9064 -44018 9130 -44013
rect 9064 -44074 9069 -44018
rect 9125 -44074 9130 -44018
rect 9064 -44079 9130 -44074
rect 9067 -47577 9127 -45220
rect 9064 -47582 9130 -47577
rect 9064 -47638 9069 -47582
rect 9125 -47638 9130 -47582
rect 9064 -47643 9130 -47638
rect 9067 -51141 9127 -48784
rect 9064 -51146 9130 -51141
rect 9064 -51202 9069 -51146
rect 9125 -51202 9130 -51146
rect 9064 -51207 9130 -51202
rect 9067 -54705 9127 -52348
rect 9064 -54710 9130 -54705
rect 9064 -54766 9069 -54710
rect 9125 -54766 9130 -54710
rect 9064 -54771 9130 -54766
rect 9067 -58269 9127 -55912
rect 9064 -58274 9130 -58269
rect 9064 -58330 9069 -58274
rect 9125 -58330 9130 -58274
rect 9064 -58335 9130 -58330
rect 9067 -61833 9127 -59476
rect 9064 -61838 9130 -61833
rect 9064 -61894 9069 -61838
rect 9125 -61894 9130 -61838
rect 9064 -61899 9130 -61894
rect 9067 -65397 9127 -63040
rect 9064 -65402 9130 -65397
rect 9064 -65458 9069 -65402
rect 9125 -65458 9130 -65402
rect 9064 -65463 9130 -65458
rect 9064 -66958 9130 -66953
rect 9064 -67014 9069 -66958
rect 9125 -67014 9130 -66958
rect 9064 -67019 9130 -67014
use D_FlipFlop  D_FlipFlop_0
timestamp 1757226713
transform 1 0 606 0 1 -9985
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_1
timestamp 1757226713
transform 1 0 606 0 1 -13549
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1757226713
transform 1 0 606 0 1 -17113
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1757226713
transform 1 0 606 0 1 -20677
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1757226713
transform 1 0 606 0 1 -24241
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1757226713
transform 1 0 606 0 1 -27805
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1757226713
transform 1 0 606 0 1 -31369
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1757226713
transform 1 0 606 0 1 -34933
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_8
timestamp 1757226713
transform 1 0 606 0 1 -38497
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_9
timestamp 1757226713
transform 1 0 606 0 1 -42061
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_10
timestamp 1757226713
transform 1 0 606 0 1 -45625
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_11
timestamp 1757226713
transform 1 0 606 0 1 -49189
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_12
timestamp 1757226713
transform 1 0 606 0 1 -52753
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_13
timestamp 1757226713
transform 1 0 606 0 1 -56317
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_14
timestamp 1757226713
transform 1 0 606 0 1 -59881
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_15
timestamp 1757226713
transform 1 0 606 0 1 -63445
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_16
timestamp 1757226713
transform 1 0 606 0 1 -67009
box 0 -1796 8762 1842
<< labels >>
flabel metal3 2920 -67272 2980 -9676 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 1863 -67272 1923 -12686 0 FreeSans 160 90 0 0 EN
port 1 nsew
flabel metal3 9067 -11942 9127 -9580 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal3 9067 -15506 9127 -13144 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal3 9067 -19070 9127 -16708 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal3 9067 -22634 9127 -20272 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal3 9067 -26198 9127 -23836 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal3 9067 -29762 9127 -27400 0 FreeSans 160 0 0 0 Q5
port 8 nsew
flabel metal3 9067 -33326 9127 -30964 0 FreeSans 160 0 0 0 Q6
port 9 nsew
flabel metal3 9067 -36890 9127 -34528 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal3 9067 -40454 9127 -38092 0 FreeSans 160 0 0 0 Q8
port 11 nsew
flabel metal3 9067 -44018 9127 -41656 0 FreeSans 160 0 0 0 Q9
port 12 nsew
flabel metal3 9067 -47582 9127 -45220 0 FreeSans 160 0 0 0 Q10
port 13 nsew
flabel metal3 9067 -51146 9127 -48784 0 FreeSans 160 0 0 0 Q11
port 14 nsew
flabel metal3 9067 -54710 9127 -52348 0 FreeSans 160 0 0 0 Q12
port 15 nsew
flabel metal3 9067 -58274 9127 -55912 0 FreeSans 160 0 0 0 Q13
port 16 nsew
flabel metal3 9067 -61838 9127 -59476 0 FreeSans 160 0 0 0 Q14
port 17 nsew
flabel metal3 9067 -65402 9127 -63040 0 FreeSans 160 0 0 0 Q15
port 18 nsew
flabel metal3 2012 -67826 2014 -13340 0 FreeSans 160 90 0 0 VDD
port 19 nsew
flabel metal3 635 -68740 695 -8212 0 FreeSans 160 90 0 0 GND
port 20 nsew
<< end >>
