** sch_path: /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-05_18-41-24/parameters/INL/run_2/sar_output.sch
**.subckt sar_output
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND DC 0.158810118
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
**** begin user architecture code

* CACE gensim simulation file sar_output_2
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/samantha/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
tran 0.5u 8.5u uic
set wr_singlescale
wrdata /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-05_18-41-24/parameters/INL/run_2/sar_output_2.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)
quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
