magic
tech sky130A
magscale 1 2
timestamp 1761392116
<< metal1 >>
rect -1558 1555 544 1635
rect -1209 414 -1163 946
rect -595 414 -549 946
rect -338 625 132 705
rect 406 302 486 1067
rect -1558 -227 544 -147
use Inverter  Inverter_0
timestamp 1761294637
transform 1 0 -1566 0 1 676
box 1366 -903 2110 959
use Nand_Gate  Nand_Gate_0
timestamp 1761392116
transform 1 0 -3464 0 1 320
box 1906 -547 3264 1315
<< labels >>
flabel metal1 -1558 1572 544 1618 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 -1209 414 -1163 946 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 -595 414 -549 946 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal1 406 302 486 1067 0 FreeSans 160 0 0 0 Vout
port 5 nsew
flabel metal1 -1558 -210 544 -164 0 FreeSans 160 0 0 0 GND
port 0 nsew
<< end >>
