magic
tech sky130A
timestamp 1756538730
<< pwell >>
rect -164 -879 164 879
<< mvnmos >>
rect -50 -750 50 750
<< mvndiff >>
rect -79 744 -50 750
rect -79 -744 -73 744
rect -56 -744 -50 744
rect -79 -750 -50 -744
rect 50 744 79 750
rect 50 -744 56 744
rect 73 -744 79 744
rect 50 -750 79 -744
<< mvndiffc >>
rect -73 -744 -56 744
rect 56 -744 73 744
<< mvpsubdiff >>
rect -146 855 146 861
rect -146 838 -92 855
rect 92 838 146 855
rect -146 832 146 838
rect -146 807 -117 832
rect -146 -807 -140 807
rect -123 -807 -117 807
rect 117 807 146 832
rect -146 -832 -117 -807
rect 117 -807 123 807
rect 140 -807 146 807
rect 117 -832 146 -807
rect -146 -838 146 -832
rect -146 -855 -92 -838
rect 92 -855 146 -838
rect -146 -861 146 -855
<< mvpsubdiffcont >>
rect -92 838 92 855
rect -140 -807 -123 807
rect 123 -807 140 807
rect -92 -855 92 -838
<< poly >>
rect -50 786 50 794
rect -50 769 -42 786
rect 42 769 50 786
rect -50 750 50 769
rect -50 -769 50 -750
rect -50 -786 -42 -769
rect 42 -786 50 -769
rect -50 -794 50 -786
<< polycont >>
rect -42 769 42 786
rect -42 -786 42 -769
<< locali >>
rect -140 838 -92 855
rect 92 838 140 855
rect -140 807 -123 838
rect 123 807 140 838
rect -50 769 -42 786
rect 42 769 50 786
rect -73 744 -56 752
rect -73 -752 -56 -744
rect 56 744 73 752
rect 56 -752 73 -744
rect -50 -786 -42 -769
rect 42 -786 50 -769
rect -140 -838 -123 -807
rect 123 -838 140 -807
rect -140 -855 -92 -838
rect 92 -855 140 -838
<< viali >>
rect -42 769 42 786
rect -73 -744 -56 744
rect 56 -744 73 744
rect -42 -786 42 -769
<< metal1 >>
rect -48 786 48 789
rect -48 769 -42 786
rect 42 769 48 786
rect -48 766 48 769
rect -76 744 -53 750
rect -76 -744 -73 744
rect -56 -744 -53 744
rect -76 -750 -53 -744
rect 53 744 76 750
rect 53 -744 56 744
rect 73 -744 76 744
rect 53 -750 76 -744
rect -48 -769 48 -766
rect -48 -786 -42 -769
rect 42 -786 48 -769
rect -48 -789 48 -786
<< properties >>
string FIXED_BBOX -131 -846 131 846
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 15 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string sky130_fd_pr__nfet_g5v0d10v5_94KJBV parameters
<< end >>
