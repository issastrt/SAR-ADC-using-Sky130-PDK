** sch_path: /home/audrey/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-08-29_17-48-37/parameters/Power/run_06/power_consumption.sch
**.subckt power_consumption
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.8
VCLK CLK GND PULSE(1.8 0 0 500p 500p 1u 2u)
VEN EN net1 PULSE(1.8 0 0 500ps 500ps 1u 0)
VVin Vin GND DC 0.6
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
R1 net1 GND 0.01 m=1
**** begin user architecture code

.control
tran 0.5u 34u uic
set wr_singlescale
wrdata /home/audrey/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-08-29_17-48-37/parameters/Power/run_06/power_consumption_6.data -I(VVDD)
quit
.endc



* CACE gensim simulation file power_consumption_6
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/audrey/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice sf

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
