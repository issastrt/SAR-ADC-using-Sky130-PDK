* NGSPICE file created from SAR-ADC-using-Sky130-PDK.ext - technology: sky130A

.subckt SAR-ADC-using-Sky130-PDK VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 GND
X0 a_49391_58825# Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t2 GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1 GND.t63 EN.t0 a_9337_55365# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X2 GND.t712 Q0.t4 CDAC_v3_0.switch_8.Z.t1 VDD.t776 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X3 a_n1355_54751# Ring_Counter_0.D_FlipFlop_15.Qbar.t4 Nand_Gate_1.A.t2 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X4 VDD.t214 VDD.t212 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X5 GND.t210 EN.t1 a_44977_59439# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X6 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t130 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X7 VDD.t1 D_FlipFlop_2.3-input-nand_2.Vout.t4 D_FlipFlop_2.Nand_Gate_0.Vout VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X8 GND.t199 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 a_48541_56723# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X9 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Inverter_1.Vout VDD.t444 VDD.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X10 a_2209_59439# Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout a_2209_58825# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X11 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t65 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X12 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t64 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X13 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.CLK.t2 VDD.t483 VDD.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X14 a_23593_60797# CLK.t0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X15 GND.t502 GND.t503 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X16 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B VDD.t897 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X17 VDD.t472 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t2 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X18 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_0.CLK.t2 VDD.t459 VDD.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X19 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B VDD.t272 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X20 GND.t94 CLK.t1 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t1 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X21 a_3059_61411# Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B a_3059_60797# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X22 a_49930_48405# FFCLR.t4 GND.t641 GND.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X23 a_6623_56723# Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X24 a_n4069_55365# Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 a_n4069_54751# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X25 GND.t518 VDD.t924 a_37849_61411# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X26 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t35 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X27 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t77 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X28 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.CLK.t2 a_33020_48405# GND.t578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X29 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t129 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X30 VDD.t211 VDD.t209 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X31 VDD.t399 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t3 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X32 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t128 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X33 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t34 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X34 a_51632_31172.t2 a_51632_31172.t1 VDD.t43 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X35 GND.t500 GND.t501 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X36 VDD.t73 Ring_Counter_0.D_FlipFlop_9.Qbar Nand_Gate_6.A.t0 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X37 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t127 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X38 VDD.t424 D_FlipFlop_2.3-input-nand_1.B D_FlipFlop_2.3-input-nand_1.Vout VDD.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X39 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t126 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X40 GND.t498 GND.t499 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X41 GND.t224 Nand_Gate_6.A.t4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X42 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.CLK.t2 VDD.t375 VDD.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X43 D_FlipFlop_3.3-input-nand_1.B D_FlipFlop_7.D.t3 VDD.t17 VDD.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X44 GND.t519 VDD.t925 a_31571_59439# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X45 GND.t520 VDD.t926 a_28007_59439# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X46 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t63 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X47 D_FlipFlop_7.Nand_Gate_1.Vout D_FlipFlop_7.Inverter_1.Vout VDD.t531 VDD.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X48 a_35135_56723# Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X49 VDD.t710 D_FlipFlop_3.nPRE.t4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X50 VDD.t208 VDD.t207 Ring_Counter_0.D_FlipFlop_2.Qbar VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X51 GND.t326 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 a_9337_56723# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X52 a_5773_58825# Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X53 GND.t212 EN.t2 a_10187_61411# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X54 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t62 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X55 D_FlipFlop_5.CLK.t1 And_Gate_3.Nand_Gate_0.Vout GND.t307 GND.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X56 VDD.t700 EN.t3 D_FlipFlop_2.nPRE.t3 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X57 GND.t496 GND.t497 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X58 a_15496_48405# D_FlipFlop_5.3-input-nand_1.B a_14882_48405# GND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X59 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t33 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X60 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t9 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X61 a_30721_56723# Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X62 VDD.t588 D_FlipFlop_4.nPRE.t4 Ring_Counter_0.D_FlipFlop_10.Qbar.t2 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X63 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t125 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X64 VDD.t251 CLK.t2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t1 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X65 VDD.t534 D_FlipFlop_2.3-input-nand_2.C.t4 D_FlipFlop_2.Nand_Gate_1.Vout VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X66 a_n11404_48405# D_FlipFlop_7.nPRE.t4 GND.t103 GND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X67 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_6.Inverter_1.Vout VDD.t443 VDD.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X68 VDD.t13 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X69 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t61 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X70 VDD.t206 VDD.t205 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X71 GND.t211 EN.t4 a_24443_61411# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X72 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.CLK.t3 VDD.t484 VDD.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X73 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout Nand_Gate_3.A.t4 VDD.t909 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X74 a_20879_61411# Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B a_20879_60797# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X75 a_41413_61411# D_FlipFlop_1.nPRE.t4 a_41413_60797# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X76 a_34285_58825# Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X77 VDD.t584 And_Gate_1.A And_Gate_1.Nand_Gate_0.Vout VDD.t583 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X78 VDD.t711 D_FlipFlop_3.nPRE.t5 Ring_Counter_0.D_FlipFlop_6.Qbar VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X79 VDD.t463 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t1 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X80 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.CLK.t2 GND.t244 GND.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X81 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 VDD.t378 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X82 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t124 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X83 VDD.t807 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X84 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t60 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X85 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 VDD.t374 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X86 VDD.t885 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_2.Vout.t3 VDD.t618 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X87 GND.t521 VDD.t927 a_13751_55365# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X88 a_43754_51119# D_FlipFlop_1.3-input-nand_0.Vout a_43140_51119# GND.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X89 a_n4919_60797# CLK.t3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X90 a_40815_52049# And_Gate_6.A GND.t218 GND.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X91 a_n7633_59439# Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 a_n7633_58825# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X92 Q6.t1 D_FlipFlop_1.Qbar a_47828_51119# GND.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X93 a_48541_58825# Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X94 Ring_Counter_0.D_FlipFlop_3.Qbar.t2 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 VDD.t52 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X95 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t59 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X96 And_Gate_1.Nand_Gate_0.Vout CLK.t4 VDD.t253 VDD.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X97 a_27157_60797# CLK.t5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X98 a_27542_45397# Q5.t4 GND.t183 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X99 CDAC_v3_0.switch_5.Z.t2 a_27542_45397# VDD.t631 VDD.t630 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X100 VDD.t593 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t1 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X101 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout FFCLR.t5 VDD.t387 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X102 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.CLK.t2 VDD.t900 VDD.t899 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X103 D_FlipFlop_0.3-input-nand_2.Vout.t2 FFCLR.t6 VDD.t389 VDD.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X104 GND.t522 VDD.t928 a_6623_59439# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X105 a_49391_60797# CLK.t6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X106 VDD.t417 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X107 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t123 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X108 VDD.t873 D_FlipFlop_0.Nand_Gate_0.Vout Q7.t3 VDD.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X109 VDD.t517 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X110 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t122 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X111 VDD.t89 D_FlipFlop_6.nPRE.t4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X112 GND.t494 GND.t495 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X113 a_41168_51119# FFCLR.t7 GND.t187 GND.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X114 a_25616_51119# D_FlipFlop_3.nPRE.t6 GND.t592 GND.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X115 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t121 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X116 D_FlipFlop_0.3-input-nand_2.Vout.t0 D_FlipFlop_0.3-input-nand_2.C.t4 VDD.t325 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X117 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t120 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X118 GND.t523 VDD.t929 a_44977_61411# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X119 a_49577_52049# And_Gate_7.A GND.t643 GND.t642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X120 a_2209_61411# Nand_Gate_0.A.t4 a_2209_60797# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X121 a_16465_54751# Ring_Counter_0.D_FlipFlop_10.Qbar.t4 D_FlipFlop_4.nPRE.t0 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X122 GND.t524 VDD.t930 a_38699_55365# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X123 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t58 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X124 a_8092_51119# D_FlipFlop_4.nPRE.t5 GND.t347 GND.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X125 VDD.t254 CLK.t7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X126 a_51773_21431.t0 Vin.t0 a_50502_29172.t0 Vbias.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X127 VDD.t533 Ring_Counter_0.D_FlipFlop_7.Qbar Nand_Gate_3.A.t1 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X128 a_20029_56723# Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X129 GND.t323 Nand_Gate_3.A.t5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X130 GND.t492 GND.t493 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X131 Q5.t0 D_FlipFlop_2.nPRE.t4 VDD.t739 VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X132 GND.t525 VDD.t931 a_35135_59439# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X133 Q7.t0 D_FlipFlop_0.Qbar VDD.t524 VDD.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X134 a_42263_56723# Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X135 VDD.t740 D_FlipFlop_2.nPRE.t5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X136 a_n56_51119# D_FlipFlop_6.3-input-nand_0.Vout a_n670_51119# GND.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X137 a_52105_59439# Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t4 a_52105_58825# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X138 VDD.t699 EN.t5 Ring_Counter_0.D_FlipFlop_0.Qbar VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X139 a_9337_58825# Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X140 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout D_FlipFlop_4.nPRE.t6 VDD.t589 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X141 VDD.t204 VDD.t203 Ring_Counter_0.D_FlipFlop_14.Qbar.t0 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X142 GND.t57 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t4 a_13751_56723# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X143 GND.t700 EN.t6 a_30721_59439# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X144 VDD.t255 CLK.t8 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t0 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X145 VDD.t619 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_0.3-input-nand_2.C.t0 VDD.t618 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X146 Ring_Counter_0.D_FlipFlop_16.Qbar Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 VDD.t846 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X147 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t119 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X148 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.CLK.t2 VDD.t837 VDD.t836 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X149 VDD.t787 D_FlipFlop_5.nPRE.t4 Ring_Counter_0.D_FlipFlop_8.Qbar.t1 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X150 VDD.t436 Nand_Gate_6.A.t5 Ring_Counter_0.D_FlipFlop_9.Qbar VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X151 VDD.t698 EN.t7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X152 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Inverter_1.Vout a_10808_51119# GND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X153 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t57 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X154 Q1.t2 D_FlipFlop_6.nPRE.t5 VDD.t91 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X155 a_45827_59439# Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 a_45827_58825# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X156 GND.t341 EN.t8 a_31571_61411# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X157 GND.t703 EN.t9 a_28007_61411# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X158 a_30304_48405# D_FlipFlop_3.Nand_Gate_1.Vout a_29690_48405# GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X159 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t118 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X160 Q1.t0 D_FlipFlop_6.Qbar VDD.t309 VDD.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X161 VDD.t256 CLK.t9 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t0 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X162 a_5773_60797# CLK.t10 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X163 a_n670_51119# D_FlipFlop_6.nPRE.t6 GND.t60 GND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X164 D_FlipFlop_4.3-input-nand_2.Vout.t0 D_FlipFlop_4.3-input-nand_2.C.t4 VDD.t826 VDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X165 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t32 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X166 D_FlipFlop_0.3-input-nand_2.C.t1 EN.t10 VDD.t697 VDD.t388 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X167 VDD.t372 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_0.Qbar VDD.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X168 a_19282_52049# D_FlipFlop_5.nPRE.t5 And_Gate_3.A GND.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X169 a_47214_48405# FFCLR.t8 GND.t189 GND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X170 D_FlipFlop_0.3-input-nand_2.C.t2 D_FlipFlop_0.3-input-nand_2.Vout.t4 VDD.t5 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X171 VDD.t19 D_FlipFlop_7.D.t4 D_FlipFlop_3.3-input-nand_0.Vout VDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X172 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t117 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X173 VDD.t239 CLK.t11 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X174 GND.t490 GND.t491 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X175 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 VDD.t414 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X176 D_FlipFlop_6.3-input-nand_1.B D_FlipFlop_7.D.t5 GND.t12 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X177 GND.t526 VDD.t932 a_17315_55365# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X178 GND.t327 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t4 a_38699_56723# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X179 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t116 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X180 GND.t488 GND.t489 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X181 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t115 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X182 a_3059_56723# Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X183 VDD.t502 D_FlipFlop_6.3-input-nand_2.Vout.t4 D_FlipFlop_6.Nand_Gate_0.Vout VDD.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X184 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t56 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X185 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_0.CLK.t3 a_50544_48405# GND.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X186 D_FlipFlop_2.3-input-nand_2.C.t3 D_FlipFlop_2.3-input-nand_2.Vout.t5 a_34992_48405# GND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X187 GND.t704 EN.t11 a_12901_55365# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X188 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t114 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X189 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t113 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X190 VDD.t555 Ring_Counter_0.D_FlipFlop_13.Qbar Nand_Gate_0.A.t0 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X191 a_34285_60797# CLK.t12 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X192 D_FlipFlop_2.Qbar FFCLR.t9 VDD.t391 VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X193 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD.t580 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X194 VDD.t696 EN.t12 D_FlipFlop_5.nPRE.t2 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X195 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t112 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X196 VDD.t602 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t3 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X197 D_FlipFlop_0.Qbar Q7.t4 VDD.t910 VDD.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X198 VDD.t695 EN.t13 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X199 VDD.t448 Q1.t4 CDAC_v3_0.switch_0.Z.t0 GND.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X200 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t55 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X201 VDD.t841 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X202 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t5 VDD.t851 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X203 CDAC_v3_0.OUT CDAC_v3_0.switch_2.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X204 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.CLK.t3 VDD.t901 VDD.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X205 VDD.t802 Nand_Gate_2.A.t4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X206 a_n7633_61411# Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B a_n7633_60797# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X207 D_FlipFlop_5.3-input-nand_1.B D_FlipFlop_7.D.t6 GND.t14 GND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X208 D_FlipFlop_7.Qbar Q0.t5 a_n4744_48405# GND.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X209 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t54 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X210 a_48541_60797# CLK.t13 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X211 a_n8818_48405# D_FlipFlop_7.3-input-nand_1.Vout a_n9432_48405# GND.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X212 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.CLK.t3 VDD.t838 VDD.t836 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X213 a_23593_54751# Ring_Counter_0.D_FlipFlop_8.Qbar.t4 D_FlipFlop_5.nPRE.t0 GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X214 a_33020_48405# D_FlipFlop_2.3-input-nand_1.B a_32406_48405# GND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X215 GND.t269 Nand_Gate_1.A.t4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X216 D_FlipFlop_6.Qbar FFCLR.t10 VDD.t392 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X217 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t53 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X218 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_2.Inverter_1.Vout a_37094_48405# GND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X219 D_FlipFlop_1.3-input-nand_1.B D_FlipFlop_7.D.t7 GND.t16 GND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X220 VDD.t835 Ring_Counter_0.D_FlipFlop_5.Qbar.t4 Nand_Gate_4.A.t1 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X221 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t5 VDD.t433 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X222 GND.t239 EN.t14 a_20029_59439# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X223 D_FlipFlop_6.Qbar Q1.t5 VDD.t449 VDD.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X224 Ring_Counter_0.D_FlipFlop_11.Qbar.t3 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 VDD.t519 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X225 GND.t593 D_FlipFlop_3.nPRE.t7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X226 GND.t205 EN.t15 a_6623_61411# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X227 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t8 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X228 GND.t527 VDD.t933 a_42263_59439# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X229 a_11766_45397# Q1.t6 GND.t247 GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X230 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t111 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X231 D_FlipFlop_4.3-input-nand_2.C.t0 D_FlipFlop_4.3-input-nand_2.Vout.t4 VDD.t75 VDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X232 CDAC_v3_0.switch_0.Z.t4 a_11766_45397# VDD.t881 VDD.t880 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X233 GND.t260 EN.t16 a_37849_55365# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X234 VDD.t694 EN.t17 Nand_Gate_7.A.t1 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X235 VDD.t576 D_FlipFlop_3.3-input-nand_1.B D_FlipFlop_3.3-input-nand_1.Vout VDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X236 GND.t192 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t4 a_17315_56723# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X237 a_13751_58825# Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t3 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X238 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_6.Inverter_1.Vout a_2046_48405# GND.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X239 a_20879_56723# Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X240 VDD.t240 CLK.t14 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t0 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X241 a_n9432_48405# FFCLR.t11 GND.t191 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X242 VDD.t241 CLK.t15 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t0 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X243 a_41413_56723# Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X244 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.CLK.t4 a_6734_48405# GND.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X245 VDD.t551 Nand_Gate_3.A.t6 Ring_Counter_0.D_FlipFlop_7.Qbar VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X246 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t31 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X247 VDD.t782 D_FlipFlop_6.3-input-nand_2.C.t4 D_FlipFlop_6.Nand_Gate_1.Vout VDD.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X248 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t110 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X249 VDD.t435 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t0 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X250 GND.t133 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 a_12901_56723# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X251 GND.t241 EN.t18 a_35135_61411# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X252 D_FlipFlop_6.CLK.t1 And_Gate_1.Nand_Gate_0.Vout GND.t345 GND.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X253 GND.t528 VDD.t934 a_10187_55365# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X254 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t52 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X255 a_n4069_59439# Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 a_n4069_58825# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X256 a_52105_61411# Ring_Counter_0.D_FlipFlop_16.Q.t4 a_52105_60797# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X257 a_9337_60797# CLK.t16 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X258 GND.t718 Q7.t5 CDAC_v3_0.switch_6.Z.t131 VDD.t911 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X259 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.CLK.t4 VDD.t258 VDD.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X260 GND.t529 VDD.t935 a_30721_61411# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X261 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t51 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X262 VDD.t202 VDD.t201 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X263 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 VDD.t515 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X264 GND.t530 VDD.t936 a_24443_55365# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X265 VDD.t693 EN.t19 Nand_Gate_2.A.t3 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X266 a_43140_51119# D_FlipFlop_1.nPRE.t5 GND.t654 GND.t653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X267 GND.t531 VDD.t937 a_3059_59439# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X268 a_45827_61411# Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B a_45827_60797# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X269 a_38699_58825# Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t1 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X270 a_47828_51119# D_FlipFlop_1.Nand_Gate_0.Vout a_47214_51119# GND.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X271 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t109 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X272 VDD.t500 Ring_Counter_0.D_FlipFlop_12.Qbar D_FlipFlop_6.nPRE.t1 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X273 GND.t349 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 a_37849_56723# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X274 GND.t486 GND.t487 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X275 a_2209_56723# Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X276 GND.t61 D_FlipFlop_6.nPRE.t7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X277 VDD.t447 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t1 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X278 VDD.t242 CLK.t17 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X279 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t4 VDD.t867 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X280 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t5 VDD.t393 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X281 Q7.t2 FFCLR.t12 VDD.t357 VDD.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X282 VDD.t814 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t2 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X283 a_n4919_54751# Ring_Counter_0.D_FlipFlop_16.Qbar Ring_Counter_0.D_FlipFlop_16.Q.t3 GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X284 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t108 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X285 GND.t484 GND.t485 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X286 a_29690_51119# D_FlipFlop_3.nPRE.t8 GND.t595 GND.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X287 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.CLK.t3 VDD.t612 VDD.t611 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X288 a_27157_54751# Ring_Counter_0.D_FlipFlop_7.Qbar Nand_Gate_3.A.t2 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X289 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t107 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X290 VDD.t380 Nand_Gate_0.A.t5 Ring_Counter_0.D_FlipFlop_13.Qbar VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X291 And_Gate_7.Nand_Gate_0.Vout CLK.t18 a_49577_52049# GND.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X292 GND.t78 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t4 a_10187_56723# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X293 D_FlipFlop_1.3-input-nand_2.Vout.t0 D_FlipFlop_1.3-input-nand_2.C.t4 VDD.t281 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X294 a_n4744_51119# D_FlipFlop_7.Nand_Gate_0.Vout a_n5358_51119# GND.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X295 a_49391_54751# FFCLR.t13 Ring_Counter_0.D_FlipFlop_0.Qbar GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X296 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t50 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X297 Q2.t1 D_FlipFlop_4.Qbar a_12780_51119# GND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X298 VDD.t379 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X299 VDD.t200 VDD.t198 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X300 And_Gate_5.Nand_Gate_0.Vout CLK.t19 a_32053_52049# GND.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X301 GND.t580 D_FlipFlop_2.nPRE.t6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X302 GND.t240 EN.t20 a_44977_55365# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X303 VDD.t338 Nand_Gate_7.A.t4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X304 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t7 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X305 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t106 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X306 GND.t532 VDD.t938 a_20879_59439# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X307 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.CLK.t4 VDD.t461 VDD.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X308 GND.t676 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t4 a_24443_56723# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X309 GND.t673 EN.t21 a_41413_59439# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X310 a_17315_58825# Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t2 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X311 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 VDD.t791 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X312 VDD.t438 D_FlipFlop_5.Nand_Gate_0.Vout Q3.t3 VDD.t400 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X313 VDD.t291 CLK.t20 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t0 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X314 GND.t161 FFCLR.t14 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X315 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 VDD.t592 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X316 VDD.t79 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.3-input-nand_2.Vout.t0 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X317 VDD.t85 Nand_Gate_4.A.t4 Ring_Counter_0.D_FlipFlop_5.Qbar.t2 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X318 VDD.t197 VDD.t196 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t2 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X319 a_10808_51119# D_FlipFlop_4.3-input-nand_2.Vout.t5 GND.t52 GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X320 GND.t533 VDD.t939 a_20029_61411# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X321 a_n5358_51119# D_FlipFlop_7.nPRE.t5 GND.t105 GND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X322 VDD.t297 And_Gate_5.A And_Gate_5.Nand_Gate_0.Vout VDD.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X323 a_12901_58825# Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X324 GND.t672 EN.t22 a_42263_61411# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X325 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t105 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X326 GND.t271 Nand_Gate_1.A.t5 a_n7004_52049# GND.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X327 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_1.nPRE.t6 VDD.t857 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X328 VDD.t902 D_FlipFlop_6.Nand_Gate_0.Vout Q1.t3 VDD.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X329 VDD.t868 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X330 VDD.t86 Nand_Gate_4.A.t5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X331 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t104 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X332 D_FlipFlop_0.3-input-nand_2.C.t3 D_FlipFlop_0.3-input-nand_2.Vout.t5 a_52516_48405# GND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X333 a_13751_60797# CLK.t21 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X334 VDD.t339 Nand_Gate_7.A.t5 Ring_Counter_0.D_FlipFlop_1.Qbar VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X335 D_FlipFlop_0.Qbar EN.t23 VDD.t692 VDD.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X336 GND.t482 GND.t483 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X337 a_14882_51119# FFCLR.t15 GND.t163 GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X338 D_FlipFlop_3.3-input-nand_2.Vout.t2 D_FlipFlop_3.3-input-nand_2.C.t4 VDD.t429 VDD.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X339 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 VDD.t473 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X340 GND.t534 VDD.t940 a_31571_55365# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X341 GND.t535 VDD.t941 a_28007_55365# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X342 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.CLK.t4 VDD.t613 VDD.t611 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X343 a_19570_51119# D_FlipFlop_5.3-input-nand_2.Vout.t4 GND.t216 GND.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X344 VDD.t7 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X345 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t49 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X346 And_Gate_2.Nand_Gate_0.Vout CLK.t22 VDD.t293 VDD.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X347 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t103 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X348 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.CLK.t2 a_15496_51119# GND.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X349 CDAC_v3_0.OUT CDAC_v3_0.switch_8.Z.t2 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X350 D_FlipFlop_4.3-input-nand_2.Vout.t2 D_FlipFlop_4.nPRE.t7 VDD.t590 VDD.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X351 a_5773_54751# Ring_Counter_0.D_FlipFlop_13.Qbar Nand_Gate_0.A.t1 GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X352 a_38452_48405# FFCLR.t16 GND.t165 GND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X353 D_FlipFlop_1.3-input-nand_2.C.t0 D_FlipFlop_1.3-input-nand_2.Vout.t4 VDD.t457 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X354 a_n4069_61411# Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B a_n4069_60797# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X355 a_34992_48405# D_FlipFlop_2.3-input-nand_1.Vout a_34378_48405# GND.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X356 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t48 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X357 a_n7633_56723# Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X358 GND.t208 EN.t24 a_2209_59439# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X359 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.CLK.t4 a_41782_51119# GND.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X360 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t30 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X361 GND.t360 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 a_44977_56723# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X362 a_37849_58825# Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X363 GND.t480 GND.t481 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X364 GND.t617 Nand_Gate_2.A.t5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X365 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 VDD.t346 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X366 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t29 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X367 VDD.t707 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X368 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t28 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X369 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t5 VDD.t882 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X370 GND.t574 EN.t25 a_3059_61411# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X371 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Inverter_1.Vout VDD.t505 VDD.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X372 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout Nand_Gate_0.A.t6 VDD.t887 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X373 CDAC_v3_0.switch_3.Z.t1 a_19654_45397# GND.t66 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X374 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Inverter_1.Vout a_19570_51119# GND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X375 VDD.t401 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_5.Qbar VDD.t400 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X376 a_38699_60797# CLK.t23 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X377 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t102 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X378 a_n505_55365# Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 a_n505_54751# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X379 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t101 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X380 VDD.t528 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.3-input-nand_2.C.t0 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X381 VDD.t21 D_FlipFlop_7.D.t8 D_FlipFlop_0.3-input-nand_0.Vout VDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X382 VDD.t294 CLK.t24 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t0 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X383 a_39066_48405# D_FlipFlop_2.Nand_Gate_1.Vout a_38452_48405# GND.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X384 a_34285_54751# Ring_Counter_0.D_FlipFlop_5.Qbar.t5 Nand_Gate_4.A.t2 GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X385 D_FlipFlop_6.Qbar Q1.t7 a_4018_48405# GND.t701 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X386 GND.t123 CLK.t25 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X387 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Inverter_1.Vout VDD.t318 VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X388 VDD.t93 D_FlipFlop_6.nPRE.t8 Ring_Counter_0.D_FlipFlop_12.Qbar VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X389 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t100 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X390 VDD.t691 EN.t26 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X391 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t99 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X392 D_FlipFlop_4.3-input-nand_2.C.t1 D_FlipFlop_4.3-input-nand_2.Vout.t6 a_8706_48405# GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X393 a_10187_58825# Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t2 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X394 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t98 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X395 VDD.t525 Ring_Counter_0.D_FlipFlop_2.Qbar D_FlipFlop_1.nPRE.t0 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X396 And_Gate_1.Nand_Gate_0.Vout CLK.t26 a_n2995_52049# GND.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X397 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t97 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X398 VDD.t419 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_6.Qbar VDD.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X399 And_Gate_5.A Nand_Gate_4.A.t6 VDD.t88 VDD.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X400 D_FlipFlop_4.nPRE.t1 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t587 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X401 a_48541_54751# Ring_Counter_0.D_FlipFlop_1.Qbar Nand_Gate_7.A.t2 GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X402 GND.t478 GND.t479 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X403 GND.t604 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t5 a_31571_56723# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X404 GND.t223 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t6 a_28007_56723# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X405 a_24443_58825# Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t3 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X406 VDD.t780 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X407 D_FlipFlop_3.3-input-nand_2.C.t2 D_FlipFlop_3.3-input-nand_2.Vout.t4 VDD.t432 VDD.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X408 VDD.t295 CLK.t27 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t0 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X409 a_52105_56723# Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t1 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X410 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 VDD.t464 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X411 VDD.t741 D_FlipFlop_2.nPRE.t7 Ring_Counter_0.D_FlipFlop_4.Qbar.t0 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X412 GND.t536 VDD.t942 a_6623_55365# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X413 VDD.t234 CLK.t28 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X414 And_Gate_1.A Nand_Gate_0.A.t7 VDD.t889 VDD.t888 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X415 D_FlipFlop_4.3-input-nand_2.C.t3 FFCLR.t17 VDD.t359 VDD.t358 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X416 VDD.t907 Ring_Counter_0.D_FlipFlop_6.Qbar D_FlipFlop_3.nPRE.t2 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X417 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t47 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X418 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.CLK.t5 a_24258_48405# GND.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X419 a_45827_56723# Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X420 VDD.t370 Nand_Gate_5.A.t4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X421 CDAC_v3_0.switch_6.Z.t0 a_35430_45397# VDD.t315 VDD.t314 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X422 VDD.t235 CLK.t29 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t0 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X423 GND.t209 EN.t27 a_20879_61411# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X424 a_17315_60797# CLK.t30 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X425 GND.t537 VDD.t943 a_41413_61411# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X426 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_3.Inverter_1.Vout VDD.t504 VDD.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X427 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t5 VDD.t33 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X428 VDD.t195 VDD.t194 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t1 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X429 VDD.t690 EN.t28 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t3 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X430 D_FlipFlop_0.3-input-nand_1.B D_FlipFlop_7.D.t9 GND.t18 GND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X431 GND.t538 VDD.t944 a_35135_55365# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X432 VDD.t289 D_FlipFlop_0.3-input-nand_1.B D_FlipFlop_0.3-input-nand_1.Vout VDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X433 a_12901_60797# CLK.t31 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X434 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 VDD.t373 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X435 a_n1355_55365# Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_n1355_54751# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X436 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_0.Inverter_1.Vout VDD.t317 VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X437 VDD.t884 a_50502_29172.t2 D_FlipFlop_7.D.t1 VDD.t883 sky130_fd_pr__pfet_g5v0d10v5 ad=17.4 pd=120.58 as=17.4 ps=120.58 w=60 l=1
X438 a_9337_54751# Ring_Counter_0.D_FlipFlop_12.Qbar D_FlipFlop_6.nPRE.t2 GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X439 D_FlipFlop_7.3-input-nand_1.B D_FlipFlop_7.D.t10 VDD.t756 VDD.t755 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X440 GND.t539 VDD.t945 a_n7633_59439# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X441 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t96 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X442 GND.t354 EN.t29 a_30721_55365# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X443 a_n2028_51119# D_FlipFlop_7.D.t11 a_n2642_51119# GND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X444 a_34378_51119# D_FlipFlop_2.nPRE.t8 GND.t582 GND.t581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X445 a_44977_58825# Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X446 a_n6716_51119# D_FlipFlop_7.3-input-nand_2.Vout.t4 GND.t130 GND.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X447 Q4.t3 D_FlipFlop_3.Qbar a_30304_51119# GND.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X448 VDD.t689 EN.t30 Nand_Gate_5.A.t3 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X449 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t6 VDD.t768 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X450 VDD.t236 CLK.t32 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X451 D_FlipFlop_7.3-input-nand_2.Vout.t2 D_FlipFlop_7.3-input-nand_2.C.t4 VDD.t617 VDD.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X452 VDD.t9 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X453 VDD.t270 D_FlipFlop_7.nPRE.t6 And_Gate_0.A VDD.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X454 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t19 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X455 a_50502_29172.t3 D_FlipFlop_7.D.t2 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X456 GND.t193 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t5 a_6623_56723# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X457 VDD.t237 CLK.t33 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t0 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X458 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t95 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X459 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t46 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X460 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t6 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X461 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t94 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X462 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Inverter_1.Vout a_n6716_51119# GND.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X463 GND.t540 VDD.t946 a_2209_61411# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X464 a_n2642_51119# FFCLR.t18 GND.t167 GND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X465 a_37849_60797# CLK.t34 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X466 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t6 VDD.t708 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X467 a_32053_52049# And_Gate_5.A GND.t126 GND.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X468 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t27 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X469 Q5.t3 D_FlipFlop_2.Qbar a_39066_51119# GND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X470 GND.t476 GND.t477 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X471 Nand_Gate_6.A.t2 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t410 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X472 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.CLK.t5 GND.t263 GND.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X473 a_n10790_48405# D_FlipFlop_7.3-input-nand_1.B a_n11404_48405# GND.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X474 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t26 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X475 GND.t474 GND.t475 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X476 GND.t472 GND.t473 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X477 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t45 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X478 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t93 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X479 GND.t42 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t6 a_35135_56723# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X480 a_31571_58825# Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X481 GND.t541 VDD.t947 a_52105_59439# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X482 a_28007_58825# Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t3 GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X483 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t25 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X484 Q3.t2 D_FlipFlop_5.nPRE.t6 VDD.t788 VDD.t635 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X485 VDD.t238 CLK.t35 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t0 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X486 a_12166_51119# D_FlipFlop_4.nPRE.t8 GND.t289 GND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X487 GND.t470 GND.t471 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X488 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t92 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X489 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t91 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X490 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t90 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X491 D_FlipFlop_3.3-input-nand_2.Vout.t1 D_FlipFlop_3.nPRE.t9 VDD.t752 VDD.t637 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X492 D_FlipFlop_7.3-input-nand_2.Vout.t3 D_FlipFlop_7.3-input-nand_2.C.t5 a_n8818_51119# GND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X493 VDD.t193 VDD.t192 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X494 a_10187_60797# CLK.t36 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X495 VDD.t853 Q2.t4 CDAC_v3_0.switch_2.Z.t6 GND.t650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X496 VDD.t858 D_FlipFlop_1.nPRE.t7 Ring_Counter_0.D_FlipFlop_2.Qbar VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X497 VDD.t688 EN.t31 D_FlipFlop_7.nPRE.t2 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X498 a_16854_51119# D_FlipFlop_5.nPRE.t7 GND.t172 GND.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X499 VDD.t266 Ring_Counter_0.D_FlipFlop_4.Qbar.t4 D_FlipFlop_2.nPRE.t0 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X500 GND.t267 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 a_30721_56723# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X501 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t89 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X502 Ring_Counter_0.D_FlipFlop_10.Qbar.t0 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 VDD.t11 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X503 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t88 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X504 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.CLK.t3 GND.t179 GND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X505 And_Gate_2.Nand_Gate_0.Vout CLK.t37 a_5767_52049# GND.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X506 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t0 Ring_Counter_0.D_FlipFlop_16.Q.t5 VDD.t219 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X507 GND.t542 VDD.t948 a_45827_59439# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X508 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t44 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X509 GND.t468 GND.t469 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X510 GND.t466 GND.t467 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X511 VDD.t595 And_Gate_4.A And_Gate_4.Nand_Gate_0.Vout VDD.t594 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X512 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t87 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X513 a_24443_60797# CLK.t38 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X514 GND.t662 EN.t32 a_20029_55365# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X515 D_FlipFlop_7.3-input-nand_2.C.t0 D_FlipFlop_7.3-input-nand_2.Vout.t5 VDD.t304 VDD.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X516 Q4.t0 D_FlipFlop_3.nPRE.t10 VDD.t753 VDD.t639 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X517 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t6 VDD.t860 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X518 a_n4069_56723# Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X519 VDD.t382 Q5.t5 CDAC_v3_0.switch_5.Z.t0 GND.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X520 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t24 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X521 Ring_Counter_0.D_FlipFlop_6.Qbar Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 VDD.t360 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X522 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t328 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X523 a_15710_45397# Q2.t5 GND.t652 GND.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X524 GND.t543 VDD.t949 a_42263_55365# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X525 D_FlipFlop_1.3-input-nand_2.C.t1 D_FlipFlop_1.3-input-nand_2.Vout.t5 a_43754_48405# GND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X526 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t86 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X527 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t85 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X528 VDD.t599 And_Gate_2.A And_Gate_2.Nand_Gate_0.Vout VDD.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X529 VDD.t743 CLK.t39 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X530 Q2.t0 D_FlipFlop_4.Qbar VDD.t412 VDD.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X531 a_13751_54751# D_FlipFlop_4.nPRE.t9 Ring_Counter_0.D_FlipFlop_10.Qbar.t3 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X532 And_Gate_4.Nand_Gate_0.Vout CLK.t40 VDD.t745 VDD.t744 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X533 a_19654_45397# Q3.t4 GND.t611 GND.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X534 a_21542_48405# D_FlipFlop_5.Nand_Gate_1.Vout a_20928_48405# GND.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X535 VDD.t687 EN.t33 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X536 VDD.t686 EN.t34 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X537 GND.t20 Nand_Gate_4.A.t7 a_36806_52049# GND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X538 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t7 VDD.t54 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X539 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t84 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X540 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 VDD.t311 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X541 D_FlipFlop_5.Qbar FFCLR.t19 VDD.t636 VDD.t635 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X542 a_6623_58825# Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t0 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X543 D_FlipFlop_3.3-input-nand_2.C.t1 FFCLR.t20 VDD.t638 VDD.t637 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X544 VDD.t216 D_FlipFlop_4.3-input-nand_2.Vout.t7 D_FlipFlop_4.Nand_Gate_0.Vout VDD.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X545 GND.t290 D_FlipFlop_4.nPRE.t10 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X546 GND.t234 EN.t35 a_n7633_61411# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X547 a_4018_48405# D_FlipFlop_6.Nand_Gate_1.Vout a_3404_48405# GND.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X548 VDD.t546 D_FlipFlop_0.3-input-nand_2.Vout.t6 D_FlipFlop_0.Nand_Gate_0.Vout VDD.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X549 VDD.t757 D_FlipFlop_7.D.t12 D_FlipFlop_5.3-input-nand_0.Vout VDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X550 a_45856_51119# D_FlipFlop_1.3-input-nand_2.Vout.t6 GND.t258 GND.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X551 a_44977_60797# CLK.t41 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X552 VDD.t552 Nand_Gate_3.A.t7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X553 GND.t464 GND.t465 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X554 a_16465_55365# Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_16465_54751# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X555 CDAC_v3_0.switch_7.Z.t0 a_31486_45397# VDD.t302 VDD.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X556 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.CLK.t5 VDD.t486 VDD.t485 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X557 GND.t679 Nand_Gate_0.A.t8 a_1758_52049# GND.t678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X558 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout Nand_Gate_1.A.t6 VDD.t467 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X559 D_FlipFlop_5.Qbar Q3.t5 a_21542_48405# GND.t612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X560 Nand_Gate_3.A.t0 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD.t522 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X561 GND.t544 VDD.t950 a_3059_55365# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X562 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t23 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X563 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t22 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X564 a_38699_54751# Nand_Gate_5.A.t5 Ring_Counter_0.D_FlipFlop_3.Qbar.t1 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X565 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t21 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X566 GND.t303 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 a_20029_56723# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X567 D_FlipFlop_3.3-input-nand_2.C.t3 D_FlipFlop_3.3-input-nand_2.Vout.t5 a_26230_48405# GND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X568 D_FlipFlop_3.Qbar FFCLR.t21 VDD.t640 VDD.t639 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X569 GND.t618 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t6 a_42263_56723# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X570 a_35135_58825# Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t2 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X571 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t18 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X572 VDD.t746 CLK.t42 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t0 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X573 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t83 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X574 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.CLK.t3 VDD.t38 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X575 VDD.t641 FFCLR.t22 Ring_Counter_0.D_FlipFlop_0.Qbar VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X576 VDD.t704 D_FlipFlop_6.nPRE.t9 And_Gate_1.A VDD.t703 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X577 VDD.t775 Q0.t6 CDAC_v3_0.switch_8.Z.t0 GND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X578 VDD.t556 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X579 D_FlipFlop_4.Qbar Q2.t6 VDD.t854 VDD.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X580 VDD.t271 D_FlipFlop_7.nPRE.t7 Ring_Counter_0.D_FlipFlop_14.Qbar.t1 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X581 a_30721_58825# Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X582 Ring_Counter_0.D_FlipFlop_8.Qbar.t3 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 VDD.t404 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X583 Ring_Counter_0.D_FlipFlop_9.Qbar Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 VDD.t575 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X584 GND.t590 Nand_Gate_5.A.t6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X585 GND.t226 Nand_Gate_6.A.t6 a_19282_52049# GND.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X586 a_24258_48405# D_FlipFlop_3.3-input-nand_1.B a_23644_48405# GND.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X587 VDD.t354 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X588 VDD.t642 FFCLR.t23 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X589 D_FlipFlop_2.3-input-nand_1.B D_FlipFlop_7.D.t13 GND.t598 GND.t597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X590 a_n505_59439# Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 a_n505_58825# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X591 GND.t545 VDD.t951 a_n4069_59439# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X592 a_31571_60797# CLK.t43 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X593 a_28007_60797# CLK.t44 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X594 GND.t355 EN.t36 a_52105_61411# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X595 a_50544_48405# D_FlipFlop_0.3-input-nand_1.B a_49930_48405# GND.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X596 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t82 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X597 D_FlipFlop_2.CLK.t1 And_Gate_5.Nand_Gate_0.Vout GND.t513 GND.t512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X598 GND.t462 GND.t463 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X599 VDD.t827 D_FlipFlop_4.3-input-nand_2.C.t5 D_FlipFlop_4.Nand_Gate_1.Vout VDD.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X600 D_FlipFlop_6.3-input-nand_2.Vout.t1 D_FlipFlop_6.3-input-nand_2.C.t5 a_n56_51119# GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X601 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B VDD.t319 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X602 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t20 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X603 VDD.t327 D_FlipFlop_0.3-input-nand_2.C.t5 D_FlipFlop_0.Nand_Gate_1.Vout VDD.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X604 VDD.t69 D_FlipFlop_5.3-input-nand_1.B D_FlipFlop_5.3-input-nand_1.Vout VDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X605 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD.t512 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X606 GND.t460 GND.t461 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X607 GND.t356 EN.t37 a_45827_61411# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X608 GND.t585 CLK.t45 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t1 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X609 GND.t546 VDD.t952 a_20879_55365# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X610 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.CLK.t4 a_n2028_51119# GND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X611 GND.t357 EN.t38 a_41413_55365# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X612 a_17315_54751# Nand_Gate_6.A.t7 Ring_Counter_0.D_FlipFlop_9.Qbar GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X613 GND.t29 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t6 a_3059_56723# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X614 a_32406_48405# D_FlipFlop_2.nPRE.t9 GND.t116 GND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X615 VDD.t191 VDD.t189 FFCLR.t0 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X616 VDD.t758 D_FlipFlop_7.D.t14 D_FlipFlop_4.3-input-nand_0.Vout VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X617 Nand_Gate_0.A.t3 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t724 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X618 VDD.t492 D_FlipFlop_4.nPRE.t11 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X619 a_12901_54751# Ring_Counter_0.D_FlipFlop_11.Qbar.t4 Nand_Gate_2.A.t1 GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X620 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t7 VDD.t803 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X621 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 VDD.t320 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X622 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t19 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X623 And_Gate_0.A Nand_Gate_1.A.t7 VDD.t469 VDD.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X624 VDD.t579 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X625 VDD.t363 Ring_Counter_0.D_FlipFlop_8.Qbar.t5 D_FlipFlop_5.nPRE.t1 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X626 VDD.t778 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X627 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.CLK.t4 VDD.t39 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X628 GND.t458 GND.t459 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X629 a_23593_55365# Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_23593_54751# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X630 GND.t91 CLK.t46 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t1 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X631 VDD.t188 VDD.t187 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X632 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t81 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X633 Nand_Gate_4.A.t0 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD.t398 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X634 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.CLK.t5 a_n10790_48405# GND.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X635 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t43 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X636 a_20029_58825# Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X637 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t42 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X638 GND.t456 GND.t457 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X639 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t80 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X640 a_n1355_59439# Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout a_n1355_58825# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X641 a_6623_60797# CLK.t47 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X642 a_42263_58825# Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t1 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X643 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t17 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X644 GND.t235 EN.t39 a_2209_55365# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X645 GND.t454 GND.t455 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X646 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t41 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X647 VDD.t248 CLK.t48 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X648 a_37849_54751# Ring_Counter_0.D_FlipFlop_4.Qbar.t5 D_FlipFlop_2.nPRE.t1 GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X649 GND.t452 GND.t453 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X650 VDD.t186 VDD.t185 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t0 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X651 CDAC_v3_0.switch_2.Z.t1 a_15710_45397# GND.t317 GND.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X652 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t79 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X653 VDD.t249 CLK.t49 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t0 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X654 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X655 GND.t635 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t6 a_20879_56723# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X656 VDD.t886 Ring_Counter_0.D_FlipFlop_1.Qbar Nand_Gate_7.A.t3 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X657 GND.t181 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 a_41413_56723# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X658 GND.t450 GND.t451 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X659 Ring_Counter_0.D_FlipFlop_7.Qbar Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 VDD.t366 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X660 GND.t155 Nand_Gate_7.A.t6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X661 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t18 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X662 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t78 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X663 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t77 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X664 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t17 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X665 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t16 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X666 VDD.t95 D_FlipFlop_4.3-input-nand_1.B D_FlipFlop_4.3-input-nand_1.Vout VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X667 D_FlipFlop_2.3-input-nand_2.Vout.t1 D_FlipFlop_2.3-input-nand_2.C.t5 VDD.t535 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X668 a_35135_60797# CLK.t50 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X669 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t76 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X670 VDD.t685 EN.t40 Ring_Counter_0.D_FlipFlop_16.Q.t1 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X671 a_10187_54751# Nand_Gate_2.A.t6 Ring_Counter_0.D_FlipFlop_11.Qbar.t2 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X672 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t40 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X673 GND.t448 GND.t449 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X674 CDAC_v3_0.switch_5.Z.t3 a_27542_45397# GND.t509 GND.t508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X675 GND.t446 GND.t447 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X676 a_30721_60797# CLK.t51 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X677 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.CLK.t5 VDD.t840 VDD.t839 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X678 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD.t806 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X679 GND.t93 CLK.t52 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t1 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X680 VDD.t499 D_FlipFlop_4.Nand_Gate_0.Vout Q2.t3 VDD.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X681 a_24443_54751# Nand_Gate_3.A.t8 Ring_Counter_0.D_FlipFlop_7.Qbar GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X682 VDD.t305 Ring_Counter_0.D_FlipFlop_11.Qbar.t5 Nand_Gate_2.A.t2 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X683 VDD.t250 CLK.t53 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X684 VDD.t908 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X685 VDD.t922 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.3-input-nand_2.Vout.t3 VDD.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X686 a_3059_58825# Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t3 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X687 a_n505_61411# Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B a_n505_60797# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X688 GND.t663 EN.t41 a_n4069_61411# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X689 a_20928_48405# FFCLR.t24 GND.t511 GND.t510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X690 D_FlipFlop_6.nPRE.t0 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t267 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X691 VDD.t759 D_FlipFlop_7.D.t15 D_FlipFlop_7.3-input-nand_0.Vout VDD.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X692 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t4 VDD.t845 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X693 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t75 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X694 GND.t629 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 a_2209_56723# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X695 VDD.t184 VDD.t183 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t0 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X696 GND.t444 GND.t445 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X697 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t5 VDD.t779 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X698 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout D_FlipFlop_7.nPRE.t8 VDD.t912 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X699 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 VDD.t279 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X700 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t15 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X701 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t74 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X702 a_n4919_55365# Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_n4919_54751# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X703 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.CLK.t6 GND.t301 GND.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X704 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t39 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X705 D_FlipFlop_5.3-input-nand_2.Vout.t2 D_FlipFlop_5.3-input-nand_2.C.t4 VDD.t737 VDD.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X706 a_49930_51119# EN.t42 GND.t237 GND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X707 a_27157_55365# Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_27157_54751# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X708 a_1758_52049# D_FlipFlop_6.nPRE.t10 And_Gate_1.A GND.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X709 VDD.t182 VDD.t181 Ring_Counter_0.D_FlipFlop_15.Qbar.t0 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X710 Ring_Counter_0.D_FlipFlop_13.Qbar Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 VDD.t727 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X711 a_49391_55365# Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout a_49391_54751# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X712 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 VDD.t445 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X713 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t73 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X714 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t38 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X715 D_FlipFlop_2.3-input-nand_2.C.t2 D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t3 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X716 D_FlipFlop_7.3-input-nand_0.Vout FFCLR.t25 VDD.t644 VDD.t643 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X717 a_26230_48405# D_FlipFlop_3.3-input-nand_1.Vout a_25616_48405# GND.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X718 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.CLK.t3 a_33020_51119# GND.t579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X719 GND.t547 VDD.t953 a_n7633_55365# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X720 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t16 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X721 a_52516_48405# D_FlipFlop_0.3-input-nand_1.Vout a_51902_48405# GND.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X722 a_44977_54751# Ring_Counter_0.D_FlipFlop_2.Qbar D_FlipFlop_1.nPRE.t1 GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X723 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t72 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X724 a_20879_58825# Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t1 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X725 CDAC_v3_0.switch_8.Z.t3 a_7822_45397# GND.t722 GND.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X726 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t37 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X727 VDD.t288 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_4.Qbar VDD.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X728 a_41413_58825# Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X729 GND.t442 GND.t443 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X730 Ring_Counter_0.D_FlipFlop_5.Qbar.t1 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 VDD.t47 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X731 VDD.t466 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.3-input-nand_2.C.t0 VDD.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X732 VDD.t760 D_FlipFlop_7.D.t16 D_FlipFlop_1.3-input-nand_0.Vout VDD.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X733 VDD.t844 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t3 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X734 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t71 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X735 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Inverter_1.Vout VDD.t397 VDD.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X736 a_20029_60797# CLK.t54 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X737 a_15496_51119# D_FlipFlop_7.D.t17 a_14882_51119# GND.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X738 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 VDD.t334 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X739 a_n1355_61411# D_FlipFlop_7.nPRE.t9 a_n1355_60797# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X740 GND.t81 CLK.t55 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t1 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X741 VDD.t629 D_FlipFlop_7.3-input-nand_1.B D_FlipFlop_7.3-input-nand_1.Vout VDD.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X742 a_42263_60797# CLK.t56 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X743 GND.t440 GND.t441 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X744 And_Gate_4.A Nand_Gate_3.A.t9 VDD.t554 VDD.t553 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X745 a_n11404_51119# FFCLR.t26 GND.t336 GND.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X746 a_54618_48405# D_FlipFlop_0.3-input-nand_2.C.t6 GND.t145 GND.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X747 Ring_Counter_0.D_FlipFlop_1.Qbar Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 VDD.t606 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X748 VDD.t684 EN.t43 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X749 a_16465_59439# Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout a_16465_58825# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X750 D_FlipFlop_3.3-input-nand_0.Vout FFCLR.t27 VDD.t564 VDD.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X751 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t582 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X752 GND.t82 CLK.t57 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t1 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X753 D_FlipFlop_5.3-input-nand_2.C.t1 D_FlipFlop_5.3-input-nand_2.Vout.t5 VDD.t421 VDD.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X754 VDD.t610 D_FlipFlop_3.3-input-nand_2.Vout.t6 D_FlipFlop_3.Nand_Gate_0.Vout VDD.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X755 VDD.t180 VDD.t179 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t0 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X756 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t14 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X757 a_31571_54751# Nand_Gate_4.A.t8 Ring_Counter_0.D_FlipFlop_5.Qbar.t0 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X758 a_28007_54751# D_FlipFlop_3.nPRE.t11 Ring_Counter_0.D_FlipFlop_6.Qbar GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X759 GND.t548 VDD.t954 a_52105_55365# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X760 VDD.t231 CLK.t58 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X761 a_5773_55365# Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_5773_54751# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X762 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.nPRE.t10 VDD.t913 VDD.t643 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X763 GND.t438 GND.t439 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X764 D_FlipFlop_4.3-input-nand_0.Vout FFCLR.t28 VDD.t565 VDD.t493 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X765 GND.t583 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t4 a_n7633_56723# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X766 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_0.Inverter_1.Vout a_54618_48405# GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X767 a_2209_58825# Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X768 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 VDD.t762 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X769 GND.t549 VDD.t955 a_45827_55365# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X770 CDAC_v3_0.switch_0.Z.t5 a_11766_45397# GND.t675 GND.t674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X771 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 VDD.t616 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X772 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 VDD.t600 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X773 GND.t23 Nand_Gate_4.A.t9 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X774 VDD.t361 Q4.t4 CDAC_v3_0.switch_4.Z.t0 GND.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X775 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t36 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X776 VDD.t232 CLK.t59 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X777 a_3059_60797# CLK.t60 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X778 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t70 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X779 D_FlipFlop_0.3-input-nand_1.B D_FlipFlop_7.D.t18 VDD.t717 VDD.t716 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X780 VDD.t859 D_FlipFlop_1.nPRE.t8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X781 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t15 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X782 VDD.t543 D_FlipFlop_1.3-input-nand_1.B D_FlipFlop_1.3-input-nand_1.Vout VDD.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X783 a_34285_55365# Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_34285_54751# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X784 VDD.t336 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.3-input-nand_2.Vout.t0 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X785 Ring_Counter_0.D_FlipFlop_12.Qbar Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 VDD.t632 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X786 D_FlipFlop_1.Nand_Gate_1.Vout D_FlipFlop_1.Inverter_1.Vout VDD.t396 VDD.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X787 a_37094_48405# D_FlipFlop_2.3-input-nand_2.C.t6 GND.t716 GND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X788 D_FlipFlop_1.nPRE.t3 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD.t923 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X789 VDD.t683 EN.t44 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X790 VDD.t742 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X791 CDAC_v3_0.switch_4.Z.t3 a_23598_45397# GND.t202 GND.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X792 VDD.t233 CLK.t61 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X793 D_FlipFlop_3.CLK.t0 And_Gate_4.Nand_Gate_0.Vout VDD.t597 VDD.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X794 VDD.t508 Q7.t6 CDAC_v3_0.switch_6.Z.t2 GND.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X795 a_48541_55365# Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_48541_54751# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X796 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t69 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X797 a_23598_45397# Q4.t5 GND.t170 GND.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X798 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 VDD.t623 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X799 CDAC_v3_0.OUT CDAC_v3_0.switch_2.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X800 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.nPRE.t12 VDD.t754 VDD.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X801 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t35 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X802 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t68 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X803 VDD.t682 EN.t45 Nand_Gate_1.A.t0 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X804 a_2046_48405# D_FlipFlop_6.3-input-nand_2.C.t6 GND.t196 GND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X805 VDD.t431 D_FlipFlop_3.3-input-nand_2.C.t5 D_FlipFlop_3.Nand_Gate_1.Vout VDD.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X806 GND.t242 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t6 a_52105_56723# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X807 D_FlipFlop_6.3-input-nand_2.Vout.t3 D_FlipFlop_6.nPRE.t11 VDD.t705 VDD.t566 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X808 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD.t581 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X809 Ring_Counter_0.D_FlipFlop_4.Qbar.t3 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 VDD.t702 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X810 a_6734_48405# D_FlipFlop_4.3-input-nand_1.B a_6120_48405# GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X811 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B VDD.t80 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X812 D_FlipFlop_3.nPRE.t0 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD.t491 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X813 a_6623_54751# D_FlipFlop_6.nPRE.t12 Ring_Counter_0.D_FlipFlop_12.Qbar GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X814 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.nPRE.t12 VDD.t494 VDD.t493 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X815 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t34 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X816 GND.t436 GND.t437 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X817 GND.t565 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t7 a_45827_56723# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X818 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t33 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X819 a_35430_45397# Q7.t7 GND.t298 GND.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X820 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t32 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X821 VDD.t890 Nand_Gate_0.A.t9 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X822 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t31 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X823 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X824 a_30304_51119# D_FlipFlop_3.Nand_Gate_0.Vout a_29690_51119# GND.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X825 a_n505_56723# Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X826 a_23593_59439# Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout a_23593_58825# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X827 a_20879_60797# CLK.t62 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X828 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t14 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X829 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.CLK.t6 GND.t516 GND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X830 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t13 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X831 a_41413_60797# CLK.t63 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X832 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t13 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X833 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t67 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X834 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t906 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X835 GND.t139 CLK.t64 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X836 GND.t141 CLK.t65 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t1 GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X837 Q2.t2 D_FlipFlop_4.nPRE.t13 VDD.t731 VDD.t568 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X838 VDD.t221 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t2 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X839 GND.t434 GND.t435 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X840 a_35135_54751# D_FlipFlop_2.nPRE.t10 Ring_Counter_0.D_FlipFlop_4.Qbar.t1 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X841 VDD.t877 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.3-input-nand_2.C.t3 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X842 VDD.t321 CLK.t66 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X843 a_47214_51119# D_FlipFlop_1.nPRE.t9 GND.t656 GND.t655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X844 a_9337_55365# Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_9337_54751# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X845 VDD.t621 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X846 GND.t173 D_FlipFlop_5.nPRE.t8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X847 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t66 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X848 a_n7633_58825# Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t3 GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X849 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t30 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X850 a_30721_54751# Ring_Counter_0.D_FlipFlop_6.Qbar D_FlipFlop_3.nPRE.t3 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X851 a_16465_61411# Nand_Gate_6.A.t8 a_16465_60797# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X852 VDD.t50 Ring_Counter_0.D_FlipFlop_3.Qbar.t4 Nand_Gate_5.A.t1 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X853 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 VDD.t284 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X854 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.CLK.t6 a_50544_51119# GND.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X855 D_FlipFlop_2.3-input-nand_2.Vout.t3 D_FlipFlop_2.3-input-nand_2.C.t7 a_34992_51119# GND.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X856 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t65 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X857 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B VDD.t437 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X858 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t29 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X859 VDD.t681 EN.t46 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X860 VDD.t322 CLK.t67 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X861 VDD.t323 CLK.t68 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X862 GND.t550 VDD.t956 a_n4069_55365# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X863 D_FlipFlop_6.3-input-nand_2.C.t2 FFCLR.t29 VDD.t567 VDD.t566 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X864 VDD.t548 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.3-input-nand_2.Vout.t3 VDD.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X865 Q0.t1 D_FlipFlop_7.Qbar a_n4744_51119# GND.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X866 a_2209_60797# CLK.t69 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X867 Q6.t0 D_FlipFlop_1.Qbar VDD.t477 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X868 a_n8818_51119# D_FlipFlop_7.3-input-nand_0.Vout a_n9432_51119# GND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X869 a_33020_51119# D_FlipFlop_7.D.t19 a_32406_51119# GND.t569 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X870 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t64 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X871 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t63 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X872 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t12 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X873 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Inverter_1.Vout a_37094_51119# GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X874 a_51902_48405# EN.t47 GND.t708 GND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X875 a_12780_48405# D_FlipFlop_4.Nand_Gate_1.Vout a_12166_48405# GND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X876 GND.t325 Nand_Gate_3.A.t10 a_28044_52049# GND.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X877 a_n1355_56723# Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X878 a_56590_48405# D_FlipFlop_0.Nand_Gate_1.Vout a_55976_48405# GND.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X879 a_17468_48405# D_FlipFlop_5.3-input-nand_1.Vout a_16854_48405# GND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X880 D_FlipFlop_4.Qbar FFCLR.t30 VDD.t569 VDD.t568 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X881 a_52105_58825# Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t0 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X882 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD.t608 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X883 Ring_Counter_0.D_FlipFlop_2.Qbar Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 VDD.t345 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X884 GND.t432 GND.t433 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X885 D_FlipFlop_1.3-input-nand_0.Vout FFCLR.t31 VDD.t570 VDD.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X886 GND.t142 CLK.t70 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t1 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X887 D_FlipFlop_2.nPRE.t2 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD.t310 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X888 VDD.t865 Ring_Counter_0.D_FlipFlop_14.Qbar.t4 D_FlipFlop_7.nPRE.t3 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X889 VDD.t324 CLK.t71 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X890 VDD.t574 D_FlipFlop_1.3-input-nand_2.Vout.t7 D_FlipFlop_1.Nand_Gate_0.Vout VDD.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X891 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t62 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X892 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Inverter_1.Vout a_2046_51119# GND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X893 a_n9432_51119# D_FlipFlop_7.nPRE.t11 GND.t720 GND.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X894 a_n4919_59439# Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout a_n4919_58825# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X895 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t61 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X896 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.CLK.t7 a_6734_51119# GND.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X897 a_55976_48405# EN.t48 GND.t711 GND.t710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X898 a_45827_58825# Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t2 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X899 GND.t551 VDD.t957 a_n505_59439# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X900 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t60 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X901 VDD.t789 Q3.t6 CDAC_v3_0.switch_3.Z.t10 GND.t613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X902 D_FlipFlop_0.Qbar Q7.t8 a_56590_48405# GND.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X903 D_FlipFlop_5.3-input-nand_2.C.t2 D_FlipFlop_5.3-input-nand_2.Vout.t6 a_17468_48405# GND.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X904 a_27157_59439# Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout a_27157_58825# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X905 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t12 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X906 GND.t106 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t4 a_n4069_56723# GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X907 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 VDD.t331 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X908 VDD.t572 FFCLR.t32 And_Gate_7.A VDD.t571 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X909 a_20029_54751# Ring_Counter_0.D_FlipFlop_9.Qbar Nand_Gate_6.A.t1 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X910 a_49391_59439# Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout a_49391_58825# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X911 GND.t143 CLK.t72 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t1 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X912 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t28 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X913 a_42263_54751# D_FlipFlop_1.nPRE.t10 Ring_Counter_0.D_FlipFlop_2.Qbar GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X914 VDD.t680 EN.t49 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X915 VDD.t243 CLK.t73 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X916 VDD.t917 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X917 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B VDD.t56 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X918 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t27 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X919 GND.t430 GND.t431 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X920 a_3404_48405# FFCLR.t33 GND.t600 GND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X921 VDD.t573 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.3-input-nand_2.C.t2 VDD.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X922 VDD.t178 VDD.t177 Ring_Counter_0.D_FlipFlop_3.Qbar.t0 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X923 a_13751_55365# Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 a_13751_54751# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X924 D_FlipFlop_1.Qbar Q6.t4 VDD.t28 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X925 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Inverter_1.Vout VDD.t441 VDD.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X926 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t11 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X927 a_23593_61411# Nand_Gate_3.A.t11 a_23593_60797# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X928 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 VDD.t849 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X929 And_Gate_7.A Nand_Gate_7.A.t7 VDD.t341 VDD.t340 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X930 VDD.t415 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X931 a_41782_48405# D_FlipFlop_1.3-input-nand_1.B a_41168_48405# GND.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X932 GND.t312 D_FlipFlop_1.nPRE.t11 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X933 D_FlipFlop_3.CLK.t1 And_Gate_4.Nand_Gate_0.Vout GND.t353 GND.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X934 VDD.t244 CLK.t74 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X935 D_FlipFlop_1.Nand_Gate_1.Vout D_FlipFlop_1.Inverter_1.Vout a_45856_48405# GND.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X936 D_FlipFlop_7.CLK.t1 And_Gate_0.Nand_Gate_0.Vout GND.t152 GND.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X937 VDD.t622 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X938 VDD.t220 Ring_Counter_0.D_FlipFlop_16.Q.t6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X939 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t59 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X940 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.nPRE.t12 VDD.t537 VDD.t536 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X941 a_n7633_60797# CLK.t75 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X942 VDD.t283 D_FlipFlop_1.3-input-nand_2.C.t5 D_FlipFlop_1.Nand_Gate_1.Vout VDD.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X943 a_8706_48405# D_FlipFlop_4.3-input-nand_1.Vout a_8092_48405# GND.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X944 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 VDD.t342 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X945 GND.t428 GND.t429 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X946 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t26 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X947 a_38699_55365# Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 a_38699_54751# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X948 a_23644_48405# D_FlipFlop_3.nPRE.t13 GND.t175 GND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X949 VDD.t274 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X950 CDAC_v3_0.switch_6.Z.t1 a_35430_45397# GND.t135 GND.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X951 Q0.t3 D_FlipFlop_7.nPRE.t12 VDD.t914 VDD.t763 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X952 a_3059_54751# Nand_Gate_0.A.t10 Ring_Counter_0.D_FlipFlop_13.Qbar GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X953 a_28332_48405# D_FlipFlop_3.3-input-nand_2.C.t6 GND.t648 GND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X954 GND.t709 EN.t50 a_n1355_59439# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X955 a_5773_59439# Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout a_5773_58825# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X956 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t25 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X957 VDD.t176 VDD.t174 Ring_Counter_0.D_FlipFlop_16.Qbar VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X958 Ring_Counter_0.D_FlipFlop_0.Qbar Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout VDD.t800 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X959 a_6120_48405# D_FlipFlop_4.nPRE.t14 GND.t577 GND.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X960 VDD.t797 And_Gate_0.A And_Gate_0.Nand_Gate_0.Vout VDD.t796 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X961 a_51632_31172.t0 CDAC_v3_0.OUT a_51773_21431.t2 Vbias.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X962 D_FlipFlop_5.3-input-nand_1.B D_FlipFlop_7.D.t20 VDD.t719 VDD.t718 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X963 Ring_Counter_0.D_FlipFlop_14.Qbar.t3 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 VDD.t834 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X964 VDD.t245 CLK.t76 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X965 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 VDD.t381 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X966 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t58 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X967 GND.t646 Nand_Gate_0.A.t11 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X968 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_4.Inverter_1.Vout VDD.t440 VDD.t439 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X969 D_FlipFlop_1.3-input-nand_1.B D_FlipFlop_7.D.t21 VDD.t721 VDD.t720 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X970 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_3.Inverter_1.Vout a_28332_48405# GND.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X971 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t57 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X972 a_34285_59439# Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout a_34285_58825# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X973 D_FlipFlop_0.CLK.t0 And_Gate_7.Nand_Gate_0.Vout VDD.t870 VDD.t869 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X974 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 VDD.t850 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X975 a_n4069_58825# Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t3 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X976 a_52105_60797# CLK.t77 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t2 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X977 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t24 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X978 GND.t426 GND.t427 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X979 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t511 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X980 D_FlipFlop_0.3-input-nand_2.Vout.t1 D_FlipFlop_0.3-input-nand_2.C.t7 a_52516_51119# GND.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X981 GND.t89 CLK.t78 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t1 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X982 VDD.t246 CLK.t79 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X983 a_16465_56723# Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X984 a_15710_45397# Q2.t7 VDD.t856 VDD.t855 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X985 VDD.t679 EN.t51 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X986 VDD.t470 Nand_Gate_1.A.t8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X987 a_n4919_61411# Nand_Gate_1.A.t9 a_n4919_60797# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X988 VDD.t264 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X989 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t56 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X990 a_48541_59439# Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout a_48541_58825# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X991 a_45827_60797# CLK.t80 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X992 a_17315_55365# Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 a_17315_54751# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X993 a_20879_54751# D_FlipFlop_5.nPRE.t9 Ring_Counter_0.D_FlipFlop_8.Qbar.t2 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X994 GND.t207 EN.t52 a_n505_61411# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X995 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t55 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X996 a_41413_54751# Ring_Counter_0.D_FlipFlop_3.Qbar.t5 Nand_Gate_5.A.t2 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X997 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t23 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X998 a_27157_61411# D_FlipFlop_3.nPRE.t14 a_27157_60797# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X999 GND.t424 GND.t425 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1000 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t22 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1001 a_38452_51119# D_FlipFlop_2.nPRE.t11 GND.t118 GND.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1002 D_FlipFlop_7.Qbar FFCLR.t34 VDD.t764 VDD.t763 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1003 VDD.t876 Ring_Counter_0.D_FlipFlop_0.Qbar FFCLR.t2 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1004 a_12901_55365# Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_12901_54751# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1005 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 VDD.t918 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1006 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t54 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1007 a_34992_51119# D_FlipFlop_2.3-input-nand_0.Vout a_34378_51119# GND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1008 a_49391_61411# Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B a_49391_60797# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1009 GND.t659 Q2.t8 CDAC_v3_0.switch_2.Z.t7 VDD.t866 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1010 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t10 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1011 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t921 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1012 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 VDD.t825 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1013 VDD.t173 VDD.t172 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t0 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1014 VDD.t171 VDD.t170 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1015 D_FlipFlop_5.nPRE.t3 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t785 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1016 VDD.t247 CLK.t81 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1017 VDD.t30 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1018 VDD.t489 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1019 GND.t422 GND.t423 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1020 And_Gate_6.Nand_Gate_0.Vout CLK.t82 VDD.t225 VDD.t224 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1021 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.CLK.t5 VDD.t41 VDD.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1022 D_FlipFlop_1.3-input-nand_2.Vout.t2 D_FlipFlop_1.nPRE.t13 VDD.t539 VDD.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1023 VDD.t532 D_FlipFlop_1.Nand_Gate_0.Vout Q6.t3 VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1024 VDD.t169 VDD.t168 Ring_Counter_0.D_FlipFlop_11.Qbar.t0 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1025 VDD.t167 VDD.t166 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t0 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1026 a_39066_51119# D_FlipFlop_2.Nand_Gate_0.Vout a_38452_51119# GND.t619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1027 GND.t79 CLK.t83 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t1 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1028 VDD.t226 CLK.t84 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1029 Q1.t1 D_FlipFlop_6.Qbar a_4018_51119# GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1030 VDD.t348 D_FlipFlop_3.Nand_Gate_0.Vout Q4.t1 VDD.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1031 D_FlipFlop_4.3-input-nand_2.Vout.t1 D_FlipFlop_4.3-input-nand_2.C.t6 a_8706_51119# GND.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1032 a_9337_59439# Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout a_9337_58825# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1033 VDD.t423 And_Gate_6.A And_Gate_6.Nand_Gate_0.Vout VDD.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1034 a_37849_55365# Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_37849_54751# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1035 a_2209_54751# Ring_Counter_0.D_FlipFlop_14.Qbar.t5 D_FlipFlop_7.nPRE.t0 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1036 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t53 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1037 Q6.t2 D_FlipFlop_1.nPRE.t14 VDD.t541 VDD.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1038 a_54330_52049# FFCLR.t35 And_Gate_7.A GND.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1039 Nand_Gate_7.A.t0 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD.t634 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1040 VDD.t268 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t2 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1041 a_n11757_52049# And_Gate_0.A GND.t616 GND.t615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1042 VDD.t25 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1043 a_5767_52049# And_Gate_2.A GND.t359 GND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1044 GND.t552 VDD.t958 a_n1355_61411# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1045 D_FlipFlop_2.3-input-nand_0.Vout FFCLR.t36 VDD.t765 VDD.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1046 a_5773_61411# D_FlipFlop_6.nPRE.t13 a_5773_60797# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1047 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t52 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1048 GND.t420 GND.t421 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1049 a_10187_55365# Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 a_10187_54751# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1050 VDD.t893 Q6.t5 CDAC_v3_0.switch_7.Z.t66 GND.t682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1051 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.CLK.t7 a_24258_51119# GND.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1052 VDD.t722 D_FlipFlop_7.D.t22 D_FlipFlop_6.3-input-nand_0.Vout VDD.t487 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1053 VDD.t871 Ring_Counter_0.D_FlipFlop_16.Qbar Ring_Counter_0.D_FlipFlop_16.Q.t2 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1054 GND.t661 EN.t53 a_16465_59439# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1055 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t51 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1056 GND.t148 Nand_Gate_7.A.t8 a_54330_52049# GND.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1057 VDD.t227 CLK.t85 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1058 a_23593_56723# Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1059 a_43754_48405# D_FlipFlop_1.3-input-nand_1.Vout a_43140_48405# GND.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1060 VDD.t678 EN.t54 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1061 VDD.t228 CLK.t86 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1062 D_FlipFlop_1.Qbar Q6.t6 a_47828_48405# GND.t683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1063 a_7822_45397# Q0.t7 VDD.t774 VDD.t773 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1064 VDD.t750 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1065 GND.t80 CLK.t87 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t1 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1066 D_FlipFlop_1.3-input-nand_2.C.t3 FFCLR.t37 VDD.t766 VDD.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1067 a_24443_55365# Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 a_24443_54751# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1068 Nand_Gate_2.A.t0 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t49 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1069 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout Nand_Gate_6.A.t9 VDD.t58 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1070 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t50 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1071 VDD.t82 D_FlipFlop_1.Nand_Gate_1.Vout D_FlipFlop_1.Qbar VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1072 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t49 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1073 CDAC_v3_0.switch_7.Z.t1 a_31486_45397# GND.t128 GND.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1074 a_34285_61411# D_FlipFlop_2.nPRE.t12 a_34285_60797# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1075 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t21 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1076 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Inverter_1.Vout VDD.t66 VDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1077 a_n4069_60797# CLK.t88 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1078 VDD.t577 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_3.Qbar VDD.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1079 CDAC_v3_0.OUT CDAC_v3_0.switch_2.Z.t3 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1080 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 VDD.t497 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1081 a_31486_45397# Q6.t7 GND.t685 GND.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1082 D_FlipFlop_6.3-input-nand_0.Vout FFCLR.t38 VDD.t767 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1083 a_36806_52049# D_FlipFlop_2.nPRE.t13 And_Gate_5.A GND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1084 a_41168_48405# D_FlipFlop_1.nPRE.t15 GND.t314 GND.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1085 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t798 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1086 a_25616_48405# FFCLR.t39 GND.t603 GND.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1087 GND.t74 Ring_Counter_0.D_FlipFlop_16.Q.t7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1088 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t20 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1089 And_Gate_3.A Nand_Gate_6.A.t10 VDD.t60 VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1090 VDD.t165 VDD.t164 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t0 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1091 VDD.t163 VDD.t162 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t0 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1092 VDD.t259 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t2 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1093 VDD.t161 VDD.t160 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1094 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t19 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1095 VDD.t229 CLK.t89 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1096 VDD.t265 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1097 VDD.t230 CLK.t90 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1098 D_FlipFlop_1.Qbar FFCLR.t40 VDD.t559 VDD.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1099 a_48541_61411# FFCLR.t41 a_48541_60797# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1100 D_FlipFlop_5.3-input-nand_0.Vout FFCLR.t42 VDD.t560 VDD.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1101 GND.t418 GND.t419 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1102 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t18 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1103 a_8092_48405# FFCLR.t43 GND.t330 GND.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1104 VDD.t307 D_FlipFlop_5.3-input-nand_2.Vout.t7 D_FlipFlop_5.Nand_Gate_0.Vout VDD.t306 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1105 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.nPRE.t14 VDD.t286 VDD.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1106 VDD.t471 Nand_Gate_1.A.t10 Ring_Counter_0.D_FlipFlop_15.Qbar.t1 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1107 VDD.t677 EN.t55 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1108 a_n56_48405# D_FlipFlop_6.3-input-nand_1.Vout a_n670_48405# GND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1109 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t48 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1110 VDD.t488 D_FlipFlop_6.3-input-nand_1.B D_FlipFlop_6.3-input-nand_1.Vout VDD.t487 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1111 a_n7633_54751# Ring_Counter_0.D_FlipFlop_16.Q.t8 Ring_Counter_0.D_FlipFlop_16.Qbar GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1112 a_44977_55365# Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_44977_54751# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1113 a_11766_45397# Q1.t8 VDD.t904 VDD.t903 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1114 a_n10790_51119# D_FlipFlop_7.D.t23 a_n11404_51119# GND.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1115 a_13751_59439# Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 a_13751_58825# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1116 D_FlipFlop_0.CLK.t1 And_Gate_7.Nand_Gate_0.Vout GND.t665 GND.t664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1117 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t17 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1118 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_4.Inverter_1.Vout a_10808_48405# GND.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1119 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Inverter_1.Vout VDD.t627 VDD.t625 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1120 VDD.t676 EN.t56 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1121 VDD.t675 EN.t57 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1122 GND.t416 GND.t417 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1123 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t7 VDD.t446 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1124 VDD.t520 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1125 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_2.Inverter_1.Vout VDD.t65 VDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1126 GND.t414 GND.t415 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1127 a_n670_48405# FFCLR.t44 GND.t332 GND.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1128 VDD.t407 D_FlipFlop_7.nPRE.t13 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1129 a_9337_61411# Nand_Gate_2.A.t7 a_9337_60797# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1130 a_n4919_56723# Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1131 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.nPRE.t14 VDD.t479 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1132 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t47 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1133 D_FlipFlop_5.CLK.t0 And_Gate_3.Nand_Gate_0.Vout VDD.t527 VDD.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1134 GND.t575 EN.t58 a_23593_59439# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1135 a_27157_56723# Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1136 VDD.t674 EN.t59 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1137 VDD.t26 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1138 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t46 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1139 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.nPRE.t10 VDD.t365 VDD.t364 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1140 a_38699_59439# Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 a_38699_58825# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1141 a_49391_56723# Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1142 VDD.t738 D_FlipFlop_5.3-input-nand_2.C.t5 D_FlipFlop_5.Nand_Gate_1.Vout VDD.t306 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1143 a_31571_55365# Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 a_31571_54751# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1144 a_28007_55365# Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 a_28007_54751# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1145 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout D_FlipFlop_5.nPRE.t11 VDD.t351 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1146 VDD.t624 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t3 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1147 D_FlipFlop_1.3-input-nand_2.Vout.t1 D_FlipFlop_1.3-input-nand_2.C.t6 a_43754_51119# GND.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1148 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t45 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1149 D_FlipFlop_4.3-input-nand_1.B D_FlipFlop_7.D.t24 GND.t249 GND.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1150 And_Gate_6.Nand_Gate_0.Vout CLK.t91 a_40815_52049# GND.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1151 a_52105_54751# Ring_Counter_0.D_FlipFlop_0.Qbar FFCLR.t3 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1152 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout VDD.t771 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1153 GND.t553 VDD.t959 a_16465_61411# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1154 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t44 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1155 CDAC_v3_0.switch_2.Z.t0 a_15710_45397# VDD.t545 VDD.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1156 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t43 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1157 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 VDD.t730 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1158 VDD.t159 VDD.t158 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t0 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1159 VDD.t809 CLK.t92 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1160 VDD.t157 VDD.t155 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1161 a_45827_54751# Nand_Gate_7.A.t9 Ring_Counter_0.D_FlipFlop_1.Qbar GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1162 VDD.t751 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1163 VDD.t810 CLK.t93 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1164 a_21542_51119# D_FlipFlop_5.Nand_Gate_0.Vout a_20928_51119# GND.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1165 GND.t554 VDD.t960 a_n505_55365# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1166 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B VDD.t490 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1167 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_5.Inverter_1.Vout VDD.t626 VDD.t625 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1168 a_23291_52049# And_Gate_4.A GND.t351 GND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1169 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t42 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1170 VDD.t811 CLK.t94 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t0 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1171 a_4018_51119# D_FlipFlop_6.Nand_Gate_0.Vout a_3404_51119# GND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1172 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 VDD.t260 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1173 VDD.t673 EN.t60 D_FlipFlop_4.nPRE.t2 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1174 VDD.t620 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1175 GND.t412 GND.t413 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1176 VDD.t672 EN.t61 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1177 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t3 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1178 VDD.t671 EN.t62 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1179 a_51773_21431.t1 a_50454_10637.t3 Vbias.t6 Vbias.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X1180 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B VDD.t729 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1181 GND.t623 CLK.t95 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t1 GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1182 a_27542_45397# Q5.t6 VDD.t384 VDD.t383 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1183 D_FlipFlop_2.3-input-nand_2.Vout.t2 D_FlipFlop_2.nPRE.t15 VDD.t792 VDD.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1184 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t16 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1185 Q4.t2 D_FlipFlop_3.Qbar VDD.t496 VDD.t495 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1186 Q3.t1 D_FlipFlop_5.Qbar a_21542_51119# GND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1187 a_17315_59439# Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 a_17315_58825# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1188 D_FlipFlop_3.3-input-nand_2.Vout.t3 D_FlipFlop_3.3-input-nand_2.C.t7 a_26230_51119# GND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1189 VDD.t843 And_Gate_7.A And_Gate_7.Nand_Gate_0.Vout VDD.t842 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1190 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t41 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1191 And_Gate_4.Nand_Gate_0.Vout CLK.t96 a_23291_52049# GND.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1192 a_5773_56723# Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1193 VDD.t670 EN.t63 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1194 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t9 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1195 VDD.t601 Ring_Counter_0.D_FlipFlop_15.Qbar.t5 Nand_Gate_1.A.t1 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1196 GND.t410 GND.t411 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1197 And_Gate_0.Nand_Gate_0.Vout CLK.t97 a_n11757_52049# GND.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1198 D_FlipFlop_4.CLK.t0 And_Gate_2.Nand_Gate_0.Vout VDD.t550 VDD.t549 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1199 a_12901_59439# Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout a_12901_58825# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1200 a_6623_55365# Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 a_6623_54751# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1201 CDAC_v3_0.OUT CDAC_v3_0.switch_2.Z.t2 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1202 D_FlipFlop_7.CLK.t0 And_Gate_0.Nand_Gate_0.Vout VDD.t333 VDD.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1203 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD.t920 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1204 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t15 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1205 GND.t266 EN.t64 a_n4919_59439# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1206 VDD.t350 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.3-input-nand_2.Vout.t0 VDD.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1207 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t40 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1208 a_13751_61411# Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B a_13751_60797# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1209 Q5.t2 D_FlipFlop_2.Qbar VDD.t847 VDD.t385 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1210 a_24258_51119# D_FlipFlop_7.D.t25 a_23644_51119# GND.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1211 GND.t232 EN.t65 a_27157_59439# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1212 GND.t38 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t7 a_n505_56723# GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1213 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t14 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1214 And_Gate_7.Nand_Gate_0.Vout CLK.t98 VDD.t813 VDD.t812 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1215 VDD.t154 VDD.t153 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t1 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1216 VDD.t152 VDD.t151 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1217 a_43140_48405# FFCLR.t45 GND.t334 GND.t333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1218 a_34285_56723# Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1219 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t8 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1220 GND.t233 EN.t66 a_49391_59439# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1221 VDD.t521 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1222 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t39 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1223 a_47828_48405# D_FlipFlop_1.Nand_Gate_1.Vout a_47214_48405# GND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1224 a_50544_51119# D_FlipFlop_7.D.t26 a_49930_51119# GND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1225 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t6 VDD.t416 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1226 GND.t670 EN.t67 a_n1355_55365# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1227 VDD.t273 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1228 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t13 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1229 GND.t408 GND.t409 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1230 a_35135_55365# Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 a_35135_54751# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1231 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_3.nPRE.t15 VDD.t367 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1232 D_FlipFlop_5.3-input-nand_2.Vout.t1 D_FlipFlop_5.nPRE.t12 VDD.t353 VDD.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1233 a_37849_59439# Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout a_37849_58825# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1234 a_48541_56723# Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1235 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t38 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1236 a_30721_55365# Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_30721_54751# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1237 GND.t555 VDD.t961 a_23593_61411# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1238 D_FlipFlop_2.3-input-nand_2.C.t1 FFCLR.t46 VDD.t562 VDD.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1239 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t37 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1240 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t313 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1241 GND.t406 GND.t407 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1242 GND.t626 CLK.t99 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1243 CDAC_v3_0.switch_8.Z.t4 a_7822_45397# VDD.t916 VDD.t915 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1244 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t36 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1245 D_FlipFlop_3.Qbar Q4.t6 VDD.t712 VDD.t495 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1246 VDD.t330 D_FlipFlop_7.3-input-nand_2.Vout.t6 D_FlipFlop_7.Nand_Gate_0.Vout VDD.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1247 VDD.t150 VDD.t149 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t0 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1248 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t35 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1249 a_29690_48405# FFCLR.t47 GND.t688 GND.t687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1250 a_32406_51119# FFCLR.t48 GND.t690 GND.t689 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1251 Nand_Gate_5.A.t0 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD.t67 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1252 VDD.t815 CLK.t100 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1253 VDD.t148 VDD.t146 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1254 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t12 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1255 VDD.t514 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1256 a_38699_61411# Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B a_38699_60797# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1257 VDD.t816 CLK.t101 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1258 VDD.t591 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1259 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B VDD.t84 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1260 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t34 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1261 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B VDD.t633 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1262 VDD.t879 D_FlipFlop_1.nPRE.t16 And_Gate_6.A VDD.t878 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1263 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t33 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1264 GND.t404 GND.t405 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1265 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t32 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1266 a_n4744_48405# D_FlipFlop_7.Nand_Gate_1.Vout a_n5358_48405# GND.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1267 a_n4069_54751# Nand_Gate_1.A.t11 Ring_Counter_0.D_FlipFlop_15.Qbar.t2 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1268 D_FlipFlop_4.Qbar Q2.t9 a_12780_48405# GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1269 a_10187_59439# Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 a_10187_58825# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1270 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t31 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1271 VDD.t145 VDD.t144 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t0 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1272 VDD.t669 EN.t68 Nand_Gate_6.A.t3 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1273 VDD.t701 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.3-input-nand_2.C.t0 VDD.t349 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1274 VDD.t668 EN.t69 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1275 D_FlipFlop_2.Qbar Q5.t7 VDD.t386 VDD.t385 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1276 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t30 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1277 GND.t702 Q1.t9 CDAC_v3_0.switch_0.Z.t1 VDD.t905 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1278 a_24443_59439# Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 a_24443_58825# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1279 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD.t872 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1280 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.CLK.t6 a_n10790_51119# GND.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1281 GND.t671 EN.t70 a_5773_59439# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1282 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t11 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1283 And_Gate_6.A Nand_Gate_5.A.t7 VDD.t748 VDD.t747 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1284 GND.t606 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 a_n1355_56723# GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1285 a_10808_48405# D_FlipFlop_4.3-input-nand_2.C.t7 GND.t608 GND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1286 a_9337_56723# Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1287 a_n5358_48405# FFCLR.t49 GND.t692 GND.t691 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1288 GND.t402 GND.t403 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1289 VDD.t143 VDD.t142 Ring_Counter_0.D_FlipFlop_10.Qbar.t1 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1290 D_FlipFlop_5.3-input-nand_2.C.t3 FFCLR.t50 VDD.t898 VDD.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1291 D_FlipFlop_7.nPRE.t1 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t609 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1292 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout D_FlipFlop_6.nPRE.t15 VDD.t480 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1293 GND.t566 Q4.t7 CDAC_v3_0.switch_4.Z.t1 VDD.t713 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1294 VDD.t817 CLK.t102 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1295 a_17315_61411# Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B a_17315_60797# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1296 VDD.t369 D_FlipFlop_3.nPRE.t16 And_Gate_4.A VDD.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1297 VDD.t223 D_FlipFlop_7.3-input-nand_2.C.t6 D_FlipFlop_7.Nand_Gate_1.Vout VDD.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1298 GND.t400 GND.t401 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1299 GND.t637 EN.t71 a_34285_59439# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1300 a_14882_48405# D_FlipFlop_5.nPRE.t13 GND.t160 GND.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1301 VDD.t141 VDD.t139 Ring_Counter_0.D_FlipFlop_6.Qbar VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1302 a_n505_58825# Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t3 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1303 VDD.t138 VDD.t137 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t2 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1304 VDD.t136 VDD.t134 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1305 a_19570_48405# D_FlipFlop_5.3-input-nand_2.C.t6 GND.t68 GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1306 VDD.t667 EN.t72 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1307 a_20029_55365# Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_20029_54751# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1308 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.CLK.t6 a_15496_48405# GND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1309 a_12901_61411# D_FlipFlop_4.nPRE.t15 a_12901_60797# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1310 a_42263_55365# Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 a_42263_54751# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1311 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_2.nPRE.t16 VDD.t793 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1312 GND.t556 VDD.t962 a_n4919_61411# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1313 GND.t398 GND.t399 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1314 VDD.t852 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1315 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.CLK.t6 a_41782_48405# GND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1316 GND.t705 EN.t73 a_48541_59439# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1317 a_44977_59439# Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout a_44977_58825# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1318 a_23598_45397# Q4.t8 VDD.t715 VDD.t714 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1319 VDD.t749 Nand_Gate_5.A.t8 Ring_Counter_0.D_FlipFlop_3.Qbar.t3 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1320 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t11 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1321 GND.t557 VDD.t963 a_27157_61411# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1322 VDD.t666 EN.t74 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1323 D_FlipFlop_2.3-input-nand_1.B D_FlipFlop_7.D.t27 VDD.t451 VDD.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1324 VDD.t133 VDD.t132 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t0 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1325 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_5.Inverter_1.Vout a_19570_48405# GND.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1326 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 VDD.t783 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1327 GND.t558 VDD.t964 a_49391_61411# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1328 VDD.t665 EN.t75 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1329 VDD.t498 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1330 VDD.t818 CLK.t103 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1331 a_20928_51119# D_FlipFlop_5.nPRE.t14 GND.t255 GND.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1332 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t29 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1333 D_FlipFlop_1.CLK.t0 And_Gate_6.Nand_Gate_0.Vout VDD.t726 VDD.t725 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1334 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t7 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1335 VDD.t516 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1336 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B VDD.t217 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1337 GND.t630 CLK.t104 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t1 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1338 D_FlipFlop_6.3-input-nand_2.Vout.t2 D_FlipFlop_6.3-input-nand_2.C.t7 VDD.t394 VDD.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1339 GND.t396 GND.t397 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1340 GND.t706 EN.t76 a_16465_55365# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1341 a_37849_61411# Nand_Gate_5.A.t9 a_37849_60797# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1342 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t28 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1343 And_Gate_0.Nand_Gate_0.Vout CLK.t105 VDD.t820 VDD.t819 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1344 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t27 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1345 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t26 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1346 VDD.t664 EN.t77 Nand_Gate_3.A.t3 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1347 D_FlipFlop_4.CLK.t1 And_Gate_2.Nand_Gate_0.Vout GND.t322 GND.t321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1348 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t25 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1349 VDD.t663 EN.t78 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1350 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t6 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1351 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t24 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1352 a_3059_55365# Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 a_3059_54751# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1353 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t10 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1354 a_31571_59439# Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 a_31571_58825# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1355 a_28007_59439# Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 a_28007_58825# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1356 GND.t206 EN.t79 a_9337_59439# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1357 a_26230_51119# D_FlipFlop_3.3-input-nand_0.Vout a_25616_51119# GND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1358 a_n1355_58825# Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1359 D_FlipFlop_6.3-input-nand_1.B D_FlipFlop_7.D.t28 VDD.t453 VDD.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1360 a_10187_61411# Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B a_10187_60797# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1361 VDD.t821 CLK.t106 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1362 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t23 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1363 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.CLK.t7 GND.t6 GND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1364 CDAC_v3_0.OUT CDAC_v3_0.switch_0.Z.t3 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1365 a_13751_56723# Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1366 VDD.t662 EN.t80 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1367 a_52516_51119# D_FlipFlop_0.3-input-nand_0.Vout a_51902_51119# GND.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1368 VDD.t131 VDD.t130 Ring_Counter_0.D_FlipFlop_8.Qbar.t0 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1369 VDD.t129 VDD.t128 Ring_Counter_0.D_FlipFlop_9.Qbar VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1370 VDD.t808 Ring_Counter_0.D_FlipFlop_16.Q.t9 Ring_Counter_0.D_FlipFlop_16.Qbar VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1371 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout Nand_Gate_2.A.t8 VDD.t405 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1372 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t9 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1373 GND.t394 GND.t395 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1374 And_Gate_5.Nand_Gate_0.Vout CLK.t107 VDD.t823 VDD.t822 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1375 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t22 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1376 D_FlipFlop_7.D.t29 Vbias.t1 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X1377 a_n7004_52049# D_FlipFlop_7.nPRE.t14 And_Gate_0.A GND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1378 VDD.t805 D_FlipFlop_2.Nand_Gate_0.Vout Q5.t1 VDD.t804 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1379 GND.t392 GND.t393 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1380 a_24443_61411# Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B a_24443_60797# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1381 GND.t559 VDD.t965 a_5773_61411# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1382 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.CLK.t4 VDD.t736 VDD.t735 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1383 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t21 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1384 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B VDD.t801 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1385 GND.t154 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 a_16465_56723# GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1386 a_54618_51119# D_FlipFlop_0.3-input-nand_2.Vout.t7 GND.t319 GND.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1387 D_FlipFlop_6.3-input-nand_2.C.t0 D_FlipFlop_6.3-input-nand_2.Vout.t5 VDD.t262 VDD.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1388 VDD.t892 And_Gate_3.A And_Gate_3.Nand_Gate_0.Vout VDD.t891 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1389 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t20 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1390 CDAC_v3_0.OUT CDAC_v3_0.switch_0.Z.t2 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1391 a_n2028_48405# D_FlipFlop_6.3-input-nand_1.B a_n2642_48405# GND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1392 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1393 a_45568_52049# D_FlipFlop_1.nPRE.t17 And_Gate_6.A GND.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1394 VDD.t919 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1395 a_34378_48405# FFCLR.t51 GND.t694 GND.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1396 a_38699_56723# Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1397 a_n6716_48405# D_FlipFlop_7.3-input-nand_2.C.t7 GND.t77 GND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1398 VDD.t824 CLK.t108 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t0 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1399 GND.t390 GND.t391 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1400 D_FlipFlop_3.Qbar Q4.t9 a_30304_48405# GND.t504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1401 VDD.t770 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.3-input-nand_2.Vout.t3 VDD.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1402 a_20879_55365# Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 a_20879_54751# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1403 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t8 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1404 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t19 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1405 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.CLK.t5 VDD.t377 VDD.t376 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1406 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t18 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1407 VDD.t661 EN.t81 Nand_Gate_0.A.t2 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1408 a_41413_55365# Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_41413_54751# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1409 GND.t560 VDD.t966 a_34285_61411# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1410 a_n505_60797# CLK.t109 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1411 VDD.t660 EN.t82 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1412 GND.t388 GND.t389 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1413 VDD.t127 VDD.t125 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t0 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1414 FFCLR.t1 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t3 VDD.t607 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1415 VDD.t124 VDD.t122 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1416 VDD.t659 EN.t83 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1417 VDD.t434 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1418 a_6623_59439# Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 a_6623_58825# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1419 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Inverter_1.Vout a_54618_51119# GND.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1420 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B VDD.t557 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1421 GND.t386 GND.t387 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1422 D_FlipFlop_7.Nand_Gate_1.Vout D_FlipFlop_7.Inverter_1.Vout a_n6716_48405# GND.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1423 VDD.t518 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1424 D_FlipFlop_7.3-input-nand_1.B D_FlipFlop_7.D.t30 GND.t253 GND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1425 And_Gate_3.Nand_Gate_0.Vout CLK.t110 VDD.t829 VDD.t828 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1426 VDD.t337 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t2 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1427 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t10 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1428 a_n2642_48405# D_FlipFlop_6.nPRE.t16 GND.t283 GND.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1429 GND.t101 Nand_Gate_5.A.t10 a_45568_52049# GND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1430 GND.t561 VDD.t967 a_48541_61411# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1431 GND.t114 EN.t84 a_23593_55365# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1432 a_44977_61411# Nand_Gate_7.A.t10 a_44977_60797# GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1433 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t9 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1434 D_FlipFlop_2.Qbar Q5.t8 a_39066_48405# GND.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1435 VDD.t658 EN.t85 Nand_Gate_4.A.t3 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1436 VDD.t657 EN.t86 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1437 VDD.t45 a_51632_31172.t3 a_50502_29172.t1 VDD.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X1438 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B VDD.t848 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1439 VDD.t875 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_2.Qbar VDD.t804 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1440 a_n2995_52049# And_Gate_1.A GND.t343 GND.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1441 VDD.t121 VDD.t120 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1442 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.CLK.t7 VDD.t615 VDD.t614 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1443 VDD.t312 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t1 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1444 VDD.t406 Nand_Gate_2.A.t9 Ring_Counter_0.D_FlipFlop_11.Qbar.t1 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1445 a_37094_51119# D_FlipFlop_2.3-input-nand_2.Vout.t7 GND.t2 GND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1446 a_35135_59439# Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 a_35135_58825# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1447 a_12166_48405# FFCLR.t52 GND.t696 GND.t695 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1448 GND.t384 GND.t385 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1449 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t17 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1450 D_FlipFlop_7.3-input-nand_2.C.t1 D_FlipFlop_7.3-input-nand_2.Vout.t7 a_n8818_48405# GND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1451 a_28044_52049# D_FlipFlop_3.nPRE.t17 And_Gate_4.A GND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1452 a_16854_48405# FFCLR.t53 GND.t698 GND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1453 GND.t562 VDD.t968 a_13751_59439# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1454 CDAC_v3_0.switch_3.Z.t0 a_19654_45397# VDD.t97 VDD.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1455 a_2209_55365# Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_2209_54751# GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1456 VDD.t830 CLK.t111 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t0 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1457 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t16 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1458 a_17315_56723# Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1459 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t15 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1460 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t7 VDD.t355 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1461 VDD.t733 D_FlipFlop_4.nPRE.t16 And_Gate_2.A VDD.t732 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1462 VDD.t119 VDD.t118 Ring_Counter_0.D_FlipFlop_7.Qbar VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1463 a_30721_59439# Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout a_30721_58825# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1464 VDD.t605 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.3-input-nand_2.C.t2 VDD.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1465 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t603 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1466 a_2046_51119# D_FlipFlop_6.3-input-nand_2.Vout.t6 GND.t98 GND.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1467 D_FlipFlop_0.3-input-nand_0.Vout EN.t87 VDD.t656 VDD.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1468 a_12901_56723# Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1469 a_6734_51119# D_FlipFlop_7.D.t31 a_6120_51119# GND.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1470 CDAC_v3_0.switch_4.Z.t2 a_23598_45397# VDD.t403 VDD.t402 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1471 a_31571_61411# Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B a_31571_60797# GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1472 a_28007_61411# Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B a_28007_60797# GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1473 GND.t563 VDD.t969 a_9337_61411# GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1474 VDD.t218 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1475 a_n1355_60797# CLK.t112 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1476 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t8 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1477 GND.t382 GND.t383 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1478 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.CLK.t5 VDD.t863 VDD.t862 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1479 Ring_Counter_0.D_FlipFlop_16.Q.t0 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t413 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1480 a_50454_10637.t2 a_50454_10637.t1 Vbias.t3 Vbias.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X1481 And_Gate_2.A Nand_Gate_2.A.t10 VDD.t32 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1482 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B VDD.t874 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1483 D_FlipFlop_3.3-input-nand_1.B D_FlipFlop_7.D.t32 GND.t109 GND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1484 VDD.t455 D_FlipFlop_5.nPRE.t15 And_Gate_3.A VDD.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1485 GND.t571 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 a_23593_56723# GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1486 a_16465_58825# Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1487 CDAC_v3_0.OUT CDAC_v3_0.switch_3.Z.t2 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1488 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t14 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1489 VDD.t728 a_50454_10637.t0 Vbias.t4 sky130_fd_pr__res_xhigh_po_5p73 l=150
X1490 D_FlipFlop_1.CLK.t1 And_Gate_6.Nand_Gate_0.Vout GND.t573 GND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1491 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout Nand_Gate_7.A.t11 VDD.t329 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1492 GND.t564 VDD.t970 a_38699_59439# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1493 VDD.t786 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1494 VDD.t655 EN.t88 D_FlipFlop_6.nPRE.t3 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1495 a_35430_45397# Q7.t9 VDD.t510 VDD.t509 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1496 VDD.t654 EN.t89 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t0 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1497 a_37849_56723# Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1498 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t6 VDD.t761 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1499 Q0.t0 D_FlipFlop_7.Qbar VDD.t426 VDD.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1500 GND.t713 EN.t90 a_n4919_55365# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1501 VDD.t117 VDD.t115 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t1 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1502 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD.t777 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1503 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t13 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1504 VDD.t462 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1505 CDAC_v3_0.OUT CDAC_v3_0.switch_4.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1506 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B VDD.t290 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1507 VDD.t63 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.3-input-nand_2.Vout.t0 VDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1508 a_45856_48405# D_FlipFlop_1.3-input-nand_2.C.t7 GND.t113 GND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1509 VDD.t723 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t3 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1510 VDD.t513 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t1 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1511 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout Nand_Gate_4.A.t10 VDD.t23 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1512 GND.t714 EN.t91 a_27157_55365# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1513 VDD.t114 VDD.t113 Ring_Counter_0.D_FlipFlop_13.Qbar VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1514 D_FlipFlop_2.CLK.t0 And_Gate_5.Nand_Gate_0.Vout VDD.t646 VDD.t645 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1515 GND.t631 EN.t92 a_49391_55365# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1516 D_FlipFlop_0.3-input-nand_1.Vout FFCLR.t54 VDD.t475 VDD.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1517 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t12 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1518 a_10187_56723# Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1519 VDD.t831 CLK.t113 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t0 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1520 VDD.t653 EN.t93 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1521 Ring_Counter_0.D_FlipFlop_15.Qbar.t3 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 VDD.t481 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1522 a_20029_59439# Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout a_20029_58825# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1523 D_FlipFlop_4.3-input-nand_1.B D_FlipFlop_7.D.t33 VDD.t276 VDD.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1524 VDD.t112 VDD.t110 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1525 a_6623_61411# Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B a_6623_60797# GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1526 GND.t380 GND.t381 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1527 VDD.t507 D_FlipFlop_7.Nand_Gate_0.Vout Q0.t2 VDD.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1528 a_42263_59439# Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 a_42263_58825# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1529 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.CLK.t6 VDD.t864 VDD.t862 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1530 D_FlipFlop_7.3-input-nand_2.Vout.t1 D_FlipFlop_7.nPRE.t15 VDD.t409 VDD.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1531 a_n7633_55365# Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 a_n7633_54751# GND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1532 GND.t586 VDD.t971 a_17315_59439# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1533 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t7 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1534 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t6 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1535 VDD.t734 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1536 a_24443_56723# Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1537 VDD.t61 Nand_Gate_6.A.t11 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1538 a_51902_51119# FFCLR.t55 GND.t274 GND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1539 a_12780_51119# D_FlipFlop_4.Nand_Gate_0.Vout a_12166_51119# GND.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1540 VDD.t109 VDD.t108 Ring_Counter_0.D_FlipFlop_5.Qbar.t3 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1541 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t11 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1542 a_56590_51119# D_FlipFlop_0.Nand_Gate_0.Vout a_55976_51119# GND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1543 a_17468_51119# D_FlipFlop_5.3-input-nand_0.Vout a_16854_51119# GND.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1544 GND.t378 GND.t379 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1545 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1546 GND.t632 EN.t94 a_12901_59439# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1547 a_14529_52049# And_Gate_3.A GND.t681 GND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1548 VDD.t34 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1549 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t10 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1550 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t9 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1551 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.CLK.t7 GND.t658 GND.t657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1552 VDD.t652 EN.t95 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1553 VDD.t832 CLK.t114 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1554 a_35135_61411# Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B a_35135_60797# GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1555 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t8 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1556 GND.t96 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 a_n4919_56723# GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1557 VDD.t107 VDD.t105 Ring_Counter_0.D_FlipFlop_1.Qbar VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1558 GND.t638 EN.t96 a_13751_61411# GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1559 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t7 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1560 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t7 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1561 D_FlipFlop_6.3-input-nand_2.C.t1 D_FlipFlop_6.3-input-nand_2.Vout.t7 a_n56_48405# GND.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1562 D_FlipFlop_7.Qbar Q0.t8 VDD.t772 VDD.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1563 a_55976_51119# FFCLR.t56 GND.t276 GND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1564 VDD.t558 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.3-input-nand_2.C.t2 VDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1565 a_30721_61411# Nand_Gate_4.A.t11 a_30721_60797# GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1566 Q3.t0 D_FlipFlop_5.Qbar VDD.t71 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1567 GND.t31 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 a_27157_56723# GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1568 a_23593_58825# Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1569 GND.t376 GND.t377 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1570 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t6 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1571 Q7.t1 D_FlipFlop_0.Qbar a_56590_51119# GND.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1572 D_FlipFlop_5.3-input-nand_2.Vout.t0 D_FlipFlop_5.3-input-nand_2.C.t7 a_17468_51119# GND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1573 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.CLK.t6 a_n2028_48405# GND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1574 And_Gate_3.Nand_Gate_0.Vout CLK.t115 a_14529_52049# GND.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1575 GND.t644 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t7 a_49391_56723# GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1576 VDD.t769 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1577 GND.t633 EN.t97 a_5773_55365# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1578 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t7 VDD.t781 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1579 a_3059_59439# Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 a_3059_58825# GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1580 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1581 GND.t374 GND.t375 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1582 CDAC_v3_0.OUT CDAC_v3_0.switch_5.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1583 a_52105_55365# Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t4 a_52105_54751# GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1584 GND.t627 EN.t98 a_37849_59439# GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1585 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1586 VDD.t578 D_FlipFlop_7.Nand_Gate_1.Vout D_FlipFlop_7.Qbar VDD.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1587 a_44977_56723# Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1588 GND.t204 D_FlipFlop_7.nPRE.t16 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1589 a_3404_51119# D_FlipFlop_6.nPRE.t17 GND.t285 GND.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1590 GND.t614 Q3.t7 CDAC_v3_0.switch_3.Z.t11 VDD.t790 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1591 VDD.t651 EN.t99 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 VDD.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1592 D_FlipFlop_7.3-input-nand_2.C.t3 FFCLR.t57 VDD.t476 VDD.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1593 a_16465_60797# CLK.t116 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1594 GND.t372 GND.t373 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1595 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B VDD.t709 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1596 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t6 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1597 GND.t221 Q5.t9 CDAC_v3_0.switch_5.Z.t1 VDD.t427 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1598 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t5 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1599 a_45827_55365# Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 a_45827_54751# GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1600 GND.t628 EN.t100 a_38699_61411# GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1601 VDD.t36 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t2 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1602 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout Nand_Gate_5.A.t11 VDD.t263 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1603 GND.t370 GND.t371 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1604 VDD.t833 CLK.t117 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1605 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.CLK.t7 GND.t35 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1606 GND.t621 EN.t101 a_34285_55365# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1607 a_n505_54751# D_FlipFlop_7.nPRE.t17 Ring_Counter_0.D_FlipFlop_14.Qbar.t2 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1608 a_41782_51119# D_FlipFlop_7.D.t34 a_41168_51119# GND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1609 VDD.t104 VDD.t103 Ring_Counter_0.D_FlipFlop_12.Qbar VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1610 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t4 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1611 GND.t587 VDD.t972 a_10187_59439# GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1612 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Inverter_1.Vout a_45856_51119# GND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1613 VDD.t650 EN.t102 D_FlipFlop_1.nPRE.t2 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1614 a_10520_52049# D_FlipFlop_4.nPRE.t17 And_Gate_2.A GND.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1615 Vbias.t8 a_50454_10637.t4 D_FlipFlop_7.D.t0 Vbias.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X1616 VDD.t102 VDD.t100 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1617 GND.t686 Q6.t8 CDAC_v3_0.switch_7.Z.t67 VDD.t894 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1618 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t3 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1619 a_19654_45397# Q3.t8 VDD.t299 VDD.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1620 VDD.t649 EN.t103 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 VDD.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1621 CDAC_v3_0.OUT CDAC_v3_0.switch_7.Z.t2 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1622 a_8706_51119# D_FlipFlop_4.3-input-nand_0.Vout a_8092_51119# GND.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1623 VDD.t706 Ring_Counter_0.D_FlipFlop_10.Qbar.t5 D_FlipFlop_4.nPRE.t3 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1624 D_FlipFlop_6.CLK.t0 And_Gate_1.Nand_Gate_0.Vout VDD.t586 VDD.t585 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1625 GND.t620 EN.t104 a_48541_55365# GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1626 GND.t588 VDD.t973 a_24443_59439# GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1627 VDD.t648 EN.t105 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1628 D_FlipFlop_5.Qbar Q3.t9 VDD.t300 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1629 a_23644_51119# FFCLR.t58 GND.t278 GND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1630 a_20879_59439# Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 a_20879_58825# GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1631 a_31571_56723# Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1632 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.CLK.t7 VDD.t784 VDD.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1633 a_28007_56723# Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 GND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1634 VDD.t456 D_FlipFlop_5.nPRE.t16 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1635 a_28332_51119# D_FlipFlop_3.3-input-nand_2.Vout.t7 GND.t363 GND.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1636 VDD.t99 VDD.t98 Ring_Counter_0.D_FlipFlop_4.Qbar.t2 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1637 GND.t10 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 a_5773_56723# GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1638 a_41413_59439# Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout a_41413_58825# GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1639 VDD.t795 D_FlipFlop_2.nPRE.t17 And_Gate_5.A VDD.t794 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1640 VDD.t647 EN.t106 D_FlipFlop_3.nPRE.t1 VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1641 GND.t27 Nand_Gate_2.A.t11 a_10520_52049# GND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1642 Nand_Gate_1.A.t3 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t799 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1643 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t5 VDD.t362 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1644 VDD.t861 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1645 a_20029_61411# D_FlipFlop_5.nPRE.t17 a_20029_60797# GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1646 a_7822_45397# Q0.t9 GND.t87 GND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1647 a_31486_45397# Q6.t9 VDD.t896 VDD.t895 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1648 CDAC_v3_0.OUT CDAC_v3_0.switch_6.Z.t3 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1649 a_6120_51119# FFCLR.t59 GND.t280 GND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1650 a_42263_61411# Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B a_42263_60797# GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1651 a_n4919_58825# Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1652 GND.t567 EN.t107 a_17315_61411# GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1653 VDD.t278 D_FlipFlop_7.D.t35 D_FlipFlop_2.3-input-nand_0.Vout VDD.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1654 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.CLK.t7 VDD.t344 VDD.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1655 GND.t368 GND.t369 sky130_fd_pr__cap_mim_m3_1 l=6.88 w=6.88
X1656 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Inverter_1.Vout a_28332_51119# GND.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1657 GND.t272 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 a_34285_56723# GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1658 a_27157_58825# Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1659 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Inverter_1.Vout VDD.t530 VDD.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1660 GND.t589 VDD.t974 a_12901_61411# GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1661 VDD.t15 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t0 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
R0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t2 169.46
R1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t1 167.809
R2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t3 167.809
R3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t5 167.227
R4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n0 151.594
R5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t7 150.273
R6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t6 74.8641
R7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t4 73.6304
R8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t0 61.84
R9 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 12.3891
R10 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n2 11.4489
R11 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n8 0.38637
R12 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n1 0.280391
R13 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n3 0.200143
R14 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.152844
R15 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.149957
R16 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n4 0.149957
R17 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.063
R18 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.063
R19 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n7 0.063
R20 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n5 0.063
R21 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.0454219
R22 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t0 169.46
R23 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t3 167.809
R24 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t1 167.809
R25 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t5 167.226
R26 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n6 150.273
R27 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t4 150.273
R28 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t6 74.951
R29 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t7 73.6304
R30 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t2 60.3943
R31 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n4 12.3891
R32 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n8 11.4489
R33 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n10 1.68257
R34 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n0 1.44615
R35 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n2 1.2342
R36 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 1.08448
R37 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.932141
R38 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n9 0.3496
R39 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n7 0.280391
R40 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.063
R41 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.063
R42 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n3 0.063
R43 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.063
R44 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n5 0.063
R45 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n1 0.063
R46 GND.n2100 GND.n2099 73717.4
R47 GND.n721 GND.n720 61368.3
R48 GND.n4363 GND.n4362 29655.4
R49 GND.n1087 GND.n1086 28217.6
R50 GND.n3998 GND.n49 22149.2
R51 GND.n1520 GND.n1519 18700
R52 GND.n3997 GND.n3996 17786.4
R53 GND.n2946 GND.n357 17283.1
R54 GND.n2393 GND.n526 16860.5
R55 GND.n2947 GND.n486 16437.9
R56 GND.n2297 GND.n599 15443.5
R57 GND.n2296 GND.n2295 14598.3
R58 GND.n4288 GND.n4287 13725.7
R59 GND.n1303 GND.n773 13604
R60 GND.n1521 GND.n823 13224.9
R61 GND.n1173 GND.n1172 12758.8
R62 GND.n2393 GND.n2392 12678
R63 GND.n2523 GND.n533 11385.3
R64 GND.n1303 GND.n802 11310.7
R65 GND.n1519 GND.n802 10838.4
R66 GND.n3995 GND.n94 9624.05
R67 GND.n2392 GND.n599 9471.19
R68 GND.n3333 GND.n3332 9120.66
R69 GND.n1173 GND.n773 8545.2
R70 GND.n3333 GND.n357 7631.64
R71 GND.n4362 GND.n10 7473.67
R72 GND.n3996 GND.n3995 7128.25
R73 GND.n4286 GND.n54 6971.5
R74 GND.n4236 GND.n54 6971.5
R75 GND.n4286 GND.n55 6971.5
R76 GND.n4236 GND.n55 6971.5
R77 GND.n4232 GND.n50 6971.5
R78 GND.n4276 GND.n4232 6971.5
R79 GND.n4235 GND.n50 6971.5
R80 GND.n4276 GND.n4235 6971.5
R81 GND.n4317 GND.n27 6971.5
R82 GND.n4321 GND.n27 6971.5
R83 GND.n4317 GND.n28 6971.5
R84 GND.n4321 GND.n28 6971.5
R85 GND.n4290 GND.n44 6971.5
R86 GND.n4294 GND.n44 6971.5
R87 GND.n4290 GND.n45 6971.5
R88 GND.n4294 GND.n45 6971.5
R89 GND.n4050 GND.n64 6971.5
R90 GND.n4064 GND.n64 6971.5
R91 GND.n4050 GND.n65 6971.5
R92 GND.n4064 GND.n65 6971.5
R93 GND.n4069 GND.n4045 6971.5
R94 GND.n4069 GND.n4046 6971.5
R95 GND.n4045 GND.n4044 6971.5
R96 GND.n4046 GND.n4044 6971.5
R97 GND.n4082 GND.n72 6971.5
R98 GND.n4082 GND.n73 6971.5
R99 GND.n72 GND.n71 6971.5
R100 GND.n73 GND.n71 6971.5
R101 GND.n86 GND.n83 6971.5
R102 GND.n91 GND.n83 6971.5
R103 GND.n87 GND.n86 6971.5
R104 GND.n91 GND.n87 6971.5
R105 GND.n4020 GND.n67 6971.5
R106 GND.n4022 GND.n67 6971.5
R107 GND.n4020 GND.n68 6971.5
R108 GND.n4022 GND.n68 6971.5
R109 GND.n4026 GND.n89 6971.5
R110 GND.n4032 GND.n89 6971.5
R111 GND.n4026 GND.n90 6971.5
R112 GND.n4032 GND.n90 6971.5
R113 GND.n3975 GND.n129 6971.5
R114 GND.n3975 GND.n3974 6971.5
R115 GND.n130 GND.n129 6971.5
R116 GND.n3974 GND.n130 6971.5
R117 GND.n3994 GND.n96 6971.5
R118 GND.n3994 GND.n97 6971.5
R119 GND.n96 GND.n95 6971.5
R120 GND.n97 GND.n95 6971.5
R121 GND.n3309 GND.n386 6971.5
R122 GND.n3309 GND.n3308 6971.5
R123 GND.n3307 GND.n386 6971.5
R124 GND.n3308 GND.n3307 6971.5
R125 GND.n3331 GND.n362 6971.5
R126 GND.n384 GND.n362 6971.5
R127 GND.n3331 GND.n363 6971.5
R128 GND.n384 GND.n363 6971.5
R129 GND.n3320 GND.n372 6971.5
R130 GND.n373 GND.n372 6971.5
R131 GND.n3320 GND.n383 6971.5
R132 GND.n383 GND.n373 6971.5
R133 GND.n374 GND.n358 6971.5
R134 GND.n374 GND.n370 6971.5
R135 GND.n377 GND.n358 6971.5
R136 GND.n377 GND.n370 6971.5
R137 GND.n445 GND.n388 6971.5
R138 GND.n437 GND.n388 6971.5
R139 GND.n445 GND.n389 6971.5
R140 GND.n437 GND.n389 6971.5
R141 GND.n432 GND.n360 6971.5
R142 GND.n443 GND.n432 6971.5
R143 GND.n442 GND.n360 6971.5
R144 GND.n443 GND.n442 6971.5
R145 GND.n3128 GND.n3049 6971.5
R146 GND.n3142 GND.n3049 6971.5
R147 GND.n3128 GND.n3050 6971.5
R148 GND.n3142 GND.n3050 6971.5
R149 GND.n3147 GND.n3123 6971.5
R150 GND.n3147 GND.n3124 6971.5
R151 GND.n3123 GND.n3122 6971.5
R152 GND.n3124 GND.n3122 6971.5
R153 GND.n3160 GND.n3057 6971.5
R154 GND.n3160 GND.n3058 6971.5
R155 GND.n3057 GND.n3056 6971.5
R156 GND.n3058 GND.n3056 6971.5
R157 GND.n3071 GND.n3068 6971.5
R158 GND.n3076 GND.n3068 6971.5
R159 GND.n3072 GND.n3071 6971.5
R160 GND.n3076 GND.n3072 6971.5
R161 GND.n3098 GND.n3052 6971.5
R162 GND.n3100 GND.n3052 6971.5
R163 GND.n3098 GND.n3053 6971.5
R164 GND.n3100 GND.n3053 6971.5
R165 GND.n3104 GND.n3074 6971.5
R166 GND.n3110 GND.n3074 6971.5
R167 GND.n3104 GND.n3075 6971.5
R168 GND.n3110 GND.n3075 6971.5
R169 GND.n3335 GND.n352 6971.5
R170 GND.n3339 GND.n352 6971.5
R171 GND.n3335 GND.n353 6971.5
R172 GND.n3339 GND.n353 6971.5
R173 GND.n2945 GND.n488 6971.5
R174 GND.n2945 GND.n489 6971.5
R175 GND.n488 GND.n487 6971.5
R176 GND.n489 GND.n487 6971.5
R177 GND.n2802 GND.n553 6971.5
R178 GND.n2802 GND.n554 6971.5
R179 GND.n2801 GND.n553 6971.5
R180 GND.n2801 GND.n554 6971.5
R181 GND.n2575 GND.n2495 6971.5
R182 GND.n2589 GND.n2495 6971.5
R183 GND.n2575 GND.n2496 6971.5
R184 GND.n2589 GND.n2496 6971.5
R185 GND.n2594 GND.n2570 6971.5
R186 GND.n2594 GND.n2571 6971.5
R187 GND.n2570 GND.n2569 6971.5
R188 GND.n2571 GND.n2569 6971.5
R189 GND.n2607 GND.n2503 6971.5
R190 GND.n2607 GND.n2504 6971.5
R191 GND.n2503 GND.n2502 6971.5
R192 GND.n2504 GND.n2502 6971.5
R193 GND.n2517 GND.n2514 6971.5
R194 GND.n2522 GND.n2514 6971.5
R195 GND.n2518 GND.n2517 6971.5
R196 GND.n2522 GND.n2518 6971.5
R197 GND.n2545 GND.n2498 6971.5
R198 GND.n2547 GND.n2498 6971.5
R199 GND.n2545 GND.n2499 6971.5
R200 GND.n2547 GND.n2499 6971.5
R201 GND.n2551 GND.n2520 6971.5
R202 GND.n2557 GND.n2520 6971.5
R203 GND.n2551 GND.n2521 6971.5
R204 GND.n2557 GND.n2521 6971.5
R205 GND.n2822 GND.n524 6971.5
R206 GND.n2822 GND.n525 6971.5
R207 GND.n2821 GND.n524 6971.5
R208 GND.n2821 GND.n525 6971.5
R209 GND.n2383 GND.n2335 6971.5
R210 GND.n2383 GND.n2336 6971.5
R211 GND.n2382 GND.n2336 6971.5
R212 GND.n2382 GND.n2335 6971.5
R213 GND.n2391 GND.n601 6971.5
R214 GND.n2391 GND.n602 6971.5
R215 GND.n601 GND.n600 6971.5
R216 GND.n602 GND.n600 6971.5
R217 GND.n1830 GND.n1752 6971.5
R218 GND.n1844 GND.n1752 6971.5
R219 GND.n1830 GND.n1753 6971.5
R220 GND.n1844 GND.n1753 6971.5
R221 GND.n1849 GND.n1825 6971.5
R222 GND.n1849 GND.n1826 6971.5
R223 GND.n1825 GND.n1824 6971.5
R224 GND.n1826 GND.n1824 6971.5
R225 GND.n1862 GND.n1760 6971.5
R226 GND.n1862 GND.n1761 6971.5
R227 GND.n1760 GND.n1759 6971.5
R228 GND.n1761 GND.n1759 6971.5
R229 GND.n1774 GND.n1771 6971.5
R230 GND.n1775 GND.n1771 6971.5
R231 GND.n1776 GND.n1774 6971.5
R232 GND.n1776 GND.n1775 6971.5
R233 GND.n1800 GND.n1755 6971.5
R234 GND.n1802 GND.n1755 6971.5
R235 GND.n1800 GND.n1756 6971.5
R236 GND.n1802 GND.n1756 6971.5
R237 GND.n1806 GND.n1778 6971.5
R238 GND.n1812 GND.n1778 6971.5
R239 GND.n1806 GND.n1779 6971.5
R240 GND.n1812 GND.n1779 6971.5
R241 GND.n621 GND.n620 6971.5
R242 GND.n2299 GND.n620 6971.5
R243 GND.n2298 GND.n621 6971.5
R244 GND.n2299 GND.n2298 6971.5
R245 GND.n2286 GND.n633 6971.5
R246 GND.n2286 GND.n634 6971.5
R247 GND.n2285 GND.n634 6971.5
R248 GND.n2285 GND.n633 6971.5
R249 GND.n1999 GND.n883 6971.5
R250 GND.n1999 GND.n884 6971.5
R251 GND.n1998 GND.n883 6971.5
R252 GND.n1998 GND.n884 6971.5
R253 GND.n1573 GND.n900 6971.5
R254 GND.n1587 GND.n900 6971.5
R255 GND.n1573 GND.n901 6971.5
R256 GND.n1587 GND.n901 6971.5
R257 GND.n1592 GND.n1568 6971.5
R258 GND.n1592 GND.n1569 6971.5
R259 GND.n1568 GND.n1567 6971.5
R260 GND.n1569 GND.n1567 6971.5
R261 GND.n1605 GND.n908 6971.5
R262 GND.n1605 GND.n909 6971.5
R263 GND.n908 GND.n907 6971.5
R264 GND.n909 GND.n907 6971.5
R265 GND.n922 GND.n919 6971.5
R266 GND.n927 GND.n919 6971.5
R267 GND.n923 GND.n922 6971.5
R268 GND.n927 GND.n923 6971.5
R269 GND.n1543 GND.n903 6971.5
R270 GND.n1545 GND.n903 6971.5
R271 GND.n1543 GND.n904 6971.5
R272 GND.n1545 GND.n904 6971.5
R273 GND.n1549 GND.n925 6971.5
R274 GND.n1555 GND.n925 6971.5
R275 GND.n1549 GND.n926 6971.5
R276 GND.n1555 GND.n926 6971.5
R277 GND.n2020 GND.n813 6971.5
R278 GND.n2016 GND.n813 6971.5
R279 GND.n2020 GND.n814 6971.5
R280 GND.n2016 GND.n814 6971.5
R281 GND.n2034 GND.n804 6971.5
R282 GND.n2030 GND.n804 6971.5
R283 GND.n2030 GND.n805 6971.5
R284 GND.n2034 GND.n805 6971.5
R285 GND.n2040 GND.n800 6971.5
R286 GND.n2040 GND.n801 6971.5
R287 GND.n2039 GND.n800 6971.5
R288 GND.n2039 GND.n801 6971.5
R289 GND.n1225 GND.n943 6971.5
R290 GND.n1239 GND.n943 6971.5
R291 GND.n1225 GND.n944 6971.5
R292 GND.n1239 GND.n944 6971.5
R293 GND.n1244 GND.n1220 6971.5
R294 GND.n1244 GND.n1221 6971.5
R295 GND.n1220 GND.n1219 6971.5
R296 GND.n1221 GND.n1219 6971.5
R297 GND.n1257 GND.n951 6971.5
R298 GND.n1257 GND.n952 6971.5
R299 GND.n951 GND.n950 6971.5
R300 GND.n952 GND.n950 6971.5
R301 GND.n965 GND.n962 6971.5
R302 GND.n970 GND.n962 6971.5
R303 GND.n966 GND.n965 6971.5
R304 GND.n970 GND.n966 6971.5
R305 GND.n1195 GND.n946 6971.5
R306 GND.n1197 GND.n946 6971.5
R307 GND.n1195 GND.n947 6971.5
R308 GND.n1197 GND.n947 6971.5
R309 GND.n1201 GND.n968 6971.5
R310 GND.n1207 GND.n968 6971.5
R311 GND.n1201 GND.n969 6971.5
R312 GND.n1207 GND.n969 6971.5
R313 GND.n1355 GND.n1275 6971.5
R314 GND.n1369 GND.n1275 6971.5
R315 GND.n1355 GND.n1276 6971.5
R316 GND.n1369 GND.n1276 6971.5
R317 GND.n1374 GND.n1350 6971.5
R318 GND.n1374 GND.n1351 6971.5
R319 GND.n1350 GND.n1349 6971.5
R320 GND.n1351 GND.n1349 6971.5
R321 GND.n1387 GND.n1283 6971.5
R322 GND.n1387 GND.n1284 6971.5
R323 GND.n1283 GND.n1282 6971.5
R324 GND.n1284 GND.n1282 6971.5
R325 GND.n1297 GND.n1294 6971.5
R326 GND.n1302 GND.n1294 6971.5
R327 GND.n1298 GND.n1297 6971.5
R328 GND.n1302 GND.n1298 6971.5
R329 GND.n1325 GND.n1278 6971.5
R330 GND.n1327 GND.n1278 6971.5
R331 GND.n1325 GND.n1279 6971.5
R332 GND.n1327 GND.n1279 6971.5
R333 GND.n1331 GND.n1300 6971.5
R334 GND.n1337 GND.n1300 6971.5
R335 GND.n1331 GND.n1301 6971.5
R336 GND.n1337 GND.n1301 6971.5
R337 GND.n1441 GND.n929 6971.5
R338 GND.n1446 GND.n1441 6971.5
R339 GND.n1442 GND.n929 6971.5
R340 GND.n1446 GND.n1442 6971.5
R341 GND.n1494 GND.n1490 6971.5
R342 GND.n1494 GND.n1408 6971.5
R343 GND.n1490 GND.n1489 6971.5
R344 GND.n1489 GND.n1408 6971.5
R345 GND.n1458 GND.n932 6971.5
R346 GND.n1463 GND.n1458 6971.5
R347 GND.n1459 GND.n932 6971.5
R348 GND.n1463 GND.n1459 6971.5
R349 GND.n1420 GND.n1419 6971.5
R350 GND.n1419 GND.n1412 6971.5
R351 GND.n1424 GND.n1420 6971.5
R352 GND.n1424 GND.n1412 6971.5
R353 GND.n1440 GND.n931 6971.5
R354 GND.n1467 GND.n1440 6971.5
R355 GND.n1468 GND.n931 6971.5
R356 GND.n1468 GND.n1467 6971.5
R357 GND.n1471 GND.n1426 6971.5
R358 GND.n1477 GND.n1426 6971.5
R359 GND.n1471 GND.n1427 6971.5
R360 GND.n1477 GND.n1427 6971.5
R361 GND.n2060 GND.n771 6971.5
R362 GND.n2060 GND.n772 6971.5
R363 GND.n2059 GND.n771 6971.5
R364 GND.n2059 GND.n772 6971.5
R365 GND.n1163 GND.n1125 6971.5
R366 GND.n1163 GND.n1126 6971.5
R367 GND.n1162 GND.n1126 6971.5
R368 GND.n1162 GND.n1125 6971.5
R369 GND.n1111 GND.n979 6971.5
R370 GND.n1111 GND.n980 6971.5
R371 GND.n1116 GND.n979 6971.5
R372 GND.n1116 GND.n980 6971.5
R373 GND.n1017 GND.n1005 6971.5
R374 GND.n1024 GND.n1005 6971.5
R375 GND.n1017 GND.n1006 6971.5
R376 GND.n1024 GND.n1006 6971.5
R377 GND.n1063 GND.n1012 6971.5
R378 GND.n1063 GND.n1013 6971.5
R379 GND.n1012 GND.n1011 6971.5
R380 GND.n1013 GND.n1011 6971.5
R381 GND.n1040 GND.n1008 6971.5
R382 GND.n1035 GND.n1008 6971.5
R383 GND.n1040 GND.n1009 6971.5
R384 GND.n1035 GND.n1009 6971.5
R385 GND.n1088 GND.n996 6971.5
R386 GND.n1092 GND.n996 6971.5
R387 GND.n1088 GND.n997 6971.5
R388 GND.n1092 GND.n997 6971.5
R389 GND.n2098 GND.n683 6971.5
R390 GND.n2098 GND.n684 6971.5
R391 GND.n683 GND.n682 6971.5
R392 GND.n684 GND.n682 6971.5
R393 GND.n3488 GND.n193 6971.5
R394 GND.n3880 GND.n193 6971.5
R395 GND.n3488 GND.n194 6971.5
R396 GND.n3880 GND.n194 6971.5
R397 GND.n3507 GND.n301 6971.5
R398 GND.n3492 GND.n301 6971.5
R399 GND.n3507 GND.n302 6971.5
R400 GND.n3492 GND.n302 6971.5
R401 GND.n3529 GND.n293 6971.5
R402 GND.n3511 GND.n293 6971.5
R403 GND.n3529 GND.n294 6971.5
R404 GND.n3511 GND.n294 6971.5
R405 GND.n3551 GND.n285 6971.5
R406 GND.n3533 GND.n285 6971.5
R407 GND.n3551 GND.n286 6971.5
R408 GND.n3533 GND.n286 6971.5
R409 GND.n3570 GND.n277 6971.5
R410 GND.n3555 GND.n277 6971.5
R411 GND.n3570 GND.n278 6971.5
R412 GND.n3555 GND.n278 6971.5
R413 GND.n3590 GND.n269 6971.5
R414 GND.n3574 GND.n269 6971.5
R415 GND.n3590 GND.n270 6971.5
R416 GND.n3574 GND.n270 6971.5
R417 GND.n3609 GND.n251 6971.5
R418 GND.n3594 GND.n251 6971.5
R419 GND.n3609 GND.n252 6971.5
R420 GND.n3594 GND.n252 6971.5
R421 GND.n3615 GND.n248 6971.5
R422 GND.n3615 GND.n249 6971.5
R423 GND.n3616 GND.n248 6971.5
R424 GND.n3616 GND.n249 6971.5
R425 GND.n3921 GND.n8 6971.5
R426 GND.n4364 GND.n8 6971.5
R427 GND.n3921 GND.n9 6971.5
R428 GND.n4364 GND.n9 6971.5
R429 GND.n3926 GND.n3911 6971.5
R430 GND.n3926 GND.n3912 6971.5
R431 GND.n3927 GND.n3911 6971.5
R432 GND.n3927 GND.n3912 6971.5
R433 GND.n3950 GND.n186 6971.5
R434 GND.n3950 GND.n187 6971.5
R435 GND.n3951 GND.n186 6971.5
R436 GND.n3951 GND.n187 6971.5
R437 GND.n3884 GND.n188 6971.5
R438 GND.n3893 GND.n188 6971.5
R439 GND.n3884 GND.n189 6971.5
R440 GND.n3893 GND.n189 6971.5
R441 GND.n3406 GND.n3399 6971.5
R442 GND.n3406 GND.n3400 6971.5
R443 GND.n3407 GND.n3399 6971.5
R444 GND.n3407 GND.n3400 6971.5
R445 GND.n3436 GND.n330 6971.5
R446 GND.n3428 GND.n330 6971.5
R447 GND.n3436 GND.n331 6971.5
R448 GND.n3428 GND.n331 6971.5
R449 GND.n3447 GND.n325 6971.5
R450 GND.n3439 GND.n325 6971.5
R451 GND.n3447 GND.n326 6971.5
R452 GND.n3439 GND.n326 6971.5
R453 GND.n4326 GND.n21 6971.5
R454 GND.n4343 GND.n21 6971.5
R455 GND.n4326 GND.n22 6971.5
R456 GND.n4343 GND.n22 6971.5
R457 GND.n3967 GND.n134 6971.5
R458 GND.n3967 GND.n135 6971.5
R459 GND.n3971 GND.n135 6971.5
R460 GND.n3971 GND.n134 6971.5
R461 GND.n3361 GND.n346 6971.5
R462 GND.n3361 GND.n347 6971.5
R463 GND.n3344 GND.n347 6971.5
R464 GND.n3344 GND.n346 6971.5
R465 GND.n2791 GND.n2739 6971.5
R466 GND.n2791 GND.n2740 6971.5
R467 GND.n2795 GND.n2740 6971.5
R468 GND.n2795 GND.n2739 6971.5
R469 GND.n719 GND.n714 6971.5
R470 GND.n719 GND.n717 6971.5
R471 GND.n714 GND.n704 6971.5
R472 GND.n717 GND.n704 6971.5
R473 GND.n722 GND.n710 6971.5
R474 GND.n723 GND.n722 6971.5
R475 GND.n710 GND.n708 6971.5
R476 GND.n723 GND.n708 6971.5
R477 GND.n2128 GND.n666 6971.5
R478 GND.n2137 GND.n666 6971.5
R479 GND.n2128 GND.n667 6971.5
R480 GND.n2137 GND.n667 6971.5
R481 GND.n2116 GND.n671 6971.5
R482 GND.n2125 GND.n671 6971.5
R483 GND.n2116 GND.n672 6971.5
R484 GND.n2125 GND.n672 6971.5
R485 GND.n2104 GND.n675 6971.5
R486 GND.n2113 GND.n675 6971.5
R487 GND.n2104 GND.n676 6971.5
R488 GND.n2113 GND.n676 6971.5
R489 GND.n762 GND.n728 6971.5
R490 GND.n762 GND.n729 6971.5
R491 GND.n763 GND.n728 6971.5
R492 GND.n763 GND.n729 6971.5
R493 GND.n3458 GND.n320 6971.5
R494 GND.n3450 GND.n320 6971.5
R495 GND.n3458 GND.n321 6971.5
R496 GND.n3450 GND.n321 6971.5
R497 GND.n2892 GND.n497 6971.5
R498 GND.n2892 GND.n498 6971.5
R499 GND.n2893 GND.n497 6971.5
R500 GND.n2893 GND.n498 6971.5
R501 GND.n2872 GND.n499 6971.5
R502 GND.n2881 GND.n499 6971.5
R503 GND.n2872 GND.n500 6971.5
R504 GND.n2881 GND.n500 6971.5
R505 GND.n2860 GND.n503 6971.5
R506 GND.n2869 GND.n503 6971.5
R507 GND.n2860 GND.n504 6971.5
R508 GND.n2869 GND.n504 6971.5
R509 GND.n2829 GND.n516 6971.5
R510 GND.n2838 GND.n516 6971.5
R511 GND.n2829 GND.n517 6971.5
R512 GND.n2838 GND.n517 6971.5
R513 GND.n2221 GND.n2205 6971.5
R514 GND.n2213 GND.n2205 6971.5
R515 GND.n2221 GND.n2206 6971.5
R516 GND.n2213 GND.n2206 6971.5
R517 GND.n2226 GND.n2203 6971.5
R518 GND.n2226 GND.n2204 6971.5
R519 GND.n2227 GND.n2203 6971.5
R520 GND.n2227 GND.n2204 6971.5
R521 GND.n2250 GND.n2183 6971.5
R522 GND.n2250 GND.n2184 6971.5
R523 GND.n2251 GND.n2183 6971.5
R524 GND.n2251 GND.n2184 6971.5
R525 GND.n2171 GND.n649 6971.5
R526 GND.n2180 GND.n649 6971.5
R527 GND.n2171 GND.n650 6971.5
R528 GND.n2180 GND.n650 6971.5
R529 GND.n2159 GND.n653 6971.5
R530 GND.n2168 GND.n653 6971.5
R531 GND.n2159 GND.n654 6971.5
R532 GND.n2168 GND.n654 6971.5
R533 GND.n1915 GND.n886 6971.5
R534 GND.n1920 GND.n1915 6971.5
R535 GND.n1916 GND.n886 6971.5
R536 GND.n1920 GND.n1916 6971.5
R537 GND.n1968 GND.n1964 6971.5
R538 GND.n1968 GND.n1882 6971.5
R539 GND.n1964 GND.n1963 6971.5
R540 GND.n1963 GND.n1882 6971.5
R541 GND.n1932 GND.n889 6971.5
R542 GND.n1937 GND.n1932 6971.5
R543 GND.n1933 GND.n889 6971.5
R544 GND.n1937 GND.n1933 6971.5
R545 GND.n1894 GND.n1893 6971.5
R546 GND.n1893 GND.n1886 6971.5
R547 GND.n1898 GND.n1894 6971.5
R548 GND.n1898 GND.n1886 6971.5
R549 GND.n1914 GND.n888 6971.5
R550 GND.n1941 GND.n1914 6971.5
R551 GND.n1942 GND.n888 6971.5
R552 GND.n1942 GND.n1941 6971.5
R553 GND.n1945 GND.n1900 6971.5
R554 GND.n1951 GND.n1900 6971.5
R555 GND.n1945 GND.n1901 6971.5
R556 GND.n1951 GND.n1901 6971.5
R557 GND.n1703 GND.n1624 6971.5
R558 GND.n1717 GND.n1624 6971.5
R559 GND.n1703 GND.n1625 6971.5
R560 GND.n1717 GND.n1625 6971.5
R561 GND.n1722 GND.n1698 6971.5
R562 GND.n1722 GND.n1699 6971.5
R563 GND.n1698 GND.n1697 6971.5
R564 GND.n1699 GND.n1697 6971.5
R565 GND.n1735 GND.n1632 6971.5
R566 GND.n1735 GND.n1633 6971.5
R567 GND.n1632 GND.n1631 6971.5
R568 GND.n1633 GND.n1631 6971.5
R569 GND.n1646 GND.n1643 6971.5
R570 GND.n1651 GND.n1643 6971.5
R571 GND.n1647 GND.n1646 6971.5
R572 GND.n1651 GND.n1647 6971.5
R573 GND.n1673 GND.n1627 6971.5
R574 GND.n1675 GND.n1627 6971.5
R575 GND.n1673 GND.n1628 6971.5
R576 GND.n1675 GND.n1628 6971.5
R577 GND.n1679 GND.n1649 6971.5
R578 GND.n1685 GND.n1649 6971.5
R579 GND.n1679 GND.n1650 6971.5
R580 GND.n1685 GND.n1650 6971.5
R581 GND.n2445 GND.n571 6971.5
R582 GND.n2459 GND.n571 6971.5
R583 GND.n2445 GND.n572 6971.5
R584 GND.n2459 GND.n572 6971.5
R585 GND.n2464 GND.n2440 6971.5
R586 GND.n2464 GND.n2441 6971.5
R587 GND.n2440 GND.n2439 6971.5
R588 GND.n2441 GND.n2439 6971.5
R589 GND.n2477 GND.n579 6971.5
R590 GND.n2477 GND.n580 6971.5
R591 GND.n579 GND.n578 6971.5
R592 GND.n580 GND.n578 6971.5
R593 GND.n593 GND.n590 6971.5
R594 GND.n598 GND.n590 6971.5
R595 GND.n594 GND.n593 6971.5
R596 GND.n598 GND.n594 6971.5
R597 GND.n2415 GND.n574 6971.5
R598 GND.n2417 GND.n574 6971.5
R599 GND.n2415 GND.n575 6971.5
R600 GND.n2417 GND.n575 6971.5
R601 GND.n2421 GND.n596 6971.5
R602 GND.n2427 GND.n596 6971.5
R603 GND.n2421 GND.n597 6971.5
R604 GND.n2427 GND.n597 6971.5
R605 GND.n2661 GND.n557 6971.5
R606 GND.n2666 GND.n2661 6971.5
R607 GND.n2662 GND.n557 6971.5
R608 GND.n2666 GND.n2662 6971.5
R609 GND.n2714 GND.n2710 6971.5
R610 GND.n2714 GND.n2628 6971.5
R611 GND.n2710 GND.n2709 6971.5
R612 GND.n2709 GND.n2628 6971.5
R613 GND.n2678 GND.n560 6971.5
R614 GND.n2683 GND.n2678 6971.5
R615 GND.n2679 GND.n560 6971.5
R616 GND.n2683 GND.n2679 6971.5
R617 GND.n2640 GND.n2639 6971.5
R618 GND.n2639 GND.n2632 6971.5
R619 GND.n2644 GND.n2640 6971.5
R620 GND.n2644 GND.n2632 6971.5
R621 GND.n2660 GND.n559 6971.5
R622 GND.n2687 GND.n2660 6971.5
R623 GND.n2688 GND.n559 6971.5
R624 GND.n2688 GND.n2687 6971.5
R625 GND.n2691 GND.n2646 6971.5
R626 GND.n2697 GND.n2646 6971.5
R627 GND.n2691 GND.n2647 6971.5
R628 GND.n2697 GND.n2647 6971.5
R629 GND.n2999 GND.n458 6971.5
R630 GND.n3013 GND.n458 6971.5
R631 GND.n2999 GND.n459 6971.5
R632 GND.n3013 GND.n459 6971.5
R633 GND.n3018 GND.n2994 6971.5
R634 GND.n3018 GND.n2995 6971.5
R635 GND.n2994 GND.n2993 6971.5
R636 GND.n2995 GND.n2993 6971.5
R637 GND.n3031 GND.n466 6971.5
R638 GND.n3031 GND.n467 6971.5
R639 GND.n466 GND.n465 6971.5
R640 GND.n467 GND.n465 6971.5
R641 GND.n480 GND.n477 6971.5
R642 GND.n485 GND.n477 6971.5
R643 GND.n481 GND.n480 6971.5
R644 GND.n485 GND.n481 6971.5
R645 GND.n2969 GND.n461 6971.5
R646 GND.n2971 GND.n461 6971.5
R647 GND.n2969 GND.n462 6971.5
R648 GND.n2971 GND.n462 6971.5
R649 GND.n2975 GND.n483 6971.5
R650 GND.n2981 GND.n483 6971.5
R651 GND.n2975 GND.n484 6971.5
R652 GND.n2981 GND.n484 6971.5
R653 GND.n3256 GND.n3178 6971.5
R654 GND.n3270 GND.n3178 6971.5
R655 GND.n3256 GND.n3179 6971.5
R656 GND.n3270 GND.n3179 6971.5
R657 GND.n3275 GND.n3251 6971.5
R658 GND.n3275 GND.n3252 6971.5
R659 GND.n3251 GND.n3250 6971.5
R660 GND.n3252 GND.n3250 6971.5
R661 GND.n3288 GND.n3186 6971.5
R662 GND.n3288 GND.n3187 6971.5
R663 GND.n3186 GND.n3185 6971.5
R664 GND.n3187 GND.n3185 6971.5
R665 GND.n3200 GND.n3197 6971.5
R666 GND.n3201 GND.n3197 6971.5
R667 GND.n3202 GND.n3200 6971.5
R668 GND.n3202 GND.n3201 6971.5
R669 GND.n3226 GND.n3181 6971.5
R670 GND.n3228 GND.n3181 6971.5
R671 GND.n3226 GND.n3182 6971.5
R672 GND.n3228 GND.n3182 6971.5
R673 GND.n3232 GND.n3204 6971.5
R674 GND.n3238 GND.n3204 6971.5
R675 GND.n3232 GND.n3205 6971.5
R676 GND.n3238 GND.n3205 6971.5
R677 GND.n4179 GND.n4100 6971.5
R678 GND.n4193 GND.n4100 6971.5
R679 GND.n4179 GND.n4101 6971.5
R680 GND.n4193 GND.n4101 6971.5
R681 GND.n4198 GND.n4174 6971.5
R682 GND.n4198 GND.n4175 6971.5
R683 GND.n4174 GND.n4173 6971.5
R684 GND.n4175 GND.n4173 6971.5
R685 GND.n4211 GND.n4108 6971.5
R686 GND.n4211 GND.n4109 6971.5
R687 GND.n4108 GND.n4107 6971.5
R688 GND.n4109 GND.n4107 6971.5
R689 GND.n4122 GND.n4119 6971.5
R690 GND.n4127 GND.n4119 6971.5
R691 GND.n4123 GND.n4122 6971.5
R692 GND.n4127 GND.n4123 6971.5
R693 GND.n4149 GND.n4103 6971.5
R694 GND.n4151 GND.n4103 6971.5
R695 GND.n4149 GND.n4104 6971.5
R696 GND.n4151 GND.n4104 6971.5
R697 GND.n4155 GND.n4125 6971.5
R698 GND.n4161 GND.n4125 6971.5
R699 GND.n4155 GND.n4126 6971.5
R700 GND.n4161 GND.n4126 6971.5
R701 GND.n4239 GND.n52 6971.5
R702 GND.n4274 GND.n4239 6971.5
R703 GND.n4240 GND.n52 6971.5
R704 GND.n4274 GND.n4240 6971.5
R705 GND.n2297 GND.n2296 6705.65
R706 GND.n2523 GND.n526 5288.7
R707 GND.n4261 GND.n51 5246.88
R708 GND.n4261 GND.n4238 5246.88
R709 GND.n4264 GND.n51 5246.88
R710 GND.n4264 GND.n4238 5246.88
R711 GND.n43 GND.n32 5246.88
R712 GND.n4314 GND.n32 5246.88
R713 GND.n43 GND.n33 5246.88
R714 GND.n4314 GND.n33 5246.88
R715 GND.n40 GND.n39 5246.88
R716 GND.n4301 GND.n39 5246.88
R717 GND.n4301 GND.n4300 5246.88
R718 GND.n4300 GND.n40 5246.88
R719 GND.n4012 GND.n66 5246.88
R720 GND.n4008 GND.n66 5246.88
R721 GND.n4012 GND.n70 5246.88
R722 GND.n4008 GND.n70 5246.88
R723 GND.n4000 GND.n88 5246.88
R724 GND.n4001 GND.n88 5246.88
R725 GND.n4042 GND.n4000 5246.88
R726 GND.n4042 GND.n4001 5246.88
R727 GND.n3983 GND.n115 5246.88
R728 GND.n3983 GND.n116 5246.88
R729 GND.n115 GND.n111 5246.88
R730 GND.n116 GND.n111 5246.88
R731 GND.n3986 GND.n106 5246.88
R732 GND.n3986 GND.n107 5246.88
R733 GND.n110 GND.n107 5246.88
R734 GND.n110 GND.n106 5246.88
R735 GND.n414 GND.n387 5246.88
R736 GND.n414 GND.n413 5246.88
R737 GND.n412 GND.n387 5246.88
R738 GND.n413 GND.n412 5246.88
R739 GND.n408 GND.n359 5246.88
R740 GND.n420 GND.n408 5246.88
R741 GND.n421 GND.n359 5246.88
R742 GND.n421 GND.n420 5246.88
R743 GND.n3090 GND.n3051 5246.88
R744 GND.n3086 GND.n3051 5246.88
R745 GND.n3090 GND.n3055 5246.88
R746 GND.n3086 GND.n3055 5246.88
R747 GND.n3078 GND.n3073 5246.88
R748 GND.n3079 GND.n3073 5246.88
R749 GND.n3120 GND.n3078 5246.88
R750 GND.n3120 GND.n3079 5246.88
R751 GND.n2934 GND.n2917 5246.88
R752 GND.n2934 GND.n2918 5246.88
R753 GND.n2917 GND.n2912 5246.88
R754 GND.n2918 GND.n2912 5246.88
R755 GND.n2937 GND.n2907 5246.88
R756 GND.n2937 GND.n2908 5246.88
R757 GND.n2911 GND.n2908 5246.88
R758 GND.n2911 GND.n2907 5246.88
R759 GND.n544 GND.n534 5246.88
R760 GND.n2809 GND.n534 5246.88
R761 GND.n544 GND.n537 5246.88
R762 GND.n2809 GND.n537 5246.88
R763 GND.n2537 GND.n2497 5246.88
R764 GND.n2533 GND.n2497 5246.88
R765 GND.n2537 GND.n2501 5246.88
R766 GND.n2533 GND.n2501 5246.88
R767 GND.n2525 GND.n2519 5246.88
R768 GND.n2526 GND.n2519 5246.88
R769 GND.n2567 GND.n2525 5246.88
R770 GND.n2567 GND.n2526 5246.88
R771 GND.n2816 GND.n528 5246.88
R772 GND.n2812 GND.n528 5246.88
R773 GND.n2812 GND.n529 5246.88
R774 GND.n2816 GND.n529 5246.88
R775 GND.n2378 GND.n2349 5246.88
R776 GND.n2369 GND.n2349 5246.88
R777 GND.n2378 GND.n2350 5246.88
R778 GND.n2369 GND.n2350 5246.88
R779 GND.n1792 GND.n1754 5246.88
R780 GND.n1788 GND.n1754 5246.88
R781 GND.n1792 GND.n1758 5246.88
R782 GND.n1788 GND.n1758 5246.88
R783 GND.n1780 GND.n1777 5246.88
R784 GND.n1781 GND.n1777 5246.88
R785 GND.n1822 GND.n1780 5246.88
R786 GND.n1822 GND.n1781 5246.88
R787 GND.n2280 GND.n637 5246.88
R788 GND.n2266 GND.n637 5246.88
R789 GND.n2280 GND.n638 5246.88
R790 GND.n2266 GND.n638 5246.88
R791 GND.n872 GND.n824 5246.88
R792 GND.n2006 GND.n824 5246.88
R793 GND.n872 GND.n827 5246.88
R794 GND.n2006 GND.n827 5246.88
R795 GND.n1535 GND.n902 5246.88
R796 GND.n1531 GND.n902 5246.88
R797 GND.n1535 GND.n906 5246.88
R798 GND.n1531 GND.n906 5246.88
R799 GND.n1523 GND.n924 5246.88
R800 GND.n1524 GND.n924 5246.88
R801 GND.n1565 GND.n1523 5246.88
R802 GND.n1565 GND.n1524 5246.88
R803 GND.n2013 GND.n818 5246.88
R804 GND.n2009 GND.n818 5246.88
R805 GND.n2009 GND.n819 5246.88
R806 GND.n2013 GND.n819 5246.88
R807 GND.n855 GND.n833 5246.88
R808 GND.n857 GND.n833 5246.88
R809 GND.n856 GND.n855 5246.88
R810 GND.n857 GND.n856 5246.88
R811 GND.n1187 GND.n945 5246.88
R812 GND.n1183 GND.n945 5246.88
R813 GND.n1187 GND.n949 5246.88
R814 GND.n1183 GND.n949 5246.88
R815 GND.n1175 GND.n967 5246.88
R816 GND.n1176 GND.n967 5246.88
R817 GND.n1217 GND.n1175 5246.88
R818 GND.n1217 GND.n1176 5246.88
R819 GND.n1317 GND.n1277 5246.88
R820 GND.n1313 GND.n1277 5246.88
R821 GND.n1317 GND.n1281 5246.88
R822 GND.n1313 GND.n1281 5246.88
R823 GND.n1305 GND.n1299 5246.88
R824 GND.n1306 GND.n1299 5246.88
R825 GND.n1347 GND.n1305 5246.88
R826 GND.n1347 GND.n1306 5246.88
R827 GND.n1447 GND.n930 5246.88
R828 GND.n1457 GND.n1447 5246.88
R829 GND.n1448 GND.n930 5246.88
R830 GND.n1457 GND.n1448 5246.88
R831 GND.n1428 GND.n1425 5246.88
R832 GND.n1429 GND.n1425 5246.88
R833 GND.n1487 GND.n1428 5246.88
R834 GND.n1487 GND.n1429 5246.88
R835 GND.n1157 GND.n1129 5246.88
R836 GND.n1143 GND.n1129 5246.88
R837 GND.n1157 GND.n1130 5246.88
R838 GND.n1143 GND.n1130 5246.88
R839 GND.n1052 GND.n1007 5246.88
R840 GND.n1048 GND.n1007 5246.88
R841 GND.n1052 GND.n1010 5246.88
R842 GND.n1048 GND.n1010 5246.88
R843 GND.n2087 GND.n693 5246.88
R844 GND.n2087 GND.n694 5246.88
R845 GND.n2089 GND.n693 5246.88
R846 GND.n2089 GND.n694 5246.88
R847 GND.n3945 GND.n3896 5246.88
R848 GND.n3938 GND.n3896 5246.88
R849 GND.n3945 GND.n3897 5246.88
R850 GND.n3938 GND.n3897 5246.88
R851 GND.n3425 GND.n3384 5246.88
R852 GND.n3418 GND.n3384 5246.88
R853 GND.n3425 GND.n3385 5246.88
R854 GND.n3418 GND.n3385 5246.88
R855 GND.n4339 GND.n14 5246.88
R856 GND.n4353 GND.n14 5246.88
R857 GND.n4339 GND.n15 5246.88
R858 GND.n4353 GND.n15 5246.88
R859 GND.n167 GND.n145 5246.88
R860 GND.n169 GND.n145 5246.88
R861 GND.n168 GND.n167 5246.88
R862 GND.n169 GND.n168 5246.88
R863 GND.n3357 GND.n339 5246.88
R864 GND.n3370 GND.n339 5246.88
R865 GND.n3357 GND.n340 5246.88
R866 GND.n3370 GND.n340 5246.88
R867 GND.n2773 GND.n2750 5246.88
R868 GND.n2775 GND.n2750 5246.88
R869 GND.n2774 GND.n2773 5246.88
R870 GND.n2775 GND.n2774 5246.88
R871 GND.n2310 GND.n607 5246.88
R872 GND.n2321 GND.n607 5246.88
R873 GND.n2310 GND.n608 5246.88
R874 GND.n2321 GND.n608 5246.88
R875 GND.n2317 GND.n609 5246.88
R876 GND.n2317 GND.n610 5246.88
R877 GND.n2313 GND.n610 5246.88
R878 GND.n2313 GND.n609 5246.88
R879 GND.n791 GND.n781 5246.88
R880 GND.n2047 GND.n781 5246.88
R881 GND.n791 GND.n784 5246.88
R882 GND.n2047 GND.n784 5246.88
R883 GND.n2050 GND.n775 5246.88
R884 GND.n2050 GND.n776 5246.88
R885 GND.n2054 GND.n776 5246.88
R886 GND.n2054 GND.n775 5246.88
R887 GND.n989 GND.n988 5246.88
R888 GND.n1104 GND.n988 5246.88
R889 GND.n1103 GND.n989 5246.88
R890 GND.n1104 GND.n1103 5246.88
R891 GND.n1100 GND.n991 5246.88
R892 GND.n1100 GND.n992 5246.88
R893 GND.n1096 GND.n992 5246.88
R894 GND.n1096 GND.n991 5246.88
R895 GND.n757 GND.n730 5246.88
R896 GND.n750 GND.n730 5246.88
R897 GND.n757 GND.n731 5246.88
R898 GND.n750 GND.n731 5246.88
R899 GND.n2887 GND.n309 5246.88
R900 GND.n3469 GND.n309 5246.88
R901 GND.n2887 GND.n310 5246.88
R902 GND.n3469 GND.n310 5246.88
R903 GND.n2842 GND.n514 5246.88
R904 GND.n2848 GND.n514 5246.88
R905 GND.n2842 GND.n515 5246.88
R906 GND.n2848 GND.n515 5246.88
R907 GND.n2245 GND.n2185 5246.88
R908 GND.n2238 GND.n2185 5246.88
R909 GND.n2245 GND.n2186 5246.88
R910 GND.n2238 GND.n2186 5246.88
R911 GND.n2141 GND.n664 5246.88
R912 GND.n2147 GND.n664 5246.88
R913 GND.n2141 GND.n665 5246.88
R914 GND.n2147 GND.n665 5246.88
R915 GND.n1921 GND.n887 5246.88
R916 GND.n1931 GND.n1921 5246.88
R917 GND.n1922 GND.n887 5246.88
R918 GND.n1931 GND.n1922 5246.88
R919 GND.n1902 GND.n1899 5246.88
R920 GND.n1903 GND.n1899 5246.88
R921 GND.n1961 GND.n1902 5246.88
R922 GND.n1961 GND.n1903 5246.88
R923 GND.n1665 GND.n1626 5246.88
R924 GND.n1661 GND.n1626 5246.88
R925 GND.n1665 GND.n1630 5246.88
R926 GND.n1661 GND.n1630 5246.88
R927 GND.n1653 GND.n1648 5246.88
R928 GND.n1654 GND.n1648 5246.88
R929 GND.n1695 GND.n1653 5246.88
R930 GND.n1695 GND.n1654 5246.88
R931 GND.n2407 GND.n573 5246.88
R932 GND.n2403 GND.n573 5246.88
R933 GND.n2407 GND.n577 5246.88
R934 GND.n2403 GND.n577 5246.88
R935 GND.n2395 GND.n595 5246.88
R936 GND.n2396 GND.n595 5246.88
R937 GND.n2437 GND.n2395 5246.88
R938 GND.n2437 GND.n2396 5246.88
R939 GND.n2667 GND.n558 5246.88
R940 GND.n2677 GND.n2667 5246.88
R941 GND.n2668 GND.n558 5246.88
R942 GND.n2677 GND.n2668 5246.88
R943 GND.n2648 GND.n2645 5246.88
R944 GND.n2649 GND.n2645 5246.88
R945 GND.n2707 GND.n2648 5246.88
R946 GND.n2707 GND.n2649 5246.88
R947 GND.n2961 GND.n460 5246.88
R948 GND.n2957 GND.n460 5246.88
R949 GND.n2961 GND.n464 5246.88
R950 GND.n2957 GND.n464 5246.88
R951 GND.n2949 GND.n482 5246.88
R952 GND.n2950 GND.n482 5246.88
R953 GND.n2991 GND.n2949 5246.88
R954 GND.n2991 GND.n2950 5246.88
R955 GND.n3218 GND.n3180 5246.88
R956 GND.n3214 GND.n3180 5246.88
R957 GND.n3218 GND.n3184 5246.88
R958 GND.n3214 GND.n3184 5246.88
R959 GND.n3206 GND.n3203 5246.88
R960 GND.n3207 GND.n3203 5246.88
R961 GND.n3248 GND.n3206 5246.88
R962 GND.n3248 GND.n3207 5246.88
R963 GND.n4141 GND.n4102 5246.88
R964 GND.n4137 GND.n4102 5246.88
R965 GND.n4141 GND.n4106 5246.88
R966 GND.n4137 GND.n4106 5246.88
R967 GND.n4129 GND.n4124 5246.88
R968 GND.n4130 GND.n4124 5246.88
R969 GND.n4171 GND.n4129 5246.88
R970 GND.n4171 GND.n4130 5246.88
R971 GND.n2947 GND.n2946 4866.1
R972 GND.n3998 GND.n3997 4362.71
R973 GND.n4249 GND.n53 3522.26
R974 GND.n4249 GND.n4237 3522.26
R975 GND.n4252 GND.n53 3522.26
R976 GND.n4252 GND.n4237 3522.26
R977 GND.n4083 GND.n60 3522.26
R978 GND.n4083 GND.n62 3522.26
R979 GND.n4084 GND.n60 3522.26
R980 GND.n4084 GND.n62 3522.26
R981 GND.n4043 GND.n81 3522.26
R982 GND.n4043 GND.n79 3522.26
R983 GND.n4070 GND.n81 3522.26
R984 GND.n4070 GND.n79 3522.26
R985 GND.n3318 GND.n446 3522.26
R986 GND.n449 GND.n446 3522.26
R987 GND.n3318 GND.n447 3522.26
R988 GND.n449 GND.n447 3522.26
R989 GND.n395 GND.n361 3522.26
R990 GND.n396 GND.n395 3522.26
R991 GND.n398 GND.n361 3522.26
R992 GND.n398 GND.n396 3522.26
R993 GND.n3161 GND.n3045 3522.26
R994 GND.n3161 GND.n3047 3522.26
R995 GND.n3162 GND.n3045 3522.26
R996 GND.n3162 GND.n3047 3522.26
R997 GND.n3121 GND.n3066 3522.26
R998 GND.n3121 GND.n3064 3522.26
R999 GND.n3148 GND.n3066 3522.26
R1000 GND.n3148 GND.n3064 3522.26
R1001 GND.n2608 GND.n2491 3522.26
R1002 GND.n2608 GND.n2493 3522.26
R1003 GND.n2609 GND.n2491 3522.26
R1004 GND.n2609 GND.n2493 3522.26
R1005 GND.n2568 GND.n2512 3522.26
R1006 GND.n2568 GND.n2510 3522.26
R1007 GND.n2595 GND.n2512 3522.26
R1008 GND.n2595 GND.n2510 3522.26
R1009 GND.n2343 GND.n2337 3522.26
R1010 GND.n2347 GND.n2337 3522.26
R1011 GND.n2343 GND.n2338 3522.26
R1012 GND.n2347 GND.n2338 3522.26
R1013 GND.n2367 GND.n2359 3522.26
R1014 GND.n2367 GND.n2360 3522.26
R1015 GND.n2360 GND.n2358 3522.26
R1016 GND.n2359 GND.n2358 3522.26
R1017 GND.n1863 GND.n1749 3522.26
R1018 GND.n1863 GND.n1751 3522.26
R1019 GND.n1864 GND.n1749 3522.26
R1020 GND.n1864 GND.n1751 3522.26
R1021 GND.n1823 GND.n1769 3522.26
R1022 GND.n1823 GND.n1767 3522.26
R1023 GND.n1850 GND.n1769 3522.26
R1024 GND.n1850 GND.n1767 3522.26
R1025 GND.n2293 GND.n625 3522.26
R1026 GND.n635 GND.n625 3522.26
R1027 GND.n2293 GND.n626 3522.26
R1028 GND.n635 GND.n626 3522.26
R1029 GND.n2264 GND.n2259 3522.26
R1030 GND.n2270 GND.n2259 3522.26
R1031 GND.n2270 GND.n2261 3522.26
R1032 GND.n2264 GND.n2261 3522.26
R1033 GND.n1606 GND.n896 3522.26
R1034 GND.n1606 GND.n898 3522.26
R1035 GND.n1607 GND.n896 3522.26
R1036 GND.n1607 GND.n898 3522.26
R1037 GND.n1566 GND.n917 3522.26
R1038 GND.n1566 GND.n915 3522.26
R1039 GND.n1593 GND.n917 3522.26
R1040 GND.n1593 GND.n915 3522.26
R1041 GND.n838 GND.n835 3522.26
R1042 GND.n852 GND.n835 3522.26
R1043 GND.n838 GND.n836 3522.26
R1044 GND.n852 GND.n836 3522.26
R1045 GND.n2027 GND.n810 3522.26
R1046 GND.n2023 GND.n810 3522.26
R1047 GND.n2023 GND.n811 3522.26
R1048 GND.n2027 GND.n811 3522.26
R1049 GND.n1258 GND.n939 3522.26
R1050 GND.n1258 GND.n941 3522.26
R1051 GND.n1259 GND.n939 3522.26
R1052 GND.n1259 GND.n941 3522.26
R1053 GND.n1218 GND.n960 3522.26
R1054 GND.n1218 GND.n958 3522.26
R1055 GND.n1245 GND.n960 3522.26
R1056 GND.n1245 GND.n958 3522.26
R1057 GND.n1388 GND.n1271 3522.26
R1058 GND.n1388 GND.n1273 3522.26
R1059 GND.n1389 GND.n1271 3522.26
R1060 GND.n1389 GND.n1273 3522.26
R1061 GND.n1348 GND.n1292 3522.26
R1062 GND.n1348 GND.n1290 3522.26
R1063 GND.n1375 GND.n1292 3522.26
R1064 GND.n1375 GND.n1290 3522.26
R1065 GND.n1517 GND.n933 3522.26
R1066 GND.n1465 GND.n933 3522.26
R1067 GND.n1517 GND.n934 3522.26
R1068 GND.n1465 GND.n934 3522.26
R1069 GND.n1488 GND.n1417 3522.26
R1070 GND.n1488 GND.n1415 3522.26
R1071 GND.n1495 GND.n1417 3522.26
R1072 GND.n1495 GND.n1415 3522.26
R1073 GND.n1170 GND.n972 3522.26
R1074 GND.n1127 GND.n972 3522.26
R1075 GND.n1170 GND.n973 3522.26
R1076 GND.n1127 GND.n973 3522.26
R1077 GND.n1141 GND.n1136 3522.26
R1078 GND.n1147 GND.n1136 3522.26
R1079 GND.n1147 GND.n1138 3522.26
R1080 GND.n1141 GND.n1138 3522.26
R1081 GND.n1064 GND.n1002 3522.26
R1082 GND.n1064 GND.n1004 3522.26
R1083 GND.n1065 GND.n1002 3522.26
R1084 GND.n1065 GND.n1004 3522.26
R1085 GND.n3935 GND.n3904 3522.26
R1086 GND.n3913 GND.n3904 3522.26
R1087 GND.n3935 GND.n3905 3522.26
R1088 GND.n3913 GND.n3905 3522.26
R1089 GND.n3415 GND.n3390 3522.26
R1090 GND.n3401 GND.n3390 3522.26
R1091 GND.n3415 GND.n3391 3522.26
R1092 GND.n3401 GND.n3391 3522.26
R1093 GND.n4323 GND.n23 3522.26
R1094 GND.n4335 GND.n23 3522.26
R1095 GND.n4323 GND.n24 3522.26
R1096 GND.n4335 GND.n24 3522.26
R1097 GND.n4356 GND.n11 3522.26
R1098 GND.n4360 GND.n11 3522.26
R1099 GND.n4356 GND.n12 3522.26
R1100 GND.n4360 GND.n12 3522.26
R1101 GND.n150 GND.n147 3522.26
R1102 GND.n164 GND.n147 3522.26
R1103 GND.n150 GND.n148 3522.26
R1104 GND.n164 GND.n148 3522.26
R1105 GND.n3964 GND.n140 3522.26
R1106 GND.n3960 GND.n140 3522.26
R1107 GND.n3960 GND.n141 3522.26
R1108 GND.n3964 GND.n141 3522.26
R1109 GND.n3341 GND.n348 3522.26
R1110 GND.n3353 GND.n348 3522.26
R1111 GND.n3341 GND.n349 3522.26
R1112 GND.n3353 GND.n349 3522.26
R1113 GND.n3376 GND.n336 3522.26
R1114 GND.n3376 GND.n337 3522.26
R1115 GND.n3375 GND.n337 3522.26
R1116 GND.n3375 GND.n336 3522.26
R1117 GND.n2756 GND.n2752 3522.26
R1118 GND.n2770 GND.n2752 3522.26
R1119 GND.n2756 GND.n2753 3522.26
R1120 GND.n2770 GND.n2753 3522.26
R1121 GND.n2788 GND.n2745 3522.26
R1122 GND.n2784 GND.n2745 3522.26
R1123 GND.n2784 GND.n2746 3522.26
R1124 GND.n2788 GND.n2746 3522.26
R1125 GND.n747 GND.n738 3522.26
R1126 GND.n741 GND.n738 3522.26
R1127 GND.n747 GND.n739 3522.26
R1128 GND.n741 GND.n739 3522.26
R1129 GND.n319 GND.n318 3522.26
R1130 GND.n3461 GND.n319 3522.26
R1131 GND.n318 GND.n316 3522.26
R1132 GND.n3461 GND.n316 3522.26
R1133 GND.n2845 GND.n507 3522.26
R1134 GND.n2857 GND.n507 3522.26
R1135 GND.n2845 GND.n508 3522.26
R1136 GND.n2857 GND.n508 3522.26
R1137 GND.n2235 GND.n2193 3522.26
R1138 GND.n2200 GND.n2193 3522.26
R1139 GND.n2235 GND.n2194 3522.26
R1140 GND.n2200 GND.n2194 3522.26
R1141 GND.n2144 GND.n657 3522.26
R1142 GND.n2156 GND.n657 3522.26
R1143 GND.n2144 GND.n658 3522.26
R1144 GND.n2156 GND.n658 3522.26
R1145 GND.n2082 GND.n697 3522.26
R1146 GND.n711 GND.n697 3522.26
R1147 GND.n2082 GND.n698 3522.26
R1148 GND.n711 GND.n698 3522.26
R1149 GND.n1991 GND.n890 3522.26
R1150 GND.n1939 GND.n890 3522.26
R1151 GND.n1991 GND.n891 3522.26
R1152 GND.n1939 GND.n891 3522.26
R1153 GND.n1962 GND.n1891 3522.26
R1154 GND.n1962 GND.n1889 3522.26
R1155 GND.n1969 GND.n1891 3522.26
R1156 GND.n1969 GND.n1889 3522.26
R1157 GND.n1736 GND.n1620 3522.26
R1158 GND.n1736 GND.n1622 3522.26
R1159 GND.n1737 GND.n1620 3522.26
R1160 GND.n1737 GND.n1622 3522.26
R1161 GND.n1696 GND.n1641 3522.26
R1162 GND.n1696 GND.n1639 3522.26
R1163 GND.n1723 GND.n1641 3522.26
R1164 GND.n1723 GND.n1639 3522.26
R1165 GND.n2478 GND.n567 3522.26
R1166 GND.n2478 GND.n569 3522.26
R1167 GND.n2479 GND.n567 3522.26
R1168 GND.n2479 GND.n569 3522.26
R1169 GND.n2438 GND.n588 3522.26
R1170 GND.n2438 GND.n586 3522.26
R1171 GND.n2465 GND.n588 3522.26
R1172 GND.n2465 GND.n586 3522.26
R1173 GND.n2737 GND.n561 3522.26
R1174 GND.n2685 GND.n561 3522.26
R1175 GND.n2737 GND.n562 3522.26
R1176 GND.n2685 GND.n562 3522.26
R1177 GND.n2708 GND.n2637 3522.26
R1178 GND.n2708 GND.n2635 3522.26
R1179 GND.n2715 GND.n2637 3522.26
R1180 GND.n2715 GND.n2635 3522.26
R1181 GND.n3032 GND.n454 3522.26
R1182 GND.n3032 GND.n456 3522.26
R1183 GND.n3033 GND.n454 3522.26
R1184 GND.n3033 GND.n456 3522.26
R1185 GND.n2992 GND.n475 3522.26
R1186 GND.n2992 GND.n473 3522.26
R1187 GND.n3019 GND.n475 3522.26
R1188 GND.n3019 GND.n473 3522.26
R1189 GND.n3289 GND.n3175 3522.26
R1190 GND.n3289 GND.n3177 3522.26
R1191 GND.n3290 GND.n3175 3522.26
R1192 GND.n3290 GND.n3177 3522.26
R1193 GND.n3249 GND.n3195 3522.26
R1194 GND.n3249 GND.n3193 3522.26
R1195 GND.n3276 GND.n3195 3522.26
R1196 GND.n3276 GND.n3193 3522.26
R1197 GND.n4212 GND.n4096 3522.26
R1198 GND.n4212 GND.n4098 3522.26
R1199 GND.n4213 GND.n4096 3522.26
R1200 GND.n4213 GND.n4098 3522.26
R1201 GND.n4172 GND.n4117 3522.26
R1202 GND.n4172 GND.n4115 3522.26
R1203 GND.n4199 GND.n4117 3522.26
R1204 GND.n4199 GND.n4115 3522.26
R1205 GND.n1521 GND.n1520 3449.15
R1206 GND.n4288 GND.n49 3026.55
R1207 GND.n3490 GND.n3471 1967.95
R1208 GND.n3509 GND.n300 1967.95
R1209 GND.n3531 GND.n292 1967.95
R1210 GND.n3553 GND.n284 1967.95
R1211 GND.n3572 GND.n276 1967.95
R1212 GND.n3592 GND.n268 1967.95
R1213 GND.n3611 GND.n250 1967.95
R1214 GND.n2182 GND.n2181 1886.95
R1215 GND.n2883 GND.n2882 1886.95
R1216 GND.n2212 GND.n284 1746.61
R1217 GND.n1113 GND.n982 1691.24
R1218 GND.t0 GND.t514 1325.61
R1219 GND.t514 GND.t693 1325.61
R1220 GND.t578 GND.t219 1325.61
R1221 GND.t219 GND.t115 1325.61
R1222 GND.t339 GND.t687 1325.61
R1223 GND.t308 GND.t602 1325.61
R1224 GND.t338 GND.t72 1325.61
R1225 GND.t174 GND.t338 1325.61
R1226 GND.t612 GND.t200 1325.61
R1227 GND.t200 GND.t510 1325.61
R1228 GND.t131 GND.t268 1325.61
R1229 GND.t268 GND.t697 1325.61
R1230 GND.t33 GND.t48 1325.61
R1231 GND.t48 GND.t159 1325.61
R1232 GND.t120 GND.t660 1325.61
R1233 GND.t120 GND.t695 1325.61
R1234 GND.t361 GND.t71 1325.61
R1235 GND.t329 GND.t361 1325.61
R1236 GND.n2127 GND.n2126 1316.99
R1237 GND.n3438 GND.n3437 1316.99
R1238 GND.n3895 GND.n3894 1316.99
R1239 GND.t504 GND.n268 1083.81
R1240 GND.n2100 GND.n680 1036.71
R1241 GND.n2320 GND.n2319 999.98
R1242 GND.n2048 GND.n780 999.98
R1243 GND.n1112 GND.n984 999.98
R1244 GND.n3334 GND.n356 999.98
R1245 GND.n128 GND.n127 999.98
R1246 GND.n4316 GND.n4315 999.98
R1247 GND.t305 GND.t666 994.698
R1248 GND.t311 GND.t655 994.698
R1249 GND.t320 GND.t653 994.698
R1250 GND.t619 GND.t117 994.698
R1251 GND.t157 GND.t594 994.698
R1252 GND.t54 GND.t591 994.698
R1253 GND.t227 GND.t254 994.698
R1254 GND.t292 GND.t288 994.698
R1255 GND.t605 GND.t346 994.698
R1256 GND.t699 GND.t284 994.698
R1257 GND.t59 GND.t153 994.698
R1258 GND.t295 GND.t104 994.698
R1259 GND.t45 GND.t719 994.698
R1260 GND.t275 GND.n982 993.078
R1261 GND.n3882 GND.n3881 987.285
R1262 GND.n1114 GND.t677 931.518
R1263 GND.t56 GND.t683 925.207
R1264 GND.t56 GND.t188 925.207
R1265 GND.t256 GND.t337 925.207
R1266 GND.t4 GND.t315 925.207
R1267 GND.t315 GND.t313 925.207
R1268 GND.t185 GND.t667 925.207
R1269 GND.t667 GND.t164 925.207
R1270 GND.t64 GND.t286 925.207
R1271 GND.t576 GND.t64 925.207
R1272 GND.t214 GND.t701 925.207
R1273 GND.t599 GND.t214 925.207
R1274 GND.t668 GND.t99 925.207
R1275 GND.t668 GND.t331 925.207
R1276 GND.t156 GND.t287 925.207
R1277 GND.t340 GND.t259 925.207
R1278 GND.t340 GND.t691 925.207
R1279 GND.t328 GND.t150 925.207
R1280 GND.t328 GND.t190 925.207
R1281 GND.t364 GND.t507 925.207
R1282 GND.t507 GND.t102 925.207
R1283 GND.t281 GND.n773 912.077
R1284 GND.n1520 GND.t645 912.077
R1285 GND.n2297 GND.t291 912.077
R1286 GND.t49 GND.n526 912.077
R1287 GND.n2946 GND.t213 912.077
R1288 GND.n3995 GND.t132 912.077
R1289 GND.t220 GND.n4288 912.077
R1290 GND.n802 GND.t111 806.775
R1291 GND.n2392 GND.t649 806.775
R1292 GND.t634 GND.n3333 806.775
R1293 GND.n3997 GND.t194 806.775
R1294 GND.t366 GND.n10 806.775
R1295 GND.t222 GND.n276 803.14
R1296 GND.t158 GND.t581 789.019
R1297 GND.t723 GND.t69 789.019
R1298 GND.n1994 GND.t717 781.308
R1299 GND.t287 GND.n3882 763.973
R1300 GND.n165 GND.t344 736.533
R1301 GND.n166 GND.t124 736.533
R1302 GND.n3354 GND.t321 736.533
R1303 GND.t584 GND.n3358 736.533
R1304 GND.n2771 GND.t306 736.533
R1305 GND.n2772 GND.t636 736.533
R1306 GND.n4336 GND.t151 736.533
R1307 GND.t625 GND.n4340 736.533
R1308 GND.n4361 GND.t252 736.533
R1309 GND.n1128 GND.t664 736.533
R1310 GND.n1158 GND.t85 736.533
R1311 GND.n853 GND.t572 736.533
R1312 GND.n854 GND.t622 736.533
R1313 GND.n636 GND.t512 736.533
R1314 GND.n2281 GND.t122 736.533
R1315 GND.n2348 GND.t352 736.533
R1316 GND.n2379 GND.t624 736.533
R1317 GND.t677 GND.n1113 701.473
R1318 GND.t293 GND.t324 690.949
R1319 GND.n616 GND.n615 690.949
R1320 GND.t362 GND.t176 690.949
R1321 GND.n2320 GND.n2318 690.949
R1322 GND.t100 GND.t197 690.949
R1323 GND.n783 GND.n782 690.949
R1324 GND.t257 GND.t669 690.949
R1325 GND.n2049 GND.n2048 690.949
R1326 GND.t136 GND.t147 690.949
R1327 GND.n1102 GND.n990 690.949
R1328 GND.t318 GND.t601 690.949
R1329 GND.n1101 GND.n984 690.949
R1330 GND.t19 GND.t46 690.949
R1331 GND.n826 GND.n825 690.949
R1332 GND.t1 GND.t119 690.949
R1333 GND.n2008 GND.n2007 690.949
R1334 GND.t225 GND.t506 690.949
R1335 GND.n536 GND.n535 690.949
R1336 GND.t215 GND.t609 690.949
R1337 GND.n2811 GND.n2810 690.949
R1338 GND.t229 GND.t26 690.949
R1339 GND.n2936 GND.n2935 690.949
R1340 GND.t51 GND.t348 690.949
R1341 GND.n2913 GND.n356 690.949
R1342 GND.t230 GND.t678 690.949
R1343 GND.n3985 GND.n3984 690.949
R1344 GND.t517 GND.t97 690.949
R1345 GND.n127 GND.n126 690.949
R1346 GND.t270 GND.t310 690.949
R1347 GND.n4299 GND.n4298 690.949
R1348 GND.t129 GND.t203 690.949
R1349 GND.n4315 GND.n31 690.949
R1350 GND.n1993 GND.n823 669.51
R1351 GND.n555 GND.n533 669.51
R1352 GND.n2146 GND.t715 662.808
R1353 GND.n2145 GND.t657 662.808
R1354 GND.n2157 GND.t657 662.808
R1355 GND.n2158 GND.t0 662.808
R1356 GND.n2170 GND.t578 662.808
R1357 GND.n2181 GND.t115 662.808
R1358 GND.n2182 GND.t504 662.808
R1359 GND.t687 GND.n2247 662.808
R1360 GND.n2246 GND.t294 662.808
R1361 GND.n2192 GND.t294 662.808
R1362 GND.t647 GND.n2192 662.808
R1363 GND.n2237 GND.t647 662.808
R1364 GND.n2236 GND.t515 662.808
R1365 GND.n2201 GND.t515 662.808
R1366 GND.n2202 GND.t222 662.808
R1367 GND.t602 GND.n2223 662.808
R1368 GND.n2222 GND.t72 662.808
R1369 GND.n2212 GND.t174 662.808
R1370 GND.n2828 GND.t612 662.808
R1371 GND.n2839 GND.t510 662.808
R1372 GND.t505 GND.n2843 662.808
R1373 GND.n2844 GND.t505 662.808
R1374 GND.t67 GND.n2844 662.808
R1375 GND.n2847 GND.t67 662.808
R1376 GND.n2846 GND.t34 662.808
R1377 GND.n2859 GND.t131 662.808
R1378 GND.n2870 GND.t697 662.808
R1379 GND.n2871 GND.t33 662.808
R1380 GND.t660 GND.n2883 662.808
R1381 GND.t695 GND.n2889 662.808
R1382 GND.n2888 GND.t228 662.808
R1383 GND.t228 GND.n2884 662.808
R1384 GND.n2884 GND.t607 662.808
R1385 GND.t300 GND.n308 662.808
R1386 GND.n3460 GND.t300 662.808
R1387 GND.n3459 GND.t71 662.808
R1388 GND.n3449 GND.t329 662.808
R1389 GND.t124 GND.t166 626.173
R1390 GND.n3966 GND.n138 626.173
R1391 GND.t279 GND.t584 626.173
R1392 GND.n3360 GND.n3359 626.173
R1393 GND.t636 GND.t162 626.173
R1394 GND.n2790 GND.n2743 626.173
R1395 GND.t335 GND.t625 626.173
R1396 GND.n4342 GND.n4341 626.173
R1397 GND.t236 GND.t85 626.173
R1398 GND.n1140 GND.n1139 626.173
R1399 GND.t622 GND.t186 626.173
R1400 GND.n2029 GND.n808 626.173
R1401 GND.t689 GND.t122 626.173
R1402 GND.n2263 GND.n2262 626.173
R1403 GND.t277 GND.t624 626.173
R1404 GND.n2354 GND.n2353 626.173
R1405 GND.n2169 GND.n250 623.946
R1406 GND.t715 GND.n2143 608.681
R1407 GND.n2102 GND.n2101 584.846
R1408 GND.n2102 GND.n2100 578.735
R1409 GND.t337 GND.n2102 568.082
R1410 GND.t344 GND.t180 535.005
R1411 GND.n3965 GND.n139 535.005
R1412 GND.t302 GND.t321 535.005
R1413 GND.n3371 GND.n338 535.005
R1414 GND.t265 GND.t306 535.005
R1415 GND.n2789 GND.n2744 535.005
R1416 GND.t365 GND.t151 535.005
R1417 GND.n4355 GND.n4354 535.005
R1418 GND.t664 GND.t264 535.005
R1419 GND.n1144 GND.n1142 535.005
R1420 GND.t572 GND.t639 535.005
R1421 GND.n2028 GND.n809 535.005
R1422 GND.t512 GND.t579 535.005
R1423 GND.n2267 GND.n2265 535.005
R1424 GND.t304 GND.t352 535.005
R1425 GND.n2368 GND.n2355 535.005
R1426 GND.t308 GND.n276 522.473
R1427 GND.t34 GND.n292 522.473
R1428 GND.t159 GND.n300 522.473
R1429 GND.n1087 GND.t305 497.349
R1430 GND.n1093 GND.t275 497.349
R1431 GND.t146 GND.n1112 497.349
R1432 GND.n1146 GND.t17 497.349
R1433 GND.n1145 GND.t281 497.349
R1434 GND.t655 GND.n2056 497.349
R1435 GND.t111 GND.n780 497.349
R1436 GND.t653 GND.n2036 497.349
R1437 GND.n2022 GND.t15 497.349
R1438 GND.n2021 GND.t645 497.349
R1439 GND.n2015 GND.t117 497.349
R1440 GND.n2269 GND.t597 497.349
R1441 GND.n2268 GND.t291 497.349
R1442 GND.t594 GND.n614 497.349
R1443 GND.n2319 GND.t649 497.349
R1444 GND.n2340 GND.t591 497.349
R1445 GND.t108 GND.n2357 497.349
R1446 GND.n2356 GND.t49 497.349
R1447 GND.t254 GND.n2818 497.349
R1448 GND.n2783 GND.t13 497.349
R1449 GND.n2782 GND.t213 497.349
R1450 GND.n2914 GND.t288 497.349
R1451 GND.n3334 GND.t634 497.349
R1452 GND.n3340 GND.t346 497.349
R1453 GND.t248 GND.n3373 497.349
R1454 GND.n3372 GND.t132 497.349
R1455 GND.n112 GND.t284 497.349
R1456 GND.n128 GND.t194 497.349
R1457 GND.n3973 GND.t59 497.349
R1458 GND.t11 GND.n48 497.349
R1459 GND.n4289 GND.t220 497.349
R1460 GND.n4295 GND.t104 497.349
R1461 GND.n4316 GND.t366 497.349
R1462 GND.n4322 GND.t719 497.349
R1463 GND.n4275 GND.n10 473.918
R1464 GND.n4285 GND.n56 467.2
R1465 GND.n4285 GND.n4284 467.2
R1466 GND.n4233 GND.n4230 467.2
R1467 GND.n4234 GND.n4233 467.2
R1468 GND.n4028 GND.n4027 467.2
R1469 GND.n4027 GND.n4025 467.2
R1470 GND.n85 GND.n75 467.2
R1471 GND.n85 GND.n84 467.2
R1472 GND.n4081 GND.n4080 467.2
R1473 GND.n4080 GND.n4079 467.2
R1474 GND.n4049 GND.n4047 467.2
R1475 GND.n4068 GND.n4047 467.2
R1476 GND.n4066 GND.n4065 467.2
R1477 GND.n4065 GND.n4063 467.2
R1478 GND.n4023 GND.n4021 467.2
R1479 GND.n4024 GND.n4023 467.2
R1480 GND.n441 GND.n433 467.2
R1481 GND.n434 GND.n433 467.2
R1482 GND.n378 GND.n376 467.2
R1483 GND.n376 GND.n375 467.2
R1484 GND.n381 GND.n380 467.2
R1485 GND.n382 GND.n381 467.2
R1486 GND.n3330 GND.n3329 467.2
R1487 GND.n3330 GND.n364 467.2
R1488 GND.n3310 GND.n3306 467.2
R1489 GND.n3306 GND.n365 467.2
R1490 GND.n438 GND.n436 467.2
R1491 GND.n439 GND.n438 467.2
R1492 GND.n3106 GND.n3105 467.2
R1493 GND.n3105 GND.n3103 467.2
R1494 GND.n3070 GND.n3060 467.2
R1495 GND.n3070 GND.n3069 467.2
R1496 GND.n3159 GND.n3158 467.2
R1497 GND.n3158 GND.n3157 467.2
R1498 GND.n3127 GND.n3125 467.2
R1499 GND.n3146 GND.n3125 467.2
R1500 GND.n3144 GND.n3143 467.2
R1501 GND.n3143 GND.n3141 467.2
R1502 GND.n3101 GND.n3099 467.2
R1503 GND.n3102 GND.n3101 467.2
R1504 GND.n2553 GND.n2552 467.2
R1505 GND.n2552 GND.n2550 467.2
R1506 GND.n2516 GND.n2506 467.2
R1507 GND.n2516 GND.n2515 467.2
R1508 GND.n2606 GND.n2605 467.2
R1509 GND.n2605 GND.n2604 467.2
R1510 GND.n2574 GND.n2572 467.2
R1511 GND.n2593 GND.n2572 467.2
R1512 GND.n2591 GND.n2590 467.2
R1513 GND.n2590 GND.n2588 467.2
R1514 GND.n2548 GND.n2546 467.2
R1515 GND.n2549 GND.n2548 467.2
R1516 GND.n1808 GND.n1807 467.2
R1517 GND.n1807 GND.n1805 467.2
R1518 GND.n1773 GND.n1763 467.2
R1519 GND.n1773 GND.n1772 467.2
R1520 GND.n1861 GND.n1860 467.2
R1521 GND.n1860 GND.n1859 467.2
R1522 GND.n1829 GND.n1827 467.2
R1523 GND.n1848 GND.n1827 467.2
R1524 GND.n1846 GND.n1845 467.2
R1525 GND.n1845 GND.n1843 467.2
R1526 GND.n1803 GND.n1801 467.2
R1527 GND.n1804 GND.n1803 467.2
R1528 GND.n1551 GND.n1550 467.2
R1529 GND.n1550 GND.n1548 467.2
R1530 GND.n921 GND.n911 467.2
R1531 GND.n921 GND.n920 467.2
R1532 GND.n1604 GND.n1603 467.2
R1533 GND.n1603 GND.n1602 467.2
R1534 GND.n1572 GND.n1570 467.2
R1535 GND.n1591 GND.n1570 467.2
R1536 GND.n1589 GND.n1588 467.2
R1537 GND.n1588 GND.n1586 467.2
R1538 GND.n1546 GND.n1544 467.2
R1539 GND.n1547 GND.n1546 467.2
R1540 GND.n1203 GND.n1202 467.2
R1541 GND.n1202 GND.n1200 467.2
R1542 GND.n964 GND.n954 467.2
R1543 GND.n964 GND.n963 467.2
R1544 GND.n1256 GND.n1255 467.2
R1545 GND.n1255 GND.n1254 467.2
R1546 GND.n1224 GND.n1222 467.2
R1547 GND.n1243 GND.n1222 467.2
R1548 GND.n1241 GND.n1240 467.2
R1549 GND.n1240 GND.n1238 467.2
R1550 GND.n1198 GND.n1196 467.2
R1551 GND.n1199 GND.n1198 467.2
R1552 GND.n1333 GND.n1332 467.2
R1553 GND.n1332 GND.n1330 467.2
R1554 GND.n1296 GND.n1286 467.2
R1555 GND.n1296 GND.n1295 467.2
R1556 GND.n1386 GND.n1385 467.2
R1557 GND.n1385 GND.n1384 467.2
R1558 GND.n1354 GND.n1352 467.2
R1559 GND.n1373 GND.n1352 467.2
R1560 GND.n1371 GND.n1370 467.2
R1561 GND.n1370 GND.n1368 467.2
R1562 GND.n1328 GND.n1326 467.2
R1563 GND.n1329 GND.n1328 467.2
R1564 GND.n1473 GND.n1472 467.2
R1565 GND.n1472 GND.n1470 467.2
R1566 GND.n1423 GND.n1422 467.2
R1567 GND.n1422 GND.n1421 467.2
R1568 GND.n1462 GND.n1460 467.2
R1569 GND.n1462 GND.n1461 467.2
R1570 GND.n1492 GND.n1491 467.2
R1571 GND.n1493 GND.n1492 467.2
R1572 GND.n1445 GND.n1443 467.2
R1573 GND.n1445 GND.n1444 467.2
R1574 GND.n1439 GND.n1438 467.2
R1575 GND.n1469 GND.n1438 467.2
R1576 GND.n1062 GND.n1061 467.2
R1577 GND.n1061 GND.n1060 467.2
R1578 GND.n1025 GND.n1023 467.2
R1579 GND.n1026 GND.n1025 467.2
R1580 GND.n1036 GND.n1034 467.2
R1581 GND.n1037 GND.n1036 467.2
R1582 GND.n4320 GND.n4319 467.2
R1583 GND.n4319 GND.n4318 467.2
R1584 GND.n4293 GND.n4292 467.2
R1585 GND.n4292 GND.n4291 467.2
R1586 GND.n3969 GND.n3968 467.2
R1587 GND.n3970 GND.n3969 467.2
R1588 GND.n132 GND.n131 467.2
R1589 GND.n131 GND.n124 467.2
R1590 GND.n102 GND.n101 467.2
R1591 GND.n101 GND.n100 467.2
R1592 GND.n3362 GND.n345 467.2
R1593 GND.n3345 GND.n345 467.2
R1594 GND.n3338 GND.n3337 467.2
R1595 GND.n3337 GND.n3336 467.2
R1596 GND.n2903 GND.n2902 467.2
R1597 GND.n2902 GND.n2901 467.2
R1598 GND.n2793 GND.n2792 467.2
R1599 GND.n2794 GND.n2793 467.2
R1600 GND.n2800 GND.n2799 467.2
R1601 GND.n2800 GND.n551 467.2
R1602 GND.n2820 GND.n2819 467.2
R1603 GND.n2820 GND.n522 467.2
R1604 GND.n2381 GND.n2380 467.2
R1605 GND.n2381 GND.n2331 467.2
R1606 GND.n2329 GND.n2328 467.2
R1607 GND.n2328 GND.n2327 467.2
R1608 GND.n2300 GND.n619 467.2
R1609 GND.n643 GND.n619 467.2
R1610 GND.n2284 GND.n2283 467.2
R1611 GND.n2284 GND.n2282 467.2
R1612 GND.n1997 GND.n1996 467.2
R1613 GND.n1997 GND.n879 467.2
R1614 GND.n2018 GND.n2017 467.2
R1615 GND.n2019 GND.n2018 467.2
R1616 GND.n2032 GND.n2031 467.2
R1617 GND.n2033 GND.n2032 467.2
R1618 GND.n2038 GND.n2037 467.2
R1619 GND.n2038 GND.n798 467.2
R1620 GND.n2058 GND.n2057 467.2
R1621 GND.n2058 GND.n769 467.2
R1622 GND.n1161 GND.n1160 467.2
R1623 GND.n1161 GND.n1159 467.2
R1624 GND.n1117 GND.n978 467.2
R1625 GND.n1110 GND.n978 467.2
R1626 GND.n1091 GND.n1090 467.2
R1627 GND.n1090 GND.n1089 467.2
R1628 GND.n3879 GND.n195 467.2
R1629 GND.n3487 GND.n195 467.2
R1630 GND.n3493 GND.n303 467.2
R1631 GND.n3506 GND.n303 467.2
R1632 GND.n3512 GND.n295 467.2
R1633 GND.n3528 GND.n295 467.2
R1634 GND.n3534 GND.n287 467.2
R1635 GND.n3550 GND.n287 467.2
R1636 GND.n3556 GND.n279 467.2
R1637 GND.n3569 GND.n279 467.2
R1638 GND.n3575 GND.n271 467.2
R1639 GND.n3589 GND.n271 467.2
R1640 GND.n3595 GND.n253 467.2
R1641 GND.n3608 GND.n253 467.2
R1642 GND.n3614 GND.n3613 467.2
R1643 GND.n3614 GND.n245 467.2
R1644 GND.n718 GND.n703 467.2
R1645 GND.n718 GND.n705 467.2
R1646 GND.n709 GND.n707 467.2
R1647 GND.n724 GND.n709 467.2
R1648 GND.n2179 GND.n651 467.2
R1649 GND.n2172 GND.n651 467.2
R1650 GND.n2167 GND.n655 467.2
R1651 GND.n2160 GND.n655 467.2
R1652 GND.n2136 GND.n668 467.2
R1653 GND.n2129 GND.n668 467.2
R1654 GND.n2214 GND.n2207 467.2
R1655 GND.n2220 GND.n2207 467.2
R1656 GND.n2225 GND.n2224 467.2
R1657 GND.n2225 GND.n2198 467.2
R1658 GND.n2249 GND.n2248 467.2
R1659 GND.n2249 GND.n647 467.2
R1660 GND.n2880 GND.n501 467.2
R1661 GND.n2873 GND.n501 467.2
R1662 GND.n2868 GND.n505 467.2
R1663 GND.n2861 GND.n505 467.2
R1664 GND.n2837 GND.n518 467.2
R1665 GND.n2830 GND.n518 467.2
R1666 GND.n3440 GND.n327 467.2
R1667 GND.n3446 GND.n327 467.2
R1668 GND.n3451 GND.n322 467.2
R1669 GND.n3457 GND.n322 467.2
R1670 GND.n2891 GND.n2890 467.2
R1671 GND.n2891 GND.n493 467.2
R1672 GND.n3892 GND.n190 467.2
R1673 GND.n3885 GND.n190 467.2
R1674 GND.n3405 GND.n3404 467.2
R1675 GND.n3405 GND.n3395 467.2
R1676 GND.n3429 GND.n332 467.2
R1677 GND.n3435 GND.n332 467.2
R1678 GND.n4365 GND.n7 467.2
R1679 GND.n3920 GND.n7 467.2
R1680 GND.n3925 GND.n3924 467.2
R1681 GND.n3925 GND.n3909 467.2
R1682 GND.n3949 GND.n3948 467.2
R1683 GND.n3949 GND.n184 467.2
R1684 GND.n2124 GND.n673 467.2
R1685 GND.n2117 GND.n673 467.2
R1686 GND.n2112 GND.n677 467.2
R1687 GND.n2105 GND.n677 467.2
R1688 GND.n761 GND.n760 467.2
R1689 GND.n761 GND.n726 467.2
R1690 GND.n2097 GND.n2096 467.2
R1691 GND.n2097 GND.n685 467.2
R1692 GND.n4327 GND.n20 467.2
R1693 GND.n4344 GND.n20 467.2
R1694 GND.n1947 GND.n1946 467.2
R1695 GND.n1946 GND.n1944 467.2
R1696 GND.n1897 GND.n1896 467.2
R1697 GND.n1896 GND.n1895 467.2
R1698 GND.n1936 GND.n1934 467.2
R1699 GND.n1936 GND.n1935 467.2
R1700 GND.n1966 GND.n1965 467.2
R1701 GND.n1967 GND.n1966 467.2
R1702 GND.n1919 GND.n1917 467.2
R1703 GND.n1919 GND.n1918 467.2
R1704 GND.n1913 GND.n1912 467.2
R1705 GND.n1943 GND.n1912 467.2
R1706 GND.n1681 GND.n1680 467.2
R1707 GND.n1680 GND.n1678 467.2
R1708 GND.n1645 GND.n1635 467.2
R1709 GND.n1645 GND.n1644 467.2
R1710 GND.n1734 GND.n1733 467.2
R1711 GND.n1733 GND.n1732 467.2
R1712 GND.n1702 GND.n1700 467.2
R1713 GND.n1721 GND.n1700 467.2
R1714 GND.n1719 GND.n1718 467.2
R1715 GND.n1718 GND.n1716 467.2
R1716 GND.n1676 GND.n1674 467.2
R1717 GND.n1677 GND.n1676 467.2
R1718 GND.n2423 GND.n2422 467.2
R1719 GND.n2422 GND.n2420 467.2
R1720 GND.n592 GND.n582 467.2
R1721 GND.n592 GND.n591 467.2
R1722 GND.n2476 GND.n2475 467.2
R1723 GND.n2475 GND.n2474 467.2
R1724 GND.n2444 GND.n2442 467.2
R1725 GND.n2463 GND.n2442 467.2
R1726 GND.n2461 GND.n2460 467.2
R1727 GND.n2460 GND.n2458 467.2
R1728 GND.n2418 GND.n2416 467.2
R1729 GND.n2419 GND.n2418 467.2
R1730 GND.n2693 GND.n2692 467.2
R1731 GND.n2692 GND.n2690 467.2
R1732 GND.n2643 GND.n2642 467.2
R1733 GND.n2642 GND.n2641 467.2
R1734 GND.n2682 GND.n2680 467.2
R1735 GND.n2682 GND.n2681 467.2
R1736 GND.n2712 GND.n2711 467.2
R1737 GND.n2713 GND.n2712 467.2
R1738 GND.n2665 GND.n2663 467.2
R1739 GND.n2665 GND.n2664 467.2
R1740 GND.n2659 GND.n2658 467.2
R1741 GND.n2689 GND.n2658 467.2
R1742 GND.n2977 GND.n2976 467.2
R1743 GND.n2976 GND.n2974 467.2
R1744 GND.n479 GND.n469 467.2
R1745 GND.n479 GND.n478 467.2
R1746 GND.n3030 GND.n3029 467.2
R1747 GND.n3029 GND.n3028 467.2
R1748 GND.n2998 GND.n2996 467.2
R1749 GND.n3017 GND.n2996 467.2
R1750 GND.n3015 GND.n3014 467.2
R1751 GND.n3014 GND.n3012 467.2
R1752 GND.n2972 GND.n2970 467.2
R1753 GND.n2973 GND.n2972 467.2
R1754 GND.n3234 GND.n3233 467.2
R1755 GND.n3233 GND.n3231 467.2
R1756 GND.n3199 GND.n3189 467.2
R1757 GND.n3199 GND.n3198 467.2
R1758 GND.n3287 GND.n3286 467.2
R1759 GND.n3286 GND.n3285 467.2
R1760 GND.n3255 GND.n3253 467.2
R1761 GND.n3274 GND.n3253 467.2
R1762 GND.n3272 GND.n3271 467.2
R1763 GND.n3271 GND.n3269 467.2
R1764 GND.n3229 GND.n3227 467.2
R1765 GND.n3230 GND.n3229 467.2
R1766 GND.n4157 GND.n4156 467.2
R1767 GND.n4156 GND.n4154 467.2
R1768 GND.n4121 GND.n4111 467.2
R1769 GND.n4121 GND.n4120 467.2
R1770 GND.n4210 GND.n4209 467.2
R1771 GND.n4209 GND.n4208 467.2
R1772 GND.n4178 GND.n4176 467.2
R1773 GND.n4197 GND.n4176 467.2
R1774 GND.n4195 GND.n4194 467.2
R1775 GND.n4194 GND.n4192 467.2
R1776 GND.n4152 GND.n4150 467.2
R1777 GND.n4153 GND.n4152 467.2
R1778 GND.n4243 GND.n4242 467.2
R1779 GND.n4244 GND.n4243 467.2
R1780 GND.t683 GND.n680 462.603
R1781 GND.t188 GND.n759 462.603
R1782 GND.n758 GND.t198 462.603
R1783 GND.n737 GND.t198 462.603
R1784 GND.t112 GND.n737 462.603
R1785 GND.n749 GND.t112 462.603
R1786 GND.n748 GND.t5 462.603
R1787 GND.t5 GND.n679 462.603
R1788 GND.n2103 GND.t256 462.603
R1789 GND.n2114 GND.t333 462.603
R1790 GND.n2115 GND.t4 462.603
R1791 GND.n2126 GND.t313 462.603
R1792 GND.n2127 GND.t185 462.603
R1793 GND.n2138 GND.t164 462.603
R1794 GND.t47 GND.n2142 462.603
R1795 GND.n2143 GND.t47 462.603
R1796 GND.n3448 GND.t286 462.603
R1797 GND.n3438 GND.t576 462.603
R1798 GND.n3437 GND.t701 462.603
R1799 GND.n3427 GND.t599 462.603
R1800 GND.n3426 GND.t231 462.603
R1801 GND.n3389 GND.t231 462.603
R1802 GND.t195 GND.n3389 462.603
R1803 GND.n3417 GND.t195 462.603
R1804 GND.n3416 GND.t178 462.603
R1805 GND.n3402 GND.t178 462.603
R1806 GND.t99 GND.n3403 462.603
R1807 GND.t331 GND.n192 462.603
R1808 GND.n3883 GND.t156 462.603
R1809 GND.n3894 GND.t282 462.603
R1810 GND.t259 GND.n3895 462.603
R1811 GND.t691 GND.n3947 462.603
R1812 GND.n3946 GND.t309 462.603
R1813 GND.n3903 GND.t309 462.603
R1814 GND.t76 GND.n3903 462.603
R1815 GND.n3937 GND.t76 462.603
R1816 GND.n3936 GND.t243 462.603
R1817 GND.n3914 GND.t243 462.603
R1818 GND.t150 GND.n3915 462.603
R1819 GND.t190 GND.n3923 462.603
R1820 GND.n3922 GND.t364 462.603
R1821 GND.n4363 GND.t102 462.603
R1822 GND.n1095 GND.n1094 424.125
R1823 GND.n2055 GND.n774 424.125
R1824 GND.n2014 GND.n817 424.125
R1825 GND.n2312 GND.n2311 424.125
R1826 GND.n2817 GND.n527 424.125
R1827 GND.n2916 GND.n2915 424.125
R1828 GND.n114 GND.n113 424.125
R1829 GND.n4297 GND.n4296 424.125
R1830 GND.n3471 GND.n3470 421.002
R1831 GND.n2798 GND.t171 416.356
R1832 GND.n3972 GND.n133 411.909
R1833 GND.n3343 GND.n3342 411.909
R1834 GND.n4325 GND.n4324 411.909
R1835 GND.n2035 GND.n803 411.909
R1836 GND.n2342 GND.n2341 411.909
R1837 GND.n1115 GND.t273 394.51
R1838 GND.t717 GND.n1993 394.51
R1839 GND.t581 GND.n1995 394.51
R1840 GND.t69 GND.n555 394.51
R1841 GND.t171 GND.n2797 394.51
R1842 GND.t177 GND.t710 388.161
R1843 GND.t723 GND.n2798 372.664
R1844 GND.t3 GND.t367 363.363
R1845 GND.t367 GND.t707 363.363
R1846 GND.t121 GND.t261 363.363
R1847 GND.n2102 GND.t333 357.123
R1848 GND.n4263 GND.n4262 351.625
R1849 GND.n4265 GND.n4263 351.625
R1850 GND.n4041 GND.n4002 351.625
R1851 GND.n4007 GND.n4002 351.625
R1852 GND.n4010 GND.n4009 351.625
R1853 GND.n4009 GND.n4003 351.625
R1854 GND.n422 GND.n407 351.625
R1855 GND.n410 GND.n407 351.625
R1856 GND.n415 GND.n411 351.625
R1857 GND.n411 GND.n406 351.625
R1858 GND.n3119 GND.n3080 351.625
R1859 GND.n3085 GND.n3080 351.625
R1860 GND.n3088 GND.n3087 351.625
R1861 GND.n3087 GND.n3081 351.625
R1862 GND.n2566 GND.n2527 351.625
R1863 GND.n2532 GND.n2527 351.625
R1864 GND.n2535 GND.n2534 351.625
R1865 GND.n2534 GND.n2528 351.625
R1866 GND.n1821 GND.n1782 351.625
R1867 GND.n1787 GND.n1782 351.625
R1868 GND.n1790 GND.n1789 351.625
R1869 GND.n1789 GND.n1783 351.625
R1870 GND.n1564 GND.n1525 351.625
R1871 GND.n1530 GND.n1525 351.625
R1872 GND.n1533 GND.n1532 351.625
R1873 GND.n1532 GND.n1526 351.625
R1874 GND.n1216 GND.n1177 351.625
R1875 GND.n1182 GND.n1177 351.625
R1876 GND.n1185 GND.n1184 351.625
R1877 GND.n1184 GND.n1178 351.625
R1878 GND.n1346 GND.n1307 351.625
R1879 GND.n1312 GND.n1307 351.625
R1880 GND.n1315 GND.n1314 351.625
R1881 GND.n1314 GND.n1308 351.625
R1882 GND.n1486 GND.n1430 351.625
R1883 GND.n1449 GND.n1430 351.625
R1884 GND.n1456 GND.n1455 351.625
R1885 GND.n1456 GND.n1431 351.625
R1886 GND.n1049 GND.n1047 351.625
R1887 GND.n1050 GND.n1049 351.625
R1888 GND.n4352 GND.n16 351.625
R1889 GND.n4338 GND.n16 351.625
R1890 GND.n4313 GND.n34 351.625
R1891 GND.n42 GND.n34 351.625
R1892 GND.n3982 GND.n3981 351.625
R1893 GND.n3982 GND.n117 351.625
R1894 GND.n2933 GND.n2932 351.625
R1895 GND.n2933 GND.n2919 351.625
R1896 GND.n2808 GND.n538 351.625
R1897 GND.n545 GND.n538 351.625
R1898 GND.n2370 GND.n2351 351.625
R1899 GND.n2377 GND.n2351 351.625
R1900 GND.n640 GND.n639 351.625
R1901 GND.n2279 GND.n639 351.625
R1902 GND.n2005 GND.n828 351.625
R1903 GND.n873 GND.n828 351.625
R1904 GND.n858 GND.n832 351.625
R1905 GND.n834 GND.n832 351.625
R1906 GND.n1132 GND.n1131 351.625
R1907 GND.n1156 GND.n1131 351.625
R1908 GND.n4302 GND.n38 351.625
R1909 GND.n175 GND.n38 351.625
R1910 GND.n146 GND.n144 351.625
R1911 GND.n170 GND.n144 351.625
R1912 GND.n109 GND.n108 351.625
R1913 GND.n109 GND.n104 351.625
R1914 GND.n3356 GND.n341 351.625
R1915 GND.n3369 GND.n341 351.625
R1916 GND.n2910 GND.n2909 351.625
R1917 GND.n2910 GND.n2905 351.625
R1918 GND.n2751 GND.n2749 351.625
R1919 GND.n2776 GND.n2749 351.625
R1920 GND.n2814 GND.n2813 351.625
R1921 GND.n2815 GND.n2814 351.625
R1922 GND.n2309 GND.n606 351.625
R1923 GND.n2322 GND.n606 351.625
R1924 GND.n2316 GND.n2315 351.625
R1925 GND.n2315 GND.n2314 351.625
R1926 GND.n2011 GND.n2010 351.625
R1927 GND.n2012 GND.n2011 351.625
R1928 GND.n792 GND.n785 351.625
R1929 GND.n2046 GND.n785 351.625
R1930 GND.n2052 GND.n2051 351.625
R1931 GND.n2053 GND.n2052 351.625
R1932 GND.n1076 GND.n987 351.625
R1933 GND.n1105 GND.n987 351.625
R1934 GND.n1099 GND.n1098 351.625
R1935 GND.n1098 GND.n1097 351.625
R1936 GND.n2239 GND.n2187 351.625
R1937 GND.n2244 GND.n2187 351.625
R1938 GND.n2849 GND.n513 351.625
R1939 GND.n2841 GND.n513 351.625
R1940 GND.n3468 GND.n311 351.625
R1941 GND.n2886 GND.n311 351.625
R1942 GND.n3419 GND.n3386 351.625
R1943 GND.n3424 GND.n3386 351.625
R1944 GND.n3939 GND.n3898 351.625
R1945 GND.n3944 GND.n3898 351.625
R1946 GND.n751 GND.n732 351.625
R1947 GND.n756 GND.n732 351.625
R1948 GND.n2140 GND.n663 351.625
R1949 GND.n2148 GND.n663 351.625
R1950 GND.n2086 GND.n2085 351.625
R1951 GND.n2086 GND.n691 351.625
R1952 GND.n1960 GND.n1904 351.625
R1953 GND.n1923 GND.n1904 351.625
R1954 GND.n1930 GND.n1929 351.625
R1955 GND.n1930 GND.n1905 351.625
R1956 GND.n1694 GND.n1655 351.625
R1957 GND.n1660 GND.n1655 351.625
R1958 GND.n1663 GND.n1662 351.625
R1959 GND.n1662 GND.n1656 351.625
R1960 GND.n2436 GND.n2397 351.625
R1961 GND.n2402 GND.n2397 351.625
R1962 GND.n2405 GND.n2404 351.625
R1963 GND.n2404 GND.n2398 351.625
R1964 GND.n2706 GND.n2650 351.625
R1965 GND.n2669 GND.n2650 351.625
R1966 GND.n2676 GND.n2675 351.625
R1967 GND.n2676 GND.n2651 351.625
R1968 GND.n2990 GND.n2951 351.625
R1969 GND.n2956 GND.n2951 351.625
R1970 GND.n2959 GND.n2958 351.625
R1971 GND.n2958 GND.n2952 351.625
R1972 GND.n3247 GND.n3208 351.625
R1973 GND.n3213 GND.n3208 351.625
R1974 GND.n3216 GND.n3215 351.625
R1975 GND.n3215 GND.n3209 351.625
R1976 GND.n4170 GND.n4131 351.625
R1977 GND.n4136 GND.n4131 351.625
R1978 GND.n4139 GND.n4138 351.625
R1979 GND.n4138 GND.n4132 351.625
R1980 GND.n1113 GND.t146 293.226
R1981 GND.n2146 GND.n2145 280.668
R1982 GND.n2158 GND.n2157 280.668
R1983 GND.n2170 GND.n2169 280.668
R1984 GND.n2247 GND.n2246 280.668
R1985 GND.n2237 GND.n2236 280.668
R1986 GND.n2202 GND.n2201 280.668
R1987 GND.n2223 GND.n2222 280.668
R1988 GND.n2843 GND.n2839 280.668
R1989 GND.n2847 GND.n2846 280.668
R1990 GND.n2859 GND.n2858 280.668
R1991 GND.n2871 GND.n2870 280.668
R1992 GND.n2889 GND.n2888 280.668
R1993 GND.n3470 GND.n308 280.668
R1994 GND.n3460 GND.n3459 280.668
R1995 GND.t339 GND.n268 241.806
R1996 GND.n3471 GND.t607 241.806
R1997 GND.n4251 GND.n4250 236.048
R1998 GND.n4253 GND.n4251 236.048
R1999 GND.n80 GND.n78 236.048
R2000 GND.n4071 GND.n80 236.048
R2001 GND.n61 GND.n59 236.048
R2002 GND.n4085 GND.n61 236.048
R2003 GND.n397 GND.n394 236.048
R2004 GND.n399 GND.n397 236.048
R2005 GND.n450 GND.n448 236.048
R2006 GND.n451 GND.n450 236.048
R2007 GND.n3065 GND.n3063 236.048
R2008 GND.n3149 GND.n3065 236.048
R2009 GND.n3046 GND.n3044 236.048
R2010 GND.n3163 GND.n3046 236.048
R2011 GND.n2511 GND.n2509 236.048
R2012 GND.n2596 GND.n2511 236.048
R2013 GND.n2492 GND.n2490 236.048
R2014 GND.n2610 GND.n2492 236.048
R2015 GND.n1768 GND.n1766 236.048
R2016 GND.n1851 GND.n1768 236.048
R2017 GND.n1750 GND.n1748 236.048
R2018 GND.n1865 GND.n1750 236.048
R2019 GND.n916 GND.n914 236.048
R2020 GND.n1594 GND.n916 236.048
R2021 GND.n897 GND.n895 236.048
R2022 GND.n1608 GND.n897 236.048
R2023 GND.n959 GND.n957 236.048
R2024 GND.n1246 GND.n959 236.048
R2025 GND.n940 GND.n938 236.048
R2026 GND.n1260 GND.n940 236.048
R2027 GND.n1291 GND.n1289 236.048
R2028 GND.n1376 GND.n1291 236.048
R2029 GND.n1272 GND.n1270 236.048
R2030 GND.n1390 GND.n1272 236.048
R2031 GND.n1416 GND.n1414 236.048
R2032 GND.n1496 GND.n1416 236.048
R2033 GND.n1464 GND.n935 236.048
R2034 GND.n1464 GND.n936 236.048
R2035 GND.n1003 GND.n1001 236.048
R2036 GND.n1066 GND.n1003 236.048
R2037 GND.n4334 GND.n25 236.048
R2038 GND.n26 GND.n25 236.048
R2039 GND.n2346 GND.n2339 236.048
R2040 GND.n2344 GND.n2339 236.048
R2041 GND.n628 GND.n627 236.048
R2042 GND.n2292 GND.n627 236.048
R2043 GND.n851 GND.n837 236.048
R2044 GND.n839 GND.n837 236.048
R2045 GND.n975 GND.n974 236.048
R2046 GND.n1169 GND.n974 236.048
R2047 GND.n4359 GND.n4358 236.048
R2048 GND.n4358 GND.n4357 236.048
R2049 GND.n151 GND.n149 236.048
R2050 GND.n163 GND.n149 236.048
R2051 GND.n3962 GND.n3961 236.048
R2052 GND.n3963 GND.n3962 236.048
R2053 GND.n351 GND.n350 236.048
R2054 GND.n3352 GND.n350 236.048
R2055 GND.n3374 GND.n335 236.048
R2056 GND.n3374 GND.n334 236.048
R2057 GND.n2757 GND.n2754 236.048
R2058 GND.n2769 GND.n2754 236.048
R2059 GND.n2786 GND.n2785 236.048
R2060 GND.n2787 GND.n2786 236.048
R2061 GND.n2363 GND.n2362 236.048
R2062 GND.n2362 GND.n2361 236.048
R2063 GND.n2271 GND.n2260 236.048
R2064 GND.n2260 GND.n2258 236.048
R2065 GND.n2025 GND.n2024 236.048
R2066 GND.n2026 GND.n2025 236.048
R2067 GND.n1148 GND.n1137 236.048
R2068 GND.n1137 GND.n1135 236.048
R2069 GND.n2155 GND.n659 236.048
R2070 GND.n660 GND.n659 236.048
R2071 GND.n2196 GND.n2195 236.048
R2072 GND.n2234 GND.n2195 236.048
R2073 GND.n2856 GND.n509 236.048
R2074 GND.n510 GND.n509 236.048
R2075 GND.n3462 GND.n317 236.048
R2076 GND.n317 GND.n315 236.048
R2077 GND.n3393 GND.n3392 236.048
R2078 GND.n3414 GND.n3392 236.048
R2079 GND.n3907 GND.n3906 236.048
R2080 GND.n3934 GND.n3906 236.048
R2081 GND.n742 GND.n740 236.048
R2082 GND.n746 GND.n740 236.048
R2083 GND.n700 GND.n699 236.048
R2084 GND.n2081 GND.n699 236.048
R2085 GND.n1890 GND.n1888 236.048
R2086 GND.n1970 GND.n1890 236.048
R2087 GND.n1938 GND.n892 236.048
R2088 GND.n1938 GND.n893 236.048
R2089 GND.n1640 GND.n1638 236.048
R2090 GND.n1724 GND.n1640 236.048
R2091 GND.n1621 GND.n1619 236.048
R2092 GND.n1738 GND.n1621 236.048
R2093 GND.n587 GND.n585 236.048
R2094 GND.n2466 GND.n587 236.048
R2095 GND.n568 GND.n566 236.048
R2096 GND.n2480 GND.n568 236.048
R2097 GND.n2636 GND.n2634 236.048
R2098 GND.n2716 GND.n2636 236.048
R2099 GND.n2684 GND.n563 236.048
R2100 GND.n2684 GND.n564 236.048
R2101 GND.n474 GND.n472 236.048
R2102 GND.n3020 GND.n474 236.048
R2103 GND.n455 GND.n453 236.048
R2104 GND.n3034 GND.n455 236.048
R2105 GND.n3194 GND.n3192 236.048
R2106 GND.n3277 GND.n3194 236.048
R2107 GND.n3176 GND.n3174 236.048
R2108 GND.n3291 GND.n3176 236.048
R2109 GND.n4116 GND.n4114 236.048
R2110 GND.n4200 GND.n4116 236.048
R2111 GND.n4097 GND.n4095 236.048
R2112 GND.n4214 GND.n4097 236.048
R2113 GND.n3449 GND.n3448 226.542
R2114 GND.n2099 GND.t299 214.944
R2115 GND.n1095 GND.n1093 210.605
R2116 GND.n1146 GND.n1145 210.605
R2117 GND.n2056 GND.n2055 210.605
R2118 GND.n2036 GND.n2035 210.605
R2119 GND.n2022 GND.n2021 210.605
R2120 GND.n2015 GND.n2014 210.605
R2121 GND.n2269 GND.n2268 210.605
R2122 GND.n2312 GND.n614 210.605
R2123 GND.n2341 GND.n2340 210.605
R2124 GND.n2357 GND.n2356 210.605
R2125 GND.n2818 GND.n2817 210.605
R2126 GND.n2783 GND.n2782 210.605
R2127 GND.n2915 GND.n2914 210.605
R2128 GND.n3343 GND.n3340 210.605
R2129 GND.n3373 GND.n3372 210.605
R2130 GND.n113 GND.n112 210.605
R2131 GND.n3973 GND.n3972 210.605
R2132 GND.n4289 GND.n48 210.605
R2133 GND.n4296 GND.n4295 210.605
R2134 GND.n4325 GND.n4322 210.605
R2135 GND.n1172 GND.n971 203.037
R2136 GND.n2295 GND.n624 203.037
R2137 GND.n2796 GND.n486 203.037
R2138 GND.t180 GND.n133 201.528
R2139 GND.t596 GND.n165 201.528
R2140 GND.t342 GND.n3965 201.528
R2141 GND.n3342 GND.t302 201.528
R2142 GND.t107 GND.n3354 201.528
R2143 GND.t358 GND.n338 201.528
R2144 GND.n2755 GND.t265 201.528
R2145 GND.t568 GND.n2771 201.528
R2146 GND.t680 GND.n2789 201.528
R2147 GND.n4324 GND.t365 201.528
R2148 GND.t570 GND.n4336 201.528
R2149 GND.n4355 GND.t615 201.528
R2150 GND.n4354 GND.t252 201.528
R2151 GND.n1171 GND.t264 201.528
R2152 GND.t251 GND.n1128 201.528
R2153 GND.n1142 GND.t642 201.528
R2154 GND.t639 GND.n803 201.528
R2155 GND.t110 GND.n853 201.528
R2156 GND.t217 GND.n2028 201.528
R2157 GND.n2294 GND.t579 201.528
R2158 GND.t569 GND.n636 201.528
R2159 GND.n2265 GND.t125 201.528
R2160 GND.n2342 GND.t304 201.528
R2161 GND.t250 GND.n2348 201.528
R2162 GND.n2355 GND.t350 201.528
R2163 GND.n759 GND.n758 195.891
R2164 GND.n749 GND.n748 195.891
R2165 GND.n2103 GND.n679 195.891
R2166 GND.n2115 GND.n2114 195.891
R2167 GND.n2142 GND.n2138 195.891
R2168 GND.n3427 GND.n3426 195.891
R2169 GND.n3417 GND.n3416 195.891
R2170 GND.n3403 GND.n3402 195.891
R2171 GND.n3883 GND.n192 195.891
R2172 GND.n3947 GND.n3946 195.891
R2173 GND.n3937 GND.n3936 195.891
R2174 GND.n3915 GND.n3914 195.891
R2175 GND.n3923 GND.n3922 195.891
R2176 GND.n1086 GND.t299 194.081
R2177 GND.n695 GND.t710 194.081
R2178 GND.t137 GND.n696 194.081
R2179 GND.n2088 GND.t137 194.081
R2180 GND.n2088 GND.t144 194.081
R2181 GND.t144 GND.n2084 194.081
R2182 GND.n2083 GND.t262 194.081
R2183 GND.n712 GND.t262 192.101
R2184 GND.t320 GND.n802 187.923
R2185 GND.n2392 GND.t54 187.923
R2186 GND.n3333 GND.t605 187.923
R2187 GND.n3997 GND.t153 187.923
R2188 GND.t45 GND.n10 187.923
R2189 GND.n716 GND.t707 181.681
R2190 GND.n715 GND.t261 181.681
R2191 GND.n3475 GND.t712 176.673
R2192 GND.n3497 GND.t702 176.673
R2193 GND.n3519 GND.t659 176.673
R2194 GND.n3538 GND.t614 176.673
R2195 GND.n3560 GND.t566 176.673
R2196 GND.n3579 GND.t221 176.673
R2197 GND.n3599 GND.t686 176.673
R2198 GND.n256 GND.t718 176.673
R2199 GND.t11 GND.n139 174.317
R2200 GND.t248 GND.n3371 174.317
R2201 GND.t13 GND.n2744 174.317
R2202 GND.t17 GND.n1144 174.317
R2203 GND.t15 GND.n809 174.317
R2204 GND.t597 GND.n2267 174.317
R2205 GND.n2368 GND.t108 174.317
R2206 GND.n2099 GND.t177 173.219
R2207 GND.n4226 GND.n56 173.012
R2208 GND.n4284 GND.n4283 173.012
R2209 GND.n4278 GND.n4230 173.012
R2210 GND.n4234 GND.n4231 173.012
R2211 GND.n4254 GND.n4250 173.012
R2212 GND.n4254 GND.n4253 173.012
R2213 GND.n4262 GND.n4260 173.012
R2214 GND.n4266 GND.n4265 173.012
R2215 GND.n4072 GND.n78 173.012
R2216 GND.n4072 GND.n4071 173.012
R2217 GND.n4086 GND.n59 173.012
R2218 GND.n4086 GND.n4085 173.012
R2219 GND.n400 GND.n394 173.012
R2220 GND.n400 GND.n399 173.012
R2221 GND.n3317 GND.n448 173.012
R2222 GND.n3317 GND.n451 173.012
R2223 GND.n3150 GND.n3063 173.012
R2224 GND.n3150 GND.n3149 173.012
R2225 GND.n3164 GND.n3044 173.012
R2226 GND.n3164 GND.n3163 173.012
R2227 GND.n2597 GND.n2509 173.012
R2228 GND.n2597 GND.n2596 173.012
R2229 GND.n2611 GND.n2490 173.012
R2230 GND.n2611 GND.n2610 173.012
R2231 GND.n1852 GND.n1766 173.012
R2232 GND.n1852 GND.n1851 173.012
R2233 GND.n1866 GND.n1748 173.012
R2234 GND.n1866 GND.n1865 173.012
R2235 GND.n1595 GND.n914 173.012
R2236 GND.n1595 GND.n1594 173.012
R2237 GND.n1609 GND.n895 173.012
R2238 GND.n1609 GND.n1608 173.012
R2239 GND.n1247 GND.n957 173.012
R2240 GND.n1247 GND.n1246 173.012
R2241 GND.n1261 GND.n938 173.012
R2242 GND.n1261 GND.n1260 173.012
R2243 GND.n1377 GND.n1289 173.012
R2244 GND.n1377 GND.n1376 173.012
R2245 GND.n1391 GND.n1270 173.012
R2246 GND.n1391 GND.n1390 173.012
R2247 GND.n1497 GND.n1414 173.012
R2248 GND.n1497 GND.n1496 173.012
R2249 GND.n1516 GND.n935 173.012
R2250 GND.n1516 GND.n936 173.012
R2251 GND.n1054 GND.n1047 173.012
R2252 GND.n1051 GND.n1050 173.012
R2253 GND.n1062 GND.n1014 173.012
R2254 GND.n1060 GND.n1059 173.012
R2255 GND.n1023 GND.n1022 173.012
R2256 GND.n1027 GND.n1026 173.012
R2257 GND.n1067 GND.n1001 173.012
R2258 GND.n1067 GND.n1066 173.012
R2259 GND.n1042 GND.n1034 173.012
R2260 GND.n1039 GND.n1037 173.012
R2261 GND.n4352 GND.n4351 173.012
R2262 GND.n4338 GND.n4337 173.012
R2263 GND.n4334 GND.n4333 173.012
R2264 GND.n4333 GND.n26 173.012
R2265 GND.n4313 GND.n4312 173.012
R2266 GND.n42 GND.n41 173.012
R2267 GND.n3981 GND.n3980 173.012
R2268 GND.n119 GND.n117 173.012
R2269 GND.n2932 GND.n2931 173.012
R2270 GND.n2921 GND.n2919 173.012
R2271 GND.n2808 GND.n2807 173.012
R2272 GND.n546 GND.n545 173.012
R2273 GND.n2371 GND.n2370 173.012
R2274 GND.n2377 GND.n2376 173.012
R2275 GND.n2346 GND.n2345 173.012
R2276 GND.n2345 GND.n2344 173.012
R2277 GND.n2276 GND.n640 173.012
R2278 GND.n2279 GND.n2278 173.012
R2279 GND.n2291 GND.n628 173.012
R2280 GND.n2292 GND.n2291 173.012
R2281 GND.n2005 GND.n2004 173.012
R2282 GND.n874 GND.n873 173.012
R2283 GND.n859 GND.n858 173.012
R2284 GND.n844 GND.n834 173.012
R2285 GND.n851 GND.n850 173.012
R2286 GND.n850 GND.n839 173.012
R2287 GND.n1153 GND.n1132 173.012
R2288 GND.n1156 GND.n1155 173.012
R2289 GND.n1168 GND.n975 173.012
R2290 GND.n1169 GND.n1168 173.012
R2291 GND.n4359 GND.n13 173.012
R2292 GND.n4357 GND.n13 173.012
R2293 GND.n4320 GND.n29 173.012
R2294 GND.n4318 GND.n30 173.012
R2295 GND.n4303 GND.n4302 173.012
R2296 GND.n176 GND.n175 173.012
R2297 GND.n4293 GND.n46 173.012
R2298 GND.n4291 GND.n47 173.012
R2299 GND.n156 GND.n146 173.012
R2300 GND.n171 GND.n170 173.012
R2301 GND.n162 GND.n151 173.012
R2302 GND.n163 GND.n162 173.012
R2303 GND.n3963 GND.n3959 173.012
R2304 GND.n3961 GND.n3959 173.012
R2305 GND.n3968 GND.n137 173.012
R2306 GND.n3970 GND.n136 173.012
R2307 GND.n132 GND.n125 173.012
R2308 GND.n3977 GND.n124 173.012
R2309 GND.n108 GND.n105 173.012
R2310 GND.n3988 GND.n104 173.012
R2311 GND.n3992 GND.n102 173.012
R2312 GND.n100 GND.n98 173.012
R2313 GND.n3356 GND.n3355 173.012
R2314 GND.n3369 GND.n3368 173.012
R2315 GND.n3351 GND.n351 173.012
R2316 GND.n3352 GND.n3351 173.012
R2317 GND.n3377 GND.n334 173.012
R2318 GND.n3377 GND.n335 173.012
R2319 GND.n3363 GND.n3362 173.012
R2320 GND.n3346 GND.n3345 173.012
R2321 GND.n3338 GND.n354 173.012
R2322 GND.n3336 GND.n355 173.012
R2323 GND.n2909 GND.n2906 173.012
R2324 GND.n2939 GND.n2905 173.012
R2325 GND.n2943 GND.n2903 173.012
R2326 GND.n2901 GND.n490 173.012
R2327 GND.n2762 GND.n2751 173.012
R2328 GND.n2777 GND.n2776 173.012
R2329 GND.n2768 GND.n2757 173.012
R2330 GND.n2769 GND.n2768 173.012
R2331 GND.n2787 GND.n2781 173.012
R2332 GND.n2785 GND.n2781 173.012
R2333 GND.n2792 GND.n2742 173.012
R2334 GND.n2794 GND.n2741 173.012
R2335 GND.n2799 GND.n552 173.012
R2336 GND.n2804 GND.n551 173.012
R2337 GND.n2813 GND.n532 173.012
R2338 GND.n2815 GND.n530 173.012
R2339 GND.n2819 GND.n523 173.012
R2340 GND.n2824 GND.n522 173.012
R2341 GND.n2366 GND.n2363 173.012
R2342 GND.n2366 GND.n2361 173.012
R2343 GND.n2380 GND.n2334 173.012
R2344 GND.n2385 GND.n2331 173.012
R2345 GND.n2389 GND.n2329 173.012
R2346 GND.n2327 GND.n603 173.012
R2347 GND.n2309 GND.n2308 173.012
R2348 GND.n2323 GND.n2322 173.012
R2349 GND.n2316 GND.n611 173.012
R2350 GND.n2314 GND.n613 173.012
R2351 GND.n2301 GND.n2300 173.012
R2352 GND.n644 GND.n643 173.012
R2353 GND.n2272 GND.n2271 173.012
R2354 GND.n2272 GND.n2258 173.012
R2355 GND.n2283 GND.n632 173.012
R2356 GND.n2282 GND.n631 173.012
R2357 GND.n1996 GND.n882 173.012
R2358 GND.n2001 GND.n879 173.012
R2359 GND.n2010 GND.n822 173.012
R2360 GND.n2012 GND.n820 173.012
R2361 GND.n2017 GND.n816 173.012
R2362 GND.n2019 GND.n815 173.012
R2363 GND.n2024 GND.n812 173.012
R2364 GND.n2026 GND.n812 173.012
R2365 GND.n2031 GND.n807 173.012
R2366 GND.n2033 GND.n806 173.012
R2367 GND.n2037 GND.n799 173.012
R2368 GND.n2042 GND.n798 173.012
R2369 GND.n793 GND.n792 173.012
R2370 GND.n2046 GND.n2045 173.012
R2371 GND.n2051 GND.n779 173.012
R2372 GND.n2053 GND.n777 173.012
R2373 GND.n2057 GND.n770 173.012
R2374 GND.n2062 GND.n769 173.012
R2375 GND.n1149 GND.n1148 173.012
R2376 GND.n1149 GND.n1135 173.012
R2377 GND.n1160 GND.n1124 173.012
R2378 GND.n1159 GND.n1123 173.012
R2379 GND.n1118 GND.n1117 173.012
R2380 GND.n1110 GND.n1109 173.012
R2381 GND.n1077 GND.n1076 173.012
R2382 GND.n1106 GND.n1105 173.012
R2383 GND.n1099 GND.n993 173.012
R2384 GND.n1097 GND.n995 173.012
R2385 GND.n1091 GND.n998 173.012
R2386 GND.n1089 GND.n1085 173.012
R2387 GND.n3879 GND.n3878 173.012
R2388 GND.n3487 GND.n3486 173.012
R2389 GND.n3494 GND.n3493 173.012
R2390 GND.n3506 GND.n3505 173.012
R2391 GND.n3513 GND.n3512 173.012
R2392 GND.n3528 GND.n3527 173.012
R2393 GND.n3535 GND.n3534 173.012
R2394 GND.n3550 GND.n3549 173.012
R2395 GND.n3557 GND.n3556 173.012
R2396 GND.n3569 GND.n3568 173.012
R2397 GND.n3576 GND.n3575 173.012
R2398 GND.n3589 GND.n3588 173.012
R2399 GND.n3596 GND.n3595 173.012
R2400 GND.n3608 GND.n3607 173.012
R2401 GND.n3613 GND.n247 173.012
R2402 GND.n3618 GND.n245 173.012
R2403 GND.n2076 GND.n703 173.012
R2404 GND.n2074 GND.n705 173.012
R2405 GND.n2070 GND.n707 173.012
R2406 GND.n2068 GND.n724 173.012
R2407 GND.n2179 GND.n2178 173.012
R2408 GND.n2173 GND.n2172 173.012
R2409 GND.n2167 GND.n2166 173.012
R2410 GND.n2161 GND.n2160 173.012
R2411 GND.n2155 GND.n2154 173.012
R2412 GND.n2154 GND.n660 173.012
R2413 GND.n2136 GND.n2135 173.012
R2414 GND.n2130 GND.n2129 173.012
R2415 GND.n2215 GND.n2214 173.012
R2416 GND.n2220 GND.n2219 173.012
R2417 GND.n2224 GND.n2199 173.012
R2418 GND.n2229 GND.n2198 173.012
R2419 GND.n2233 GND.n2196 173.012
R2420 GND.n2234 GND.n2233 173.012
R2421 GND.n2240 GND.n2239 173.012
R2422 GND.n2244 GND.n2243 173.012
R2423 GND.n2248 GND.n648 173.012
R2424 GND.n2253 GND.n647 173.012
R2425 GND.n2880 GND.n2879 173.012
R2426 GND.n2874 GND.n2873 173.012
R2427 GND.n2868 GND.n2867 173.012
R2428 GND.n2862 GND.n2861 173.012
R2429 GND.n2856 GND.n2855 173.012
R2430 GND.n2855 GND.n510 173.012
R2431 GND.n2850 GND.n2849 173.012
R2432 GND.n2841 GND.n2840 173.012
R2433 GND.n2837 GND.n2836 173.012
R2434 GND.n2831 GND.n2830 173.012
R2435 GND.n3441 GND.n3440 173.012
R2436 GND.n3446 GND.n3445 173.012
R2437 GND.n3452 GND.n3451 173.012
R2438 GND.n3457 GND.n3456 173.012
R2439 GND.n3463 GND.n3462 173.012
R2440 GND.n3463 GND.n315 173.012
R2441 GND.n3468 GND.n3467 173.012
R2442 GND.n2886 GND.n2885 173.012
R2443 GND.n2890 GND.n496 173.012
R2444 GND.n2895 GND.n493 173.012
R2445 GND.n3892 GND.n3891 173.012
R2446 GND.n3886 GND.n3885 173.012
R2447 GND.n3404 GND.n3398 173.012
R2448 GND.n3409 GND.n3395 173.012
R2449 GND.n3413 GND.n3393 173.012
R2450 GND.n3414 GND.n3413 173.012
R2451 GND.n3420 GND.n3419 173.012
R2452 GND.n3424 GND.n3423 173.012
R2453 GND.n3430 GND.n3429 173.012
R2454 GND.n3435 GND.n3434 173.012
R2455 GND.n4366 GND.n4365 173.012
R2456 GND.n3920 GND.n3919 173.012
R2457 GND.n3924 GND.n3910 173.012
R2458 GND.n3929 GND.n3909 173.012
R2459 GND.n3933 GND.n3907 173.012
R2460 GND.n3934 GND.n3933 173.012
R2461 GND.n3940 GND.n3939 173.012
R2462 GND.n3944 GND.n3943 173.012
R2463 GND.n3948 GND.n185 173.012
R2464 GND.n3953 GND.n184 173.012
R2465 GND.n2124 GND.n2123 173.012
R2466 GND.n2118 GND.n2117 173.012
R2467 GND.n2112 GND.n2111 173.012
R2468 GND.n2106 GND.n2105 173.012
R2469 GND.n745 GND.n742 173.012
R2470 GND.n746 GND.n745 173.012
R2471 GND.n752 GND.n751 173.012
R2472 GND.n756 GND.n755 173.012
R2473 GND.n760 GND.n727 173.012
R2474 GND.n765 GND.n726 173.012
R2475 GND.n2140 GND.n2139 173.012
R2476 GND.n2149 GND.n2148 173.012
R2477 GND.n2080 GND.n700 173.012
R2478 GND.n2081 GND.n2080 173.012
R2479 GND.n2085 GND.n692 173.012
R2480 GND.n2091 GND.n691 173.012
R2481 GND.n2096 GND.n2095 173.012
R2482 GND.n687 GND.n685 173.012
R2483 GND.n4345 GND.n4344 173.012
R2484 GND.n4328 GND.n4327 173.012
R2485 GND.n1971 GND.n1888 173.012
R2486 GND.n1971 GND.n1970 173.012
R2487 GND.n1990 GND.n892 173.012
R2488 GND.n1990 GND.n893 173.012
R2489 GND.n1725 GND.n1638 173.012
R2490 GND.n1725 GND.n1724 173.012
R2491 GND.n1739 GND.n1619 173.012
R2492 GND.n1739 GND.n1738 173.012
R2493 GND.n2467 GND.n585 173.012
R2494 GND.n2467 GND.n2466 173.012
R2495 GND.n2481 GND.n566 173.012
R2496 GND.n2481 GND.n2480 173.012
R2497 GND.n2717 GND.n2634 173.012
R2498 GND.n2717 GND.n2716 173.012
R2499 GND.n2736 GND.n563 173.012
R2500 GND.n2736 GND.n564 173.012
R2501 GND.n3021 GND.n472 173.012
R2502 GND.n3021 GND.n3020 173.012
R2503 GND.n3035 GND.n453 173.012
R2504 GND.n3035 GND.n3034 173.012
R2505 GND.n3278 GND.n3192 173.012
R2506 GND.n3278 GND.n3277 173.012
R2507 GND.n3292 GND.n3174 173.012
R2508 GND.n3292 GND.n3291 173.012
R2509 GND.n4201 GND.n4114 173.012
R2510 GND.n4201 GND.n4200 173.012
R2511 GND.n4215 GND.n4095 173.012
R2512 GND.n4215 GND.n4214 173.012
R2513 GND.n4242 GND.n4241 173.012
R2514 GND.n4245 GND.n4244 173.012
R2515 GND.t37 GND.n82 169.232
R2516 GND.t37 GND.n3999 169.232
R2517 GND.t138 GND.n63 169.232
R2518 GND.t138 GND.n69 169.232
R2519 GND.t43 GND.n3067 169.232
R2520 GND.t43 GND.n3077 169.232
R2521 GND.t62 GND.n3048 169.232
R2522 GND.t62 GND.n3054 169.232
R2523 GND.t25 GND.n2513 169.232
R2524 GND.t25 GND.n2524 169.232
R2525 GND.t50 GND.n2494 169.232
R2526 GND.t50 GND.n2500 169.232
R2527 GND.t21 GND.n1770 169.232
R2528 GND.t21 GND.n622 169.232
R2529 GND.t22 GND.n623 169.232
R2530 GND.t22 GND.n1757 169.232
R2531 GND.t55 GND.n918 169.232
R2532 GND.t55 GND.n1522 169.232
R2533 GND.t40 GND.n899 169.232
R2534 GND.t40 GND.n905 169.232
R2535 GND.t95 GND.n961 169.232
R2536 GND.t95 GND.n1174 169.232
R2537 GND.t84 GND.n942 169.232
R2538 GND.t84 GND.n948 169.232
R2539 GND.t90 GND.n1293 169.232
R2540 GND.t90 GND.n1304 169.232
R2541 GND.t149 GND.n1274 169.232
R2542 GND.t149 GND.n1280 169.232
R2543 GND.t70 GND.n1418 169.232
R2544 GND.t70 GND.n928 169.232
R2545 GND.n1518 GND.t28 169.232
R2546 GND.n1466 GND.t28 169.232
R2547 GND.t41 GND.n1892 169.232
R2548 GND.t41 GND.n885 169.232
R2549 GND.n1992 GND.t83 169.232
R2550 GND.n1940 GND.t83 169.232
R2551 GND.t140 GND.n1642 169.232
R2552 GND.t140 GND.n1652 169.232
R2553 GND.t30 GND.n1623 169.232
R2554 GND.t30 GND.n1629 169.232
R2555 GND.t73 GND.n589 169.232
R2556 GND.t73 GND.n2394 169.232
R2557 GND.t8 GND.n570 169.232
R2558 GND.t8 GND.n576 169.232
R2559 GND.t44 GND.n2638 169.232
R2560 GND.t44 GND.n556 169.232
R2561 GND.n2738 GND.t32 169.232
R2562 GND.n2686 GND.t32 169.232
R2563 GND.t7 GND.n476 169.232
R2564 GND.t7 GND.n2948 169.232
R2565 GND.t39 GND.n457 169.232
R2566 GND.t39 GND.n463 169.232
R2567 GND.t24 GND.n3196 169.232
R2568 GND.t24 GND.n92 169.232
R2569 GND.t36 GND.n93 169.232
R2570 GND.t36 GND.n3183 169.232
R2571 GND.t75 GND.n4118 169.232
R2572 GND.t75 GND.n4128 169.232
R2573 GND.t53 GND.n4099 169.232
R2574 GND.t53 GND.n4105 169.232
R2575 GND.n1115 GND.n971 167.056
R2576 GND.n1995 GND.n624 167.056
R2577 GND.n2797 GND.n2796 167.056
R2578 GND.n3882 GND.t282 161.233
R2579 GND.t58 GND.n983 156.579
R2580 GND.t58 GND.n981 156.579
R2581 GND.n3332 GND.t92 156.579
R2582 GND.n385 GND.t92 156.579
R2583 GND.n3319 GND.t9 156.579
R2584 GND.t9 GND.n94 156.579
R2585 GND.n4287 GND.t88 156.579
R2586 GND.n4275 GND.t88 156.579
R2587 GND.n2755 GND.n486 155.944
R2588 GND.n1172 GND.n1171 155.944
R2589 GND.n2007 GND.n823 155.944
R2590 GND.n2295 GND.n2294 155.944
R2591 GND.n2810 GND.n533 155.944
R2592 GND.n4029 GND.n4028 150.213
R2593 GND.n4025 GND.n4019 150.213
R2594 GND.n4041 GND.n4040 150.213
R2595 GND.n4011 GND.n4007 150.213
R2596 GND.n4011 GND.n4010 150.213
R2597 GND.n4040 GND.n4003 150.213
R2598 GND.n4078 GND.n75 150.213
R2599 GND.n84 GND.n74 150.213
R2600 GND.n4081 GND.n74 150.213
R2601 GND.n4079 GND.n4078 150.213
R2602 GND.n4062 GND.n4049 150.213
R2603 GND.n4068 GND.n4067 150.213
R2604 GND.n4067 GND.n4066 150.213
R2605 GND.n4063 GND.n4062 150.213
R2606 GND.n4021 GND.n4019 150.213
R2607 GND.n4029 GND.n4024 150.213
R2608 GND.n441 GND.n440 150.213
R2609 GND.n435 GND.n434 150.213
R2610 GND.n423 GND.n422 150.213
R2611 GND.n416 GND.n410 150.213
R2612 GND.n416 GND.n415 150.213
R2613 GND.n423 GND.n406 150.213
R2614 GND.n379 GND.n378 150.213
R2615 GND.n375 GND.n369 150.213
R2616 GND.n380 GND.n369 150.213
R2617 GND.n382 GND.n379 150.213
R2618 GND.n3329 GND.n3328 150.213
R2619 GND.n3311 GND.n364 150.213
R2620 GND.n3311 GND.n3310 150.213
R2621 GND.n3328 GND.n365 150.213
R2622 GND.n436 GND.n435 150.213
R2623 GND.n440 GND.n439 150.213
R2624 GND.n3107 GND.n3106 150.213
R2625 GND.n3103 GND.n3097 150.213
R2626 GND.n3119 GND.n3118 150.213
R2627 GND.n3089 GND.n3085 150.213
R2628 GND.n3089 GND.n3088 150.213
R2629 GND.n3118 GND.n3081 150.213
R2630 GND.n3156 GND.n3060 150.213
R2631 GND.n3069 GND.n3059 150.213
R2632 GND.n3159 GND.n3059 150.213
R2633 GND.n3157 GND.n3156 150.213
R2634 GND.n3140 GND.n3127 150.213
R2635 GND.n3146 GND.n3145 150.213
R2636 GND.n3145 GND.n3144 150.213
R2637 GND.n3141 GND.n3140 150.213
R2638 GND.n3099 GND.n3097 150.213
R2639 GND.n3107 GND.n3102 150.213
R2640 GND.n2554 GND.n2553 150.213
R2641 GND.n2550 GND.n2544 150.213
R2642 GND.n2566 GND.n2565 150.213
R2643 GND.n2536 GND.n2532 150.213
R2644 GND.n2536 GND.n2535 150.213
R2645 GND.n2565 GND.n2528 150.213
R2646 GND.n2603 GND.n2506 150.213
R2647 GND.n2515 GND.n2505 150.213
R2648 GND.n2606 GND.n2505 150.213
R2649 GND.n2604 GND.n2603 150.213
R2650 GND.n2587 GND.n2574 150.213
R2651 GND.n2593 GND.n2592 150.213
R2652 GND.n2592 GND.n2591 150.213
R2653 GND.n2588 GND.n2587 150.213
R2654 GND.n2546 GND.n2544 150.213
R2655 GND.n2554 GND.n2549 150.213
R2656 GND.n1809 GND.n1808 150.213
R2657 GND.n1805 GND.n1799 150.213
R2658 GND.n1821 GND.n1820 150.213
R2659 GND.n1791 GND.n1787 150.213
R2660 GND.n1791 GND.n1790 150.213
R2661 GND.n1820 GND.n1783 150.213
R2662 GND.n1858 GND.n1763 150.213
R2663 GND.n1772 GND.n1762 150.213
R2664 GND.n1861 GND.n1762 150.213
R2665 GND.n1859 GND.n1858 150.213
R2666 GND.n1842 GND.n1829 150.213
R2667 GND.n1848 GND.n1847 150.213
R2668 GND.n1847 GND.n1846 150.213
R2669 GND.n1843 GND.n1842 150.213
R2670 GND.n1801 GND.n1799 150.213
R2671 GND.n1809 GND.n1804 150.213
R2672 GND.n1552 GND.n1551 150.213
R2673 GND.n1548 GND.n1542 150.213
R2674 GND.n1564 GND.n1563 150.213
R2675 GND.n1534 GND.n1530 150.213
R2676 GND.n1534 GND.n1533 150.213
R2677 GND.n1563 GND.n1526 150.213
R2678 GND.n1601 GND.n911 150.213
R2679 GND.n920 GND.n910 150.213
R2680 GND.n1604 GND.n910 150.213
R2681 GND.n1602 GND.n1601 150.213
R2682 GND.n1585 GND.n1572 150.213
R2683 GND.n1591 GND.n1590 150.213
R2684 GND.n1590 GND.n1589 150.213
R2685 GND.n1586 GND.n1585 150.213
R2686 GND.n1544 GND.n1542 150.213
R2687 GND.n1552 GND.n1547 150.213
R2688 GND.n1204 GND.n1203 150.213
R2689 GND.n1200 GND.n1194 150.213
R2690 GND.n1216 GND.n1215 150.213
R2691 GND.n1186 GND.n1182 150.213
R2692 GND.n1186 GND.n1185 150.213
R2693 GND.n1215 GND.n1178 150.213
R2694 GND.n1253 GND.n954 150.213
R2695 GND.n963 GND.n953 150.213
R2696 GND.n1256 GND.n953 150.213
R2697 GND.n1254 GND.n1253 150.213
R2698 GND.n1237 GND.n1224 150.213
R2699 GND.n1243 GND.n1242 150.213
R2700 GND.n1242 GND.n1241 150.213
R2701 GND.n1238 GND.n1237 150.213
R2702 GND.n1196 GND.n1194 150.213
R2703 GND.n1204 GND.n1199 150.213
R2704 GND.n1334 GND.n1333 150.213
R2705 GND.n1330 GND.n1324 150.213
R2706 GND.n1346 GND.n1345 150.213
R2707 GND.n1316 GND.n1312 150.213
R2708 GND.n1316 GND.n1315 150.213
R2709 GND.n1345 GND.n1308 150.213
R2710 GND.n1383 GND.n1286 150.213
R2711 GND.n1295 GND.n1285 150.213
R2712 GND.n1386 GND.n1285 150.213
R2713 GND.n1384 GND.n1383 150.213
R2714 GND.n1367 GND.n1354 150.213
R2715 GND.n1373 GND.n1372 150.213
R2716 GND.n1372 GND.n1371 150.213
R2717 GND.n1368 GND.n1367 150.213
R2718 GND.n1326 GND.n1324 150.213
R2719 GND.n1334 GND.n1329 150.213
R2720 GND.n1474 GND.n1473 150.213
R2721 GND.n1470 GND.n1437 150.213
R2722 GND.n1486 GND.n1485 150.213
R2723 GND.n1454 GND.n1449 150.213
R2724 GND.n1455 GND.n1454 150.213
R2725 GND.n1485 GND.n1431 150.213
R2726 GND.n1423 GND.n1413 150.213
R2727 GND.n1421 GND.n1411 150.213
R2728 GND.n1460 GND.n1411 150.213
R2729 GND.n1461 GND.n1413 150.213
R2730 GND.n1491 GND.n1409 150.213
R2731 GND.n1493 GND.n1407 150.213
R2732 GND.n1443 GND.n1407 150.213
R2733 GND.n1444 GND.n1409 150.213
R2734 GND.n1439 GND.n1437 150.213
R2735 GND.n1474 GND.n1469 150.213
R2736 GND.n1948 GND.n1947 150.213
R2737 GND.n1944 GND.n1911 150.213
R2738 GND.n1960 GND.n1959 150.213
R2739 GND.n1928 GND.n1923 150.213
R2740 GND.n1929 GND.n1928 150.213
R2741 GND.n1959 GND.n1905 150.213
R2742 GND.n1897 GND.n1887 150.213
R2743 GND.n1895 GND.n1885 150.213
R2744 GND.n1934 GND.n1885 150.213
R2745 GND.n1935 GND.n1887 150.213
R2746 GND.n1965 GND.n1883 150.213
R2747 GND.n1967 GND.n1881 150.213
R2748 GND.n1917 GND.n1881 150.213
R2749 GND.n1918 GND.n1883 150.213
R2750 GND.n1913 GND.n1911 150.213
R2751 GND.n1948 GND.n1943 150.213
R2752 GND.n1682 GND.n1681 150.213
R2753 GND.n1678 GND.n1672 150.213
R2754 GND.n1694 GND.n1693 150.213
R2755 GND.n1664 GND.n1660 150.213
R2756 GND.n1664 GND.n1663 150.213
R2757 GND.n1693 GND.n1656 150.213
R2758 GND.n1731 GND.n1635 150.213
R2759 GND.n1644 GND.n1634 150.213
R2760 GND.n1734 GND.n1634 150.213
R2761 GND.n1732 GND.n1731 150.213
R2762 GND.n1715 GND.n1702 150.213
R2763 GND.n1721 GND.n1720 150.213
R2764 GND.n1720 GND.n1719 150.213
R2765 GND.n1716 GND.n1715 150.213
R2766 GND.n1674 GND.n1672 150.213
R2767 GND.n1682 GND.n1677 150.213
R2768 GND.n2424 GND.n2423 150.213
R2769 GND.n2420 GND.n2414 150.213
R2770 GND.n2436 GND.n2435 150.213
R2771 GND.n2406 GND.n2402 150.213
R2772 GND.n2406 GND.n2405 150.213
R2773 GND.n2435 GND.n2398 150.213
R2774 GND.n2473 GND.n582 150.213
R2775 GND.n591 GND.n581 150.213
R2776 GND.n2476 GND.n581 150.213
R2777 GND.n2474 GND.n2473 150.213
R2778 GND.n2457 GND.n2444 150.213
R2779 GND.n2463 GND.n2462 150.213
R2780 GND.n2462 GND.n2461 150.213
R2781 GND.n2458 GND.n2457 150.213
R2782 GND.n2416 GND.n2414 150.213
R2783 GND.n2424 GND.n2419 150.213
R2784 GND.n2694 GND.n2693 150.213
R2785 GND.n2690 GND.n2657 150.213
R2786 GND.n2706 GND.n2705 150.213
R2787 GND.n2674 GND.n2669 150.213
R2788 GND.n2675 GND.n2674 150.213
R2789 GND.n2705 GND.n2651 150.213
R2790 GND.n2643 GND.n2633 150.213
R2791 GND.n2641 GND.n2631 150.213
R2792 GND.n2680 GND.n2631 150.213
R2793 GND.n2681 GND.n2633 150.213
R2794 GND.n2711 GND.n2629 150.213
R2795 GND.n2713 GND.n2627 150.213
R2796 GND.n2663 GND.n2627 150.213
R2797 GND.n2664 GND.n2629 150.213
R2798 GND.n2659 GND.n2657 150.213
R2799 GND.n2694 GND.n2689 150.213
R2800 GND.n2978 GND.n2977 150.213
R2801 GND.n2974 GND.n2968 150.213
R2802 GND.n2990 GND.n2989 150.213
R2803 GND.n2960 GND.n2956 150.213
R2804 GND.n2960 GND.n2959 150.213
R2805 GND.n2989 GND.n2952 150.213
R2806 GND.n3027 GND.n469 150.213
R2807 GND.n478 GND.n468 150.213
R2808 GND.n3030 GND.n468 150.213
R2809 GND.n3028 GND.n3027 150.213
R2810 GND.n3011 GND.n2998 150.213
R2811 GND.n3017 GND.n3016 150.213
R2812 GND.n3016 GND.n3015 150.213
R2813 GND.n3012 GND.n3011 150.213
R2814 GND.n2970 GND.n2968 150.213
R2815 GND.n2978 GND.n2973 150.213
R2816 GND.n3235 GND.n3234 150.213
R2817 GND.n3231 GND.n3225 150.213
R2818 GND.n3247 GND.n3246 150.213
R2819 GND.n3217 GND.n3213 150.213
R2820 GND.n3217 GND.n3216 150.213
R2821 GND.n3246 GND.n3209 150.213
R2822 GND.n3284 GND.n3189 150.213
R2823 GND.n3198 GND.n3188 150.213
R2824 GND.n3287 GND.n3188 150.213
R2825 GND.n3285 GND.n3284 150.213
R2826 GND.n3268 GND.n3255 150.213
R2827 GND.n3274 GND.n3273 150.213
R2828 GND.n3273 GND.n3272 150.213
R2829 GND.n3269 GND.n3268 150.213
R2830 GND.n3227 GND.n3225 150.213
R2831 GND.n3235 GND.n3230 150.213
R2832 GND.n4158 GND.n4157 150.213
R2833 GND.n4154 GND.n4148 150.213
R2834 GND.n4170 GND.n4169 150.213
R2835 GND.n4140 GND.n4136 150.213
R2836 GND.n4140 GND.n4139 150.213
R2837 GND.n4169 GND.n4132 150.213
R2838 GND.n4207 GND.n4111 150.213
R2839 GND.n4120 GND.n4110 150.213
R2840 GND.n4210 GND.n4110 150.213
R2841 GND.n4208 GND.n4207 150.213
R2842 GND.n4191 GND.n4178 150.213
R2843 GND.n4197 GND.n4196 150.213
R2844 GND.n4196 GND.n4195 150.213
R2845 GND.n4192 GND.n4191 150.213
R2846 GND.n4150 GND.n4148 150.213
R2847 GND.n4158 GND.n4153 150.213
R2848 GND.n720 GND.n713 147.357
R2849 GND.n2828 GND.n284 140.334
R2850 GND.n2858 GND.n292 140.334
R2851 GND.n2882 GND.n300 140.334
R2852 GND.n166 GND.t596 110.361
R2853 GND.t166 GND.n138 110.361
R2854 GND.n3966 GND.t342 110.361
R2855 GND.n3358 GND.t107 110.361
R2856 GND.n3359 GND.t279 110.361
R2857 GND.n3360 GND.t358 110.361
R2858 GND.n2772 GND.t568 110.361
R2859 GND.t162 GND.n2743 110.361
R2860 GND.n2790 GND.t680 110.361
R2861 GND.n4340 GND.t570 110.361
R2862 GND.n4341 GND.t335 110.361
R2863 GND.n4342 GND.t615 110.361
R2864 GND.t251 GND.n1158 110.361
R2865 GND.n1139 GND.t236 110.361
R2866 GND.t642 GND.n1140 110.361
R2867 GND.n854 GND.t110 110.361
R2868 GND.t186 GND.n808 110.361
R2869 GND.n2029 GND.t217 110.361
R2870 GND.t569 GND.n2281 110.361
R2871 GND.n2262 GND.t689 110.361
R2872 GND.t125 GND.n2263 110.361
R2873 GND.t250 GND.n2379 110.361
R2874 GND.n2353 GND.t277 110.361
R2875 GND.t350 GND.n2354 110.361
R2876 GND.n3625 GND 105.755
R2877 GND.n4226 GND.n57 105.082
R2878 GND.n4283 GND.n57 105.082
R2879 GND.n4278 GND.n4277 105.082
R2880 GND.n4277 GND.n4231 105.082
R2881 GND.n1059 GND.n1015 105.082
R2882 GND.n1015 GND.n1014 105.082
R2883 GND.n1027 GND.n1018 105.082
R2884 GND.n1022 GND.n1018 105.082
R2885 GND.n1042 GND.n1041 105.082
R2886 GND.n1041 GND.n1039 105.082
R2887 GND.n4308 GND.n30 105.082
R2888 GND.n4308 GND.n29 105.082
R2889 GND.n180 GND.n47 105.082
R2890 GND.n180 GND.n46 105.082
R2891 GND.n158 GND.n136 105.082
R2892 GND.n158 GND.n137 105.082
R2893 GND.n3977 GND.n3976 105.082
R2894 GND.n3976 GND.n125 105.082
R2895 GND.n3993 GND.n98 105.082
R2896 GND.n3993 GND.n3992 105.082
R2897 GND.n3346 GND.n344 105.082
R2898 GND.n3363 GND.n344 105.082
R2899 GND.n2927 GND.n355 105.082
R2900 GND.n2927 GND.n354 105.082
R2901 GND.n2944 GND.n490 105.082
R2902 GND.n2944 GND.n2943 105.082
R2903 GND.n2764 GND.n2741 105.082
R2904 GND.n2764 GND.n2742 105.082
R2905 GND.n2804 GND.n2803 105.082
R2906 GND.n2803 GND.n552 105.082
R2907 GND.n2824 GND.n2823 105.082
R2908 GND.n2823 GND.n523 105.082
R2909 GND.n2385 GND.n2384 105.082
R2910 GND.n2384 GND.n2334 105.082
R2911 GND.n2390 GND.n603 105.082
R2912 GND.n2390 GND.n2389 105.082
R2913 GND.n644 GND.n618 105.082
R2914 GND.n2301 GND.n618 105.082
R2915 GND.n2287 GND.n631 105.082
R2916 GND.n2287 GND.n632 105.082
R2917 GND.n2001 GND.n2000 105.082
R2918 GND.n2000 GND.n882 105.082
R2919 GND.n866 GND.n815 105.082
R2920 GND.n866 GND.n816 105.082
R2921 GND.n846 GND.n806 105.082
R2922 GND.n846 GND.n807 105.082
R2923 GND.n2042 GND.n2041 105.082
R2924 GND.n2041 GND.n799 105.082
R2925 GND.n2062 GND.n2061 105.082
R2926 GND.n2061 GND.n770 105.082
R2927 GND.n1164 GND.n1123 105.082
R2928 GND.n1164 GND.n1124 105.082
R2929 GND.n1109 GND.n977 105.082
R2930 GND.n1118 GND.n977 105.082
R2931 GND.n1085 GND.n999 105.082
R2932 GND.n999 GND.n998 105.082
R2933 GND.n3486 GND.n196 105.082
R2934 GND.n3878 GND.n196 105.082
R2935 GND.n3505 GND.n304 105.082
R2936 GND.n3494 GND.n304 105.082
R2937 GND.n3527 GND.n296 105.082
R2938 GND.n3513 GND.n296 105.082
R2939 GND.n3549 GND.n288 105.082
R2940 GND.n3535 GND.n288 105.082
R2941 GND.n3568 GND.n280 105.082
R2942 GND.n3557 GND.n280 105.082
R2943 GND.n3588 GND.n272 105.082
R2944 GND.n3576 GND.n272 105.082
R2945 GND.n3607 GND.n254 105.082
R2946 GND.n3596 GND.n254 105.082
R2947 GND.n3618 GND.n3617 105.082
R2948 GND.n3617 GND.n247 105.082
R2949 GND.n2076 GND.n2075 105.082
R2950 GND.n2075 GND.n2074 105.082
R2951 GND.n2070 GND.n2069 105.082
R2952 GND.n2069 GND.n2068 105.082
R2953 GND.n2173 GND.n652 105.082
R2954 GND.n2178 GND.n652 105.082
R2955 GND.n2161 GND.n656 105.082
R2956 GND.n2166 GND.n656 105.082
R2957 GND.n2130 GND.n669 105.082
R2958 GND.n2135 GND.n669 105.082
R2959 GND.n2219 GND.n2208 105.082
R2960 GND.n2215 GND.n2208 105.082
R2961 GND.n2229 GND.n2228 105.082
R2962 GND.n2228 GND.n2199 105.082
R2963 GND.n2253 GND.n2252 105.082
R2964 GND.n2252 GND.n648 105.082
R2965 GND.n2874 GND.n502 105.082
R2966 GND.n2879 GND.n502 105.082
R2967 GND.n2862 GND.n506 105.082
R2968 GND.n2867 GND.n506 105.082
R2969 GND.n2831 GND.n519 105.082
R2970 GND.n2836 GND.n519 105.082
R2971 GND.n3445 GND.n328 105.082
R2972 GND.n3441 GND.n328 105.082
R2973 GND.n3456 GND.n323 105.082
R2974 GND.n3452 GND.n323 105.082
R2975 GND.n2895 GND.n2894 105.082
R2976 GND.n2894 GND.n496 105.082
R2977 GND.n3886 GND.n191 105.082
R2978 GND.n3891 GND.n191 105.082
R2979 GND.n3409 GND.n3408 105.082
R2980 GND.n3408 GND.n3398 105.082
R2981 GND.n3434 GND.n333 105.082
R2982 GND.n3430 GND.n333 105.082
R2983 GND.n3919 GND.n6 105.082
R2984 GND.n4366 GND.n6 105.082
R2985 GND.n3929 GND.n3928 105.082
R2986 GND.n3928 GND.n3910 105.082
R2987 GND.n3953 GND.n3952 105.082
R2988 GND.n3952 GND.n185 105.082
R2989 GND.n2118 GND.n674 105.082
R2990 GND.n2123 GND.n674 105.082
R2991 GND.n2106 GND.n678 105.082
R2992 GND.n2111 GND.n678 105.082
R2993 GND.n765 GND.n764 105.082
R2994 GND.n764 GND.n727 105.082
R2995 GND.n687 GND.n686 105.082
R2996 GND.n2095 GND.n686 105.082
R2997 GND.n4345 GND.n19 105.082
R2998 GND.n4328 GND.n19 105.082
R2999 GND.n4273 GND.n4245 105.082
R3000 GND.n4273 GND.n4241 105.082
R3001 GND.n1113 GND.n983 101.754
R3002 GND.n3612 GND.n3611 100.371
R3003 GND.n3611 GND.n3610 100.371
R3004 GND.n3593 GND.n3592 100.371
R3005 GND.n3592 GND.n3591 100.371
R3006 GND.n3573 GND.n3572 100.371
R3007 GND.n3572 GND.n3571 100.371
R3008 GND.n3554 GND.n3553 100.371
R3009 GND.n3553 GND.n3552 100.371
R3010 GND.n3532 GND.n3531 100.371
R3011 GND.n3531 GND.n3530 100.371
R3012 GND.n3510 GND.n3509 100.371
R3013 GND.n3509 GND.n3508 100.371
R3014 GND.n3491 GND.n3490 100.371
R3015 GND.n3490 GND.n3489 100.371
R3016 GND.n3622 GND 99.1472
R3017 GND.t121 GND.n721 92.3206
R3018 GND.n721 GND.t640 89.9046
R3019 GND.n2311 GND.n2310 86.0562
R3020 GND.n791 GND.n774 86.0562
R3021 GND.n1094 GND.n989 86.0562
R3022 GND.n872 GND.n817 86.0562
R3023 GND.n544 GND.n527 86.0562
R3024 GND.n2917 GND.n2916 86.0562
R3025 GND.n115 GND.n114 86.0562
R3026 GND.n4297 GND.n43 86.0562
R3027 GND.t311 GND.n773 82.622
R3028 GND.n1520 GND.t619 82.622
R3029 GND.t157 GND.n2297 82.622
R3030 GND.t227 GND.n526 82.622
R3031 GND.n2946 GND.t292 82.622
R3032 GND.n3995 GND.t699 82.622
R3033 GND.n4288 GND.t295 82.622
R3034 GND.n696 GND.n695 82.1844
R3035 GND.n2084 GND.n2083 82.1844
R3036 GND.n3319 GND.n385 81.7745
R3037 GND.n273 GND 79.3211
R3038 GND.n713 GND.n712 76.9339
R3039 GND.n716 GND.n715 76.9339
R3040 GND.n3623 GND 75.8872
R3041 GND.n4072 GND.n79 73.1255
R3042 GND.n3999 GND.n79 73.1255
R3043 GND.n81 GND.n80 73.1255
R3044 GND.n82 GND.n81 73.1255
R3045 GND.n62 GND.n61 73.1255
R3046 GND.n69 GND.n62 73.1255
R3047 GND.n4086 GND.n60 73.1255
R3048 GND.n63 GND.n60 73.1255
R3049 GND.n3150 GND.n3064 73.1255
R3050 GND.n3077 GND.n3064 73.1255
R3051 GND.n3066 GND.n3065 73.1255
R3052 GND.n3067 GND.n3066 73.1255
R3053 GND.n3047 GND.n3046 73.1255
R3054 GND.n3054 GND.n3047 73.1255
R3055 GND.n3164 GND.n3045 73.1255
R3056 GND.n3048 GND.n3045 73.1255
R3057 GND.n2597 GND.n2510 73.1255
R3058 GND.n2524 GND.n2510 73.1255
R3059 GND.n2512 GND.n2511 73.1255
R3060 GND.n2513 GND.n2512 73.1255
R3061 GND.n2493 GND.n2492 73.1255
R3062 GND.n2500 GND.n2493 73.1255
R3063 GND.n2611 GND.n2491 73.1255
R3064 GND.n2494 GND.n2491 73.1255
R3065 GND.n1852 GND.n1767 73.1255
R3066 GND.n1767 GND.n622 73.1255
R3067 GND.n1769 GND.n1768 73.1255
R3068 GND.n1770 GND.n1769 73.1255
R3069 GND.n1751 GND.n1750 73.1255
R3070 GND.n1757 GND.n1751 73.1255
R3071 GND.n1866 GND.n1749 73.1255
R3072 GND.n1749 GND.n623 73.1255
R3073 GND.n1595 GND.n915 73.1255
R3074 GND.n1522 GND.n915 73.1255
R3075 GND.n917 GND.n916 73.1255
R3076 GND.n918 GND.n917 73.1255
R3077 GND.n898 GND.n897 73.1255
R3078 GND.n905 GND.n898 73.1255
R3079 GND.n1609 GND.n896 73.1255
R3080 GND.n899 GND.n896 73.1255
R3081 GND.n1247 GND.n958 73.1255
R3082 GND.n1174 GND.n958 73.1255
R3083 GND.n960 GND.n959 73.1255
R3084 GND.n961 GND.n960 73.1255
R3085 GND.n941 GND.n940 73.1255
R3086 GND.n948 GND.n941 73.1255
R3087 GND.n1261 GND.n939 73.1255
R3088 GND.n942 GND.n939 73.1255
R3089 GND.n1377 GND.n1290 73.1255
R3090 GND.n1304 GND.n1290 73.1255
R3091 GND.n1292 GND.n1291 73.1255
R3092 GND.n1293 GND.n1292 73.1255
R3093 GND.n1273 GND.n1272 73.1255
R3094 GND.n1280 GND.n1273 73.1255
R3095 GND.n1391 GND.n1271 73.1255
R3096 GND.n1274 GND.n1271 73.1255
R3097 GND.n1497 GND.n1415 73.1255
R3098 GND.n1415 GND.n928 73.1255
R3099 GND.n1417 GND.n1416 73.1255
R3100 GND.n1418 GND.n1417 73.1255
R3101 GND.n1465 GND.n1464 73.1255
R3102 GND.n1466 GND.n1465 73.1255
R3103 GND.n1517 GND.n1516 73.1255
R3104 GND.n1518 GND.n1517 73.1255
R3105 GND.n162 GND.n148 73.1255
R3106 GND.n148 GND.t344 73.1255
R3107 GND.n149 GND.n147 73.1255
R3108 GND.n147 GND.t344 73.1255
R3109 GND.n3351 GND.n349 73.1255
R3110 GND.n349 GND.t321 73.1255
R3111 GND.n350 GND.n348 73.1255
R3112 GND.n348 GND.t321 73.1255
R3113 GND.n2768 GND.n2753 73.1255
R3114 GND.n2753 GND.t306 73.1255
R3115 GND.n2754 GND.n2752 73.1255
R3116 GND.n2752 GND.t306 73.1255
R3117 GND.n2154 GND.n658 73.1255
R3118 GND.n658 GND.t657 73.1255
R3119 GND.n659 GND.n657 73.1255
R3120 GND.n657 GND.t657 73.1255
R3121 GND.n2233 GND.n2194 73.1255
R3122 GND.n2194 GND.t515 73.1255
R3123 GND.n2195 GND.n2193 73.1255
R3124 GND.n2193 GND.t515 73.1255
R3125 GND.n2855 GND.n508 73.1255
R3126 GND.t34 GND.n508 73.1255
R3127 GND.n509 GND.n507 73.1255
R3128 GND.t34 GND.n507 73.1255
R3129 GND.n3463 GND.n316 73.1255
R3130 GND.t300 GND.n316 73.1255
R3131 GND.n319 GND.n317 73.1255
R3132 GND.t300 GND.n319 73.1255
R3133 GND.n745 GND.n739 73.1255
R3134 GND.n739 GND.t5 73.1255
R3135 GND.n740 GND.n738 73.1255
R3136 GND.n738 GND.t5 73.1255
R3137 GND.n4358 GND.n12 73.1255
R3138 GND.n12 GND.t252 73.1255
R3139 GND.n13 GND.n11 73.1255
R3140 GND.n11 GND.t252 73.1255
R3141 GND.n4333 GND.n24 73.1255
R3142 GND.n24 GND.t151 73.1255
R3143 GND.n25 GND.n23 73.1255
R3144 GND.n23 GND.t151 73.1255
R3145 GND.n3413 GND.n3391 73.1255
R3146 GND.n3391 GND.t178 73.1255
R3147 GND.n3392 GND.n3390 73.1255
R3148 GND.n3390 GND.t178 73.1255
R3149 GND.n3933 GND.n3905 73.1255
R3150 GND.n3905 GND.t243 73.1255
R3151 GND.n3906 GND.n3904 73.1255
R3152 GND.n3904 GND.t243 73.1255
R3153 GND.n2080 GND.n698 73.1255
R3154 GND.n698 GND.t262 73.1255
R3155 GND.n699 GND.n697 73.1255
R3156 GND.n697 GND.t262 73.1255
R3157 GND.n1004 GND.n1003 73.1255
R3158 GND.n1004 GND.n981 73.1255
R3159 GND.n1067 GND.n1002 73.1255
R3160 GND.n1002 GND.n983 73.1255
R3161 GND.n1168 GND.n973 73.1255
R3162 GND.t664 GND.n973 73.1255
R3163 GND.n974 GND.n972 73.1255
R3164 GND.t664 GND.n972 73.1255
R3165 GND.n1138 GND.n1137 73.1255
R3166 GND.t17 GND.n1138 73.1255
R3167 GND.n1149 GND.n1136 73.1255
R3168 GND.t17 GND.n1136 73.1255
R3169 GND.n850 GND.n836 73.1255
R3170 GND.n836 GND.t572 73.1255
R3171 GND.n837 GND.n835 73.1255
R3172 GND.n835 GND.t572 73.1255
R3173 GND.n2025 GND.n811 73.1255
R3174 GND.t15 GND.n811 73.1255
R3175 GND.n812 GND.n810 73.1255
R3176 GND.t15 GND.n810 73.1255
R3177 GND.n1971 GND.n1889 73.1255
R3178 GND.n1889 GND.n885 73.1255
R3179 GND.n1891 GND.n1890 73.1255
R3180 GND.n1892 GND.n1891 73.1255
R3181 GND.n1939 GND.n1938 73.1255
R3182 GND.n1940 GND.n1939 73.1255
R3183 GND.n1991 GND.n1990 73.1255
R3184 GND.n1992 GND.n1991 73.1255
R3185 GND.n2291 GND.n626 73.1255
R3186 GND.t512 GND.n626 73.1255
R3187 GND.n627 GND.n625 73.1255
R3188 GND.t512 GND.n625 73.1255
R3189 GND.n2261 GND.n2260 73.1255
R3190 GND.t597 GND.n2261 73.1255
R3191 GND.n2272 GND.n2259 73.1255
R3192 GND.t597 GND.n2259 73.1255
R3193 GND.n1725 GND.n1639 73.1255
R3194 GND.n1652 GND.n1639 73.1255
R3195 GND.n1641 GND.n1640 73.1255
R3196 GND.n1642 GND.n1641 73.1255
R3197 GND.n1622 GND.n1621 73.1255
R3198 GND.n1629 GND.n1622 73.1255
R3199 GND.n1739 GND.n1620 73.1255
R3200 GND.n1623 GND.n1620 73.1255
R3201 GND.n2467 GND.n586 73.1255
R3202 GND.n2394 GND.n586 73.1255
R3203 GND.n588 GND.n587 73.1255
R3204 GND.n589 GND.n588 73.1255
R3205 GND.n569 GND.n568 73.1255
R3206 GND.n576 GND.n569 73.1255
R3207 GND.n2481 GND.n567 73.1255
R3208 GND.n570 GND.n567 73.1255
R3209 GND.n2345 GND.n2338 73.1255
R3210 GND.n2338 GND.t352 73.1255
R3211 GND.n2339 GND.n2337 73.1255
R3212 GND.n2337 GND.t352 73.1255
R3213 GND.n2362 GND.n2358 73.1255
R3214 GND.t108 GND.n2358 73.1255
R3215 GND.n2367 GND.n2366 73.1255
R3216 GND.t108 GND.n2367 73.1255
R3217 GND.n2717 GND.n2635 73.1255
R3218 GND.n2635 GND.n556 73.1255
R3219 GND.n2637 GND.n2636 73.1255
R3220 GND.n2638 GND.n2637 73.1255
R3221 GND.n2685 GND.n2684 73.1255
R3222 GND.n2686 GND.n2685 73.1255
R3223 GND.n2737 GND.n2736 73.1255
R3224 GND.n2738 GND.n2737 73.1255
R3225 GND.n3021 GND.n473 73.1255
R3226 GND.n2948 GND.n473 73.1255
R3227 GND.n475 GND.n474 73.1255
R3228 GND.n476 GND.n475 73.1255
R3229 GND.n456 GND.n455 73.1255
R3230 GND.n463 GND.n456 73.1255
R3231 GND.n3035 GND.n454 73.1255
R3232 GND.n457 GND.n454 73.1255
R3233 GND.n2786 GND.n2746 73.1255
R3234 GND.t13 GND.n2746 73.1255
R3235 GND.n2781 GND.n2745 73.1255
R3236 GND.t13 GND.n2745 73.1255
R3237 GND.n400 GND.n396 73.1255
R3238 GND.n396 GND.n385 73.1255
R3239 GND.n397 GND.n361 73.1255
R3240 GND.n3332 GND.n361 73.1255
R3241 GND.n450 GND.n449 73.1255
R3242 GND.n449 GND.n94 73.1255
R3243 GND.n3318 GND.n3317 73.1255
R3244 GND.n3319 GND.n3318 73.1255
R3245 GND.n3278 GND.n3193 73.1255
R3246 GND.n3193 GND.n92 73.1255
R3247 GND.n3195 GND.n3194 73.1255
R3248 GND.n3196 GND.n3195 73.1255
R3249 GND.n3177 GND.n3176 73.1255
R3250 GND.n3183 GND.n3177 73.1255
R3251 GND.n3292 GND.n3175 73.1255
R3252 GND.n3175 GND.n93 73.1255
R3253 GND.n3375 GND.n3374 73.1255
R3254 GND.t248 GND.n3375 73.1255
R3255 GND.n3377 GND.n3376 73.1255
R3256 GND.n3376 GND.t248 73.1255
R3257 GND.n4201 GND.n4115 73.1255
R3258 GND.n4128 GND.n4115 73.1255
R3259 GND.n4117 GND.n4116 73.1255
R3260 GND.n4118 GND.n4117 73.1255
R3261 GND.n4098 GND.n4097 73.1255
R3262 GND.n4105 GND.n4098 73.1255
R3263 GND.n4215 GND.n4096 73.1255
R3264 GND.n4099 GND.n4096 73.1255
R3265 GND.n3962 GND.n141 73.1255
R3266 GND.n141 GND.t11 73.1255
R3267 GND.n3959 GND.n140 73.1255
R3268 GND.t11 GND.n140 73.1255
R3269 GND.n4254 GND.n4237 73.1255
R3270 GND.n4275 GND.n4237 73.1255
R3271 GND.n4251 GND.n53 73.1255
R3272 GND.n4287 GND.n53 73.1255
R3273 GND.n3620 GND 71.1372
R3274 GND.n3477 GND.t722 69.8913
R3275 GND.n3499 GND.t675 69.8913
R3276 GND.n3521 GND.t317 69.8913
R3277 GND.n3540 GND.t66 69.8913
R3278 GND.n3562 GND.t202 69.8913
R3279 GND.n3581 GND.t509 69.8913
R3280 GND.n3601 GND.t128 69.8913
R3281 GND.n258 GND.t135 69.8913
R3282 GND.n281 GND 66.1038
R3283 GND.n4028 GND.n90 65.0005
R3284 GND.t37 GND.n90 65.0005
R3285 GND.n4025 GND.n89 65.0005
R3286 GND.t37 GND.n89 65.0005
R3287 GND.n4024 GND.n68 65.0005
R3288 GND.t138 GND.n68 65.0005
R3289 GND.n4021 GND.n67 65.0005
R3290 GND.t138 GND.n67 65.0005
R3291 GND.n4042 GND.n4041 65.0005
R3292 GND.t37 GND.n4042 65.0005
R3293 GND.n4007 GND.n88 65.0005
R3294 GND.t37 GND.n88 65.0005
R3295 GND.n4003 GND.n70 65.0005
R3296 GND.t138 GND.n70 65.0005
R3297 GND.n4010 GND.n66 65.0005
R3298 GND.t138 GND.n66 65.0005
R3299 GND.n4071 GND.n4070 65.0005
R3300 GND.n4070 GND.t37 65.0005
R3301 GND.n4043 GND.n78 65.0005
R3302 GND.t37 GND.n4043 65.0005
R3303 GND.n87 GND.n75 65.0005
R3304 GND.t37 GND.n87 65.0005
R3305 GND.n84 GND.n83 65.0005
R3306 GND.t37 GND.n83 65.0005
R3307 GND.n4079 GND.n71 65.0005
R3308 GND.t138 GND.n71 65.0005
R3309 GND.n4082 GND.n4081 65.0005
R3310 GND.t138 GND.n4082 65.0005
R3311 GND.n4049 GND.n4044 65.0005
R3312 GND.t37 GND.n4044 65.0005
R3313 GND.n4069 GND.n4068 65.0005
R3314 GND.t37 GND.n4069 65.0005
R3315 GND.n4063 GND.n65 65.0005
R3316 GND.t138 GND.n65 65.0005
R3317 GND.n4066 GND.n64 65.0005
R3318 GND.t138 GND.n64 65.0005
R3319 GND.n4085 GND.n4084 65.0005
R3320 GND.n4084 GND.t138 65.0005
R3321 GND.n4083 GND.n59 65.0005
R3322 GND.t138 GND.n4083 65.0005
R3323 GND.n3106 GND.n3075 65.0005
R3324 GND.t43 GND.n3075 65.0005
R3325 GND.n3103 GND.n3074 65.0005
R3326 GND.t43 GND.n3074 65.0005
R3327 GND.n3102 GND.n3053 65.0005
R3328 GND.t62 GND.n3053 65.0005
R3329 GND.n3099 GND.n3052 65.0005
R3330 GND.t62 GND.n3052 65.0005
R3331 GND.n3120 GND.n3119 65.0005
R3332 GND.t43 GND.n3120 65.0005
R3333 GND.n3085 GND.n3073 65.0005
R3334 GND.t43 GND.n3073 65.0005
R3335 GND.n3081 GND.n3055 65.0005
R3336 GND.t62 GND.n3055 65.0005
R3337 GND.n3088 GND.n3051 65.0005
R3338 GND.t62 GND.n3051 65.0005
R3339 GND.n3149 GND.n3148 65.0005
R3340 GND.n3148 GND.t43 65.0005
R3341 GND.n3121 GND.n3063 65.0005
R3342 GND.t43 GND.n3121 65.0005
R3343 GND.n3072 GND.n3060 65.0005
R3344 GND.t43 GND.n3072 65.0005
R3345 GND.n3069 GND.n3068 65.0005
R3346 GND.t43 GND.n3068 65.0005
R3347 GND.n3157 GND.n3056 65.0005
R3348 GND.t62 GND.n3056 65.0005
R3349 GND.n3160 GND.n3159 65.0005
R3350 GND.t62 GND.n3160 65.0005
R3351 GND.n3127 GND.n3122 65.0005
R3352 GND.t43 GND.n3122 65.0005
R3353 GND.n3147 GND.n3146 65.0005
R3354 GND.t43 GND.n3147 65.0005
R3355 GND.n3141 GND.n3050 65.0005
R3356 GND.t62 GND.n3050 65.0005
R3357 GND.n3144 GND.n3049 65.0005
R3358 GND.t62 GND.n3049 65.0005
R3359 GND.n3163 GND.n3162 65.0005
R3360 GND.n3162 GND.t62 65.0005
R3361 GND.n3161 GND.n3044 65.0005
R3362 GND.t62 GND.n3161 65.0005
R3363 GND.n2553 GND.n2521 65.0005
R3364 GND.t25 GND.n2521 65.0005
R3365 GND.n2550 GND.n2520 65.0005
R3366 GND.t25 GND.n2520 65.0005
R3367 GND.n2549 GND.n2499 65.0005
R3368 GND.t50 GND.n2499 65.0005
R3369 GND.n2546 GND.n2498 65.0005
R3370 GND.t50 GND.n2498 65.0005
R3371 GND.n2567 GND.n2566 65.0005
R3372 GND.t25 GND.n2567 65.0005
R3373 GND.n2532 GND.n2519 65.0005
R3374 GND.t25 GND.n2519 65.0005
R3375 GND.n2528 GND.n2501 65.0005
R3376 GND.t50 GND.n2501 65.0005
R3377 GND.n2535 GND.n2497 65.0005
R3378 GND.t50 GND.n2497 65.0005
R3379 GND.n2596 GND.n2595 65.0005
R3380 GND.n2595 GND.t25 65.0005
R3381 GND.n2568 GND.n2509 65.0005
R3382 GND.t25 GND.n2568 65.0005
R3383 GND.n2518 GND.n2506 65.0005
R3384 GND.t25 GND.n2518 65.0005
R3385 GND.n2515 GND.n2514 65.0005
R3386 GND.t25 GND.n2514 65.0005
R3387 GND.n2604 GND.n2502 65.0005
R3388 GND.t50 GND.n2502 65.0005
R3389 GND.n2607 GND.n2606 65.0005
R3390 GND.t50 GND.n2607 65.0005
R3391 GND.n2574 GND.n2569 65.0005
R3392 GND.t25 GND.n2569 65.0005
R3393 GND.n2594 GND.n2593 65.0005
R3394 GND.t25 GND.n2594 65.0005
R3395 GND.n2588 GND.n2496 65.0005
R3396 GND.t50 GND.n2496 65.0005
R3397 GND.n2591 GND.n2495 65.0005
R3398 GND.t50 GND.n2495 65.0005
R3399 GND.n2610 GND.n2609 65.0005
R3400 GND.n2609 GND.t50 65.0005
R3401 GND.n2608 GND.n2490 65.0005
R3402 GND.t50 GND.n2608 65.0005
R3403 GND.n1808 GND.n1779 65.0005
R3404 GND.t21 GND.n1779 65.0005
R3405 GND.n1805 GND.n1778 65.0005
R3406 GND.t21 GND.n1778 65.0005
R3407 GND.n1804 GND.n1756 65.0005
R3408 GND.t22 GND.n1756 65.0005
R3409 GND.n1801 GND.n1755 65.0005
R3410 GND.t22 GND.n1755 65.0005
R3411 GND.n1822 GND.n1821 65.0005
R3412 GND.t21 GND.n1822 65.0005
R3413 GND.n1787 GND.n1777 65.0005
R3414 GND.t21 GND.n1777 65.0005
R3415 GND.n1783 GND.n1758 65.0005
R3416 GND.t22 GND.n1758 65.0005
R3417 GND.n1790 GND.n1754 65.0005
R3418 GND.t22 GND.n1754 65.0005
R3419 GND.n1851 GND.n1850 65.0005
R3420 GND.n1850 GND.t21 65.0005
R3421 GND.n1823 GND.n1766 65.0005
R3422 GND.t21 GND.n1823 65.0005
R3423 GND.n1776 GND.n1763 65.0005
R3424 GND.t21 GND.n1776 65.0005
R3425 GND.n1772 GND.n1771 65.0005
R3426 GND.t21 GND.n1771 65.0005
R3427 GND.n1859 GND.n1759 65.0005
R3428 GND.t22 GND.n1759 65.0005
R3429 GND.n1862 GND.n1861 65.0005
R3430 GND.t22 GND.n1862 65.0005
R3431 GND.n1829 GND.n1824 65.0005
R3432 GND.t21 GND.n1824 65.0005
R3433 GND.n1849 GND.n1848 65.0005
R3434 GND.t21 GND.n1849 65.0005
R3435 GND.n1843 GND.n1753 65.0005
R3436 GND.t22 GND.n1753 65.0005
R3437 GND.n1846 GND.n1752 65.0005
R3438 GND.t22 GND.n1752 65.0005
R3439 GND.n1865 GND.n1864 65.0005
R3440 GND.n1864 GND.t22 65.0005
R3441 GND.n1863 GND.n1748 65.0005
R3442 GND.t22 GND.n1863 65.0005
R3443 GND.n1551 GND.n926 65.0005
R3444 GND.t55 GND.n926 65.0005
R3445 GND.n1548 GND.n925 65.0005
R3446 GND.t55 GND.n925 65.0005
R3447 GND.n1547 GND.n904 65.0005
R3448 GND.t40 GND.n904 65.0005
R3449 GND.n1544 GND.n903 65.0005
R3450 GND.t40 GND.n903 65.0005
R3451 GND.n1565 GND.n1564 65.0005
R3452 GND.t55 GND.n1565 65.0005
R3453 GND.n1530 GND.n924 65.0005
R3454 GND.t55 GND.n924 65.0005
R3455 GND.n1526 GND.n906 65.0005
R3456 GND.t40 GND.n906 65.0005
R3457 GND.n1533 GND.n902 65.0005
R3458 GND.t40 GND.n902 65.0005
R3459 GND.n1594 GND.n1593 65.0005
R3460 GND.n1593 GND.t55 65.0005
R3461 GND.n1566 GND.n914 65.0005
R3462 GND.t55 GND.n1566 65.0005
R3463 GND.n923 GND.n911 65.0005
R3464 GND.t55 GND.n923 65.0005
R3465 GND.n920 GND.n919 65.0005
R3466 GND.t55 GND.n919 65.0005
R3467 GND.n1602 GND.n907 65.0005
R3468 GND.t40 GND.n907 65.0005
R3469 GND.n1605 GND.n1604 65.0005
R3470 GND.t40 GND.n1605 65.0005
R3471 GND.n1572 GND.n1567 65.0005
R3472 GND.t55 GND.n1567 65.0005
R3473 GND.n1592 GND.n1591 65.0005
R3474 GND.t55 GND.n1592 65.0005
R3475 GND.n1586 GND.n901 65.0005
R3476 GND.t40 GND.n901 65.0005
R3477 GND.n1589 GND.n900 65.0005
R3478 GND.t40 GND.n900 65.0005
R3479 GND.n1608 GND.n1607 65.0005
R3480 GND.n1607 GND.t40 65.0005
R3481 GND.n1606 GND.n895 65.0005
R3482 GND.t40 GND.n1606 65.0005
R3483 GND.n1203 GND.n969 65.0005
R3484 GND.t95 GND.n969 65.0005
R3485 GND.n1200 GND.n968 65.0005
R3486 GND.t95 GND.n968 65.0005
R3487 GND.n1199 GND.n947 65.0005
R3488 GND.t84 GND.n947 65.0005
R3489 GND.n1196 GND.n946 65.0005
R3490 GND.t84 GND.n946 65.0005
R3491 GND.n1217 GND.n1216 65.0005
R3492 GND.t95 GND.n1217 65.0005
R3493 GND.n1182 GND.n967 65.0005
R3494 GND.t95 GND.n967 65.0005
R3495 GND.n1178 GND.n949 65.0005
R3496 GND.t84 GND.n949 65.0005
R3497 GND.n1185 GND.n945 65.0005
R3498 GND.t84 GND.n945 65.0005
R3499 GND.n1246 GND.n1245 65.0005
R3500 GND.n1245 GND.t95 65.0005
R3501 GND.n1218 GND.n957 65.0005
R3502 GND.t95 GND.n1218 65.0005
R3503 GND.n966 GND.n954 65.0005
R3504 GND.t95 GND.n966 65.0005
R3505 GND.n963 GND.n962 65.0005
R3506 GND.t95 GND.n962 65.0005
R3507 GND.n1254 GND.n950 65.0005
R3508 GND.t84 GND.n950 65.0005
R3509 GND.n1257 GND.n1256 65.0005
R3510 GND.t84 GND.n1257 65.0005
R3511 GND.n1224 GND.n1219 65.0005
R3512 GND.t95 GND.n1219 65.0005
R3513 GND.n1244 GND.n1243 65.0005
R3514 GND.t95 GND.n1244 65.0005
R3515 GND.n1238 GND.n944 65.0005
R3516 GND.t84 GND.n944 65.0005
R3517 GND.n1241 GND.n943 65.0005
R3518 GND.t84 GND.n943 65.0005
R3519 GND.n1260 GND.n1259 65.0005
R3520 GND.n1259 GND.t84 65.0005
R3521 GND.n1258 GND.n938 65.0005
R3522 GND.t84 GND.n1258 65.0005
R3523 GND.n1333 GND.n1301 65.0005
R3524 GND.t90 GND.n1301 65.0005
R3525 GND.n1330 GND.n1300 65.0005
R3526 GND.t90 GND.n1300 65.0005
R3527 GND.n1329 GND.n1279 65.0005
R3528 GND.t149 GND.n1279 65.0005
R3529 GND.n1326 GND.n1278 65.0005
R3530 GND.t149 GND.n1278 65.0005
R3531 GND.n1347 GND.n1346 65.0005
R3532 GND.t90 GND.n1347 65.0005
R3533 GND.n1312 GND.n1299 65.0005
R3534 GND.t90 GND.n1299 65.0005
R3535 GND.n1308 GND.n1281 65.0005
R3536 GND.t149 GND.n1281 65.0005
R3537 GND.n1315 GND.n1277 65.0005
R3538 GND.t149 GND.n1277 65.0005
R3539 GND.n1376 GND.n1375 65.0005
R3540 GND.n1375 GND.t90 65.0005
R3541 GND.n1348 GND.n1289 65.0005
R3542 GND.t90 GND.n1348 65.0005
R3543 GND.n1298 GND.n1286 65.0005
R3544 GND.t90 GND.n1298 65.0005
R3545 GND.n1295 GND.n1294 65.0005
R3546 GND.t90 GND.n1294 65.0005
R3547 GND.n1384 GND.n1282 65.0005
R3548 GND.t149 GND.n1282 65.0005
R3549 GND.n1387 GND.n1386 65.0005
R3550 GND.t149 GND.n1387 65.0005
R3551 GND.n1354 GND.n1349 65.0005
R3552 GND.t90 GND.n1349 65.0005
R3553 GND.n1374 GND.n1373 65.0005
R3554 GND.t90 GND.n1374 65.0005
R3555 GND.n1368 GND.n1276 65.0005
R3556 GND.t149 GND.n1276 65.0005
R3557 GND.n1371 GND.n1275 65.0005
R3558 GND.t149 GND.n1275 65.0005
R3559 GND.n1390 GND.n1389 65.0005
R3560 GND.n1389 GND.t149 65.0005
R3561 GND.n1388 GND.n1270 65.0005
R3562 GND.t149 GND.n1388 65.0005
R3563 GND.n1473 GND.n1427 65.0005
R3564 GND.t70 GND.n1427 65.0005
R3565 GND.n1470 GND.n1426 65.0005
R3566 GND.t70 GND.n1426 65.0005
R3567 GND.n1469 GND.n1468 65.0005
R3568 GND.n1468 GND.t28 65.0005
R3569 GND.n1440 GND.n1439 65.0005
R3570 GND.n1440 GND.t28 65.0005
R3571 GND.n1487 GND.n1486 65.0005
R3572 GND.t70 GND.n1487 65.0005
R3573 GND.n1449 GND.n1425 65.0005
R3574 GND.t70 GND.n1425 65.0005
R3575 GND.n1448 GND.n1431 65.0005
R3576 GND.n1448 GND.t28 65.0005
R3577 GND.n1455 GND.n1447 65.0005
R3578 GND.n1447 GND.t28 65.0005
R3579 GND.n1496 GND.n1495 65.0005
R3580 GND.n1495 GND.t70 65.0005
R3581 GND.n1488 GND.n1414 65.0005
R3582 GND.t70 GND.n1488 65.0005
R3583 GND.n1424 GND.n1423 65.0005
R3584 GND.t70 GND.n1424 65.0005
R3585 GND.n1421 GND.n1419 65.0005
R3586 GND.t70 GND.n1419 65.0005
R3587 GND.n1461 GND.n1459 65.0005
R3588 GND.n1459 GND.t28 65.0005
R3589 GND.n1460 GND.n1458 65.0005
R3590 GND.n1458 GND.t28 65.0005
R3591 GND.n1491 GND.n1489 65.0005
R3592 GND.t70 GND.n1489 65.0005
R3593 GND.n1494 GND.n1493 65.0005
R3594 GND.t70 GND.n1494 65.0005
R3595 GND.n1444 GND.n1442 65.0005
R3596 GND.n1442 GND.t28 65.0005
R3597 GND.n1443 GND.n1441 65.0005
R3598 GND.n1441 GND.t28 65.0005
R3599 GND.n936 GND.n934 65.0005
R3600 GND.n934 GND.t28 65.0005
R3601 GND.n935 GND.n933 65.0005
R3602 GND.n933 GND.t28 65.0005
R3603 GND.n3964 GND.n3963 65.0005
R3604 GND.n3965 GND.n3964 65.0005
R3605 GND.n164 GND.n163 65.0005
R3606 GND.n165 GND.n164 65.0005
R3607 GND.n151 GND.n150 65.0005
R3608 GND.n150 GND.n133 65.0005
R3609 GND.n170 GND.n169 65.0005
R3610 GND.n169 GND.n139 65.0005
R3611 GND.n167 GND.n146 65.0005
R3612 GND.n167 GND.n166 65.0005
R3613 GND.n3968 GND.n3967 65.0005
R3614 GND.n3967 GND.n3966 65.0005
R3615 GND.n336 GND.n334 65.0005
R3616 GND.n338 GND.n336 65.0005
R3617 GND.n3353 GND.n3352 65.0005
R3618 GND.n3354 GND.n3353 65.0005
R3619 GND.n3341 GND.n351 65.0005
R3620 GND.n3342 GND.n3341 65.0005
R3621 GND.n3370 GND.n3369 65.0005
R3622 GND.n3371 GND.n3370 65.0005
R3623 GND.n3357 GND.n3356 65.0005
R3624 GND.n3358 GND.n3357 65.0005
R3625 GND.n3362 GND.n3361 65.0005
R3626 GND.n3361 GND.n3360 65.0005
R3627 GND.n2788 GND.n2787 65.0005
R3628 GND.n2789 GND.n2788 65.0005
R3629 GND.n2770 GND.n2769 65.0005
R3630 GND.n2771 GND.n2770 65.0005
R3631 GND.n2757 GND.n2756 65.0005
R3632 GND.n2756 GND.n2755 65.0005
R3633 GND.n2776 GND.n2775 65.0005
R3634 GND.n2775 GND.n2744 65.0005
R3635 GND.n2773 GND.n2751 65.0005
R3636 GND.n2773 GND.n2772 65.0005
R3637 GND.n2792 GND.n2791 65.0005
R3638 GND.n2791 GND.n2790 65.0005
R3639 GND.n2322 GND.n2321 65.0005
R3640 GND.n2321 GND.n2320 65.0005
R3641 GND.n2310 GND.n2309 65.0005
R3642 GND.n2317 GND.n2316 65.0005
R3643 GND.n2318 GND.n2317 65.0005
R3644 GND.n2047 GND.n2046 65.0005
R3645 GND.n2048 GND.n2047 65.0005
R3646 GND.n792 GND.n791 65.0005
R3647 GND.n2051 GND.n2050 65.0005
R3648 GND.n2050 GND.n2049 65.0005
R3649 GND.n1105 GND.n1104 65.0005
R3650 GND.n1104 GND.n984 65.0005
R3651 GND.n1076 GND.n989 65.0005
R3652 GND.n1100 GND.n1099 65.0005
R3653 GND.n1101 GND.n1100 65.0005
R3654 GND.n2148 GND.n2147 65.0005
R3655 GND.n2147 GND.n2146 65.0005
R3656 GND.n2156 GND.n2155 65.0005
R3657 GND.n2157 GND.n2156 65.0005
R3658 GND.n2144 GND.n660 65.0005
R3659 GND.n2145 GND.n2144 65.0005
R3660 GND.n2168 GND.n2167 65.0005
R3661 GND.n2169 GND.n2168 65.0005
R3662 GND.n2160 GND.n2159 65.0005
R3663 GND.n2159 GND.n2158 65.0005
R3664 GND.n2180 GND.n2179 65.0005
R3665 GND.n2181 GND.n2180 65.0005
R3666 GND.n2172 GND.n2171 65.0005
R3667 GND.n2171 GND.n2170 65.0005
R3668 GND.n2248 GND.n2184 65.0005
R3669 GND.n2247 GND.n2184 65.0005
R3670 GND.n2183 GND.n647 65.0005
R3671 GND.n2183 GND.n2182 65.0005
R3672 GND.n2239 GND.n2238 65.0005
R3673 GND.n2238 GND.n2237 65.0005
R3674 GND.n2245 GND.n2244 65.0005
R3675 GND.n2246 GND.n2245 65.0005
R3676 GND.n2200 GND.n2196 65.0005
R3677 GND.n2201 GND.n2200 65.0005
R3678 GND.n2235 GND.n2234 65.0005
R3679 GND.n2236 GND.n2235 65.0005
R3680 GND.n2224 GND.n2204 65.0005
R3681 GND.n2223 GND.n2204 65.0005
R3682 GND.n2203 GND.n2198 65.0005
R3683 GND.n2203 GND.n2202 65.0005
R3684 GND.n2214 GND.n2213 65.0005
R3685 GND.n2213 GND.n2212 65.0005
R3686 GND.n2221 GND.n2220 65.0005
R3687 GND.n2222 GND.n2221 65.0005
R3688 GND.n2838 GND.n2837 65.0005
R3689 GND.n2839 GND.n2838 65.0005
R3690 GND.n2830 GND.n2829 65.0005
R3691 GND.n2829 GND.n2828 65.0005
R3692 GND.n2849 GND.n2848 65.0005
R3693 GND.n2848 GND.n2847 65.0005
R3694 GND.n2842 GND.n2841 65.0005
R3695 GND.n2843 GND.n2842 65.0005
R3696 GND.n2857 GND.n2856 65.0005
R3697 GND.n2858 GND.n2857 65.0005
R3698 GND.n2845 GND.n510 65.0005
R3699 GND.n2846 GND.n2845 65.0005
R3700 GND.n2869 GND.n2868 65.0005
R3701 GND.n2870 GND.n2869 65.0005
R3702 GND.n2861 GND.n2860 65.0005
R3703 GND.n2860 GND.n2859 65.0005
R3704 GND.n2881 GND.n2880 65.0005
R3705 GND.n2882 GND.n2881 65.0005
R3706 GND.n2873 GND.n2872 65.0005
R3707 GND.n2872 GND.n2871 65.0005
R3708 GND.n2890 GND.n498 65.0005
R3709 GND.n2889 GND.n498 65.0005
R3710 GND.n497 GND.n493 65.0005
R3711 GND.n2883 GND.n497 65.0005
R3712 GND.n3469 GND.n3468 65.0005
R3713 GND.n3470 GND.n3469 65.0005
R3714 GND.n2887 GND.n2886 65.0005
R3715 GND.n2888 GND.n2887 65.0005
R3716 GND.n3462 GND.n3461 65.0005
R3717 GND.n3461 GND.n3460 65.0005
R3718 GND.n318 GND.n315 65.0005
R3719 GND.n318 GND.n308 65.0005
R3720 GND.n3451 GND.n3450 65.0005
R3721 GND.n3450 GND.n3449 65.0005
R3722 GND.n3458 GND.n3457 65.0005
R3723 GND.n3459 GND.n3458 65.0005
R3724 GND.n760 GND.n729 65.0005
R3725 GND.n759 GND.n729 65.0005
R3726 GND.n728 GND.n726 65.0005
R3727 GND.n728 GND.n680 65.0005
R3728 GND.n751 GND.n750 65.0005
R3729 GND.n750 GND.n749 65.0005
R3730 GND.n757 GND.n756 65.0005
R3731 GND.n758 GND.n757 65.0005
R3732 GND.n742 GND.n741 65.0005
R3733 GND.n741 GND.n679 65.0005
R3734 GND.n747 GND.n746 65.0005
R3735 GND.n748 GND.n747 65.0005
R3736 GND.n2113 GND.n2112 65.0005
R3737 GND.n2114 GND.n2113 65.0005
R3738 GND.n2105 GND.n2104 65.0005
R3739 GND.n2104 GND.n2103 65.0005
R3740 GND.n2125 GND.n2124 65.0005
R3741 GND.n2126 GND.n2125 65.0005
R3742 GND.n2117 GND.n2116 65.0005
R3743 GND.n2116 GND.n2115 65.0005
R3744 GND.n2137 GND.n2136 65.0005
R3745 GND.n2138 GND.n2137 65.0005
R3746 GND.n2129 GND.n2128 65.0005
R3747 GND.n2128 GND.n2127 65.0005
R3748 GND.n2141 GND.n2140 65.0005
R3749 GND.n2142 GND.n2141 65.0005
R3750 GND.n724 GND.n723 65.0005
R3751 GND.n723 GND.n681 65.0005
R3752 GND.n717 GND.n705 65.0005
R3753 GND.n717 GND.n716 65.0005
R3754 GND.n714 GND.n703 65.0005
R3755 GND.n714 GND.n713 65.0005
R3756 GND.n710 GND.n707 65.0005
R3757 GND.n715 GND.n710 65.0005
R3758 GND.n711 GND.n700 65.0005
R3759 GND.n712 GND.n711 65.0005
R3760 GND.n4344 GND.n4343 65.0005
R3761 GND.n4343 GND.n4342 65.0005
R3762 GND.n4360 GND.n4359 65.0005
R3763 GND.n4361 GND.n4360 65.0005
R3764 GND.n4357 GND.n4356 65.0005
R3765 GND.n4356 GND.n4355 65.0005
R3766 GND.n4335 GND.n4334 65.0005
R3767 GND.n4336 GND.n4335 65.0005
R3768 GND.n4323 GND.n26 65.0005
R3769 GND.n4324 GND.n4323 65.0005
R3770 GND.n4353 GND.n4352 65.0005
R3771 GND.n4354 GND.n4353 65.0005
R3772 GND.n4339 GND.n4338 65.0005
R3773 GND.n4340 GND.n4339 65.0005
R3774 GND.n3440 GND.n3439 65.0005
R3775 GND.n3439 GND.n3438 65.0005
R3776 GND.n3447 GND.n3446 65.0005
R3777 GND.n3448 GND.n3447 65.0005
R3778 GND.n3429 GND.n3428 65.0005
R3779 GND.n3428 GND.n3427 65.0005
R3780 GND.n3436 GND.n3435 65.0005
R3781 GND.n3437 GND.n3436 65.0005
R3782 GND.n3419 GND.n3418 65.0005
R3783 GND.n3418 GND.n3417 65.0005
R3784 GND.n3425 GND.n3424 65.0005
R3785 GND.n3426 GND.n3425 65.0005
R3786 GND.n3401 GND.n3393 65.0005
R3787 GND.n3402 GND.n3401 65.0005
R3788 GND.n3415 GND.n3414 65.0005
R3789 GND.n3416 GND.n3415 65.0005
R3790 GND.n3404 GND.n3400 65.0005
R3791 GND.n3400 GND.n192 65.0005
R3792 GND.n3399 GND.n3395 65.0005
R3793 GND.n3403 GND.n3399 65.0005
R3794 GND.n3893 GND.n3892 65.0005
R3795 GND.n3894 GND.n3893 65.0005
R3796 GND.n3885 GND.n3884 65.0005
R3797 GND.n3884 GND.n3883 65.0005
R3798 GND.n3948 GND.n187 65.0005
R3799 GND.n3947 GND.n187 65.0005
R3800 GND.n186 GND.n184 65.0005
R3801 GND.n3895 GND.n186 65.0005
R3802 GND.n3939 GND.n3938 65.0005
R3803 GND.n3938 GND.n3937 65.0005
R3804 GND.n3945 GND.n3944 65.0005
R3805 GND.n3946 GND.n3945 65.0005
R3806 GND.n3913 GND.n3907 65.0005
R3807 GND.n3914 GND.n3913 65.0005
R3808 GND.n3935 GND.n3934 65.0005
R3809 GND.n3936 GND.n3935 65.0005
R3810 GND.n3924 GND.n3912 65.0005
R3811 GND.n3923 GND.n3912 65.0005
R3812 GND.n3911 GND.n3909 65.0005
R3813 GND.n3915 GND.n3911 65.0005
R3814 GND.n4365 GND.n4364 65.0005
R3815 GND.n4364 GND.n4363 65.0005
R3816 GND.n3921 GND.n3920 65.0005
R3817 GND.n3922 GND.n3921 65.0005
R3818 GND.n3613 GND.n249 65.0005
R3819 GND.n3612 GND.n249 65.0005
R3820 GND.n248 GND.n245 65.0005
R3821 GND.n2101 GND.n248 65.0005
R3822 GND.n3595 GND.n3594 65.0005
R3823 GND.n3594 GND.n3593 65.0005
R3824 GND.n3609 GND.n3608 65.0005
R3825 GND.n3610 GND.n3609 65.0005
R3826 GND.n3575 GND.n3574 65.0005
R3827 GND.n3574 GND.n3573 65.0005
R3828 GND.n3590 GND.n3589 65.0005
R3829 GND.n3591 GND.n3590 65.0005
R3830 GND.n3556 GND.n3555 65.0005
R3831 GND.n3555 GND.n3554 65.0005
R3832 GND.n3570 GND.n3569 65.0005
R3833 GND.n3571 GND.n3570 65.0005
R3834 GND.n3534 GND.n3533 65.0005
R3835 GND.n3533 GND.n3532 65.0005
R3836 GND.n3551 GND.n3550 65.0005
R3837 GND.n3552 GND.n3551 65.0005
R3838 GND.n3512 GND.n3511 65.0005
R3839 GND.n3511 GND.n3510 65.0005
R3840 GND.n3529 GND.n3528 65.0005
R3841 GND.n3530 GND.n3529 65.0005
R3842 GND.n3493 GND.n3492 65.0005
R3843 GND.n3492 GND.n3491 65.0005
R3844 GND.n3507 GND.n3506 65.0005
R3845 GND.n3508 GND.n3507 65.0005
R3846 GND.n3880 GND.n3879 65.0005
R3847 GND.n3881 GND.n3880 65.0005
R3848 GND.n3488 GND.n3487 65.0005
R3849 GND.n3489 GND.n3488 65.0005
R3850 GND.n2096 GND.n684 65.0005
R3851 GND.n695 GND.n684 65.0005
R3852 GND.n685 GND.n683 65.0005
R3853 GND.n1086 GND.n683 65.0005
R3854 GND.n2085 GND.n694 65.0005
R3855 GND.n2084 GND.n694 65.0005
R3856 GND.n693 GND.n691 65.0005
R3857 GND.n696 GND.n693 65.0005
R3858 GND.n2082 GND.n2081 65.0005
R3859 GND.n2083 GND.n2082 65.0005
R3860 GND.n1092 GND.n1091 65.0005
R3861 GND.n1093 GND.n1092 65.0005
R3862 GND.n1089 GND.n1088 65.0005
R3863 GND.n1088 GND.n1087 65.0005
R3864 GND.n1097 GND.n1096 65.0005
R3865 GND.n1096 GND.n1095 65.0005
R3866 GND.n1037 GND.n1009 65.0005
R3867 GND.t58 GND.n1009 65.0005
R3868 GND.n1034 GND.n1008 65.0005
R3869 GND.t58 GND.n1008 65.0005
R3870 GND.n1050 GND.n1010 65.0005
R3871 GND.t58 GND.n1010 65.0005
R3872 GND.n1047 GND.n1007 65.0005
R3873 GND.t58 GND.n1007 65.0005
R3874 GND.n1060 GND.n1011 65.0005
R3875 GND.t58 GND.n1011 65.0005
R3876 GND.n1063 GND.n1062 65.0005
R3877 GND.t58 GND.n1063 65.0005
R3878 GND.n1026 GND.n1006 65.0005
R3879 GND.t58 GND.n1006 65.0005
R3880 GND.n1023 GND.n1005 65.0005
R3881 GND.t58 GND.n1005 65.0005
R3882 GND.n1066 GND.n1065 65.0005
R3883 GND.n1065 GND.t58 65.0005
R3884 GND.n1064 GND.n1001 65.0005
R3885 GND.t58 GND.n1064 65.0005
R3886 GND.n1111 GND.n1110 65.0005
R3887 GND.n1112 GND.n1111 65.0005
R3888 GND.n1117 GND.n1116 65.0005
R3889 GND.n1116 GND.n1115 65.0005
R3890 GND.n1159 GND.n1125 65.0005
R3891 GND.n1125 GND.n971 65.0005
R3892 GND.n1160 GND.n1126 65.0005
R3893 GND.n1140 GND.n1126 65.0005
R3894 GND.n1141 GND.n1135 65.0005
R3895 GND.n1142 GND.n1141 65.0005
R3896 GND.n1127 GND.n975 65.0005
R3897 GND.n1128 GND.n1127 65.0005
R3898 GND.n1170 GND.n1169 65.0005
R3899 GND.n1171 GND.n1170 65.0005
R3900 GND.n1143 GND.n1132 65.0005
R3901 GND.n1144 GND.n1143 65.0005
R3902 GND.n1157 GND.n1156 65.0005
R3903 GND.n1158 GND.n1157 65.0005
R3904 GND.n1148 GND.n1147 65.0005
R3905 GND.n1147 GND.n1146 65.0005
R3906 GND.n2057 GND.n772 65.0005
R3907 GND.n2056 GND.n772 65.0005
R3908 GND.n771 GND.n769 65.0005
R3909 GND.n1145 GND.n771 65.0005
R3910 GND.n2054 GND.n2053 65.0005
R3911 GND.n2055 GND.n2054 65.0005
R3912 GND.n2037 GND.n801 65.0005
R3913 GND.n2036 GND.n801 65.0005
R3914 GND.n800 GND.n798 65.0005
R3915 GND.n800 GND.n780 65.0005
R3916 GND.n2034 GND.n2033 65.0005
R3917 GND.n2035 GND.n2034 65.0005
R3918 GND.n2031 GND.n2030 65.0005
R3919 GND.n2030 GND.n2029 65.0005
R3920 GND.n2027 GND.n2026 65.0005
R3921 GND.n2028 GND.n2027 65.0005
R3922 GND.n852 GND.n851 65.0005
R3923 GND.n853 GND.n852 65.0005
R3924 GND.n839 GND.n838 65.0005
R3925 GND.n838 GND.n803 65.0005
R3926 GND.n858 GND.n857 65.0005
R3927 GND.n857 GND.n809 65.0005
R3928 GND.n855 GND.n834 65.0005
R3929 GND.n855 GND.n854 65.0005
R3930 GND.n2024 GND.n2023 65.0005
R3931 GND.n2023 GND.n2022 65.0005
R3932 GND.n2017 GND.n2016 65.0005
R3933 GND.n2016 GND.n2015 65.0005
R3934 GND.n2020 GND.n2019 65.0005
R3935 GND.n2021 GND.n2020 65.0005
R3936 GND.n2013 GND.n2012 65.0005
R3937 GND.n2014 GND.n2013 65.0005
R3938 GND.n2010 GND.n2009 65.0005
R3939 GND.n2009 GND.n2008 65.0005
R3940 GND.n2006 GND.n2005 65.0005
R3941 GND.n2007 GND.n2006 65.0005
R3942 GND.n873 GND.n872 65.0005
R3943 GND.n1947 GND.n1901 65.0005
R3944 GND.t41 GND.n1901 65.0005
R3945 GND.n1944 GND.n1900 65.0005
R3946 GND.t41 GND.n1900 65.0005
R3947 GND.n1943 GND.n1942 65.0005
R3948 GND.n1942 GND.t83 65.0005
R3949 GND.n1914 GND.n1913 65.0005
R3950 GND.n1914 GND.t83 65.0005
R3951 GND.n1961 GND.n1960 65.0005
R3952 GND.t41 GND.n1961 65.0005
R3953 GND.n1923 GND.n1899 65.0005
R3954 GND.t41 GND.n1899 65.0005
R3955 GND.n1922 GND.n1905 65.0005
R3956 GND.n1922 GND.t83 65.0005
R3957 GND.n1929 GND.n1921 65.0005
R3958 GND.n1921 GND.t83 65.0005
R3959 GND.n1970 GND.n1969 65.0005
R3960 GND.n1969 GND.t41 65.0005
R3961 GND.n1962 GND.n1888 65.0005
R3962 GND.t41 GND.n1962 65.0005
R3963 GND.n1898 GND.n1897 65.0005
R3964 GND.t41 GND.n1898 65.0005
R3965 GND.n1895 GND.n1893 65.0005
R3966 GND.t41 GND.n1893 65.0005
R3967 GND.n1935 GND.n1933 65.0005
R3968 GND.n1933 GND.t83 65.0005
R3969 GND.n1934 GND.n1932 65.0005
R3970 GND.n1932 GND.t83 65.0005
R3971 GND.n1965 GND.n1963 65.0005
R3972 GND.t41 GND.n1963 65.0005
R3973 GND.n1968 GND.n1967 65.0005
R3974 GND.t41 GND.n1968 65.0005
R3975 GND.n1918 GND.n1916 65.0005
R3976 GND.n1916 GND.t83 65.0005
R3977 GND.n1917 GND.n1915 65.0005
R3978 GND.n1915 GND.t83 65.0005
R3979 GND.n893 GND.n891 65.0005
R3980 GND.n891 GND.t83 65.0005
R3981 GND.n892 GND.n890 65.0005
R3982 GND.n890 GND.t83 65.0005
R3983 GND.n1996 GND.n884 65.0005
R3984 GND.n1995 GND.n884 65.0005
R3985 GND.n883 GND.n879 65.0005
R3986 GND.n1993 GND.n883 65.0005
R3987 GND.n2282 GND.n633 65.0005
R3988 GND.n633 GND.n624 65.0005
R3989 GND.n2283 GND.n634 65.0005
R3990 GND.n2263 GND.n634 65.0005
R3991 GND.n2264 GND.n2258 65.0005
R3992 GND.n2265 GND.n2264 65.0005
R3993 GND.n635 GND.n628 65.0005
R3994 GND.n636 GND.n635 65.0005
R3995 GND.n2293 GND.n2292 65.0005
R3996 GND.n2294 GND.n2293 65.0005
R3997 GND.n2266 GND.n640 65.0005
R3998 GND.n2267 GND.n2266 65.0005
R3999 GND.n2280 GND.n2279 65.0005
R4000 GND.n2281 GND.n2280 65.0005
R4001 GND.n2271 GND.n2270 65.0005
R4002 GND.n2270 GND.n2269 65.0005
R4003 GND.n2300 GND.n2299 65.0005
R4004 GND.n2299 GND.n614 65.0005
R4005 GND.n643 GND.n621 65.0005
R4006 GND.n2268 GND.n621 65.0005
R4007 GND.n2314 GND.n2313 65.0005
R4008 GND.n2313 GND.n2312 65.0005
R4009 GND.n1681 GND.n1650 65.0005
R4010 GND.t140 GND.n1650 65.0005
R4011 GND.n1678 GND.n1649 65.0005
R4012 GND.t140 GND.n1649 65.0005
R4013 GND.n1677 GND.n1628 65.0005
R4014 GND.t30 GND.n1628 65.0005
R4015 GND.n1674 GND.n1627 65.0005
R4016 GND.t30 GND.n1627 65.0005
R4017 GND.n1695 GND.n1694 65.0005
R4018 GND.t140 GND.n1695 65.0005
R4019 GND.n1660 GND.n1648 65.0005
R4020 GND.t140 GND.n1648 65.0005
R4021 GND.n1656 GND.n1630 65.0005
R4022 GND.t30 GND.n1630 65.0005
R4023 GND.n1663 GND.n1626 65.0005
R4024 GND.t30 GND.n1626 65.0005
R4025 GND.n1724 GND.n1723 65.0005
R4026 GND.n1723 GND.t140 65.0005
R4027 GND.n1696 GND.n1638 65.0005
R4028 GND.t140 GND.n1696 65.0005
R4029 GND.n1647 GND.n1635 65.0005
R4030 GND.t140 GND.n1647 65.0005
R4031 GND.n1644 GND.n1643 65.0005
R4032 GND.t140 GND.n1643 65.0005
R4033 GND.n1732 GND.n1631 65.0005
R4034 GND.t30 GND.n1631 65.0005
R4035 GND.n1735 GND.n1734 65.0005
R4036 GND.t30 GND.n1735 65.0005
R4037 GND.n1702 GND.n1697 65.0005
R4038 GND.t140 GND.n1697 65.0005
R4039 GND.n1722 GND.n1721 65.0005
R4040 GND.t140 GND.n1722 65.0005
R4041 GND.n1716 GND.n1625 65.0005
R4042 GND.t30 GND.n1625 65.0005
R4043 GND.n1719 GND.n1624 65.0005
R4044 GND.t30 GND.n1624 65.0005
R4045 GND.n1738 GND.n1737 65.0005
R4046 GND.n1737 GND.t30 65.0005
R4047 GND.n1736 GND.n1619 65.0005
R4048 GND.t30 GND.n1736 65.0005
R4049 GND.n2423 GND.n597 65.0005
R4050 GND.t73 GND.n597 65.0005
R4051 GND.n2420 GND.n596 65.0005
R4052 GND.t73 GND.n596 65.0005
R4053 GND.n2419 GND.n575 65.0005
R4054 GND.t8 GND.n575 65.0005
R4055 GND.n2416 GND.n574 65.0005
R4056 GND.t8 GND.n574 65.0005
R4057 GND.n2437 GND.n2436 65.0005
R4058 GND.t73 GND.n2437 65.0005
R4059 GND.n2402 GND.n595 65.0005
R4060 GND.t73 GND.n595 65.0005
R4061 GND.n2398 GND.n577 65.0005
R4062 GND.t8 GND.n577 65.0005
R4063 GND.n2405 GND.n573 65.0005
R4064 GND.t8 GND.n573 65.0005
R4065 GND.n2466 GND.n2465 65.0005
R4066 GND.n2465 GND.t73 65.0005
R4067 GND.n2438 GND.n585 65.0005
R4068 GND.t73 GND.n2438 65.0005
R4069 GND.n594 GND.n582 65.0005
R4070 GND.t73 GND.n594 65.0005
R4071 GND.n591 GND.n590 65.0005
R4072 GND.t73 GND.n590 65.0005
R4073 GND.n2474 GND.n578 65.0005
R4074 GND.t8 GND.n578 65.0005
R4075 GND.n2477 GND.n2476 65.0005
R4076 GND.t8 GND.n2477 65.0005
R4077 GND.n2444 GND.n2439 65.0005
R4078 GND.t73 GND.n2439 65.0005
R4079 GND.n2464 GND.n2463 65.0005
R4080 GND.t73 GND.n2464 65.0005
R4081 GND.n2458 GND.n572 65.0005
R4082 GND.t8 GND.n572 65.0005
R4083 GND.n2461 GND.n571 65.0005
R4084 GND.t8 GND.n571 65.0005
R4085 GND.n2480 GND.n2479 65.0005
R4086 GND.n2479 GND.t8 65.0005
R4087 GND.n2478 GND.n566 65.0005
R4088 GND.t8 GND.n2478 65.0005
R4089 GND.n2329 GND.n602 65.0005
R4090 GND.n2340 GND.n602 65.0005
R4091 GND.n2327 GND.n601 65.0005
R4092 GND.n2319 GND.n601 65.0005
R4093 GND.n2335 GND.n2331 65.0005
R4094 GND.n2341 GND.n2335 65.0005
R4095 GND.n2380 GND.n2336 65.0005
R4096 GND.n2354 GND.n2336 65.0005
R4097 GND.n2361 GND.n2359 65.0005
R4098 GND.n2359 GND.n2355 65.0005
R4099 GND.n2347 GND.n2346 65.0005
R4100 GND.n2348 GND.n2347 65.0005
R4101 GND.n2344 GND.n2343 65.0005
R4102 GND.n2343 GND.n2342 65.0005
R4103 GND.n2370 GND.n2369 65.0005
R4104 GND.n2369 GND.n2368 65.0005
R4105 GND.n2378 GND.n2377 65.0005
R4106 GND.n2379 GND.n2378 65.0005
R4107 GND.n2363 GND.n2360 65.0005
R4108 GND.n2360 GND.n2357 65.0005
R4109 GND.n2819 GND.n525 65.0005
R4110 GND.n2818 GND.n525 65.0005
R4111 GND.n524 GND.n522 65.0005
R4112 GND.n2356 GND.n524 65.0005
R4113 GND.n2816 GND.n2815 65.0005
R4114 GND.n2817 GND.n2816 65.0005
R4115 GND.n2813 GND.n2812 65.0005
R4116 GND.n2812 GND.n2811 65.0005
R4117 GND.n2809 GND.n2808 65.0005
R4118 GND.n2810 GND.n2809 65.0005
R4119 GND.n545 GND.n544 65.0005
R4120 GND.n2693 GND.n2647 65.0005
R4121 GND.t44 GND.n2647 65.0005
R4122 GND.n2690 GND.n2646 65.0005
R4123 GND.t44 GND.n2646 65.0005
R4124 GND.n2689 GND.n2688 65.0005
R4125 GND.n2688 GND.t32 65.0005
R4126 GND.n2660 GND.n2659 65.0005
R4127 GND.n2660 GND.t32 65.0005
R4128 GND.n2707 GND.n2706 65.0005
R4129 GND.t44 GND.n2707 65.0005
R4130 GND.n2669 GND.n2645 65.0005
R4131 GND.t44 GND.n2645 65.0005
R4132 GND.n2668 GND.n2651 65.0005
R4133 GND.n2668 GND.t32 65.0005
R4134 GND.n2675 GND.n2667 65.0005
R4135 GND.n2667 GND.t32 65.0005
R4136 GND.n2716 GND.n2715 65.0005
R4137 GND.n2715 GND.t44 65.0005
R4138 GND.n2708 GND.n2634 65.0005
R4139 GND.t44 GND.n2708 65.0005
R4140 GND.n2644 GND.n2643 65.0005
R4141 GND.t44 GND.n2644 65.0005
R4142 GND.n2641 GND.n2639 65.0005
R4143 GND.t44 GND.n2639 65.0005
R4144 GND.n2681 GND.n2679 65.0005
R4145 GND.n2679 GND.t32 65.0005
R4146 GND.n2680 GND.n2678 65.0005
R4147 GND.n2678 GND.t32 65.0005
R4148 GND.n2711 GND.n2709 65.0005
R4149 GND.t44 GND.n2709 65.0005
R4150 GND.n2714 GND.n2713 65.0005
R4151 GND.t44 GND.n2714 65.0005
R4152 GND.n2664 GND.n2662 65.0005
R4153 GND.n2662 GND.t32 65.0005
R4154 GND.n2663 GND.n2661 65.0005
R4155 GND.n2661 GND.t32 65.0005
R4156 GND.n564 GND.n562 65.0005
R4157 GND.n562 GND.t32 65.0005
R4158 GND.n563 GND.n561 65.0005
R4159 GND.n561 GND.t32 65.0005
R4160 GND.n2799 GND.n554 65.0005
R4161 GND.n2797 GND.n554 65.0005
R4162 GND.n553 GND.n551 65.0005
R4163 GND.n555 GND.n553 65.0005
R4164 GND.n2795 GND.n2794 65.0005
R4165 GND.n2796 GND.n2795 65.0005
R4166 GND.n2977 GND.n484 65.0005
R4167 GND.t7 GND.n484 65.0005
R4168 GND.n2974 GND.n483 65.0005
R4169 GND.t7 GND.n483 65.0005
R4170 GND.n2973 GND.n462 65.0005
R4171 GND.t39 GND.n462 65.0005
R4172 GND.n2970 GND.n461 65.0005
R4173 GND.t39 GND.n461 65.0005
R4174 GND.n2991 GND.n2990 65.0005
R4175 GND.t7 GND.n2991 65.0005
R4176 GND.n2956 GND.n482 65.0005
R4177 GND.t7 GND.n482 65.0005
R4178 GND.n2952 GND.n464 65.0005
R4179 GND.t39 GND.n464 65.0005
R4180 GND.n2959 GND.n460 65.0005
R4181 GND.t39 GND.n460 65.0005
R4182 GND.n3020 GND.n3019 65.0005
R4183 GND.n3019 GND.t7 65.0005
R4184 GND.n2992 GND.n472 65.0005
R4185 GND.t7 GND.n2992 65.0005
R4186 GND.n481 GND.n469 65.0005
R4187 GND.t7 GND.n481 65.0005
R4188 GND.n478 GND.n477 65.0005
R4189 GND.t7 GND.n477 65.0005
R4190 GND.n3028 GND.n465 65.0005
R4191 GND.t39 GND.n465 65.0005
R4192 GND.n3031 GND.n3030 65.0005
R4193 GND.t39 GND.n3031 65.0005
R4194 GND.n2998 GND.n2993 65.0005
R4195 GND.t7 GND.n2993 65.0005
R4196 GND.n3018 GND.n3017 65.0005
R4197 GND.t7 GND.n3018 65.0005
R4198 GND.n3012 GND.n459 65.0005
R4199 GND.t39 GND.n459 65.0005
R4200 GND.n3015 GND.n458 65.0005
R4201 GND.t39 GND.n458 65.0005
R4202 GND.n3034 GND.n3033 65.0005
R4203 GND.n3033 GND.t39 65.0005
R4204 GND.n3032 GND.n453 65.0005
R4205 GND.t39 GND.n3032 65.0005
R4206 GND.n2785 GND.n2784 65.0005
R4207 GND.n2784 GND.n2783 65.0005
R4208 GND.n2903 GND.n489 65.0005
R4209 GND.n2914 GND.n489 65.0005
R4210 GND.n2901 GND.n488 65.0005
R4211 GND.n2782 GND.n488 65.0005
R4212 GND.n2907 GND.n2905 65.0005
R4213 GND.n2915 GND.n2907 65.0005
R4214 GND.n2909 GND.n2908 65.0005
R4215 GND.n2913 GND.n2908 65.0005
R4216 GND.n2932 GND.n2918 65.0005
R4217 GND.n2918 GND.n356 65.0005
R4218 GND.n2919 GND.n2917 65.0005
R4219 GND.n3339 GND.n3338 65.0005
R4220 GND.n3340 GND.n3339 65.0005
R4221 GND.n3336 GND.n3335 65.0005
R4222 GND.n3335 GND.n3334 65.0005
R4223 GND.n3345 GND.n3344 65.0005
R4224 GND.n3344 GND.n3343 65.0005
R4225 GND.n442 GND.n441 65.0005
R4226 GND.n442 GND.t92 65.0005
R4227 GND.n434 GND.n432 65.0005
R4228 GND.n432 GND.t92 65.0005
R4229 GND.n439 GND.n389 65.0005
R4230 GND.n389 GND.t9 65.0005
R4231 GND.n436 GND.n388 65.0005
R4232 GND.n388 GND.t9 65.0005
R4233 GND.n422 GND.n421 65.0005
R4234 GND.n421 GND.t92 65.0005
R4235 GND.n410 GND.n408 65.0005
R4236 GND.n408 GND.t92 65.0005
R4237 GND.n412 GND.n406 65.0005
R4238 GND.n412 GND.t9 65.0005
R4239 GND.n415 GND.n414 65.0005
R4240 GND.n414 GND.t9 65.0005
R4241 GND.n399 GND.n398 65.0005
R4242 GND.n398 GND.t92 65.0005
R4243 GND.n395 GND.n394 65.0005
R4244 GND.n395 GND.t92 65.0005
R4245 GND.n378 GND.n377 65.0005
R4246 GND.n377 GND.t92 65.0005
R4247 GND.n375 GND.n374 65.0005
R4248 GND.n374 GND.t92 65.0005
R4249 GND.n383 GND.n382 65.0005
R4250 GND.t9 GND.n383 65.0005
R4251 GND.n380 GND.n372 65.0005
R4252 GND.t9 GND.n372 65.0005
R4253 GND.n3329 GND.n363 65.0005
R4254 GND.n363 GND.t92 65.0005
R4255 GND.n364 GND.n362 65.0005
R4256 GND.n362 GND.t92 65.0005
R4257 GND.n3307 GND.n365 65.0005
R4258 GND.n3307 GND.t9 65.0005
R4259 GND.n3310 GND.n3309 65.0005
R4260 GND.n3309 GND.t9 65.0005
R4261 GND.n451 GND.n447 65.0005
R4262 GND.n447 GND.t9 65.0005
R4263 GND.n448 GND.n446 65.0005
R4264 GND.n446 GND.t9 65.0005
R4265 GND.n3234 GND.n3205 65.0005
R4266 GND.t24 GND.n3205 65.0005
R4267 GND.n3231 GND.n3204 65.0005
R4268 GND.t24 GND.n3204 65.0005
R4269 GND.n3230 GND.n3182 65.0005
R4270 GND.t36 GND.n3182 65.0005
R4271 GND.n3227 GND.n3181 65.0005
R4272 GND.t36 GND.n3181 65.0005
R4273 GND.n3248 GND.n3247 65.0005
R4274 GND.t24 GND.n3248 65.0005
R4275 GND.n3213 GND.n3203 65.0005
R4276 GND.t24 GND.n3203 65.0005
R4277 GND.n3209 GND.n3184 65.0005
R4278 GND.t36 GND.n3184 65.0005
R4279 GND.n3216 GND.n3180 65.0005
R4280 GND.t36 GND.n3180 65.0005
R4281 GND.n3277 GND.n3276 65.0005
R4282 GND.n3276 GND.t24 65.0005
R4283 GND.n3249 GND.n3192 65.0005
R4284 GND.t24 GND.n3249 65.0005
R4285 GND.n3202 GND.n3189 65.0005
R4286 GND.t24 GND.n3202 65.0005
R4287 GND.n3198 GND.n3197 65.0005
R4288 GND.t24 GND.n3197 65.0005
R4289 GND.n3285 GND.n3185 65.0005
R4290 GND.t36 GND.n3185 65.0005
R4291 GND.n3288 GND.n3287 65.0005
R4292 GND.t36 GND.n3288 65.0005
R4293 GND.n3255 GND.n3250 65.0005
R4294 GND.t24 GND.n3250 65.0005
R4295 GND.n3275 GND.n3274 65.0005
R4296 GND.t24 GND.n3275 65.0005
R4297 GND.n3269 GND.n3179 65.0005
R4298 GND.t36 GND.n3179 65.0005
R4299 GND.n3272 GND.n3178 65.0005
R4300 GND.t36 GND.n3178 65.0005
R4301 GND.n3291 GND.n3290 65.0005
R4302 GND.n3290 GND.t36 65.0005
R4303 GND.n3289 GND.n3174 65.0005
R4304 GND.t36 GND.n3289 65.0005
R4305 GND.n337 GND.n335 65.0005
R4306 GND.n3373 GND.n337 65.0005
R4307 GND.n102 GND.n97 65.0005
R4308 GND.n112 GND.n97 65.0005
R4309 GND.n100 GND.n96 65.0005
R4310 GND.n3372 GND.n96 65.0005
R4311 GND.n106 GND.n104 65.0005
R4312 GND.n113 GND.n106 65.0005
R4313 GND.n108 GND.n107 65.0005
R4314 GND.n126 GND.n107 65.0005
R4315 GND.n3981 GND.n116 65.0005
R4316 GND.n127 GND.n116 65.0005
R4317 GND.n117 GND.n115 65.0005
R4318 GND.n3974 GND.n132 65.0005
R4319 GND.n3974 GND.n3973 65.0005
R4320 GND.n129 GND.n124 65.0005
R4321 GND.n129 GND.n128 65.0005
R4322 GND.n3971 GND.n3970 65.0005
R4323 GND.n3972 GND.n3971 65.0005
R4324 GND.n4157 GND.n4126 65.0005
R4325 GND.t75 GND.n4126 65.0005
R4326 GND.n4154 GND.n4125 65.0005
R4327 GND.t75 GND.n4125 65.0005
R4328 GND.n4153 GND.n4104 65.0005
R4329 GND.t53 GND.n4104 65.0005
R4330 GND.n4150 GND.n4103 65.0005
R4331 GND.t53 GND.n4103 65.0005
R4332 GND.n4171 GND.n4170 65.0005
R4333 GND.t75 GND.n4171 65.0005
R4334 GND.n4136 GND.n4124 65.0005
R4335 GND.t75 GND.n4124 65.0005
R4336 GND.n4132 GND.n4106 65.0005
R4337 GND.t53 GND.n4106 65.0005
R4338 GND.n4139 GND.n4102 65.0005
R4339 GND.t53 GND.n4102 65.0005
R4340 GND.n4200 GND.n4199 65.0005
R4341 GND.n4199 GND.t75 65.0005
R4342 GND.n4172 GND.n4114 65.0005
R4343 GND.t75 GND.n4172 65.0005
R4344 GND.n4123 GND.n4111 65.0005
R4345 GND.t75 GND.n4123 65.0005
R4346 GND.n4120 GND.n4119 65.0005
R4347 GND.t75 GND.n4119 65.0005
R4348 GND.n4208 GND.n4107 65.0005
R4349 GND.t53 GND.n4107 65.0005
R4350 GND.n4211 GND.n4210 65.0005
R4351 GND.t53 GND.n4211 65.0005
R4352 GND.n4178 GND.n4173 65.0005
R4353 GND.t75 GND.n4173 65.0005
R4354 GND.n4198 GND.n4197 65.0005
R4355 GND.t75 GND.n4198 65.0005
R4356 GND.n4192 GND.n4101 65.0005
R4357 GND.t53 GND.n4101 65.0005
R4358 GND.n4195 GND.n4100 65.0005
R4359 GND.t53 GND.n4100 65.0005
R4360 GND.n4214 GND.n4213 65.0005
R4361 GND.n4213 GND.t53 65.0005
R4362 GND.n4212 GND.n4095 65.0005
R4363 GND.t53 GND.n4212 65.0005
R4364 GND.n3961 GND.n3960 65.0005
R4365 GND.n3960 GND.n48 65.0005
R4366 GND.n4294 GND.n4293 65.0005
R4367 GND.n4295 GND.n4294 65.0005
R4368 GND.n4291 GND.n4290 65.0005
R4369 GND.n4290 GND.n4289 65.0005
R4370 GND.n175 GND.n40 65.0005
R4371 GND.n4296 GND.n40 65.0005
R4372 GND.n4302 GND.n4301 65.0005
R4373 GND.n4301 GND.n31 65.0005
R4374 GND.n4314 GND.n4313 65.0005
R4375 GND.n4315 GND.n4314 65.0005
R4376 GND.n43 GND.n42 65.0005
R4377 GND.n4321 GND.n4320 65.0005
R4378 GND.n4322 GND.n4321 65.0005
R4379 GND.n4318 GND.n4317 65.0005
R4380 GND.n4317 GND.n4316 65.0005
R4381 GND.n4327 GND.n4326 65.0005
R4382 GND.n4326 GND.n4325 65.0005
R4383 GND.n4265 GND.n4264 65.0005
R4384 GND.n4264 GND.t88 65.0005
R4385 GND.n4262 GND.n4261 65.0005
R4386 GND.n4261 GND.t88 65.0005
R4387 GND.n4253 GND.n4252 65.0005
R4388 GND.n4252 GND.t88 65.0005
R4389 GND.n4250 GND.n4249 65.0005
R4390 GND.n4249 GND.t88 65.0005
R4391 GND.n4235 GND.n4234 65.0005
R4392 GND.n4235 GND.t88 65.0005
R4393 GND.n4232 GND.n4230 65.0005
R4394 GND.n4232 GND.t88 65.0005
R4395 GND.n4284 GND.n55 65.0005
R4396 GND.n55 GND.t88 65.0005
R4397 GND.n56 GND.n54 65.0005
R4398 GND.n54 GND.t88 65.0005
R4399 GND.n4242 GND.n4239 65.0005
R4400 GND.n4239 GND.t88 65.0005
R4401 GND.n4244 GND.n4240 65.0005
R4402 GND.n4240 GND.t88 65.0005
R4403 GND.n3901 GND.t692 61.1579
R4404 GND.n3902 GND.t77 61.1579
R4405 GND.n3931 GND.t244 61.1579
R4406 GND.n3917 GND.t191 61.1579
R4407 GND.n4368 GND.t103 61.1579
R4408 GND.n3383 GND.t600 61.1579
R4409 GND.n3388 GND.t196 61.1579
R4410 GND.n3411 GND.t179 61.1579
R4411 GND.n3396 GND.t332 61.1579
R4412 GND.n3889 GND.t283 61.1579
R4413 GND.n494 GND.t696 61.1579
R4414 GND.n3465 GND.t608 61.1579
R4415 GND.n314 GND.t301 61.1579
R4416 GND.n324 GND.t330 61.1579
R4417 GND.n329 GND.t577 61.1579
R4418 GND.n2834 GND.t511 61.1579
R4419 GND.n2852 GND.t68 61.1579
R4420 GND.n2853 GND.t35 61.1579
R4421 GND.n2865 GND.t698 61.1579
R4422 GND.n2877 GND.t160 61.1579
R4423 GND.n2190 GND.t688 61.1579
R4424 GND.n2191 GND.t648 61.1579
R4425 GND.n2231 GND.t516 61.1579
R4426 GND.n2210 GND.t603 61.1579
R4427 GND.n2211 GND.t175 61.1579
R4428 GND.n735 GND.t189 61.1579
R4429 GND.n736 GND.t113 61.1579
R4430 GND.n743 GND.t6 61.1579
R4431 GND.n2109 GND.t334 61.1579
R4432 GND.n2121 GND.t314 61.1579
R4433 GND.n2133 GND.t165 61.1579
R4434 GND.n2151 GND.t716 61.1579
R4435 GND.n2152 GND.t658 61.1579
R4436 GND.n2164 GND.t694 61.1579
R4437 GND.n2176 GND.t116 61.1579
R4438 GND.n2093 GND.t711 61.1579
R4439 GND.n701 GND.t145 61.1579
R4440 GND.n2078 GND.t263 61.1579
R4441 GND.n2072 GND.t708 61.1579
R4442 GND.n2066 GND.t641 61.1579
R4443 GND.n1079 GND.t148 61.1579
R4444 GND.n1166 GND.t665 61.1579
R4445 GND.n1151 GND.t643 61.1579
R4446 GND.n790 GND.t101 61.1579
R4447 GND.n848 GND.t573 61.1579
R4448 GND.n861 GND.t218 61.1579
R4449 GND.n871 GND.t20 61.1579
R4450 GND.n2289 GND.t513 61.1579
R4451 GND.n2274 GND.t126 61.1579
R4452 GND.n2305 GND.t325 61.1579
R4453 GND.n2332 GND.t353 61.1579
R4454 GND.n2364 GND.t351 61.1579
R4455 GND.n543 GND.t226 61.1579
R4456 GND.n2766 GND.t307 61.1579
R4457 GND.n2779 GND.t681 61.1579
R4458 GND.n2904 GND.t27 61.1579
R4459 GND.n3349 GND.t322 61.1579
R4460 GND.n3366 GND.t359 61.1579
R4461 GND.n103 GND.t679 61.1579
R4462 GND.n160 GND.t345 61.1579
R4463 GND.n173 GND.t343 61.1579
R4464 GND.n174 GND.t271 61.1579
R4465 GND.n4331 GND.t152 61.1579
R4466 GND.n4349 GND.t616 61.1579
R4467 GND.n4 GND.t253 61.1579
R4468 GND.n4347 GND.t336 61.1579
R4469 GND.n4306 GND.t720 61.1579
R4470 GND.n4305 GND.t130 61.1579
R4471 GND.n178 GND.t105 61.1579
R4472 GND.n3957 GND.t12 61.1579
R4473 GND.n142 GND.t167 61.1579
R4474 GND.n153 GND.t60 61.1579
R4475 GND.n122 GND.t98 61.1579
R4476 GND.n3990 GND.t285 61.1579
R4477 GND.n3379 GND.t249 61.1579
R4478 GND.n3365 GND.t280 61.1579
R4479 GND.n2925 GND.t347 61.1579
R4480 GND.n2924 GND.t52 61.1579
R4481 GND.n2941 GND.t289 61.1579
R4482 GND.n491 GND.t14 61.1579
R4483 GND.n2747 GND.t163 61.1579
R4484 GND.n2759 GND.t172 61.1579
R4485 GND.n549 GND.t216 61.1579
R4486 GND.n541 GND.t255 61.1579
R4487 GND.n520 GND.t109 61.1579
R4488 GND.n2373 GND.t278 61.1579
R4489 GND.n2387 GND.t592 61.1579
R4490 GND.n604 GND.t363 61.1579
R4491 GND.n2303 GND.t595 61.1579
R4492 GND.n2257 GND.t598 61.1579
R4493 GND.n642 GND.t690 61.1579
R4494 GND.n880 GND.t582 61.1579
R4495 GND.n877 GND.t2 61.1579
R4496 GND.n869 GND.t118 61.1579
R4497 GND.n863 GND.t16 61.1579
R4498 GND.n830 GND.t187 61.1579
R4499 GND.n841 GND.t654 61.1579
R4500 GND.n796 GND.t258 61.1579
R4501 GND.n788 GND.t656 61.1579
R4502 GND.n767 GND.t18 61.1579
R4503 GND.n1134 GND.t237 61.1579
R4504 GND.n1120 GND.t274 61.1579
R4505 GND.n985 GND.t319 61.1579
R4506 GND.n1081 GND.t276 61.1579
R4507 GND.n244 GND.t298 61.1525
R4508 GND.n3605 GND.t685 61.1525
R4509 GND.n3586 GND.t183 61.1525
R4510 GND.n3566 GND.t170 61.1525
R4511 GND.n3525 GND.t652 61.1525
R4512 GND.n3503 GND.t247 61.1525
R4513 GND.n3484 GND.t87 61.1525
R4514 GND.n3545 GND.t611 61.128
R4515 GND.n4225 GND.t234 60.3943
R4516 GND.n4280 GND.t539 60.3943
R4517 GND.n4248 GND.t623 60.3943
R4518 GND.n4257 GND.t583 60.3943
R4519 GND.n4269 GND.t547 60.3943
R4520 GND.n4036 GND.t670 60.3943
R4521 GND.n4036 GND.t554 60.3943
R4522 GND.n4006 GND.t606 60.3943
R4523 GND.n4006 GND.t38 60.3943
R4524 GND.n4074 GND.t94 60.3943
R4525 GND.n4058 GND.t709 60.3943
R4526 GND.n4058 GND.t551 60.3943
R4527 GND.n4053 GND.t552 60.3943
R4528 GND.n4053 GND.t207 60.3943
R4529 GND.n4088 GND.t204 60.3943
R4530 GND.n427 GND.t633 60.3943
R4531 GND.n427 GND.t536 60.3943
R4532 GND.n403 GND.t10 60.3943
R4533 GND.n403 GND.t193 60.3943
R4534 GND.n393 GND.t142 60.3943
R4535 GND.n3324 GND.t671 60.3943
R4536 GND.n3324 GND.t522 60.3943
R4537 GND.n3314 GND.t559 60.3943
R4538 GND.n3314 GND.t205 60.3943
R4539 GND.n3305 GND.t61 60.3943
R4540 GND.n3114 GND.t63 60.3943
R4541 GND.n3114 GND.t528 60.3943
R4542 GND.n3084 GND.t326 60.3943
R4543 GND.n3084 GND.t78 60.3943
R4544 GND.n3152 GND.t81 60.3943
R4545 GND.n3136 GND.t206 60.3943
R4546 GND.n3136 GND.t587 60.3943
R4547 GND.n3131 GND.t563 60.3943
R4548 GND.n3131 GND.t212 60.3943
R4549 GND.n3166 GND.t617 60.3943
R4550 GND.n2561 GND.t662 60.3943
R4551 GND.n2561 GND.t546 60.3943
R4552 GND.n2531 GND.t303 60.3943
R4553 GND.n2531 GND.t635 60.3943
R4554 GND.n2599 GND.t80 60.3943
R4555 GND.n2583 GND.t239 60.3943
R4556 GND.n2583 GND.t532 60.3943
R4557 GND.n2578 GND.t533 60.3943
R4558 GND.n2578 GND.t209 60.3943
R4559 GND.n2613 GND.t173 60.3943
R4560 GND.n1816 GND.t354 60.3943
R4561 GND.n1816 GND.t534 60.3943
R4562 GND.n1786 GND.t267 60.3943
R4563 GND.n1786 GND.t604 60.3943
R4564 GND.n1854 GND.t139 60.3943
R4565 GND.n1838 GND.t700 60.3943
R4566 GND.n1838 GND.t519 60.3943
R4567 GND.n1833 GND.t529 60.3943
R4568 GND.n1833 GND.t341 60.3943
R4569 GND.n1868 GND.t23 60.3943
R4570 GND.n1559 GND.t260 60.3943
R4571 GND.n1559 GND.t524 60.3943
R4572 GND.n1529 GND.t349 60.3943
R4573 GND.n1529 GND.t327 60.3943
R4574 GND.n1597 GND.t91 60.3943
R4575 GND.n1581 GND.t627 60.3943
R4576 GND.n1581 GND.t564 60.3943
R4577 GND.n1576 GND.t518 60.3943
R4578 GND.n1576 GND.t628 60.3943
R4579 GND.n1611 GND.t590 60.3943
R4580 GND.n1211 GND.t620 60.3943
R4581 GND.n1211 GND.t631 60.3943
R4582 GND.n1181 GND.t199 60.3943
R4583 GND.n1181 GND.t644 60.3943
R4584 GND.n1249 GND.t123 60.3943
R4585 GND.n1233 GND.t705 60.3943
R4586 GND.n1233 GND.t233 60.3943
R4587 GND.n1228 GND.t561 60.3943
R4588 GND.n1228 GND.t558 60.3943
R4589 GND.n1263 GND.t161 60.3943
R4590 GND.n1341 GND.t240 60.3943
R4591 GND.n1341 GND.t549 60.3943
R4592 GND.n1311 GND.t360 60.3943
R4593 GND.n1311 GND.t565 60.3943
R4594 GND.n1379 GND.t626 60.3943
R4595 GND.n1363 GND.t210 60.3943
R4596 GND.n1363 GND.t542 60.3943
R4597 GND.n1358 GND.t523 60.3943
R4598 GND.n1358 GND.t356 60.3943
R4599 GND.n1393 GND.t155 60.3943
R4600 GND.n1481 GND.t357 60.3943
R4601 GND.n1481 GND.t543 60.3943
R4602 GND.n1434 GND.t181 60.3943
R4603 GND.n1434 GND.t618 60.3943
R4604 GND.n1499 GND.t89 60.3943
R4605 GND.n1506 GND.t673 60.3943
R4606 GND.n1506 GND.t527 60.3943
R4607 GND.n1513 GND.t537 60.3943
R4608 GND.n1513 GND.t672 60.3943
R4609 GND.n1405 GND.t312 60.3943
R4610 GND.n1044 GND.t548 60.3943
R4611 GND.n1056 GND.t242 60.3943
R4612 GND.n1030 GND.t541 60.3943
R4613 GND.n1020 GND.t355 60.3943
R4614 GND.n1069 GND.t74 60.3943
R4615 GND.n1955 GND.t621 60.3943
R4616 GND.n1955 GND.t538 60.3943
R4617 GND.n1908 GND.t272 60.3943
R4618 GND.n1908 GND.t42 60.3943
R4619 GND.n1973 GND.t143 60.3943
R4620 GND.n1980 GND.t637 60.3943
R4621 GND.n1980 GND.t525 60.3943
R4622 GND.n1987 GND.t560 60.3943
R4623 GND.n1987 GND.t241 60.3943
R4624 GND.n1879 GND.t580 60.3943
R4625 GND.n1689 GND.t714 60.3943
R4626 GND.n1689 GND.t535 60.3943
R4627 GND.n1659 GND.t31 60.3943
R4628 GND.n1659 GND.t223 60.3943
R4629 GND.n1727 GND.t141 60.3943
R4630 GND.n1711 GND.t232 60.3943
R4631 GND.n1711 GND.t520 60.3943
R4632 GND.n1706 GND.t557 60.3943
R4633 GND.n1706 GND.t703 60.3943
R4634 GND.n1741 GND.t593 60.3943
R4635 GND.n2431 GND.t114 60.3943
R4636 GND.n2431 GND.t530 60.3943
R4637 GND.n2401 GND.t571 60.3943
R4638 GND.n2401 GND.t676 60.3943
R4639 GND.n2469 GND.t82 60.3943
R4640 GND.n2453 GND.t575 60.3943
R4641 GND.n2453 GND.t588 60.3943
R4642 GND.n2448 GND.t555 60.3943
R4643 GND.n2448 GND.t211 60.3943
R4644 GND.n2483 GND.t323 60.3943
R4645 GND.n2701 GND.t706 60.3943
R4646 GND.n2701 GND.t526 60.3943
R4647 GND.n2654 GND.t154 60.3943
R4648 GND.n2654 GND.t192 60.3943
R4649 GND.n2719 GND.t93 60.3943
R4650 GND.n2726 GND.t661 60.3943
R4651 GND.n2726 GND.t586 60.3943
R4652 GND.n2733 GND.t553 60.3943
R4653 GND.n2733 GND.t567 60.3943
R4654 GND.n2625 GND.t224 60.3943
R4655 GND.n2985 GND.t704 60.3943
R4656 GND.n2985 GND.t521 60.3943
R4657 GND.n2955 GND.t133 60.3943
R4658 GND.n2955 GND.t57 60.3943
R4659 GND.n3023 GND.t585 60.3943
R4660 GND.n3007 GND.t632 60.3943
R4661 GND.n3007 GND.t562 60.3943
R4662 GND.n3002 GND.t589 60.3943
R4663 GND.n3002 GND.t638 60.3943
R4664 GND.n3037 GND.t290 60.3943
R4665 GND.n3242 GND.t235 60.3943
R4666 GND.n3242 GND.t544 60.3943
R4667 GND.n3212 GND.t629 60.3943
R4668 GND.n3212 GND.t29 60.3943
R4669 GND.n3280 GND.t79 60.3943
R4670 GND.n3264 GND.t208 60.3943
R4671 GND.n3264 GND.t531 60.3943
R4672 GND.n3259 GND.t540 60.3943
R4673 GND.n3259 GND.t574 60.3943
R4674 GND.n3294 GND.t646 60.3943
R4675 GND.n4165 GND.t713 60.3943
R4676 GND.n4165 GND.t550 60.3943
R4677 GND.n4135 GND.t96 60.3943
R4678 GND.n4135 GND.t106 60.3943
R4679 GND.n4203 GND.t630 60.3943
R4680 GND.n4187 GND.t266 60.3943
R4681 GND.n4187 GND.t545 60.3943
R4682 GND.n4182 GND.t556 60.3943
R4683 GND.n4182 GND.t663 60.3943
R4684 GND.n4217 GND.t269 60.3943
R4685 GND.t640 GND.n681 60.2637
R4686 GND.n4370 GND 59.8971
R4687 GND.n289 GND 59.4951
R4688 GND.t296 GND.t297 58.6379
R4689 GND.t296 GND.t134 58.6379
R4690 GND.t682 GND.t684 58.6379
R4691 GND.t127 GND.t682 58.6379
R4692 GND.t184 GND.t182 58.6379
R4693 GND.t508 GND.t184 58.6379
R4694 GND.t168 GND.t169 58.6379
R4695 GND.t201 GND.t168 58.6379
R4696 GND.t613 GND.t610 58.6379
R4697 GND.t65 GND.t613 58.6379
R4698 GND.t650 GND.t651 58.6379
R4699 GND.t316 GND.t650 58.6379
R4700 GND.t245 GND.t246 58.6379
R4701 GND.t674 GND.t245 58.6379
R4702 GND.t86 GND.t238 58.6379
R4703 GND.t238 GND.t721 58.6379
R4704 GND.n4077 GND.n76 57.536
R4705 GND.n4056 GND.n76 57.536
R4706 GND.n4061 GND.n4051 57.536
R4707 GND.n4051 GND.n4048 57.536
R4708 GND.n4034 GND.n4033 57.536
R4709 GND.n4033 GND.n4031 57.536
R4710 GND.n3321 GND.n371 57.536
R4711 GND.n3322 GND.n3321 57.536
R4712 GND.n3327 GND.n366 57.536
R4713 GND.n3312 GND.n366 57.536
R4714 GND.n444 GND.n390 57.536
R4715 GND.n444 GND.n431 57.536
R4716 GND.n3155 GND.n3061 57.536
R4717 GND.n3134 GND.n3061 57.536
R4718 GND.n3139 GND.n3129 57.536
R4719 GND.n3129 GND.n3126 57.536
R4720 GND.n3112 GND.n3111 57.536
R4721 GND.n3111 GND.n3109 57.536
R4722 GND.n2602 GND.n2507 57.536
R4723 GND.n2581 GND.n2507 57.536
R4724 GND.n2586 GND.n2576 57.536
R4725 GND.n2576 GND.n2573 57.536
R4726 GND.n2559 GND.n2558 57.536
R4727 GND.n2558 GND.n2556 57.536
R4728 GND.n1857 GND.n1764 57.536
R4729 GND.n1836 GND.n1764 57.536
R4730 GND.n1841 GND.n1831 57.536
R4731 GND.n1831 GND.n1828 57.536
R4732 GND.n1814 GND.n1813 57.536
R4733 GND.n1813 GND.n1811 57.536
R4734 GND.n1600 GND.n912 57.536
R4735 GND.n1579 GND.n912 57.536
R4736 GND.n1584 GND.n1574 57.536
R4737 GND.n1574 GND.n1571 57.536
R4738 GND.n1557 GND.n1556 57.536
R4739 GND.n1556 GND.n1554 57.536
R4740 GND.n1252 GND.n955 57.536
R4741 GND.n1231 GND.n955 57.536
R4742 GND.n1236 GND.n1226 57.536
R4743 GND.n1226 GND.n1223 57.536
R4744 GND.n1209 GND.n1208 57.536
R4745 GND.n1208 GND.n1206 57.536
R4746 GND.n1382 GND.n1287 57.536
R4747 GND.n1361 GND.n1287 57.536
R4748 GND.n1366 GND.n1356 57.536
R4749 GND.n1356 GND.n1353 57.536
R4750 GND.n1339 GND.n1338 57.536
R4751 GND.n1338 GND.n1336 57.536
R4752 GND.n1503 GND.n1502 57.536
R4753 GND.n1504 GND.n1503 57.536
R4754 GND.n1510 GND.n1509 57.536
R4755 GND.n1511 GND.n1510 57.536
R4756 GND.n1479 GND.n1478 57.536
R4757 GND.n1478 GND.n1476 57.536
R4758 GND.n1977 GND.n1976 57.536
R4759 GND.n1978 GND.n1977 57.536
R4760 GND.n1984 GND.n1983 57.536
R4761 GND.n1985 GND.n1984 57.536
R4762 GND.n1953 GND.n1952 57.536
R4763 GND.n1952 GND.n1950 57.536
R4764 GND.n1730 GND.n1636 57.536
R4765 GND.n1709 GND.n1636 57.536
R4766 GND.n1714 GND.n1704 57.536
R4767 GND.n1704 GND.n1701 57.536
R4768 GND.n1687 GND.n1686 57.536
R4769 GND.n1686 GND.n1684 57.536
R4770 GND.n2472 GND.n583 57.536
R4771 GND.n2451 GND.n583 57.536
R4772 GND.n2456 GND.n2446 57.536
R4773 GND.n2446 GND.n2443 57.536
R4774 GND.n2429 GND.n2428 57.536
R4775 GND.n2428 GND.n2426 57.536
R4776 GND.n2723 GND.n2722 57.536
R4777 GND.n2724 GND.n2723 57.536
R4778 GND.n2730 GND.n2729 57.536
R4779 GND.n2731 GND.n2730 57.536
R4780 GND.n2699 GND.n2698 57.536
R4781 GND.n2698 GND.n2696 57.536
R4782 GND.n3026 GND.n470 57.536
R4783 GND.n3005 GND.n470 57.536
R4784 GND.n3010 GND.n3000 57.536
R4785 GND.n3000 GND.n2997 57.536
R4786 GND.n2983 GND.n2982 57.536
R4787 GND.n2982 GND.n2980 57.536
R4788 GND.n3283 GND.n3190 57.536
R4789 GND.n3262 GND.n3190 57.536
R4790 GND.n3267 GND.n3257 57.536
R4791 GND.n3257 GND.n3254 57.536
R4792 GND.n3240 GND.n3239 57.536
R4793 GND.n3239 GND.n3237 57.536
R4794 GND.n4206 GND.n4112 57.536
R4795 GND.n4185 GND.n4112 57.536
R4796 GND.n4190 GND.n4180 57.536
R4797 GND.n4180 GND.n4177 57.536
R4798 GND.n4163 GND.n4162 57.536
R4799 GND.n4162 GND.n4160 57.536
R4800 GND.n275 GND 56.8872
R4801 GND.n1114 GND.n981 53.4324
R4802 GND.n4260 GND.n4259 52.5417
R4803 GND.n4266 GND.n4259 52.5417
R4804 GND.n1054 GND.n1053 52.5417
R4805 GND.n1053 GND.n1051 52.5417
R4806 GND.n4337 GND.n17 52.5417
R4807 GND.n4351 GND.n17 52.5417
R4808 GND.n41 GND.n35 52.5417
R4809 GND.n4312 GND.n35 52.5417
R4810 GND.n119 GND.n118 52.5417
R4811 GND.n3980 GND.n118 52.5417
R4812 GND.n2921 GND.n2920 52.5417
R4813 GND.n2931 GND.n2920 52.5417
R4814 GND.n546 GND.n539 52.5417
R4815 GND.n2807 GND.n539 52.5417
R4816 GND.n2376 GND.n2352 52.5417
R4817 GND.n2371 GND.n2352 52.5417
R4818 GND.n2278 GND.n2277 52.5417
R4819 GND.n2277 GND.n2276 52.5417
R4820 GND.n874 GND.n829 52.5417
R4821 GND.n2004 GND.n829 52.5417
R4822 GND.n844 GND.n831 52.5417
R4823 GND.n859 GND.n831 52.5417
R4824 GND.n1155 GND.n1154 52.5417
R4825 GND.n1154 GND.n1153 52.5417
R4826 GND.n176 GND.n37 52.5417
R4827 GND.n4303 GND.n37 52.5417
R4828 GND.n156 GND.n143 52.5417
R4829 GND.n171 GND.n143 52.5417
R4830 GND.n3988 GND.n3987 52.5417
R4831 GND.n3987 GND.n105 52.5417
R4832 GND.n3355 GND.n342 52.5417
R4833 GND.n3368 GND.n342 52.5417
R4834 GND.n2939 GND.n2938 52.5417
R4835 GND.n2938 GND.n2906 52.5417
R4836 GND.n2762 GND.n2748 52.5417
R4837 GND.n2777 GND.n2748 52.5417
R4838 GND.n531 GND.n530 52.5417
R4839 GND.n532 GND.n531 52.5417
R4840 GND.n2308 GND.n605 52.5417
R4841 GND.n2323 GND.n605 52.5417
R4842 GND.n613 GND.n612 52.5417
R4843 GND.n612 GND.n611 52.5417
R4844 GND.n821 GND.n820 52.5417
R4845 GND.n822 GND.n821 52.5417
R4846 GND.n793 GND.n786 52.5417
R4847 GND.n2045 GND.n786 52.5417
R4848 GND.n778 GND.n777 52.5417
R4849 GND.n779 GND.n778 52.5417
R4850 GND.n1077 GND.n986 52.5417
R4851 GND.n1106 GND.n986 52.5417
R4852 GND.n995 GND.n994 52.5417
R4853 GND.n994 GND.n993 52.5417
R4854 GND.n2243 GND.n2188 52.5417
R4855 GND.n2240 GND.n2188 52.5417
R4856 GND.n2840 GND.n512 52.5417
R4857 GND.n2850 GND.n512 52.5417
R4858 GND.n2885 GND.n312 52.5417
R4859 GND.n3467 GND.n312 52.5417
R4860 GND.n3423 GND.n3387 52.5417
R4861 GND.n3420 GND.n3387 52.5417
R4862 GND.n3943 GND.n3899 52.5417
R4863 GND.n3940 GND.n3899 52.5417
R4864 GND.n755 GND.n733 52.5417
R4865 GND.n752 GND.n733 52.5417
R4866 GND.n2139 GND.n662 52.5417
R4867 GND.n2149 GND.n662 52.5417
R4868 GND.n2091 GND.n2090 52.5417
R4869 GND.n2090 GND.n692 52.5417
R4870 GND.n3626 GND.n243 50.4812
R4871 GND.n283 GND 47.3872
R4872 GND.n297 GND 46.2777
R4873 GND.t324 GND.n616 45.5839
R4874 GND.n615 GND.t362 45.5839
R4875 GND.n2318 GND.t176 45.5839
R4876 GND.n782 GND.t100 45.5839
R4877 GND.n783 GND.t257 45.5839
R4878 GND.n2049 GND.t669 45.5839
R4879 GND.t147 GND.n990 45.5839
R4880 GND.n1102 GND.t318 45.5839
R4881 GND.t601 GND.n1101 45.5839
R4882 GND.n825 GND.t19 45.5839
R4883 GND.n826 GND.t1 45.5839
R4884 GND.n2008 GND.t119 45.5839
R4885 GND.n535 GND.t225 45.5839
R4886 GND.n536 GND.t215 45.5839
R4887 GND.n2811 GND.t609 45.5839
R4888 GND.n2936 GND.t26 45.5839
R4889 GND.n2935 GND.t51 45.5839
R4890 GND.t348 GND.n2913 45.5839
R4891 GND.n3985 GND.t678 45.5839
R4892 GND.n3984 GND.t97 45.5839
R4893 GND.n126 GND.t517 45.5839
R4894 GND.n4299 GND.t270 45.5839
R4895 GND.n4298 GND.t129 45.5839
R4896 GND.t203 GND.n31 45.5839
R4897 GND.n937 GND 44.6732
R4898 GND.n3999 GND.n3998 44.1913
R4899 GND.n3998 GND.n63 44.1913
R4900 GND.n3077 GND.n357 44.1913
R4901 GND.n3048 GND.n357 44.1913
R4902 GND.n2524 GND.n2523 44.1913
R4903 GND.n2523 GND.n2494 44.1913
R4904 GND.n2296 GND.n622 44.1913
R4905 GND.n2296 GND.n623 44.1913
R4906 GND.n1522 GND.n1521 44.1913
R4907 GND.n1521 GND.n899 44.1913
R4908 GND.n1174 GND.n1173 44.1913
R4909 GND.n1173 GND.n942 44.1913
R4910 GND.n1304 GND.n1303 44.1913
R4911 GND.n1303 GND.n1274 44.1913
R4912 GND.n1519 GND.n928 44.1913
R4913 GND.n1519 GND.n1518 44.1913
R4914 GND.n1994 GND.n885 44.1913
R4915 GND.n1994 GND.n1992 44.1913
R4916 GND.n1652 GND.n599 44.1913
R4917 GND.n1623 GND.n599 44.1913
R4918 GND.n2394 GND.n2393 44.1913
R4919 GND.n2393 GND.n570 44.1913
R4920 GND.n2798 GND.n556 44.1913
R4921 GND.n2798 GND.n2738 44.1913
R4922 GND.n2948 GND.n2947 44.1913
R4923 GND.n2947 GND.n457 44.1913
R4924 GND.n3996 GND.n92 44.1913
R4925 GND.n3996 GND.n93 44.1913
R4926 GND.n4128 GND.n49 44.1913
R4927 GND.n4099 GND.n49 44.1913
R4928 GND.n1000 GND 43.1031
R4929 GND.n291 GND 42.6372
R4930 GND.n1269 GND 41.8814
R4931 GND.n1268 GND 40.5651
R4932 GND.n1399 GND 39.0896
R4933 GND.t693 GND.n250 38.8621
R4934 GND.n1398 GND 38.0271
R4935 GND.n2100 GND.n681 36.5118
R4936 GND.n894 GND 36.2978
R4937 GND.n1400 GND 35.4891
R4938 GND.n4014 GND.n4001 34.4123
R4939 GND.n4001 GND.n3999 34.4123
R4940 GND.n4002 GND.n4000 34.4123
R4941 GND.n4000 GND.n82 34.4123
R4942 GND.n4009 GND.n4008 34.4123
R4943 GND.n4008 GND.n69 34.4123
R4944 GND.n4013 GND.n4012 34.4123
R4945 GND.n4012 GND.n63 34.4123
R4946 GND.n3092 GND.n3079 34.4123
R4947 GND.n3079 GND.n3077 34.4123
R4948 GND.n3080 GND.n3078 34.4123
R4949 GND.n3078 GND.n3067 34.4123
R4950 GND.n3087 GND.n3086 34.4123
R4951 GND.n3086 GND.n3054 34.4123
R4952 GND.n3091 GND.n3090 34.4123
R4953 GND.n3090 GND.n3048 34.4123
R4954 GND.n2539 GND.n2526 34.4123
R4955 GND.n2526 GND.n2524 34.4123
R4956 GND.n2527 GND.n2525 34.4123
R4957 GND.n2525 GND.n2513 34.4123
R4958 GND.n2534 GND.n2533 34.4123
R4959 GND.n2533 GND.n2500 34.4123
R4960 GND.n2538 GND.n2537 34.4123
R4961 GND.n2537 GND.n2494 34.4123
R4962 GND.n1794 GND.n1781 34.4123
R4963 GND.n1781 GND.n622 34.4123
R4964 GND.n1782 GND.n1780 34.4123
R4965 GND.n1780 GND.n1770 34.4123
R4966 GND.n1789 GND.n1788 34.4123
R4967 GND.n1788 GND.n1757 34.4123
R4968 GND.n1793 GND.n1792 34.4123
R4969 GND.n1792 GND.n623 34.4123
R4970 GND.n1537 GND.n1524 34.4123
R4971 GND.n1524 GND.n1522 34.4123
R4972 GND.n1525 GND.n1523 34.4123
R4973 GND.n1523 GND.n918 34.4123
R4974 GND.n1532 GND.n1531 34.4123
R4975 GND.n1531 GND.n905 34.4123
R4976 GND.n1536 GND.n1535 34.4123
R4977 GND.n1535 GND.n899 34.4123
R4978 GND.n1189 GND.n1176 34.4123
R4979 GND.n1176 GND.n1174 34.4123
R4980 GND.n1177 GND.n1175 34.4123
R4981 GND.n1175 GND.n961 34.4123
R4982 GND.n1184 GND.n1183 34.4123
R4983 GND.n1183 GND.n948 34.4123
R4984 GND.n1188 GND.n1187 34.4123
R4985 GND.n1187 GND.n942 34.4123
R4986 GND.n1319 GND.n1306 34.4123
R4987 GND.n1306 GND.n1304 34.4123
R4988 GND.n1307 GND.n1305 34.4123
R4989 GND.n1305 GND.n1293 34.4123
R4990 GND.n1314 GND.n1313 34.4123
R4991 GND.n1313 GND.n1280 34.4123
R4992 GND.n1318 GND.n1317 34.4123
R4993 GND.n1317 GND.n1274 34.4123
R4994 GND.n1451 GND.n1429 34.4123
R4995 GND.n1429 GND.n928 34.4123
R4996 GND.n1430 GND.n1428 34.4123
R4997 GND.n1428 GND.n1418 34.4123
R4998 GND.n1457 GND.n1456 34.4123
R4999 GND.n1466 GND.n1457 34.4123
R5000 GND.n1450 GND.n930 34.4123
R5001 GND.n1518 GND.n930 34.4123
R5002 GND.n168 GND.n143 34.4123
R5003 GND.n168 GND.n138 34.4123
R5004 GND.n145 GND.n144 34.4123
R5005 GND.n145 GND.n138 34.4123
R5006 GND.n342 GND.n340 34.4123
R5007 GND.n3359 GND.n340 34.4123
R5008 GND.n341 GND.n339 34.4123
R5009 GND.n3359 GND.n339 34.4123
R5010 GND.n2774 GND.n2748 34.4123
R5011 GND.n2774 GND.n2743 34.4123
R5012 GND.n2750 GND.n2749 34.4123
R5013 GND.n2750 GND.n2743 34.4123
R5014 GND.n608 GND.n605 34.4123
R5015 GND.n615 GND.n608 34.4123
R5016 GND.n607 GND.n606 34.4123
R5017 GND.n615 GND.n607 34.4123
R5018 GND.n612 GND.n609 34.4123
R5019 GND.n616 GND.n609 34.4123
R5020 GND.n2315 GND.n610 34.4123
R5021 GND.n616 GND.n610 34.4123
R5022 GND.n786 GND.n784 34.4123
R5023 GND.n784 GND.n783 34.4123
R5024 GND.n785 GND.n781 34.4123
R5025 GND.n783 GND.n781 34.4123
R5026 GND.n778 GND.n775 34.4123
R5027 GND.n782 GND.n775 34.4123
R5028 GND.n2052 GND.n776 34.4123
R5029 GND.n782 GND.n776 34.4123
R5030 GND.n1103 GND.n986 34.4123
R5031 GND.n1103 GND.n1102 34.4123
R5032 GND.n988 GND.n987 34.4123
R5033 GND.n1102 GND.n988 34.4123
R5034 GND.n994 GND.n991 34.4123
R5035 GND.n991 GND.n990 34.4123
R5036 GND.n1098 GND.n992 34.4123
R5037 GND.n992 GND.n990 34.4123
R5038 GND.n2188 GND.n2186 34.4123
R5039 GND.n2192 GND.n2186 34.4123
R5040 GND.n2187 GND.n2185 34.4123
R5041 GND.n2192 GND.n2185 34.4123
R5042 GND.n515 GND.n512 34.4123
R5043 GND.n2844 GND.n515 34.4123
R5044 GND.n514 GND.n513 34.4123
R5045 GND.n2844 GND.n514 34.4123
R5046 GND.n312 GND.n310 34.4123
R5047 GND.n2884 GND.n310 34.4123
R5048 GND.n311 GND.n309 34.4123
R5049 GND.n2884 GND.n309 34.4123
R5050 GND.n733 GND.n731 34.4123
R5051 GND.n737 GND.n731 34.4123
R5052 GND.n732 GND.n730 34.4123
R5053 GND.n737 GND.n730 34.4123
R5054 GND.n665 GND.n662 34.4123
R5055 GND.n2143 GND.n665 34.4123
R5056 GND.n664 GND.n663 34.4123
R5057 GND.n2143 GND.n664 34.4123
R5058 GND.n17 GND.n15 34.4123
R5059 GND.n4341 GND.n15 34.4123
R5060 GND.n16 GND.n14 34.4123
R5061 GND.n4341 GND.n14 34.4123
R5062 GND.n3387 GND.n3385 34.4123
R5063 GND.n3389 GND.n3385 34.4123
R5064 GND.n3386 GND.n3384 34.4123
R5065 GND.n3389 GND.n3384 34.4123
R5066 GND.n3899 GND.n3897 34.4123
R5067 GND.n3903 GND.n3897 34.4123
R5068 GND.n3898 GND.n3896 34.4123
R5069 GND.n3903 GND.n3896 34.4123
R5070 GND.n2090 GND.n2089 34.4123
R5071 GND.n2089 GND.n2088 34.4123
R5072 GND.n2087 GND.n2086 34.4123
R5073 GND.n2088 GND.n2087 34.4123
R5074 GND.n1049 GND.n1048 34.4123
R5075 GND.n1048 GND.n981 34.4123
R5076 GND.n1053 GND.n1052 34.4123
R5077 GND.n1052 GND.n983 34.4123
R5078 GND.n1154 GND.n1130 34.4123
R5079 GND.n1139 GND.n1130 34.4123
R5080 GND.n1131 GND.n1129 34.4123
R5081 GND.n1139 GND.n1129 34.4123
R5082 GND.n856 GND.n831 34.4123
R5083 GND.n856 GND.n808 34.4123
R5084 GND.n833 GND.n832 34.4123
R5085 GND.n833 GND.n808 34.4123
R5086 GND.n2011 GND.n819 34.4123
R5087 GND.n825 GND.n819 34.4123
R5088 GND.n821 GND.n818 34.4123
R5089 GND.n825 GND.n818 34.4123
R5090 GND.n829 GND.n827 34.4123
R5091 GND.n827 GND.n826 34.4123
R5092 GND.n828 GND.n824 34.4123
R5093 GND.n826 GND.n824 34.4123
R5094 GND.n1925 GND.n1903 34.4123
R5095 GND.n1903 GND.n885 34.4123
R5096 GND.n1904 GND.n1902 34.4123
R5097 GND.n1902 GND.n1892 34.4123
R5098 GND.n1931 GND.n1930 34.4123
R5099 GND.n1940 GND.n1931 34.4123
R5100 GND.n1924 GND.n887 34.4123
R5101 GND.n1992 GND.n887 34.4123
R5102 GND.n2277 GND.n638 34.4123
R5103 GND.n2262 GND.n638 34.4123
R5104 GND.n639 GND.n637 34.4123
R5105 GND.n2262 GND.n637 34.4123
R5106 GND.n1667 GND.n1654 34.4123
R5107 GND.n1654 GND.n1652 34.4123
R5108 GND.n1655 GND.n1653 34.4123
R5109 GND.n1653 GND.n1642 34.4123
R5110 GND.n1662 GND.n1661 34.4123
R5111 GND.n1661 GND.n1629 34.4123
R5112 GND.n1666 GND.n1665 34.4123
R5113 GND.n1665 GND.n1623 34.4123
R5114 GND.n2409 GND.n2396 34.4123
R5115 GND.n2396 GND.n2394 34.4123
R5116 GND.n2397 GND.n2395 34.4123
R5117 GND.n2395 GND.n589 34.4123
R5118 GND.n2404 GND.n2403 34.4123
R5119 GND.n2403 GND.n576 34.4123
R5120 GND.n2408 GND.n2407 34.4123
R5121 GND.n2407 GND.n570 34.4123
R5122 GND.n2352 GND.n2350 34.4123
R5123 GND.n2353 GND.n2350 34.4123
R5124 GND.n2351 GND.n2349 34.4123
R5125 GND.n2353 GND.n2349 34.4123
R5126 GND.n2814 GND.n529 34.4123
R5127 GND.n535 GND.n529 34.4123
R5128 GND.n531 GND.n528 34.4123
R5129 GND.n535 GND.n528 34.4123
R5130 GND.n539 GND.n537 34.4123
R5131 GND.n537 GND.n536 34.4123
R5132 GND.n538 GND.n534 34.4123
R5133 GND.n536 GND.n534 34.4123
R5134 GND.n2671 GND.n2649 34.4123
R5135 GND.n2649 GND.n556 34.4123
R5136 GND.n2650 GND.n2648 34.4123
R5137 GND.n2648 GND.n2638 34.4123
R5138 GND.n2677 GND.n2676 34.4123
R5139 GND.n2686 GND.n2677 34.4123
R5140 GND.n2670 GND.n558 34.4123
R5141 GND.n2738 GND.n558 34.4123
R5142 GND.n2963 GND.n2950 34.4123
R5143 GND.n2950 GND.n2948 34.4123
R5144 GND.n2951 GND.n2949 34.4123
R5145 GND.n2949 GND.n476 34.4123
R5146 GND.n2958 GND.n2957 34.4123
R5147 GND.n2957 GND.n463 34.4123
R5148 GND.n2962 GND.n2961 34.4123
R5149 GND.n2961 GND.n457 34.4123
R5150 GND.n2911 GND.n2910 34.4123
R5151 GND.n2936 GND.n2911 34.4123
R5152 GND.n2938 GND.n2937 34.4123
R5153 GND.n2937 GND.n2936 34.4123
R5154 GND.n2920 GND.n2912 34.4123
R5155 GND.n2935 GND.n2912 34.4123
R5156 GND.n2934 GND.n2933 34.4123
R5157 GND.n2935 GND.n2934 34.4123
R5158 GND.n420 GND.n419 34.4123
R5159 GND.n420 GND.n385 34.4123
R5160 GND.n407 GND.n359 34.4123
R5161 GND.n3332 GND.n359 34.4123
R5162 GND.n413 GND.n411 34.4123
R5163 GND.n413 GND.n94 34.4123
R5164 GND.n409 GND.n387 34.4123
R5165 GND.n3319 GND.n387 34.4123
R5166 GND.n3220 GND.n3207 34.4123
R5167 GND.n3207 GND.n92 34.4123
R5168 GND.n3208 GND.n3206 34.4123
R5169 GND.n3206 GND.n3196 34.4123
R5170 GND.n3215 GND.n3214 34.4123
R5171 GND.n3214 GND.n3183 34.4123
R5172 GND.n3219 GND.n3218 34.4123
R5173 GND.n3218 GND.n93 34.4123
R5174 GND.n110 GND.n109 34.4123
R5175 GND.n3985 GND.n110 34.4123
R5176 GND.n3987 GND.n3986 34.4123
R5177 GND.n3986 GND.n3985 34.4123
R5178 GND.n118 GND.n111 34.4123
R5179 GND.n3984 GND.n111 34.4123
R5180 GND.n3983 GND.n3982 34.4123
R5181 GND.n3984 GND.n3983 34.4123
R5182 GND.n4143 GND.n4130 34.4123
R5183 GND.n4130 GND.n4128 34.4123
R5184 GND.n4131 GND.n4129 34.4123
R5185 GND.n4129 GND.n4118 34.4123
R5186 GND.n4138 GND.n4137 34.4123
R5187 GND.n4137 GND.n4105 34.4123
R5188 GND.n4142 GND.n4141 34.4123
R5189 GND.n4141 GND.n4099 34.4123
R5190 GND.n4300 GND.n38 34.4123
R5191 GND.n4300 GND.n4299 34.4123
R5192 GND.n39 GND.n37 34.4123
R5193 GND.n4299 GND.n39 34.4123
R5194 GND.n35 GND.n33 34.4123
R5195 GND.n4298 GND.n33 34.4123
R5196 GND.n34 GND.n32 34.4123
R5197 GND.n4298 GND.n32 34.4123
R5198 GND.n4259 GND.n4238 34.4123
R5199 GND.n4275 GND.n4238 34.4123
R5200 GND.n4263 GND.n51 34.4123
R5201 GND.n4287 GND.n51 34.4123
R5202 GND.n720 GND.t3 34.3246
R5203 GND.n3628 GND 33.6971
R5204 GND.n1617 GND 33.506
R5205 GND.n299 GND 33.1372
R5206 GND.n305 GND 33.0603
R5207 GND.n1616 GND 32.9511
R5208 GND.n3787 GND 31.7921
R5209 GND.n4362 GND.n4361 31.1892
R5210 GND.n1873 GND 30.7142
R5211 GND.n1874 GND 30.4131
R5212 GND.n3792 GND 29.887
R5213 GND.n4015 GND.n4013 29.7417
R5214 GND.n4013 GND.n4004 29.7417
R5215 GND.n4015 GND.n4014 29.7417
R5216 GND.n4014 GND.n4004 29.7417
R5217 GND.n418 GND.n409 29.7417
R5218 GND.n409 GND.n405 29.7417
R5219 GND.n419 GND.n418 29.7417
R5220 GND.n419 GND.n405 29.7417
R5221 GND.n3093 GND.n3091 29.7417
R5222 GND.n3091 GND.n3082 29.7417
R5223 GND.n3093 GND.n3092 29.7417
R5224 GND.n3092 GND.n3082 29.7417
R5225 GND.n2540 GND.n2538 29.7417
R5226 GND.n2538 GND.n2529 29.7417
R5227 GND.n2540 GND.n2539 29.7417
R5228 GND.n2539 GND.n2529 29.7417
R5229 GND.n1795 GND.n1793 29.7417
R5230 GND.n1793 GND.n1784 29.7417
R5231 GND.n1795 GND.n1794 29.7417
R5232 GND.n1794 GND.n1784 29.7417
R5233 GND.n1538 GND.n1536 29.7417
R5234 GND.n1536 GND.n1527 29.7417
R5235 GND.n1538 GND.n1537 29.7417
R5236 GND.n1537 GND.n1527 29.7417
R5237 GND.n1190 GND.n1188 29.7417
R5238 GND.n1188 GND.n1179 29.7417
R5239 GND.n1190 GND.n1189 29.7417
R5240 GND.n1189 GND.n1179 29.7417
R5241 GND.n1320 GND.n1318 29.7417
R5242 GND.n1318 GND.n1309 29.7417
R5243 GND.n1320 GND.n1319 29.7417
R5244 GND.n1319 GND.n1309 29.7417
R5245 GND.n1452 GND.n1450 29.7417
R5246 GND.n1450 GND.n1432 29.7417
R5247 GND.n1452 GND.n1451 29.7417
R5248 GND.n1451 GND.n1432 29.7417
R5249 GND.n1926 GND.n1924 29.7417
R5250 GND.n1924 GND.n1906 29.7417
R5251 GND.n1926 GND.n1925 29.7417
R5252 GND.n1925 GND.n1906 29.7417
R5253 GND.n1668 GND.n1666 29.7417
R5254 GND.n1666 GND.n1657 29.7417
R5255 GND.n1668 GND.n1667 29.7417
R5256 GND.n1667 GND.n1657 29.7417
R5257 GND.n2410 GND.n2408 29.7417
R5258 GND.n2408 GND.n2399 29.7417
R5259 GND.n2410 GND.n2409 29.7417
R5260 GND.n2409 GND.n2399 29.7417
R5261 GND.n2672 GND.n2670 29.7417
R5262 GND.n2670 GND.n2652 29.7417
R5263 GND.n2672 GND.n2671 29.7417
R5264 GND.n2671 GND.n2652 29.7417
R5265 GND.n2964 GND.n2962 29.7417
R5266 GND.n2962 GND.n2953 29.7417
R5267 GND.n2964 GND.n2963 29.7417
R5268 GND.n2963 GND.n2953 29.7417
R5269 GND.n3221 GND.n3219 29.7417
R5270 GND.n3219 GND.n3210 29.7417
R5271 GND.n3221 GND.n3220 29.7417
R5272 GND.n3220 GND.n3210 29.7417
R5273 GND.n4144 GND.n4142 29.7417
R5274 GND.n4142 GND.n4133 29.7417
R5275 GND.n4144 GND.n4143 29.7417
R5276 GND.n4143 GND.n4133 29.7417
R5277 GND.n2101 GND.t297 29.3192
R5278 GND.t134 GND.n3612 29.3192
R5279 GND.n3610 GND.t684 29.3192
R5280 GND.n3593 GND.t127 29.3192
R5281 GND.n3591 GND.t182 29.3192
R5282 GND.n3573 GND.t508 29.3192
R5283 GND.n3571 GND.t169 29.3192
R5284 GND.n3554 GND.t201 29.3192
R5285 GND.n3552 GND.t610 29.3192
R5286 GND.n3532 GND.t65 29.3192
R5287 GND.n3530 GND.t651 29.3192
R5288 GND.n3510 GND.t316 29.3192
R5289 GND.n3508 GND.t246 29.3192
R5290 GND.n3491 GND.t674 29.3192
R5291 GND.n3489 GND.t86 29.3192
R5292 GND.n3881 GND.t721 29.3192
R5293 GND.n3797 GND 27.9819
R5294 GND.t273 GND.n1114 27.9484
R5295 GND.n1746 GND 27.9224
R5296 GND.n1747 GND 27.8751
R5297 GND.n3472 GND 26.4516
R5298 GND.n3802 GND 26.0769
R5299 GND.n1618 GND 25.3371
R5300 GND.n565 GND 25.1306
R5301 GND.n3807 GND 24.1718
R5302 GND.n2488 GND 22.7991
R5303 GND.n4033 GND.n4032 22.5005
R5304 GND.n4032 GND.n3999 22.5005
R5305 GND.n4027 GND.n4026 22.5005
R5306 GND.n4026 GND.n82 22.5005
R5307 GND.n4023 GND.n4022 22.5005
R5308 GND.n4022 GND.n69 22.5005
R5309 GND.n4033 GND.n4020 22.5005
R5310 GND.n4020 GND.n63 22.5005
R5311 GND.n91 GND.n76 22.5005
R5312 GND.n3999 GND.n91 22.5005
R5313 GND.n86 GND.n85 22.5005
R5314 GND.n86 GND.n82 22.5005
R5315 GND.n4080 GND.n73 22.5005
R5316 GND.n73 GND.n69 22.5005
R5317 GND.n76 GND.n72 22.5005
R5318 GND.n72 GND.n63 22.5005
R5319 GND.n4051 GND.n4046 22.5005
R5320 GND.n4046 GND.n3999 22.5005
R5321 GND.n4047 GND.n4045 22.5005
R5322 GND.n4045 GND.n82 22.5005
R5323 GND.n4065 GND.n4064 22.5005
R5324 GND.n4064 GND.n69 22.5005
R5325 GND.n4051 GND.n4050 22.5005
R5326 GND.n4050 GND.n63 22.5005
R5327 GND.n3111 GND.n3110 22.5005
R5328 GND.n3110 GND.n3077 22.5005
R5329 GND.n3105 GND.n3104 22.5005
R5330 GND.n3104 GND.n3067 22.5005
R5331 GND.n3101 GND.n3100 22.5005
R5332 GND.n3100 GND.n3054 22.5005
R5333 GND.n3111 GND.n3098 22.5005
R5334 GND.n3098 GND.n3048 22.5005
R5335 GND.n3076 GND.n3061 22.5005
R5336 GND.n3077 GND.n3076 22.5005
R5337 GND.n3071 GND.n3070 22.5005
R5338 GND.n3071 GND.n3067 22.5005
R5339 GND.n3158 GND.n3058 22.5005
R5340 GND.n3058 GND.n3054 22.5005
R5341 GND.n3061 GND.n3057 22.5005
R5342 GND.n3057 GND.n3048 22.5005
R5343 GND.n3129 GND.n3124 22.5005
R5344 GND.n3124 GND.n3077 22.5005
R5345 GND.n3125 GND.n3123 22.5005
R5346 GND.n3123 GND.n3067 22.5005
R5347 GND.n3143 GND.n3142 22.5005
R5348 GND.n3142 GND.n3054 22.5005
R5349 GND.n3129 GND.n3128 22.5005
R5350 GND.n3128 GND.n3048 22.5005
R5351 GND.n2558 GND.n2557 22.5005
R5352 GND.n2557 GND.n2524 22.5005
R5353 GND.n2552 GND.n2551 22.5005
R5354 GND.n2551 GND.n2513 22.5005
R5355 GND.n2548 GND.n2547 22.5005
R5356 GND.n2547 GND.n2500 22.5005
R5357 GND.n2558 GND.n2545 22.5005
R5358 GND.n2545 GND.n2494 22.5005
R5359 GND.n2522 GND.n2507 22.5005
R5360 GND.n2524 GND.n2522 22.5005
R5361 GND.n2517 GND.n2516 22.5005
R5362 GND.n2517 GND.n2513 22.5005
R5363 GND.n2605 GND.n2504 22.5005
R5364 GND.n2504 GND.n2500 22.5005
R5365 GND.n2507 GND.n2503 22.5005
R5366 GND.n2503 GND.n2494 22.5005
R5367 GND.n2576 GND.n2571 22.5005
R5368 GND.n2571 GND.n2524 22.5005
R5369 GND.n2572 GND.n2570 22.5005
R5370 GND.n2570 GND.n2513 22.5005
R5371 GND.n2590 GND.n2589 22.5005
R5372 GND.n2589 GND.n2500 22.5005
R5373 GND.n2576 GND.n2575 22.5005
R5374 GND.n2575 GND.n2494 22.5005
R5375 GND.n1813 GND.n1812 22.5005
R5376 GND.n1812 GND.n622 22.5005
R5377 GND.n1807 GND.n1806 22.5005
R5378 GND.n1806 GND.n1770 22.5005
R5379 GND.n1803 GND.n1802 22.5005
R5380 GND.n1802 GND.n1757 22.5005
R5381 GND.n1813 GND.n1800 22.5005
R5382 GND.n1800 GND.n623 22.5005
R5383 GND.n1775 GND.n1764 22.5005
R5384 GND.n1775 GND.n622 22.5005
R5385 GND.n1774 GND.n1773 22.5005
R5386 GND.n1774 GND.n1770 22.5005
R5387 GND.n1860 GND.n1761 22.5005
R5388 GND.n1761 GND.n1757 22.5005
R5389 GND.n1764 GND.n1760 22.5005
R5390 GND.n1760 GND.n623 22.5005
R5391 GND.n1831 GND.n1826 22.5005
R5392 GND.n1826 GND.n622 22.5005
R5393 GND.n1827 GND.n1825 22.5005
R5394 GND.n1825 GND.n1770 22.5005
R5395 GND.n1845 GND.n1844 22.5005
R5396 GND.n1844 GND.n1757 22.5005
R5397 GND.n1831 GND.n1830 22.5005
R5398 GND.n1830 GND.n623 22.5005
R5399 GND.n1556 GND.n1555 22.5005
R5400 GND.n1555 GND.n1522 22.5005
R5401 GND.n1550 GND.n1549 22.5005
R5402 GND.n1549 GND.n918 22.5005
R5403 GND.n1546 GND.n1545 22.5005
R5404 GND.n1545 GND.n905 22.5005
R5405 GND.n1556 GND.n1543 22.5005
R5406 GND.n1543 GND.n899 22.5005
R5407 GND.n927 GND.n912 22.5005
R5408 GND.n1522 GND.n927 22.5005
R5409 GND.n922 GND.n921 22.5005
R5410 GND.n922 GND.n918 22.5005
R5411 GND.n1603 GND.n909 22.5005
R5412 GND.n909 GND.n905 22.5005
R5413 GND.n912 GND.n908 22.5005
R5414 GND.n908 GND.n899 22.5005
R5415 GND.n1574 GND.n1569 22.5005
R5416 GND.n1569 GND.n1522 22.5005
R5417 GND.n1570 GND.n1568 22.5005
R5418 GND.n1568 GND.n918 22.5005
R5419 GND.n1588 GND.n1587 22.5005
R5420 GND.n1587 GND.n905 22.5005
R5421 GND.n1574 GND.n1573 22.5005
R5422 GND.n1573 GND.n899 22.5005
R5423 GND.n1208 GND.n1207 22.5005
R5424 GND.n1207 GND.n1174 22.5005
R5425 GND.n1202 GND.n1201 22.5005
R5426 GND.n1201 GND.n961 22.5005
R5427 GND.n1198 GND.n1197 22.5005
R5428 GND.n1197 GND.n948 22.5005
R5429 GND.n1208 GND.n1195 22.5005
R5430 GND.n1195 GND.n942 22.5005
R5431 GND.n970 GND.n955 22.5005
R5432 GND.n1174 GND.n970 22.5005
R5433 GND.n965 GND.n964 22.5005
R5434 GND.n965 GND.n961 22.5005
R5435 GND.n1255 GND.n952 22.5005
R5436 GND.n952 GND.n948 22.5005
R5437 GND.n955 GND.n951 22.5005
R5438 GND.n951 GND.n942 22.5005
R5439 GND.n1226 GND.n1221 22.5005
R5440 GND.n1221 GND.n1174 22.5005
R5441 GND.n1222 GND.n1220 22.5005
R5442 GND.n1220 GND.n961 22.5005
R5443 GND.n1240 GND.n1239 22.5005
R5444 GND.n1239 GND.n948 22.5005
R5445 GND.n1226 GND.n1225 22.5005
R5446 GND.n1225 GND.n942 22.5005
R5447 GND.n1338 GND.n1337 22.5005
R5448 GND.n1337 GND.n1304 22.5005
R5449 GND.n1332 GND.n1331 22.5005
R5450 GND.n1331 GND.n1293 22.5005
R5451 GND.n1328 GND.n1327 22.5005
R5452 GND.n1327 GND.n1280 22.5005
R5453 GND.n1338 GND.n1325 22.5005
R5454 GND.n1325 GND.n1274 22.5005
R5455 GND.n1302 GND.n1287 22.5005
R5456 GND.n1304 GND.n1302 22.5005
R5457 GND.n1297 GND.n1296 22.5005
R5458 GND.n1297 GND.n1293 22.5005
R5459 GND.n1385 GND.n1284 22.5005
R5460 GND.n1284 GND.n1280 22.5005
R5461 GND.n1287 GND.n1283 22.5005
R5462 GND.n1283 GND.n1274 22.5005
R5463 GND.n1356 GND.n1351 22.5005
R5464 GND.n1351 GND.n1304 22.5005
R5465 GND.n1352 GND.n1350 22.5005
R5466 GND.n1350 GND.n1293 22.5005
R5467 GND.n1370 GND.n1369 22.5005
R5468 GND.n1369 GND.n1280 22.5005
R5469 GND.n1356 GND.n1355 22.5005
R5470 GND.n1355 GND.n1274 22.5005
R5471 GND.n1478 GND.n1477 22.5005
R5472 GND.n1477 GND.n928 22.5005
R5473 GND.n1472 GND.n1471 22.5005
R5474 GND.n1471 GND.n1418 22.5005
R5475 GND.n1467 GND.n1438 22.5005
R5476 GND.n1467 GND.n1466 22.5005
R5477 GND.n1478 GND.n931 22.5005
R5478 GND.n1518 GND.n931 22.5005
R5479 GND.n1503 GND.n1412 22.5005
R5480 GND.n1412 GND.n928 22.5005
R5481 GND.n1422 GND.n1420 22.5005
R5482 GND.n1420 GND.n1418 22.5005
R5483 GND.n1463 GND.n1462 22.5005
R5484 GND.n1466 GND.n1463 22.5005
R5485 GND.n1503 GND.n932 22.5005
R5486 GND.n1518 GND.n932 22.5005
R5487 GND.n1510 GND.n1408 22.5005
R5488 GND.n1408 GND.n928 22.5005
R5489 GND.n1492 GND.n1490 22.5005
R5490 GND.n1490 GND.n1418 22.5005
R5491 GND.n1446 GND.n1445 22.5005
R5492 GND.n1466 GND.n1446 22.5005
R5493 GND.n1510 GND.n929 22.5005
R5494 GND.n1518 GND.n929 22.5005
R5495 GND.n158 GND.n134 22.5005
R5496 GND.t596 GND.n134 22.5005
R5497 GND.n3969 GND.n135 22.5005
R5498 GND.t596 GND.n135 22.5005
R5499 GND.n346 GND.n344 22.5005
R5500 GND.t107 GND.n346 22.5005
R5501 GND.n347 GND.n345 22.5005
R5502 GND.t107 GND.n347 22.5005
R5503 GND.n2764 GND.n2739 22.5005
R5504 GND.t568 GND.n2739 22.5005
R5505 GND.n2793 GND.n2740 22.5005
R5506 GND.t568 GND.n2740 22.5005
R5507 GND.n656 GND.n654 22.5005
R5508 GND.t514 GND.n654 22.5005
R5509 GND.n655 GND.n653 22.5005
R5510 GND.t514 GND.n653 22.5005
R5511 GND.n652 GND.n650 22.5005
R5512 GND.t219 GND.n650 22.5005
R5513 GND.n651 GND.n649 22.5005
R5514 GND.t219 GND.n649 22.5005
R5515 GND.n2252 GND.n2251 22.5005
R5516 GND.n2251 GND.t339 22.5005
R5517 GND.n2250 GND.n2249 22.5005
R5518 GND.t339 GND.n2250 22.5005
R5519 GND.n2228 GND.n2227 22.5005
R5520 GND.n2227 GND.t308 22.5005
R5521 GND.n2226 GND.n2225 22.5005
R5522 GND.t308 GND.n2226 22.5005
R5523 GND.n2208 GND.n2206 22.5005
R5524 GND.t338 GND.n2206 22.5005
R5525 GND.n2207 GND.n2205 22.5005
R5526 GND.t338 GND.n2205 22.5005
R5527 GND.n519 GND.n517 22.5005
R5528 GND.t200 GND.n517 22.5005
R5529 GND.n518 GND.n516 22.5005
R5530 GND.t200 GND.n516 22.5005
R5531 GND.n506 GND.n504 22.5005
R5532 GND.t268 GND.n504 22.5005
R5533 GND.n505 GND.n503 22.5005
R5534 GND.t268 GND.n503 22.5005
R5535 GND.n502 GND.n500 22.5005
R5536 GND.t48 GND.n500 22.5005
R5537 GND.n501 GND.n499 22.5005
R5538 GND.t48 GND.n499 22.5005
R5539 GND.n2894 GND.n2893 22.5005
R5540 GND.n2893 GND.t120 22.5005
R5541 GND.n2892 GND.n2891 22.5005
R5542 GND.t120 GND.n2892 22.5005
R5543 GND.n323 GND.n321 22.5005
R5544 GND.t361 GND.n321 22.5005
R5545 GND.n322 GND.n320 22.5005
R5546 GND.t361 GND.n320 22.5005
R5547 GND.n764 GND.n763 22.5005
R5548 GND.n763 GND.t56 22.5005
R5549 GND.n762 GND.n761 22.5005
R5550 GND.t56 GND.n762 22.5005
R5551 GND.n678 GND.n676 22.5005
R5552 GND.t337 GND.n676 22.5005
R5553 GND.n677 GND.n675 22.5005
R5554 GND.t337 GND.n675 22.5005
R5555 GND.n674 GND.n672 22.5005
R5556 GND.t315 GND.n672 22.5005
R5557 GND.n673 GND.n671 22.5005
R5558 GND.t315 GND.n671 22.5005
R5559 GND.n669 GND.n667 22.5005
R5560 GND.t667 GND.n667 22.5005
R5561 GND.n668 GND.n666 22.5005
R5562 GND.t667 GND.n666 22.5005
R5563 GND.n2075 GND.n704 22.5005
R5564 GND.t367 GND.n704 22.5005
R5565 GND.n719 GND.n718 22.5005
R5566 GND.t367 GND.n719 22.5005
R5567 GND.n2069 GND.n708 22.5005
R5568 GND.t121 GND.n708 22.5005
R5569 GND.n722 GND.n709 22.5005
R5570 GND.n722 GND.t121 22.5005
R5571 GND.n22 GND.n20 22.5005
R5572 GND.t570 GND.n22 22.5005
R5573 GND.n21 GND.n19 22.5005
R5574 GND.t570 GND.n21 22.5005
R5575 GND.n328 GND.n326 22.5005
R5576 GND.t64 GND.n326 22.5005
R5577 GND.n327 GND.n325 22.5005
R5578 GND.t64 GND.n325 22.5005
R5579 GND.n333 GND.n331 22.5005
R5580 GND.t214 GND.n331 22.5005
R5581 GND.n332 GND.n330 22.5005
R5582 GND.t214 GND.n330 22.5005
R5583 GND.n3408 GND.n3407 22.5005
R5584 GND.n3407 GND.t668 22.5005
R5585 GND.n3406 GND.n3405 22.5005
R5586 GND.t668 GND.n3406 22.5005
R5587 GND.n191 GND.n189 22.5005
R5588 GND.t287 GND.n189 22.5005
R5589 GND.n190 GND.n188 22.5005
R5590 GND.t287 GND.n188 22.5005
R5591 GND.n3952 GND.n3951 22.5005
R5592 GND.n3951 GND.t340 22.5005
R5593 GND.n3950 GND.n3949 22.5005
R5594 GND.t340 GND.n3950 22.5005
R5595 GND.n3928 GND.n3927 22.5005
R5596 GND.n3927 GND.t328 22.5005
R5597 GND.n3926 GND.n3925 22.5005
R5598 GND.t328 GND.n3926 22.5005
R5599 GND.n9 GND.n6 22.5005
R5600 GND.t507 GND.n9 22.5005
R5601 GND.n8 GND.n7 22.5005
R5602 GND.t507 GND.n8 22.5005
R5603 GND.n3617 GND.n3616 22.5005
R5604 GND.n3616 GND.t296 22.5005
R5605 GND.n3615 GND.n3614 22.5005
R5606 GND.t296 GND.n3615 22.5005
R5607 GND.n254 GND.n252 22.5005
R5608 GND.t682 GND.n252 22.5005
R5609 GND.n253 GND.n251 22.5005
R5610 GND.t682 GND.n251 22.5005
R5611 GND.n272 GND.n270 22.5005
R5612 GND.t184 GND.n270 22.5005
R5613 GND.n271 GND.n269 22.5005
R5614 GND.t184 GND.n269 22.5005
R5615 GND.n280 GND.n278 22.5005
R5616 GND.t168 GND.n278 22.5005
R5617 GND.n279 GND.n277 22.5005
R5618 GND.t168 GND.n277 22.5005
R5619 GND.n288 GND.n286 22.5005
R5620 GND.t613 GND.n286 22.5005
R5621 GND.n287 GND.n285 22.5005
R5622 GND.t613 GND.n285 22.5005
R5623 GND.n296 GND.n294 22.5005
R5624 GND.t650 GND.n294 22.5005
R5625 GND.n295 GND.n293 22.5005
R5626 GND.t650 GND.n293 22.5005
R5627 GND.n304 GND.n302 22.5005
R5628 GND.t245 GND.n302 22.5005
R5629 GND.n303 GND.n301 22.5005
R5630 GND.t245 GND.n301 22.5005
R5631 GND.n196 GND.n194 22.5005
R5632 GND.t238 GND.n194 22.5005
R5633 GND.n195 GND.n193 22.5005
R5634 GND.t238 GND.n193 22.5005
R5635 GND.n686 GND.n682 22.5005
R5636 GND.t177 GND.n682 22.5005
R5637 GND.n2098 GND.n2097 22.5005
R5638 GND.t177 GND.n2098 22.5005
R5639 GND.n1090 GND.n997 22.5005
R5640 GND.t666 GND.n997 22.5005
R5641 GND.n999 GND.n996 22.5005
R5642 GND.t666 GND.n996 22.5005
R5643 GND.n1036 GND.n1035 22.5005
R5644 GND.n1035 GND.n981 22.5005
R5645 GND.n1041 GND.n1040 22.5005
R5646 GND.n1040 GND.n983 22.5005
R5647 GND.n1061 GND.n1013 22.5005
R5648 GND.n1013 GND.n981 22.5005
R5649 GND.n1015 GND.n1012 22.5005
R5650 GND.n1012 GND.n983 22.5005
R5651 GND.n1025 GND.n1024 22.5005
R5652 GND.n1024 GND.n981 22.5005
R5653 GND.n1018 GND.n1017 22.5005
R5654 GND.n1017 GND.n983 22.5005
R5655 GND.n980 GND.n978 22.5005
R5656 GND.t677 GND.n980 22.5005
R5657 GND.n979 GND.n977 22.5005
R5658 GND.t677 GND.n979 22.5005
R5659 GND.n1162 GND.n1161 22.5005
R5660 GND.t251 GND.n1162 22.5005
R5661 GND.n1164 GND.n1163 22.5005
R5662 GND.n1163 GND.t251 22.5005
R5663 GND.n2059 GND.n2058 22.5005
R5664 GND.t311 GND.n2059 22.5005
R5665 GND.n2061 GND.n2060 22.5005
R5666 GND.n2060 GND.t311 22.5005
R5667 GND.n2039 GND.n2038 22.5005
R5668 GND.t320 GND.n2039 22.5005
R5669 GND.n2041 GND.n2040 22.5005
R5670 GND.n2040 GND.t320 22.5005
R5671 GND.n2032 GND.n805 22.5005
R5672 GND.t110 GND.n805 22.5005
R5673 GND.n846 GND.n804 22.5005
R5674 GND.t110 GND.n804 22.5005
R5675 GND.n2018 GND.n814 22.5005
R5676 GND.t619 GND.n814 22.5005
R5677 GND.n866 GND.n813 22.5005
R5678 GND.t619 GND.n813 22.5005
R5679 GND.n1952 GND.n1951 22.5005
R5680 GND.n1951 GND.n885 22.5005
R5681 GND.n1946 GND.n1945 22.5005
R5682 GND.n1945 GND.n1892 22.5005
R5683 GND.n1941 GND.n1912 22.5005
R5684 GND.n1941 GND.n1940 22.5005
R5685 GND.n1952 GND.n888 22.5005
R5686 GND.n1992 GND.n888 22.5005
R5687 GND.n1977 GND.n1886 22.5005
R5688 GND.n1886 GND.n885 22.5005
R5689 GND.n1896 GND.n1894 22.5005
R5690 GND.n1894 GND.n1892 22.5005
R5691 GND.n1937 GND.n1936 22.5005
R5692 GND.n1940 GND.n1937 22.5005
R5693 GND.n1977 GND.n889 22.5005
R5694 GND.n1992 GND.n889 22.5005
R5695 GND.n1984 GND.n1882 22.5005
R5696 GND.n1882 GND.n885 22.5005
R5697 GND.n1966 GND.n1964 22.5005
R5698 GND.n1964 GND.n1892 22.5005
R5699 GND.n1920 GND.n1919 22.5005
R5700 GND.n1940 GND.n1920 22.5005
R5701 GND.n1984 GND.n886 22.5005
R5702 GND.n1992 GND.n886 22.5005
R5703 GND.n1998 GND.n1997 22.5005
R5704 GND.t158 GND.n1998 22.5005
R5705 GND.n2000 GND.n1999 22.5005
R5706 GND.n1999 GND.t158 22.5005
R5707 GND.n2285 GND.n2284 22.5005
R5708 GND.t569 GND.n2285 22.5005
R5709 GND.n2287 GND.n2286 22.5005
R5710 GND.n2286 GND.t569 22.5005
R5711 GND.n2298 GND.n619 22.5005
R5712 GND.n2298 GND.t157 22.5005
R5713 GND.n620 GND.n618 22.5005
R5714 GND.t157 GND.n620 22.5005
R5715 GND.n1686 GND.n1685 22.5005
R5716 GND.n1685 GND.n1652 22.5005
R5717 GND.n1680 GND.n1679 22.5005
R5718 GND.n1679 GND.n1642 22.5005
R5719 GND.n1676 GND.n1675 22.5005
R5720 GND.n1675 GND.n1629 22.5005
R5721 GND.n1686 GND.n1673 22.5005
R5722 GND.n1673 GND.n1623 22.5005
R5723 GND.n1651 GND.n1636 22.5005
R5724 GND.n1652 GND.n1651 22.5005
R5725 GND.n1646 GND.n1645 22.5005
R5726 GND.n1646 GND.n1642 22.5005
R5727 GND.n1733 GND.n1633 22.5005
R5728 GND.n1633 GND.n1629 22.5005
R5729 GND.n1636 GND.n1632 22.5005
R5730 GND.n1632 GND.n1623 22.5005
R5731 GND.n1704 GND.n1699 22.5005
R5732 GND.n1699 GND.n1652 22.5005
R5733 GND.n1700 GND.n1698 22.5005
R5734 GND.n1698 GND.n1642 22.5005
R5735 GND.n1718 GND.n1717 22.5005
R5736 GND.n1717 GND.n1629 22.5005
R5737 GND.n1704 GND.n1703 22.5005
R5738 GND.n1703 GND.n1623 22.5005
R5739 GND.n2428 GND.n2427 22.5005
R5740 GND.n2427 GND.n2394 22.5005
R5741 GND.n2422 GND.n2421 22.5005
R5742 GND.n2421 GND.n589 22.5005
R5743 GND.n2418 GND.n2417 22.5005
R5744 GND.n2417 GND.n576 22.5005
R5745 GND.n2428 GND.n2415 22.5005
R5746 GND.n2415 GND.n570 22.5005
R5747 GND.n598 GND.n583 22.5005
R5748 GND.n2394 GND.n598 22.5005
R5749 GND.n593 GND.n592 22.5005
R5750 GND.n593 GND.n589 22.5005
R5751 GND.n2475 GND.n580 22.5005
R5752 GND.n580 GND.n576 22.5005
R5753 GND.n583 GND.n579 22.5005
R5754 GND.n579 GND.n570 22.5005
R5755 GND.n2446 GND.n2441 22.5005
R5756 GND.n2441 GND.n2394 22.5005
R5757 GND.n2442 GND.n2440 22.5005
R5758 GND.n2440 GND.n589 22.5005
R5759 GND.n2460 GND.n2459 22.5005
R5760 GND.n2459 GND.n576 22.5005
R5761 GND.n2446 GND.n2445 22.5005
R5762 GND.n2445 GND.n570 22.5005
R5763 GND.n2328 GND.n600 22.5005
R5764 GND.t54 GND.n600 22.5005
R5765 GND.n2391 GND.n2390 22.5005
R5766 GND.t54 GND.n2391 22.5005
R5767 GND.n2382 GND.n2381 22.5005
R5768 GND.t250 GND.n2382 22.5005
R5769 GND.n2384 GND.n2383 22.5005
R5770 GND.n2383 GND.t250 22.5005
R5771 GND.n2821 GND.n2820 22.5005
R5772 GND.t227 GND.n2821 22.5005
R5773 GND.n2823 GND.n2822 22.5005
R5774 GND.n2822 GND.t227 22.5005
R5775 GND.n2698 GND.n2697 22.5005
R5776 GND.n2697 GND.n556 22.5005
R5777 GND.n2692 GND.n2691 22.5005
R5778 GND.n2691 GND.n2638 22.5005
R5779 GND.n2687 GND.n2658 22.5005
R5780 GND.n2687 GND.n2686 22.5005
R5781 GND.n2698 GND.n559 22.5005
R5782 GND.n2738 GND.n559 22.5005
R5783 GND.n2723 GND.n2632 22.5005
R5784 GND.n2632 GND.n556 22.5005
R5785 GND.n2642 GND.n2640 22.5005
R5786 GND.n2640 GND.n2638 22.5005
R5787 GND.n2683 GND.n2682 22.5005
R5788 GND.n2686 GND.n2683 22.5005
R5789 GND.n2723 GND.n560 22.5005
R5790 GND.n2738 GND.n560 22.5005
R5791 GND.n2730 GND.n2628 22.5005
R5792 GND.n2628 GND.n556 22.5005
R5793 GND.n2712 GND.n2710 22.5005
R5794 GND.n2710 GND.n2638 22.5005
R5795 GND.n2666 GND.n2665 22.5005
R5796 GND.n2686 GND.n2666 22.5005
R5797 GND.n2730 GND.n557 22.5005
R5798 GND.n2738 GND.n557 22.5005
R5799 GND.n2801 GND.n2800 22.5005
R5800 GND.t723 GND.n2801 22.5005
R5801 GND.n2803 GND.n2802 22.5005
R5802 GND.n2802 GND.t723 22.5005
R5803 GND.n2982 GND.n2981 22.5005
R5804 GND.n2981 GND.n2948 22.5005
R5805 GND.n2976 GND.n2975 22.5005
R5806 GND.n2975 GND.n476 22.5005
R5807 GND.n2972 GND.n2971 22.5005
R5808 GND.n2971 GND.n463 22.5005
R5809 GND.n2982 GND.n2969 22.5005
R5810 GND.n2969 GND.n457 22.5005
R5811 GND.n485 GND.n470 22.5005
R5812 GND.n2948 GND.n485 22.5005
R5813 GND.n480 GND.n479 22.5005
R5814 GND.n480 GND.n476 22.5005
R5815 GND.n3029 GND.n467 22.5005
R5816 GND.n467 GND.n463 22.5005
R5817 GND.n470 GND.n466 22.5005
R5818 GND.n466 GND.n457 22.5005
R5819 GND.n3000 GND.n2995 22.5005
R5820 GND.n2995 GND.n2948 22.5005
R5821 GND.n2996 GND.n2994 22.5005
R5822 GND.n2994 GND.n476 22.5005
R5823 GND.n3014 GND.n3013 22.5005
R5824 GND.n3013 GND.n463 22.5005
R5825 GND.n3000 GND.n2999 22.5005
R5826 GND.n2999 GND.n457 22.5005
R5827 GND.n2902 GND.n487 22.5005
R5828 GND.t292 GND.n487 22.5005
R5829 GND.n2945 GND.n2944 22.5005
R5830 GND.t292 GND.n2945 22.5005
R5831 GND.n3337 GND.n353 22.5005
R5832 GND.t605 GND.n353 22.5005
R5833 GND.n2927 GND.n352 22.5005
R5834 GND.t605 GND.n352 22.5005
R5835 GND.n444 GND.n443 22.5005
R5836 GND.n443 GND.n385 22.5005
R5837 GND.n433 GND.n360 22.5005
R5838 GND.n3332 GND.n360 22.5005
R5839 GND.n438 GND.n437 22.5005
R5840 GND.n437 GND.n94 22.5005
R5841 GND.n445 GND.n444 22.5005
R5842 GND.n3319 GND.n445 22.5005
R5843 GND.n3321 GND.n370 22.5005
R5844 GND.n385 GND.n370 22.5005
R5845 GND.n376 GND.n358 22.5005
R5846 GND.n3332 GND.n358 22.5005
R5847 GND.n381 GND.n373 22.5005
R5848 GND.n373 GND.n94 22.5005
R5849 GND.n3321 GND.n3320 22.5005
R5850 GND.n3320 GND.n3319 22.5005
R5851 GND.n384 GND.n366 22.5005
R5852 GND.n385 GND.n384 22.5005
R5853 GND.n3331 GND.n3330 22.5005
R5854 GND.n3332 GND.n3331 22.5005
R5855 GND.n3308 GND.n3306 22.5005
R5856 GND.n3308 GND.n94 22.5005
R5857 GND.n386 GND.n366 22.5005
R5858 GND.n3319 GND.n386 22.5005
R5859 GND.n3239 GND.n3238 22.5005
R5860 GND.n3238 GND.n92 22.5005
R5861 GND.n3233 GND.n3232 22.5005
R5862 GND.n3232 GND.n3196 22.5005
R5863 GND.n3229 GND.n3228 22.5005
R5864 GND.n3228 GND.n3183 22.5005
R5865 GND.n3239 GND.n3226 22.5005
R5866 GND.n3226 GND.n93 22.5005
R5867 GND.n3201 GND.n3190 22.5005
R5868 GND.n3201 GND.n92 22.5005
R5869 GND.n3200 GND.n3199 22.5005
R5870 GND.n3200 GND.n3196 22.5005
R5871 GND.n3286 GND.n3187 22.5005
R5872 GND.n3187 GND.n3183 22.5005
R5873 GND.n3190 GND.n3186 22.5005
R5874 GND.n3186 GND.n93 22.5005
R5875 GND.n3257 GND.n3252 22.5005
R5876 GND.n3252 GND.n92 22.5005
R5877 GND.n3253 GND.n3251 22.5005
R5878 GND.n3251 GND.n3196 22.5005
R5879 GND.n3271 GND.n3270 22.5005
R5880 GND.n3270 GND.n3183 22.5005
R5881 GND.n3257 GND.n3256 22.5005
R5882 GND.n3256 GND.n93 22.5005
R5883 GND.n101 GND.n95 22.5005
R5884 GND.t699 GND.n95 22.5005
R5885 GND.n3994 GND.n3993 22.5005
R5886 GND.t699 GND.n3994 22.5005
R5887 GND.n131 GND.n130 22.5005
R5888 GND.n130 GND.t153 22.5005
R5889 GND.n3976 GND.n3975 22.5005
R5890 GND.n3975 GND.t153 22.5005
R5891 GND.n4162 GND.n4161 22.5005
R5892 GND.n4161 GND.n4128 22.5005
R5893 GND.n4156 GND.n4155 22.5005
R5894 GND.n4155 GND.n4118 22.5005
R5895 GND.n4152 GND.n4151 22.5005
R5896 GND.n4151 GND.n4105 22.5005
R5897 GND.n4162 GND.n4149 22.5005
R5898 GND.n4149 GND.n4099 22.5005
R5899 GND.n4127 GND.n4112 22.5005
R5900 GND.n4128 GND.n4127 22.5005
R5901 GND.n4122 GND.n4121 22.5005
R5902 GND.n4122 GND.n4118 22.5005
R5903 GND.n4209 GND.n4109 22.5005
R5904 GND.n4109 GND.n4105 22.5005
R5905 GND.n4112 GND.n4108 22.5005
R5906 GND.n4108 GND.n4099 22.5005
R5907 GND.n4180 GND.n4175 22.5005
R5908 GND.n4175 GND.n4128 22.5005
R5909 GND.n4176 GND.n4174 22.5005
R5910 GND.n4174 GND.n4118 22.5005
R5911 GND.n4194 GND.n4193 22.5005
R5912 GND.n4193 GND.n4105 22.5005
R5913 GND.n4180 GND.n4179 22.5005
R5914 GND.n4179 GND.n4099 22.5005
R5915 GND.n4292 GND.n45 22.5005
R5916 GND.t295 GND.n45 22.5005
R5917 GND.n180 GND.n44 22.5005
R5918 GND.t295 GND.n44 22.5005
R5919 GND.n4319 GND.n28 22.5005
R5920 GND.n28 GND.t45 22.5005
R5921 GND.n4308 GND.n27 22.5005
R5922 GND.t45 GND.n27 22.5005
R5923 GND.n4277 GND.n4276 22.5005
R5924 GND.n4276 GND.n4275 22.5005
R5925 GND.n4233 GND.n50 22.5005
R5926 GND.n4287 GND.n50 22.5005
R5927 GND.n4236 GND.n57 22.5005
R5928 GND.n4275 GND.n4236 22.5005
R5929 GND.n4286 GND.n4285 22.5005
R5930 GND.n4287 GND.n4286 22.5005
R5931 GND.n4274 GND.n4273 22.5005
R5932 GND.n4275 GND.n4274 22.5005
R5933 GND.n4243 GND.n52 22.5005
R5934 GND.n4287 GND.n52 22.5005
R5935 GND.n2489 GND 22.3388
R5936 GND.n3812 GND 22.2668
R5937 GND.n4369 GND 20.4446
R5938 GND.n3817 GND 20.3617
R5939 GND.n2618 GND 20.2611
R5940 GND.n2619 GND 19.547
R5941 GND.n3474 GND 18.8872
R5942 GND.n2065 GND.n2064 18.6076
R5943 GND.n864 GND.n670 18.6076
R5944 GND.n2256 GND.n2255 18.6076
R5945 GND.n2827 GND.n2826 18.6076
R5946 GND.n2898 GND.n2897 18.6076
R5947 GND.n3382 GND.n3381 18.6076
R5948 GND.n3956 GND.n3955 18.6076
R5949 GND.n3822 GND 18.4566
R5950 GND.n2311 GND.t293 18.3746
R5951 GND.t197 GND.n774 18.3746
R5952 GND.n1094 GND.t136 18.3746
R5953 GND.t46 GND.n817 18.3746
R5954 GND.t506 GND.n527 18.3746
R5955 GND.n2916 GND.t229 18.3746
R5956 GND.n114 GND.t230 18.3746
R5957 GND.t310 GND.n4297 18.3746
R5958 GND.n2620 GND 17.7231
R5959 GND.n452 GND 16.7552
R5960 GND.n3827 GND 16.5516
R5961 GND.n3042 GND 15.1851
R5962 GND.n3832 GND 14.6465
R5963 GND.n3043 GND 13.9634
R5964 GND.n4016 GND.n4011 13.8976
R5965 GND.n4016 GND.n4015 13.8976
R5966 GND.n4039 GND.n4004 13.8976
R5967 GND.n4040 GND.n4039 13.8976
R5968 GND.n4056 GND.n74 13.8976
R5969 GND.n4078 GND.n4077 13.8976
R5970 GND.n4067 GND.n4048 13.8976
R5971 GND.n4062 GND.n4061 13.8976
R5972 GND.n4034 GND.n4019 13.8976
R5973 GND.n4031 GND.n4029 13.8976
R5974 GND.n417 GND.n416 13.8976
R5975 GND.n418 GND.n417 13.8976
R5976 GND.n424 GND.n405 13.8976
R5977 GND.n424 GND.n423 13.8976
R5978 GND.n3322 GND.n369 13.8976
R5979 GND.n379 GND.n371 13.8976
R5980 GND.n3312 GND.n3311 13.8976
R5981 GND.n3328 GND.n3327 13.8976
R5982 GND.n435 GND.n390 13.8976
R5983 GND.n440 GND.n431 13.8976
R5984 GND.n3094 GND.n3089 13.8976
R5985 GND.n3094 GND.n3093 13.8976
R5986 GND.n3117 GND.n3082 13.8976
R5987 GND.n3118 GND.n3117 13.8976
R5988 GND.n3134 GND.n3059 13.8976
R5989 GND.n3156 GND.n3155 13.8976
R5990 GND.n3145 GND.n3126 13.8976
R5991 GND.n3140 GND.n3139 13.8976
R5992 GND.n3112 GND.n3097 13.8976
R5993 GND.n3109 GND.n3107 13.8976
R5994 GND.n2541 GND.n2536 13.8976
R5995 GND.n2541 GND.n2540 13.8976
R5996 GND.n2564 GND.n2529 13.8976
R5997 GND.n2565 GND.n2564 13.8976
R5998 GND.n2581 GND.n2505 13.8976
R5999 GND.n2603 GND.n2602 13.8976
R6000 GND.n2592 GND.n2573 13.8976
R6001 GND.n2587 GND.n2586 13.8976
R6002 GND.n2559 GND.n2544 13.8976
R6003 GND.n2556 GND.n2554 13.8976
R6004 GND.n1796 GND.n1791 13.8976
R6005 GND.n1796 GND.n1795 13.8976
R6006 GND.n1819 GND.n1784 13.8976
R6007 GND.n1820 GND.n1819 13.8976
R6008 GND.n1836 GND.n1762 13.8976
R6009 GND.n1858 GND.n1857 13.8976
R6010 GND.n1847 GND.n1828 13.8976
R6011 GND.n1842 GND.n1841 13.8976
R6012 GND.n1814 GND.n1799 13.8976
R6013 GND.n1811 GND.n1809 13.8976
R6014 GND.n1539 GND.n1534 13.8976
R6015 GND.n1539 GND.n1538 13.8976
R6016 GND.n1562 GND.n1527 13.8976
R6017 GND.n1563 GND.n1562 13.8976
R6018 GND.n1579 GND.n910 13.8976
R6019 GND.n1601 GND.n1600 13.8976
R6020 GND.n1590 GND.n1571 13.8976
R6021 GND.n1585 GND.n1584 13.8976
R6022 GND.n1557 GND.n1542 13.8976
R6023 GND.n1554 GND.n1552 13.8976
R6024 GND.n1191 GND.n1186 13.8976
R6025 GND.n1191 GND.n1190 13.8976
R6026 GND.n1214 GND.n1179 13.8976
R6027 GND.n1215 GND.n1214 13.8976
R6028 GND.n1231 GND.n953 13.8976
R6029 GND.n1253 GND.n1252 13.8976
R6030 GND.n1242 GND.n1223 13.8976
R6031 GND.n1237 GND.n1236 13.8976
R6032 GND.n1209 GND.n1194 13.8976
R6033 GND.n1206 GND.n1204 13.8976
R6034 GND.n1321 GND.n1316 13.8976
R6035 GND.n1321 GND.n1320 13.8976
R6036 GND.n1344 GND.n1309 13.8976
R6037 GND.n1345 GND.n1344 13.8976
R6038 GND.n1361 GND.n1285 13.8976
R6039 GND.n1383 GND.n1382 13.8976
R6040 GND.n1372 GND.n1353 13.8976
R6041 GND.n1367 GND.n1366 13.8976
R6042 GND.n1339 GND.n1324 13.8976
R6043 GND.n1336 GND.n1334 13.8976
R6044 GND.n1454 GND.n1453 13.8976
R6045 GND.n1453 GND.n1452 13.8976
R6046 GND.n1484 GND.n1432 13.8976
R6047 GND.n1485 GND.n1484 13.8976
R6048 GND.n1504 GND.n1411 13.8976
R6049 GND.n1502 GND.n1413 13.8976
R6050 GND.n1511 GND.n1407 13.8976
R6051 GND.n1509 GND.n1409 13.8976
R6052 GND.n1479 GND.n1437 13.8976
R6053 GND.n1476 GND.n1474 13.8976
R6054 GND.n1928 GND.n1927 13.8976
R6055 GND.n1927 GND.n1926 13.8976
R6056 GND.n1958 GND.n1906 13.8976
R6057 GND.n1959 GND.n1958 13.8976
R6058 GND.n1978 GND.n1885 13.8976
R6059 GND.n1976 GND.n1887 13.8976
R6060 GND.n1985 GND.n1881 13.8976
R6061 GND.n1983 GND.n1883 13.8976
R6062 GND.n1953 GND.n1911 13.8976
R6063 GND.n1950 GND.n1948 13.8976
R6064 GND.n1669 GND.n1664 13.8976
R6065 GND.n1669 GND.n1668 13.8976
R6066 GND.n1692 GND.n1657 13.8976
R6067 GND.n1693 GND.n1692 13.8976
R6068 GND.n1709 GND.n1634 13.8976
R6069 GND.n1731 GND.n1730 13.8976
R6070 GND.n1720 GND.n1701 13.8976
R6071 GND.n1715 GND.n1714 13.8976
R6072 GND.n1687 GND.n1672 13.8976
R6073 GND.n1684 GND.n1682 13.8976
R6074 GND.n2411 GND.n2406 13.8976
R6075 GND.n2411 GND.n2410 13.8976
R6076 GND.n2434 GND.n2399 13.8976
R6077 GND.n2435 GND.n2434 13.8976
R6078 GND.n2451 GND.n581 13.8976
R6079 GND.n2473 GND.n2472 13.8976
R6080 GND.n2462 GND.n2443 13.8976
R6081 GND.n2457 GND.n2456 13.8976
R6082 GND.n2429 GND.n2414 13.8976
R6083 GND.n2426 GND.n2424 13.8976
R6084 GND.n2674 GND.n2673 13.8976
R6085 GND.n2673 GND.n2672 13.8976
R6086 GND.n2704 GND.n2652 13.8976
R6087 GND.n2705 GND.n2704 13.8976
R6088 GND.n2724 GND.n2631 13.8976
R6089 GND.n2722 GND.n2633 13.8976
R6090 GND.n2731 GND.n2627 13.8976
R6091 GND.n2729 GND.n2629 13.8976
R6092 GND.n2699 GND.n2657 13.8976
R6093 GND.n2696 GND.n2694 13.8976
R6094 GND.n2965 GND.n2960 13.8976
R6095 GND.n2965 GND.n2964 13.8976
R6096 GND.n2988 GND.n2953 13.8976
R6097 GND.n2989 GND.n2988 13.8976
R6098 GND.n3005 GND.n468 13.8976
R6099 GND.n3027 GND.n3026 13.8976
R6100 GND.n3016 GND.n2997 13.8976
R6101 GND.n3011 GND.n3010 13.8976
R6102 GND.n2983 GND.n2968 13.8976
R6103 GND.n2980 GND.n2978 13.8976
R6104 GND.n3222 GND.n3217 13.8976
R6105 GND.n3222 GND.n3221 13.8976
R6106 GND.n3245 GND.n3210 13.8976
R6107 GND.n3246 GND.n3245 13.8976
R6108 GND.n3262 GND.n3188 13.8976
R6109 GND.n3284 GND.n3283 13.8976
R6110 GND.n3273 GND.n3254 13.8976
R6111 GND.n3268 GND.n3267 13.8976
R6112 GND.n3240 GND.n3225 13.8976
R6113 GND.n3237 GND.n3235 13.8976
R6114 GND.n4145 GND.n4140 13.8976
R6115 GND.n4145 GND.n4144 13.8976
R6116 GND.n4168 GND.n4133 13.8976
R6117 GND.n4169 GND.n4168 13.8976
R6118 GND.n4185 GND.n4110 13.8976
R6119 GND.n4207 GND.n4206 13.8976
R6120 GND.n4196 GND.n4177 13.8976
R6121 GND.n4191 GND.n4190 13.8976
R6122 GND.n4163 GND.n4148 13.8976
R6123 GND.n4160 GND.n4158 13.8976
R6124 GND.n3876 GND 13.2342
R6125 GND.n3837 GND 12.7414
R6126 GND.n3171 GND 12.6471
R6127 GND.n1074 GND.n1073 12.5667
R6128 GND.n3172 GND 11.1716
R6129 GND.n3842 GND 10.8363
R6130 GND.n4224 GND 10.1098
R6131 GND.n3300 GND 10.1091
R6132 GND.n198 GND 9.38722
R6133 GND.n688 GND.n243 9.19583
R6134 GND.n3627 GND.n3626 9.18625
R6135 GND.n4371 GND.n4370 9.18624
R6136 GND.n3864 GND.n3863 9.18624
R6137 GND.n3875 GND.n3874 9.18624
R6138 GND.n3482 GND.n201 9.18624
R6139 GND.n3473 GND.n204 9.18624
R6140 GND.n306 GND.n207 9.18624
R6141 GND.n3516 GND.n210 9.18624
R6142 GND.n298 GND.n213 9.18624
R6143 GND.n3546 GND.n216 9.18624
R6144 GND.n290 GND.n219 9.18624
R6145 GND.n282 GND.n222 9.18624
R6146 GND.n274 GND.n228 9.18624
R6147 GND.n266 GND.n231 9.18624
R6148 GND.n263 GND.n234 9.18624
R6149 GND.n3621 GND.n237 9.18624
R6150 GND.n3624 GND.n240 9.18624
R6151 GND.n3847 GND 8.93128
R6152 GND.n1084 GND.n1074 8.38868
R6153 GND.n3299 GND 8.37982
R6154 GND.n3478 GND.n3477 8.32958
R6155 GND.n3500 GND.n3499 8.32958
R6156 GND.n3522 GND.n3521 8.32958
R6157 GND.n3541 GND.n3540 8.32958
R6158 GND.n3563 GND.n3562 8.32958
R6159 GND.n3602 GND.n3601 8.32958
R6160 GND.n259 GND.n258 8.32958
R6161 GND.n3583 GND.n3582 7.9105
R6162 GND.n4221 GND.n4220 7.9105
R6163 GND.n4092 GND.n4091 7.9105
R6164 GND.n3298 GND.n3297 7.9105
R6165 GND.n3302 GND.n3301 7.9105
R6166 GND.n3170 GND.n3169 7.9105
R6167 GND.n3041 GND.n3040 7.9105
R6168 GND.n2622 GND.n2621 7.9105
R6169 GND.n2617 GND.n2616 7.9105
R6170 GND.n2487 GND.n2486 7.9105
R6171 GND.n1745 GND.n1744 7.9105
R6172 GND.n1872 GND.n1871 7.9105
R6173 GND.n1876 GND.n1875 7.9105
R6174 GND.n1615 GND.n1614 7.9105
R6175 GND.n1402 GND.n1401 7.9105
R6176 GND.n1397 GND.n1396 7.9105
R6177 GND.n1267 GND.n1266 7.9105
R6178 GND.n1073 GND.n1072 7.9105
R6179 GND.t158 GND.n1994 7.71078
R6180 GND.n3173 GND 7.57106
R6181 GND.n3852 GND 7.02622
R6182 GND.n3860 GND 6.6255
R6183 GND.n3626 GND.n3625 6.49778
R6184 GND.n3623 GND.n3622 6.43528
R6185 GND.n3860 GND.n198 6.43528
R6186 GND.n3862 GND.n3861 6.43528
R6187 GND.n265 GND 5.97876
R6188 GND.n3548 GND.n291 5.93528
R6189 GND.n58 GND 5.58802
R6190 GND.n305 GND 5.26137
R6191 GND.n3857 GND 5.12115
R6192 GND.n3485 GND.n3474 5.04398
R6193 GND.n4093 GND 5.03306
R6194 GND.n4052 GND 5.0168
R6195 GND.n4059 GND 5.0168
R6196 GND.n4037 GND 5.0168
R6197 GND.n3315 GND 5.0168
R6198 GND.n3325 GND 5.0168
R6199 GND.n426 GND 5.0168
R6200 GND.n3130 GND 5.0168
R6201 GND.n3137 GND 5.0168
R6202 GND.n3115 GND 5.0168
R6203 GND.n2577 GND 5.0168
R6204 GND.n2584 GND 5.0168
R6205 GND.n2562 GND 5.0168
R6206 GND.n1832 GND 5.0168
R6207 GND.n1839 GND 5.0168
R6208 GND.n1817 GND 5.0168
R6209 GND.n1575 GND 5.0168
R6210 GND.n1582 GND 5.0168
R6211 GND.n1560 GND 5.0168
R6212 GND.n1227 GND 5.0168
R6213 GND.n1234 GND 5.0168
R6214 GND.n1212 GND 5.0168
R6215 GND.n1357 GND 5.0168
R6216 GND.n1364 GND 5.0168
R6217 GND.n1342 GND 5.0168
R6218 GND.n1514 GND 5.0168
R6219 GND.n1507 GND 5.0168
R6220 GND.n1482 GND 5.0168
R6221 GND.n1019 GND 5.0168
R6222 GND.n1029 GND 5.0168
R6223 GND.n1045 GND 5.0168
R6224 GND.n1988 GND 5.0168
R6225 GND.n1981 GND 5.0168
R6226 GND.n1956 GND 5.0168
R6227 GND.n1705 GND 5.0168
R6228 GND.n1712 GND 5.0168
R6229 GND.n1690 GND 5.0168
R6230 GND.n2447 GND 5.0168
R6231 GND.n2454 GND 5.0168
R6232 GND.n2432 GND 5.0168
R6233 GND.n2734 GND 5.0168
R6234 GND.n2727 GND 5.0168
R6235 GND.n2702 GND 5.0168
R6236 GND.n3001 GND 5.0168
R6237 GND.n3008 GND 5.0168
R6238 GND.n2986 GND 5.0168
R6239 GND.n3258 GND 5.0168
R6240 GND.n3265 GND 5.0168
R6241 GND.n3243 GND 5.0168
R6242 GND.n4181 GND 5.0168
R6243 GND.n4188 GND 5.0168
R6244 GND.n4166 GND 5.0168
R6245 GND.n4268 GND 5.0168
R6246 GND.n4281 GND 5.0168
R6247 GND.n4224 GND 5.0168
R6248 GND.n265 GND 4.73963
R6249 GND.n3862 GND 4.63722
R6250 GND.n281 GND 4.37007
R6251 GND.n3587 GND.n275 4.32659
R6252 GND.n3788 GND.n239 4.15831
R6253 GND.n3793 GND.n236 4.15831
R6254 GND.n3798 GND.n233 4.15831
R6255 GND.n3803 GND.n230 4.15831
R6256 GND.n3808 GND.n227 4.15831
R6257 GND.n3813 GND.n224 4.15831
R6258 GND.n3818 GND.n221 4.15831
R6259 GND.n3823 GND.n218 4.15831
R6260 GND.n3828 GND.n215 4.15831
R6261 GND.n3833 GND.n212 4.15831
R6262 GND.n3838 GND.n209 4.15831
R6263 GND.n3843 GND.n206 4.15831
R6264 GND.n3848 GND.n203 4.15831
R6265 GND.n3853 GND.n200 4.15831
R6266 GND.n3873 GND.n3872 4.15831
R6267 GND.n3868 GND.n3867 4.15831
R6268 GND.n3781 GND.n3628 4.15828
R6269 GND.n4371 GND.n0 3.93605
R6270 GND.n3868 GND.n3864 3.93605
R6271 GND.n3874 GND.n3873 3.93605
R6272 GND.n3853 GND.n201 3.93605
R6273 GND.n3848 GND.n204 3.93605
R6274 GND.n3843 GND.n207 3.93605
R6275 GND.n3838 GND.n210 3.93605
R6276 GND.n3833 GND.n213 3.93605
R6277 GND.n3828 GND.n216 3.93605
R6278 GND.n3823 GND.n219 3.93605
R6279 GND.n3818 GND.n222 3.93605
R6280 GND.n3813 GND.n225 3.93605
R6281 GND.n3808 GND.n228 3.93605
R6282 GND.n3803 GND.n231 3.93605
R6283 GND.n3798 GND.n234 3.93605
R6284 GND.n3793 GND.n237 3.93605
R6285 GND.n3788 GND.n240 3.93605
R6286 GND.n3783 GND.n3627 3.93605
R6287 GND.n3679 GND.n3630 3.91224
R6288 GND.n4373 GND.n1 3.91156
R6289 GND.n3732 GND.n3731 3.90049
R6290 GND.n3782 GND.n3781 3.89978
R6291 GND.n3731 GND.n3730 3.88874
R6292 GND.n3785 GND.n242 3.88874
R6293 GND.n3681 GND.n3630 3.87628
R6294 GND.n4372 GND.n3 3.87628
R6295 GND.n3870 GND.n3859 3.87628
R6296 GND.n3856 GND.n199 3.87628
R6297 GND.n3851 GND.n202 3.87628
R6298 GND.n3846 GND.n205 3.87628
R6299 GND.n3841 GND.n208 3.87628
R6300 GND.n3836 GND.n211 3.87628
R6301 GND.n3831 GND.n214 3.87628
R6302 GND.n3826 GND.n217 3.87628
R6303 GND.n3821 GND.n220 3.87628
R6304 GND.n3816 GND.n223 3.87628
R6305 GND.n3811 GND.n226 3.87628
R6306 GND.n3806 GND.n229 3.87628
R6307 GND.n3801 GND.n232 3.87628
R6308 GND.n3796 GND.n235 3.87628
R6309 GND.n3791 GND.n238 3.87628
R6310 GND.n3786 GND.n241 3.87628
R6311 GND.n3547 GND 3.84833
R6312 GND.n307 GND 3.79738
R6313 GND.n3790 GND.n239 3.66653
R6314 GND.n3795 GND.n236 3.66653
R6315 GND.n3800 GND.n233 3.66653
R6316 GND.n3805 GND.n230 3.66653
R6317 GND.n3810 GND.n227 3.66653
R6318 GND.n3815 GND.n224 3.66653
R6319 GND.n3820 GND.n221 3.66653
R6320 GND.n3825 GND.n218 3.66653
R6321 GND.n3830 GND.n215 3.66653
R6322 GND.n3835 GND.n212 3.66653
R6323 GND.n3840 GND.n209 3.66653
R6324 GND.n3845 GND.n206 3.66653
R6325 GND.n3850 GND.n203 3.66653
R6326 GND.n3855 GND.n200 3.66653
R6327 GND.n3872 GND.n3871 3.66653
R6328 GND.n3867 GND.n3866 3.66653
R6329 GND.n4374 GND.n4373 3.66653
R6330 GND GND.n3876 3.65267
R6331 GND.n3526 GND.n299 3.43528
R6332 GND.n4005 GND 3.34833
R6333 GND.n402 GND 3.34833
R6334 GND.n3083 GND 3.34833
R6335 GND.n2530 GND 3.34833
R6336 GND.n1785 GND 3.34833
R6337 GND.n1528 GND 3.34833
R6338 GND.n1180 GND 3.34833
R6339 GND.n1310 GND 3.34833
R6340 GND.n1433 GND 3.34833
R6341 GND.n1057 GND 3.34833
R6342 GND.n1907 GND 3.34833
R6343 GND.n1658 GND 3.34833
R6344 GND.n2400 GND 3.34833
R6345 GND.n2653 GND 3.34833
R6346 GND.n2954 GND 3.34833
R6347 GND.n3211 GND 3.34833
R6348 GND.n4134 GND 3.34833
R6349 GND.n4256 GND 3.34833
R6350 GND.n267 GND 3.28175
R6351 GND.n3869 GND 3.21608
R6352 GND.n3483 GND 2.95702
R6353 GND.n1074 GND.n243 2.81893
R6354 GND.n4094 GND 2.79622
R6355 GND.n297 GND 2.76137
R6356 GND.n4223 GND.n4222 2.7406
R6357 GND.n4094 GND.n4093 2.7406
R6358 GND.n3173 GND.n58 2.7406
R6359 GND.n3300 GND.n3299 2.7406
R6360 GND.n3172 GND.n3171 2.7406
R6361 GND.n3043 GND.n3042 2.7406
R6362 GND.n2620 GND.n452 2.7406
R6363 GND.n2619 GND.n2618 2.7406
R6364 GND.n2489 GND.n2488 2.7406
R6365 GND.n1618 GND.n565 2.7406
R6366 GND.n1747 GND.n1746 2.7406
R6367 GND.n1874 GND.n1873 2.7406
R6368 GND.n1617 GND.n1616 2.7406
R6369 GND.n1400 GND.n894 2.7406
R6370 GND.n1399 GND.n1398 2.7406
R6371 GND.n1269 GND.n1268 2.7406
R6372 GND.n1000 GND.n937 2.7406
R6373 GND.n3620 GND.n3619 2.71789
R6374 GND.n3544 GND 2.64112
R6375 GND.n4222 GND 2.49506
R6376 GND GND.n1057 2.36463
R6377 GND.n255 GND 2.32659
R6378 GND.n3603 GND 2.32659
R6379 GND.n3584 GND 2.32659
R6380 GND.n3564 GND 2.32659
R6381 GND.n3542 GND 2.32659
R6382 GND.n3523 GND 2.32659
R6383 GND.n3501 GND 2.32659
R6384 GND.n3479 GND 2.32659
R6385 GND.t375 GND.n3629 2.09504
R6386 GND.n3680 GND.t487 2.03299
R6387 GND.n4091 GND 2.01137
R6388 GND.n3302 GND 2.01137
R6389 GND.n3169 GND 2.01137
R6390 GND.n2616 GND 2.01137
R6391 GND.n1871 GND 2.01137
R6392 GND.n1614 GND 2.01137
R6393 GND.n1266 GND 2.01137
R6394 GND.n1396 GND 2.01137
R6395 GND.n1402 GND 2.01137
R6396 GND.n1072 GND 2.01137
R6397 GND.n1876 GND 2.01137
R6398 GND.n1744 GND 2.01137
R6399 GND.n2486 GND 2.01137
R6400 GND.n2622 GND 2.01137
R6401 GND.n3040 GND 2.01137
R6402 GND.n3297 GND 2.01137
R6403 GND.n4220 GND 2.01137
R6404 GND.n3481 GND 2.0005
R6405 GND.t435 GND.n3677 1.97121
R6406 GND.t407 GND.n3675 1.97121
R6407 GND.t443 GND.n3673 1.97121
R6408 GND.t405 GND.n3671 1.97121
R6409 GND.t437 GND.n3669 1.97121
R6410 GND.t485 GND.n3667 1.97121
R6411 GND.t457 GND.n3665 1.97121
R6412 GND.t491 GND.n3663 1.97121
R6413 GND.t411 GND.n3661 1.97121
R6414 GND.t445 GND.n3659 1.97121
R6415 GND.t455 GND.n3657 1.97121
R6416 GND.t489 GND.n3655 1.97121
R6417 GND.t477 GND.n3653 1.97121
R6418 GND.t377 GND.n3651 1.97121
R6419 GND.t481 GND.n3649 1.97121
R6420 GND.t421 GND.n3647 1.97121
R6421 GND.n3735 GND.t423 1.971
R6422 GND.n3738 GND.t385 1.971
R6423 GND.n3741 GND.t431 1.971
R6424 GND.n3744 GND.t461 1.971
R6425 GND.n3747 GND.t493 1.971
R6426 GND.n3750 GND.t409 1.971
R6427 GND.n3753 GND.t373 1.971
R6428 GND.n3756 GND.t417 1.971
R6429 GND.n3759 GND.t465 1.971
R6430 GND.n3762 GND.t369 1.971
R6431 GND.n3765 GND.t371 1.971
R6432 GND.n3768 GND.t415 1.971
R6433 GND.n3771 GND.t389 1.971
R6434 GND.n3774 GND.t433 1.971
R6435 GND.n3777 GND.t401 1.971
R6436 GND.n3780 GND.t479 1.971
R6437 GND.n3733 GND.t423 1.97064
R6438 GND.n3736 GND.t385 1.97064
R6439 GND.n3739 GND.t431 1.97064
R6440 GND.n3742 GND.t461 1.97064
R6441 GND.n3745 GND.t493 1.97064
R6442 GND.n3748 GND.t409 1.97064
R6443 GND.n3751 GND.t373 1.97064
R6444 GND.n3754 GND.t417 1.97064
R6445 GND.n3757 GND.t465 1.97064
R6446 GND.n3760 GND.t369 1.97064
R6447 GND.n3763 GND.t371 1.97064
R6448 GND.n3766 GND.t415 1.97064
R6449 GND.n3769 GND.t389 1.97064
R6450 GND.n3772 GND.t433 1.97064
R6451 GND.n3775 GND.t401 1.97064
R6452 GND.n3778 GND.t479 1.97064
R6453 GND.n3684 GND.t427 1.94807
R6454 GND.n3687 GND.t497 1.94807
R6455 GND.n3690 GND.t397 1.94807
R6456 GND.n3693 GND.t495 1.94807
R6457 GND.n3696 GND.t393 1.94807
R6458 GND.n3699 GND.t499 1.94807
R6459 GND.n3702 GND.t399 1.94807
R6460 GND.n3705 GND.t451 1.94807
R6461 GND.n3708 GND.t429 1.94807
R6462 GND.n3711 GND.t463 1.94807
R6463 GND.n3714 GND.t403 1.94807
R6464 GND.n3717 GND.t483 1.94807
R6465 GND.n3720 GND.t383 1.94807
R6466 GND.n3723 GND.t419 1.94807
R6467 GND.n3726 GND.t391 1.94807
R6468 GND.n3729 GND.t469 1.94807
R6469 GND.n3648 GND.t421 1.91309
R6470 GND.n3650 GND.t481 1.91309
R6471 GND.n3652 GND.t377 1.91309
R6472 GND.n3654 GND.t477 1.91309
R6473 GND.n3656 GND.t489 1.91309
R6474 GND.n3658 GND.t455 1.91309
R6475 GND.n3660 GND.t445 1.91309
R6476 GND.n3662 GND.t411 1.91309
R6477 GND.n3664 GND.t491 1.91309
R6478 GND.n3666 GND.t457 1.91309
R6479 GND.n3668 GND.t485 1.91309
R6480 GND.n3670 GND.t437 1.91309
R6481 GND.n3672 GND.t405 1.91309
R6482 GND.n3674 GND.t443 1.91309
R6483 GND.n3676 GND.t407 1.91309
R6484 GND.n3678 GND.t435 1.91309
R6485 GND.n3682 GND.t427 1.883
R6486 GND.n3685 GND.t497 1.883
R6487 GND.n3688 GND.t397 1.883
R6488 GND.n3691 GND.t495 1.883
R6489 GND.n3694 GND.t393 1.883
R6490 GND.n3697 GND.t499 1.883
R6491 GND.n3700 GND.t399 1.883
R6492 GND.n3703 GND.t451 1.883
R6493 GND.n3706 GND.t429 1.883
R6494 GND.n3709 GND.t463 1.883
R6495 GND.n3712 GND.t403 1.883
R6496 GND.n3715 GND.t483 1.883
R6497 GND.n3718 GND.t383 1.883
R6498 GND.n3721 GND.t419 1.883
R6499 GND.n3724 GND.t391 1.883
R6500 GND.n3727 GND.t469 1.883
R6501 GND.n273 GND 1.87007
R6502 GND.n3955 GND 1.83746
R6503 GND.n3382 GND 1.83746
R6504 GND.n2897 GND 1.83746
R6505 GND.n2827 GND 1.83746
R6506 GND.n2255 GND 1.83746
R6507 GND GND.n670 1.83746
R6508 GND GND.n2065 1.83746
R6509 GND.n3567 GND.n283 1.82659
R6510 GND.n4089 GND 1.67985
R6511 GND.n4075 GND 1.67985
R6512 GND.n3304 GND 1.67985
R6513 GND.n392 GND 1.67985
R6514 GND.n3167 GND 1.67985
R6515 GND.n3153 GND 1.67985
R6516 GND.n2614 GND 1.67985
R6517 GND.n2600 GND 1.67985
R6518 GND.n1869 GND 1.67985
R6519 GND.n1855 GND 1.67985
R6520 GND.n1612 GND 1.67985
R6521 GND.n1598 GND 1.67985
R6522 GND.n1264 GND 1.67985
R6523 GND.n1250 GND 1.67985
R6524 GND.n1394 GND 1.67985
R6525 GND.n1380 GND 1.67985
R6526 GND.n1404 GND 1.67985
R6527 GND.n1500 GND 1.67985
R6528 GND.n1070 GND 1.67985
R6529 GND.n1878 GND 1.67985
R6530 GND.n1974 GND 1.67985
R6531 GND.n1742 GND 1.67985
R6532 GND.n1728 GND 1.67985
R6533 GND.n2484 GND 1.67985
R6534 GND.n2470 GND 1.67985
R6535 GND.n2624 GND 1.67985
R6536 GND.n2720 GND 1.67985
R6537 GND.n3038 GND 1.67985
R6538 GND.n3024 GND 1.67985
R6539 GND.n3295 GND 1.67985
R6540 GND.n3281 GND 1.67985
R6541 GND.n4218 GND 1.67985
R6542 GND.n4204 GND 1.67985
R6543 GND.n4247 GND 1.67985
R6544 GND.n4055 GND.n4054 1.66898
R6545 GND.n4060 GND.n4055 1.66898
R6546 GND.n4057 GND.n77 1.66898
R6547 GND.n4076 GND.n77 1.66898
R6548 GND.n4038 GND.n4017 1.66898
R6549 GND.n4035 GND.n4018 1.66898
R6550 GND.n4030 GND.n4018 1.66898
R6551 GND.n3313 GND.n367 1.66898
R6552 GND.n3326 GND.n367 1.66898
R6553 GND.n3323 GND.n368 1.66898
R6554 GND.n391 GND.n368 1.66898
R6555 GND.n425 GND.n404 1.66898
R6556 GND.n429 GND.n428 1.66898
R6557 GND.n430 GND.n429 1.66898
R6558 GND.n3133 GND.n3132 1.66898
R6559 GND.n3138 GND.n3133 1.66898
R6560 GND.n3135 GND.n3062 1.66898
R6561 GND.n3154 GND.n3062 1.66898
R6562 GND.n3116 GND.n3095 1.66898
R6563 GND.n3113 GND.n3096 1.66898
R6564 GND.n3108 GND.n3096 1.66898
R6565 GND.n2580 GND.n2579 1.66898
R6566 GND.n2585 GND.n2580 1.66898
R6567 GND.n2582 GND.n2508 1.66898
R6568 GND.n2601 GND.n2508 1.66898
R6569 GND.n2563 GND.n2542 1.66898
R6570 GND.n2560 GND.n2543 1.66898
R6571 GND.n2555 GND.n2543 1.66898
R6572 GND.n1835 GND.n1834 1.66898
R6573 GND.n1840 GND.n1835 1.66898
R6574 GND.n1837 GND.n1765 1.66898
R6575 GND.n1856 GND.n1765 1.66898
R6576 GND.n1818 GND.n1797 1.66898
R6577 GND.n1815 GND.n1798 1.66898
R6578 GND.n1810 GND.n1798 1.66898
R6579 GND.n1578 GND.n1577 1.66898
R6580 GND.n1583 GND.n1578 1.66898
R6581 GND.n1580 GND.n913 1.66898
R6582 GND.n1599 GND.n913 1.66898
R6583 GND.n1561 GND.n1540 1.66898
R6584 GND.n1558 GND.n1541 1.66898
R6585 GND.n1553 GND.n1541 1.66898
R6586 GND.n1230 GND.n1229 1.66898
R6587 GND.n1235 GND.n1230 1.66898
R6588 GND.n1232 GND.n956 1.66898
R6589 GND.n1251 GND.n956 1.66898
R6590 GND.n1213 GND.n1192 1.66898
R6591 GND.n1210 GND.n1193 1.66898
R6592 GND.n1205 GND.n1193 1.66898
R6593 GND.n1360 GND.n1359 1.66898
R6594 GND.n1365 GND.n1360 1.66898
R6595 GND.n1362 GND.n1288 1.66898
R6596 GND.n1381 GND.n1288 1.66898
R6597 GND.n1343 GND.n1322 1.66898
R6598 GND.n1340 GND.n1323 1.66898
R6599 GND.n1335 GND.n1323 1.66898
R6600 GND.n1512 GND.n1406 1.66898
R6601 GND.n1508 GND.n1406 1.66898
R6602 GND.n1505 GND.n1410 1.66898
R6603 GND.n1501 GND.n1410 1.66898
R6604 GND.n1483 GND.n1435 1.66898
R6605 GND.n1480 GND.n1436 1.66898
R6606 GND.n1475 GND.n1436 1.66898
R6607 GND.n1021 GND.n1016 1.66898
R6608 GND.n1028 GND.n1016 1.66898
R6609 GND.n1032 GND.n1031 1.66898
R6610 GND.n1058 GND.n1032 1.66898
R6611 GND.n1055 GND.n1046 1.66898
R6612 GND.n1043 GND.n1033 1.66898
R6613 GND.n1038 GND.n1033 1.66898
R6614 GND.n3954 GND.n183 1.66898
R6615 GND.n3900 GND.n183 1.66898
R6616 GND.n3942 GND.n3941 1.66898
R6617 GND.n3930 GND.n3908 1.66898
R6618 GND.n3916 GND.n3908 1.66898
R6619 GND.n3918 GND.n5 1.66898
R6620 GND.n4367 GND.n5 1.66898
R6621 GND.n3433 GND.n3432 1.66898
R6622 GND.n3432 GND.n3431 1.66898
R6623 GND.n3422 GND.n3421 1.66898
R6624 GND.n3410 GND.n3394 1.66898
R6625 GND.n3397 GND.n3394 1.66898
R6626 GND.n3888 GND.n3887 1.66898
R6627 GND.n3890 GND.n3888 1.66898
R6628 GND.n2896 GND.n492 1.66898
R6629 GND.n495 GND.n492 1.66898
R6630 GND.n3466 GND.n313 1.66898
R6631 GND.n3455 GND.n3454 1.66898
R6632 GND.n3454 GND.n3453 1.66898
R6633 GND.n3444 GND.n3443 1.66898
R6634 GND.n3443 GND.n3442 1.66898
R6635 GND.n2833 GND.n2832 1.66898
R6636 GND.n2835 GND.n2833 1.66898
R6637 GND.n2851 GND.n511 1.66898
R6638 GND.n2864 GND.n2863 1.66898
R6639 GND.n2866 GND.n2864 1.66898
R6640 GND.n2876 GND.n2875 1.66898
R6641 GND.n2878 GND.n2876 1.66898
R6642 GND.n2254 GND.n646 1.66898
R6643 GND.n2189 GND.n646 1.66898
R6644 GND.n2242 GND.n2241 1.66898
R6645 GND.n2230 GND.n2197 1.66898
R6646 GND.n2209 GND.n2197 1.66898
R6647 GND.n2218 GND.n2217 1.66898
R6648 GND.n2217 GND.n2216 1.66898
R6649 GND.n766 GND.n725 1.66898
R6650 GND.n734 GND.n725 1.66898
R6651 GND.n754 GND.n753 1.66898
R6652 GND.n2108 GND.n2107 1.66898
R6653 GND.n2110 GND.n2108 1.66898
R6654 GND.n2120 GND.n2119 1.66898
R6655 GND.n2122 GND.n2120 1.66898
R6656 GND.n2132 GND.n2131 1.66898
R6657 GND.n2134 GND.n2132 1.66898
R6658 GND.n2150 GND.n661 1.66898
R6659 GND.n2163 GND.n2162 1.66898
R6660 GND.n2165 GND.n2163 1.66898
R6661 GND.n2175 GND.n2174 1.66898
R6662 GND.n2177 GND.n2175 1.66898
R6663 GND.n689 GND.n688 1.66898
R6664 GND.n2094 GND.n689 1.66898
R6665 GND.n2092 GND.n690 1.66898
R6666 GND.n2077 GND.n702 1.66898
R6667 GND.n2073 GND.n702 1.66898
R6668 GND.n2071 GND.n706 1.66898
R6669 GND.n2067 GND.n706 1.66898
R6670 GND.n1986 GND.n1880 1.66898
R6671 GND.n1982 GND.n1880 1.66898
R6672 GND.n1979 GND.n1884 1.66898
R6673 GND.n1975 GND.n1884 1.66898
R6674 GND.n1957 GND.n1909 1.66898
R6675 GND.n1954 GND.n1910 1.66898
R6676 GND.n1949 GND.n1910 1.66898
R6677 GND.n1708 GND.n1707 1.66898
R6678 GND.n1713 GND.n1708 1.66898
R6679 GND.n1710 GND.n1637 1.66898
R6680 GND.n1729 GND.n1637 1.66898
R6681 GND.n1691 GND.n1670 1.66898
R6682 GND.n1688 GND.n1671 1.66898
R6683 GND.n1683 GND.n1671 1.66898
R6684 GND.n2450 GND.n2449 1.66898
R6685 GND.n2455 GND.n2450 1.66898
R6686 GND.n2452 GND.n584 1.66898
R6687 GND.n2471 GND.n584 1.66898
R6688 GND.n2433 GND.n2412 1.66898
R6689 GND.n2430 GND.n2413 1.66898
R6690 GND.n2425 GND.n2413 1.66898
R6691 GND.n2732 GND.n2626 1.66898
R6692 GND.n2728 GND.n2626 1.66898
R6693 GND.n2725 GND.n2630 1.66898
R6694 GND.n2721 GND.n2630 1.66898
R6695 GND.n2703 GND.n2655 1.66898
R6696 GND.n2700 GND.n2656 1.66898
R6697 GND.n2695 GND.n2656 1.66898
R6698 GND.n3004 GND.n3003 1.66898
R6699 GND.n3009 GND.n3004 1.66898
R6700 GND.n3006 GND.n471 1.66898
R6701 GND.n3025 GND.n471 1.66898
R6702 GND.n2987 GND.n2966 1.66898
R6703 GND.n2984 GND.n2967 1.66898
R6704 GND.n2979 GND.n2967 1.66898
R6705 GND.n3261 GND.n3260 1.66898
R6706 GND.n3266 GND.n3261 1.66898
R6707 GND.n3263 GND.n3191 1.66898
R6708 GND.n3282 GND.n3191 1.66898
R6709 GND.n3244 GND.n3223 1.66898
R6710 GND.n3241 GND.n3224 1.66898
R6711 GND.n3236 GND.n3224 1.66898
R6712 GND.n4184 GND.n4183 1.66898
R6713 GND.n4189 GND.n4184 1.66898
R6714 GND.n4186 GND.n4113 1.66898
R6715 GND.n4205 GND.n4113 1.66898
R6716 GND.n4167 GND.n4146 1.66898
R6717 GND.n4164 GND.n4147 1.66898
R6718 GND.n4159 GND.n4147 1.66898
R6719 GND.n4272 GND.n4270 1.66898
R6720 GND.n4272 GND.n4271 1.66898
R6721 GND.n4267 GND.n4258 1.66898
R6722 GND.n4279 GND.n4229 1.66898
R6723 GND.n4246 GND.n4229 1.66898
R6724 GND.n4228 GND.n4227 1.66898
R6725 GND.n4282 GND.n4228 1.66898
R6726 GND.t666 GND.n982 1.62053
R6727 GND.n4087 GND.n4086 1.5505
R6728 GND.n4061 GND.n4060 1.5505
R6729 GND.n4055 GND.n4051 1.5505
R6730 GND.n4054 GND.n4048 1.5505
R6731 GND.n4077 GND.n4076 1.5505
R6732 GND.n77 GND.n76 1.5505
R6733 GND.n4057 GND.n4056 1.5505
R6734 GND.n4073 GND.n4072 1.5505
R6735 GND.n4039 GND.n4038 1.5505
R6736 GND.n4017 GND.n4016 1.5505
R6737 GND.n4035 GND.n4034 1.5505
R6738 GND.n4031 GND.n4030 1.5505
R6739 GND.n4033 GND.n4018 1.5505
R6740 GND.n3317 GND.n3316 1.5505
R6741 GND.n3327 GND.n3326 1.5505
R6742 GND.n367 GND.n366 1.5505
R6743 GND.n3313 GND.n3312 1.5505
R6744 GND.n391 GND.n371 1.5505
R6745 GND.n3321 GND.n368 1.5505
R6746 GND.n3323 GND.n3322 1.5505
R6747 GND.n401 GND.n400 1.5505
R6748 GND.n425 GND.n424 1.5505
R6749 GND.n417 GND.n404 1.5505
R6750 GND.n428 GND.n390 1.5505
R6751 GND.n431 GND.n430 1.5505
R6752 GND.n444 GND.n429 1.5505
R6753 GND.n3165 GND.n3164 1.5505
R6754 GND.n3139 GND.n3138 1.5505
R6755 GND.n3133 GND.n3129 1.5505
R6756 GND.n3132 GND.n3126 1.5505
R6757 GND.n3155 GND.n3154 1.5505
R6758 GND.n3062 GND.n3061 1.5505
R6759 GND.n3135 GND.n3134 1.5505
R6760 GND.n3151 GND.n3150 1.5505
R6761 GND.n3117 GND.n3116 1.5505
R6762 GND.n3095 GND.n3094 1.5505
R6763 GND.n3113 GND.n3112 1.5505
R6764 GND.n3109 GND.n3108 1.5505
R6765 GND.n3111 GND.n3096 1.5505
R6766 GND.n2612 GND.n2611 1.5505
R6767 GND.n2586 GND.n2585 1.5505
R6768 GND.n2580 GND.n2576 1.5505
R6769 GND.n2579 GND.n2573 1.5505
R6770 GND.n2602 GND.n2601 1.5505
R6771 GND.n2508 GND.n2507 1.5505
R6772 GND.n2582 GND.n2581 1.5505
R6773 GND.n2598 GND.n2597 1.5505
R6774 GND.n2564 GND.n2563 1.5505
R6775 GND.n2542 GND.n2541 1.5505
R6776 GND.n2560 GND.n2559 1.5505
R6777 GND.n2556 GND.n2555 1.5505
R6778 GND.n2558 GND.n2543 1.5505
R6779 GND.n1867 GND.n1866 1.5505
R6780 GND.n1841 GND.n1840 1.5505
R6781 GND.n1835 GND.n1831 1.5505
R6782 GND.n1834 GND.n1828 1.5505
R6783 GND.n1857 GND.n1856 1.5505
R6784 GND.n1765 GND.n1764 1.5505
R6785 GND.n1837 GND.n1836 1.5505
R6786 GND.n1853 GND.n1852 1.5505
R6787 GND.n1819 GND.n1818 1.5505
R6788 GND.n1797 GND.n1796 1.5505
R6789 GND.n1815 GND.n1814 1.5505
R6790 GND.n1811 GND.n1810 1.5505
R6791 GND.n1813 GND.n1798 1.5505
R6792 GND.n1610 GND.n1609 1.5505
R6793 GND.n1584 GND.n1583 1.5505
R6794 GND.n1578 GND.n1574 1.5505
R6795 GND.n1577 GND.n1571 1.5505
R6796 GND.n1600 GND.n1599 1.5505
R6797 GND.n913 GND.n912 1.5505
R6798 GND.n1580 GND.n1579 1.5505
R6799 GND.n1596 GND.n1595 1.5505
R6800 GND.n1562 GND.n1561 1.5505
R6801 GND.n1540 GND.n1539 1.5505
R6802 GND.n1558 GND.n1557 1.5505
R6803 GND.n1554 GND.n1553 1.5505
R6804 GND.n1556 GND.n1541 1.5505
R6805 GND.n1262 GND.n1261 1.5505
R6806 GND.n1236 GND.n1235 1.5505
R6807 GND.n1230 GND.n1226 1.5505
R6808 GND.n1229 GND.n1223 1.5505
R6809 GND.n1252 GND.n1251 1.5505
R6810 GND.n956 GND.n955 1.5505
R6811 GND.n1232 GND.n1231 1.5505
R6812 GND.n1248 GND.n1247 1.5505
R6813 GND.n1214 GND.n1213 1.5505
R6814 GND.n1192 GND.n1191 1.5505
R6815 GND.n1210 GND.n1209 1.5505
R6816 GND.n1206 GND.n1205 1.5505
R6817 GND.n1208 GND.n1193 1.5505
R6818 GND.n1392 GND.n1391 1.5505
R6819 GND.n1366 GND.n1365 1.5505
R6820 GND.n1360 GND.n1356 1.5505
R6821 GND.n1359 GND.n1353 1.5505
R6822 GND.n1382 GND.n1381 1.5505
R6823 GND.n1288 GND.n1287 1.5505
R6824 GND.n1362 GND.n1361 1.5505
R6825 GND.n1378 GND.n1377 1.5505
R6826 GND.n1344 GND.n1343 1.5505
R6827 GND.n1322 GND.n1321 1.5505
R6828 GND.n1340 GND.n1339 1.5505
R6829 GND.n1336 GND.n1335 1.5505
R6830 GND.n1338 GND.n1323 1.5505
R6831 GND.n1516 GND.n1515 1.5505
R6832 GND.n1509 GND.n1508 1.5505
R6833 GND.n1510 GND.n1406 1.5505
R6834 GND.n1512 GND.n1511 1.5505
R6835 GND.n1502 GND.n1501 1.5505
R6836 GND.n1503 GND.n1410 1.5505
R6837 GND.n1505 GND.n1504 1.5505
R6838 GND.n1498 GND.n1497 1.5505
R6839 GND.n1484 GND.n1483 1.5505
R6840 GND.n1453 GND.n1435 1.5505
R6841 GND.n1480 GND.n1479 1.5505
R6842 GND.n1476 GND.n1475 1.5505
R6843 GND.n1478 GND.n1436 1.5505
R6844 GND.n1068 GND.n1067 1.5505
R6845 GND.n1028 GND.n1027 1.5505
R6846 GND.n1018 GND.n1016 1.5505
R6847 GND.n1022 GND.n1021 1.5505
R6848 GND.n1059 GND.n1058 1.5505
R6849 GND.n1032 GND.n1015 1.5505
R6850 GND.n1031 GND.n1014 1.5505
R6851 GND.n1051 GND.n1046 1.5505
R6852 GND.n1055 GND.n1054 1.5505
R6853 GND.n1043 GND.n1042 1.5505
R6854 GND.n1041 GND.n1033 1.5505
R6855 GND.n1039 GND.n1038 1.5505
R6856 GND.n3619 GND.n3618 1.5505
R6857 GND.n3617 GND.n246 1.5505
R6858 GND.n261 GND.n247 1.5505
R6859 GND.n3607 GND.n3606 1.5505
R6860 GND.n3604 GND.n254 1.5505
R6861 GND.n3597 GND.n3596 1.5505
R6862 GND.n3588 GND.n3587 1.5505
R6863 GND.n3585 GND.n272 1.5505
R6864 GND.n3577 GND.n3576 1.5505
R6865 GND.n3568 GND.n3567 1.5505
R6866 GND.n3565 GND.n280 1.5505
R6867 GND.n3558 GND.n3557 1.5505
R6868 GND.n3549 GND.n3548 1.5505
R6869 GND.n3543 GND.n288 1.5505
R6870 GND.n3536 GND.n3535 1.5505
R6871 GND.n3527 GND.n3526 1.5505
R6872 GND.n3524 GND.n296 1.5505
R6873 GND.n3514 GND.n3513 1.5505
R6874 GND.n3505 GND.n3504 1.5505
R6875 GND.n3502 GND.n304 1.5505
R6876 GND.n3495 GND.n3494 1.5505
R6877 GND.n3486 GND.n3485 1.5505
R6878 GND.n3480 GND.n196 1.5505
R6879 GND.n3878 GND.n3877 1.5505
R6880 GND.n3954 GND.n3953 1.5505
R6881 GND.n3952 GND.n183 1.5505
R6882 GND.n3900 GND.n185 1.5505
R6883 GND.n3943 GND.n3942 1.5505
R6884 GND.n3941 GND.n3940 1.5505
R6885 GND.n3933 GND.n3932 1.5505
R6886 GND.n3930 GND.n3929 1.5505
R6887 GND.n3928 GND.n3908 1.5505
R6888 GND.n3916 GND.n3910 1.5505
R6889 GND.n3919 GND.n3918 1.5505
R6890 GND.n6 GND.n5 1.5505
R6891 GND.n4367 GND.n4366 1.5505
R6892 GND.n3434 GND.n3433 1.5505
R6893 GND.n3432 GND.n333 1.5505
R6894 GND.n3431 GND.n3430 1.5505
R6895 GND.n3423 GND.n3422 1.5505
R6896 GND.n3421 GND.n3420 1.5505
R6897 GND.n3413 GND.n3412 1.5505
R6898 GND.n3410 GND.n3409 1.5505
R6899 GND.n3408 GND.n3394 1.5505
R6900 GND.n3398 GND.n3397 1.5505
R6901 GND.n3887 GND.n3886 1.5505
R6902 GND.n3888 GND.n191 1.5505
R6903 GND.n3891 GND.n3890 1.5505
R6904 GND.n2896 GND.n2895 1.5505
R6905 GND.n2894 GND.n492 1.5505
R6906 GND.n496 GND.n495 1.5505
R6907 GND.n2885 GND.n313 1.5505
R6908 GND.n3467 GND.n3466 1.5505
R6909 GND.n3464 GND.n3463 1.5505
R6910 GND.n3456 GND.n3455 1.5505
R6911 GND.n3454 GND.n323 1.5505
R6912 GND.n3453 GND.n3452 1.5505
R6913 GND.n3445 GND.n3444 1.5505
R6914 GND.n3443 GND.n328 1.5505
R6915 GND.n3442 GND.n3441 1.5505
R6916 GND.n2832 GND.n2831 1.5505
R6917 GND.n2833 GND.n519 1.5505
R6918 GND.n2836 GND.n2835 1.5505
R6919 GND.n2840 GND.n511 1.5505
R6920 GND.n2851 GND.n2850 1.5505
R6921 GND.n2855 GND.n2854 1.5505
R6922 GND.n2863 GND.n2862 1.5505
R6923 GND.n2864 GND.n506 1.5505
R6924 GND.n2867 GND.n2866 1.5505
R6925 GND.n2875 GND.n2874 1.5505
R6926 GND.n2876 GND.n502 1.5505
R6927 GND.n2879 GND.n2878 1.5505
R6928 GND.n2254 GND.n2253 1.5505
R6929 GND.n2252 GND.n646 1.5505
R6930 GND.n2189 GND.n648 1.5505
R6931 GND.n2243 GND.n2242 1.5505
R6932 GND.n2241 GND.n2240 1.5505
R6933 GND.n2233 GND.n2232 1.5505
R6934 GND.n2230 GND.n2229 1.5505
R6935 GND.n2228 GND.n2197 1.5505
R6936 GND.n2209 GND.n2199 1.5505
R6937 GND.n2219 GND.n2218 1.5505
R6938 GND.n2217 GND.n2208 1.5505
R6939 GND.n2216 GND.n2215 1.5505
R6940 GND.n766 GND.n765 1.5505
R6941 GND.n764 GND.n725 1.5505
R6942 GND.n734 GND.n727 1.5505
R6943 GND.n755 GND.n754 1.5505
R6944 GND.n753 GND.n752 1.5505
R6945 GND.n745 GND.n744 1.5505
R6946 GND.n2107 GND.n2106 1.5505
R6947 GND.n2108 GND.n678 1.5505
R6948 GND.n2111 GND.n2110 1.5505
R6949 GND.n2119 GND.n2118 1.5505
R6950 GND.n2120 GND.n674 1.5505
R6951 GND.n2123 GND.n2122 1.5505
R6952 GND.n2131 GND.n2130 1.5505
R6953 GND.n2132 GND.n669 1.5505
R6954 GND.n2135 GND.n2134 1.5505
R6955 GND.n2154 GND.n2153 1.5505
R6956 GND.n2162 GND.n2161 1.5505
R6957 GND.n2163 GND.n656 1.5505
R6958 GND.n2166 GND.n2165 1.5505
R6959 GND.n2174 GND.n2173 1.5505
R6960 GND.n2175 GND.n652 1.5505
R6961 GND.n2178 GND.n2177 1.5505
R6962 GND.n2139 GND.n661 1.5505
R6963 GND.n2150 GND.n2149 1.5505
R6964 GND.n688 GND.n687 1.5505
R6965 GND.n689 GND.n686 1.5505
R6966 GND.n2095 GND.n2094 1.5505
R6967 GND.n2092 GND.n2091 1.5505
R6968 GND.n692 GND.n690 1.5505
R6969 GND.n2080 GND.n2079 1.5505
R6970 GND.n2077 GND.n2076 1.5505
R6971 GND.n2075 GND.n702 1.5505
R6972 GND.n2074 GND.n2073 1.5505
R6973 GND.n2071 GND.n2070 1.5505
R6974 GND.n2069 GND.n706 1.5505
R6975 GND.n2068 GND.n2067 1.5505
R6976 GND.n1085 GND.n1084 1.5505
R6977 GND.n1083 GND.n999 1.5505
R6978 GND.n1082 GND.n998 1.5505
R6979 GND.n1080 GND.n995 1.5505
R6980 GND.n1075 GND.n993 1.5505
R6981 GND.n1109 GND.n1108 1.5505
R6982 GND.n977 GND.n976 1.5505
R6983 GND.n1119 GND.n1118 1.5505
R6984 GND.n1123 GND.n1121 1.5505
R6985 GND.n1165 GND.n1164 1.5505
R6986 GND.n1133 GND.n1124 1.5505
R6987 GND.n1150 GND.n1149 1.5505
R6988 GND.n2063 GND.n2062 1.5505
R6989 GND.n2061 GND.n768 1.5505
R6990 GND.n787 GND.n770 1.5505
R6991 GND.n789 GND.n777 1.5505
R6992 GND.n795 GND.n779 1.5505
R6993 GND.n2043 GND.n2042 1.5505
R6994 GND.n2041 GND.n797 1.5505
R6995 GND.n840 GND.n799 1.5505
R6996 GND.n842 GND.n806 1.5505
R6997 GND.n847 GND.n846 1.5505
R6998 GND.n843 GND.n807 1.5505
R6999 GND.n862 GND.n812 1.5505
R7000 GND.n865 GND.n815 1.5505
R7001 GND.n867 GND.n866 1.5505
R7002 GND.n868 GND.n816 1.5505
R7003 GND.n870 GND.n820 1.5505
R7004 GND.n876 GND.n822 1.5505
R7005 GND.n2002 GND.n2001 1.5505
R7006 GND.n2000 GND.n878 1.5505
R7007 GND.n882 GND.n881 1.5505
R7008 GND.n631 GND.n629 1.5505
R7009 GND.n2288 GND.n2287 1.5505
R7010 GND.n641 GND.n632 1.5505
R7011 GND.n2273 GND.n2272 1.5505
R7012 GND.n645 GND.n644 1.5505
R7013 GND.n618 GND.n617 1.5505
R7014 GND.n2302 GND.n2301 1.5505
R7015 GND.n2304 GND.n613 1.5505
R7016 GND.n2306 GND.n611 1.5505
R7017 GND.n2325 GND.n603 1.5505
R7018 GND.n2390 GND.n2326 1.5505
R7019 GND.n2389 GND.n2388 1.5505
R7020 GND.n2386 GND.n2385 1.5505
R7021 GND.n2384 GND.n2333 1.5505
R7022 GND.n2374 GND.n2334 1.5505
R7023 GND.n2366 GND.n2365 1.5505
R7024 GND.n2825 GND.n2824 1.5505
R7025 GND.n2823 GND.n521 1.5505
R7026 GND.n540 GND.n523 1.5505
R7027 GND.n542 GND.n530 1.5505
R7028 GND.n548 GND.n532 1.5505
R7029 GND.n2805 GND.n2804 1.5505
R7030 GND.n2803 GND.n550 1.5505
R7031 GND.n2758 GND.n552 1.5505
R7032 GND.n2760 GND.n2741 1.5505
R7033 GND.n2765 GND.n2764 1.5505
R7034 GND.n2761 GND.n2742 1.5505
R7035 GND.n2781 GND.n2780 1.5505
R7036 GND.n2899 GND.n490 1.5505
R7037 GND.n2944 GND.n2900 1.5505
R7038 GND.n2943 GND.n2942 1.5505
R7039 GND.n2940 GND.n2939 1.5505
R7040 GND.n2923 GND.n2906 1.5505
R7041 GND.n2929 GND.n355 1.5505
R7042 GND.n2928 GND.n2927 1.5505
R7043 GND.n2926 GND.n354 1.5505
R7044 GND.n3347 GND.n3346 1.5505
R7045 GND.n3348 GND.n344 1.5505
R7046 GND.n3364 GND.n3363 1.5505
R7047 GND.n3378 GND.n3377 1.5505
R7048 GND.n3380 GND.n98 1.5505
R7049 GND.n3993 GND.n99 1.5505
R7050 GND.n3992 GND.n3991 1.5505
R7051 GND.n3989 GND.n3988 1.5505
R7052 GND.n121 GND.n105 1.5505
R7053 GND.n3978 GND.n3977 1.5505
R7054 GND.n3976 GND.n123 1.5505
R7055 GND.n152 GND.n125 1.5505
R7056 GND.n154 GND.n136 1.5505
R7057 GND.n159 GND.n158 1.5505
R7058 GND.n155 GND.n137 1.5505
R7059 GND.n3959 GND.n3958 1.5505
R7060 GND.n182 GND.n47 1.5505
R7061 GND.n181 GND.n180 1.5505
R7062 GND.n179 GND.n46 1.5505
R7063 GND.n177 GND.n176 1.5505
R7064 GND.n4304 GND.n4303 1.5505
R7065 GND.n4310 GND.n30 1.5505
R7066 GND.n4309 GND.n4308 1.5505
R7067 GND.n4307 GND.n29 1.5505
R7068 GND.n4348 GND.n13 1.5505
R7069 GND.n1078 GND.n1077 1.5505
R7070 GND.n1107 GND.n1106 1.5505
R7071 GND.n1168 GND.n1167 1.5505
R7072 GND.n1155 GND.n1122 1.5505
R7073 GND.n1153 GND.n1152 1.5505
R7074 GND.n794 GND.n793 1.5505
R7075 GND.n2045 GND.n2044 1.5505
R7076 GND.n850 GND.n849 1.5505
R7077 GND.n845 GND.n844 1.5505
R7078 GND.n860 GND.n859 1.5505
R7079 GND.n875 GND.n874 1.5505
R7080 GND.n2004 GND.n2003 1.5505
R7081 GND.n2291 GND.n2290 1.5505
R7082 GND.n2278 GND.n630 1.5505
R7083 GND.n2276 GND.n2275 1.5505
R7084 GND.n2308 GND.n2307 1.5505
R7085 GND.n2324 GND.n2323 1.5505
R7086 GND.n2345 GND.n2330 1.5505
R7087 GND.n2376 GND.n2375 1.5505
R7088 GND.n2372 GND.n2371 1.5505
R7089 GND.n547 GND.n546 1.5505
R7090 GND.n2807 GND.n2806 1.5505
R7091 GND.n2768 GND.n2767 1.5505
R7092 GND.n2763 GND.n2762 1.5505
R7093 GND.n2778 GND.n2777 1.5505
R7094 GND.n2922 GND.n2921 1.5505
R7095 GND.n2931 GND.n2930 1.5505
R7096 GND.n3351 GND.n3350 1.5505
R7097 GND.n3355 GND.n343 1.5505
R7098 GND.n3368 GND.n3367 1.5505
R7099 GND.n120 GND.n119 1.5505
R7100 GND.n3980 GND.n3979 1.5505
R7101 GND.n162 GND.n161 1.5505
R7102 GND.n157 GND.n156 1.5505
R7103 GND.n172 GND.n171 1.5505
R7104 GND.n41 GND.n36 1.5505
R7105 GND.n4312 GND.n4311 1.5505
R7106 GND.n4333 GND.n4332 1.5505
R7107 GND.n4337 GND.n18 1.5505
R7108 GND.n4351 GND.n4350 1.5505
R7109 GND.n4346 GND.n4345 1.5505
R7110 GND.n4330 GND.n19 1.5505
R7111 GND.n4329 GND.n4328 1.5505
R7112 GND.n1990 GND.n1989 1.5505
R7113 GND.n1983 GND.n1982 1.5505
R7114 GND.n1984 GND.n1880 1.5505
R7115 GND.n1986 GND.n1985 1.5505
R7116 GND.n1976 GND.n1975 1.5505
R7117 GND.n1977 GND.n1884 1.5505
R7118 GND.n1979 GND.n1978 1.5505
R7119 GND.n1972 GND.n1971 1.5505
R7120 GND.n1958 GND.n1957 1.5505
R7121 GND.n1927 GND.n1909 1.5505
R7122 GND.n1954 GND.n1953 1.5505
R7123 GND.n1950 GND.n1949 1.5505
R7124 GND.n1952 GND.n1910 1.5505
R7125 GND.n1740 GND.n1739 1.5505
R7126 GND.n1714 GND.n1713 1.5505
R7127 GND.n1708 GND.n1704 1.5505
R7128 GND.n1707 GND.n1701 1.5505
R7129 GND.n1730 GND.n1729 1.5505
R7130 GND.n1637 GND.n1636 1.5505
R7131 GND.n1710 GND.n1709 1.5505
R7132 GND.n1726 GND.n1725 1.5505
R7133 GND.n1692 GND.n1691 1.5505
R7134 GND.n1670 GND.n1669 1.5505
R7135 GND.n1688 GND.n1687 1.5505
R7136 GND.n1684 GND.n1683 1.5505
R7137 GND.n1686 GND.n1671 1.5505
R7138 GND.n2482 GND.n2481 1.5505
R7139 GND.n2456 GND.n2455 1.5505
R7140 GND.n2450 GND.n2446 1.5505
R7141 GND.n2449 GND.n2443 1.5505
R7142 GND.n2472 GND.n2471 1.5505
R7143 GND.n584 GND.n583 1.5505
R7144 GND.n2452 GND.n2451 1.5505
R7145 GND.n2468 GND.n2467 1.5505
R7146 GND.n2434 GND.n2433 1.5505
R7147 GND.n2412 GND.n2411 1.5505
R7148 GND.n2430 GND.n2429 1.5505
R7149 GND.n2426 GND.n2425 1.5505
R7150 GND.n2428 GND.n2413 1.5505
R7151 GND.n2736 GND.n2735 1.5505
R7152 GND.n2729 GND.n2728 1.5505
R7153 GND.n2730 GND.n2626 1.5505
R7154 GND.n2732 GND.n2731 1.5505
R7155 GND.n2722 GND.n2721 1.5505
R7156 GND.n2723 GND.n2630 1.5505
R7157 GND.n2725 GND.n2724 1.5505
R7158 GND.n2718 GND.n2717 1.5505
R7159 GND.n2704 GND.n2703 1.5505
R7160 GND.n2673 GND.n2655 1.5505
R7161 GND.n2700 GND.n2699 1.5505
R7162 GND.n2696 GND.n2695 1.5505
R7163 GND.n2698 GND.n2656 1.5505
R7164 GND.n3036 GND.n3035 1.5505
R7165 GND.n3010 GND.n3009 1.5505
R7166 GND.n3004 GND.n3000 1.5505
R7167 GND.n3003 GND.n2997 1.5505
R7168 GND.n3026 GND.n3025 1.5505
R7169 GND.n471 GND.n470 1.5505
R7170 GND.n3006 GND.n3005 1.5505
R7171 GND.n3022 GND.n3021 1.5505
R7172 GND.n2988 GND.n2987 1.5505
R7173 GND.n2966 GND.n2965 1.5505
R7174 GND.n2984 GND.n2983 1.5505
R7175 GND.n2980 GND.n2979 1.5505
R7176 GND.n2982 GND.n2967 1.5505
R7177 GND.n3293 GND.n3292 1.5505
R7178 GND.n3267 GND.n3266 1.5505
R7179 GND.n3261 GND.n3257 1.5505
R7180 GND.n3260 GND.n3254 1.5505
R7181 GND.n3283 GND.n3282 1.5505
R7182 GND.n3191 GND.n3190 1.5505
R7183 GND.n3263 GND.n3262 1.5505
R7184 GND.n3279 GND.n3278 1.5505
R7185 GND.n3245 GND.n3244 1.5505
R7186 GND.n3223 GND.n3222 1.5505
R7187 GND.n3241 GND.n3240 1.5505
R7188 GND.n3237 GND.n3236 1.5505
R7189 GND.n3239 GND.n3224 1.5505
R7190 GND.n4216 GND.n4215 1.5505
R7191 GND.n4190 GND.n4189 1.5505
R7192 GND.n4184 GND.n4180 1.5505
R7193 GND.n4183 GND.n4177 1.5505
R7194 GND.n4206 GND.n4205 1.5505
R7195 GND.n4113 GND.n4112 1.5505
R7196 GND.n4186 GND.n4185 1.5505
R7197 GND.n4202 GND.n4201 1.5505
R7198 GND.n4168 GND.n4167 1.5505
R7199 GND.n4146 GND.n4145 1.5505
R7200 GND.n4164 GND.n4163 1.5505
R7201 GND.n4160 GND.n4159 1.5505
R7202 GND.n4162 GND.n4147 1.5505
R7203 GND.n4271 GND.n4245 1.5505
R7204 GND.n4273 GND.n4272 1.5505
R7205 GND.n4270 GND.n4241 1.5505
R7206 GND.n4267 GND.n4266 1.5505
R7207 GND.n4260 GND.n4258 1.5505
R7208 GND.n4255 GND.n4254 1.5505
R7209 GND.n4246 GND.n4231 1.5505
R7210 GND.n4277 GND.n4229 1.5505
R7211 GND.n4279 GND.n4278 1.5505
R7212 GND.n4283 GND.n4282 1.5505
R7213 GND.n4228 GND.n57 1.5505
R7214 GND.n4227 GND.n4226 1.5505
R7215 GND.n260 GND 1.54738
R7216 GND.n3598 GND 1.54738
R7217 GND.n3578 GND 1.54738
R7218 GND.n3559 GND 1.54738
R7219 GND.n3537 GND 1.54738
R7220 GND.n3518 GND 1.54738
R7221 GND.n3496 GND 1.54738
R7222 GND.n197 GND 1.54738
R7223 GND.n3784 GND 1.51113
R7224 GND.n3789 GND 1.42306
R7225 GND.n3517 GND 1.34833
R7226 GND.n3794 GND 1.335
R7227 GND.n2 GND 1.31102
R7228 GND.n4090 GND 1.27589
R7229 GND.n3303 GND 1.27589
R7230 GND.n3168 GND 1.27589
R7231 GND.n2615 GND 1.27589
R7232 GND.n1870 GND 1.27589
R7233 GND.n1613 GND 1.27589
R7234 GND.n1265 GND 1.27589
R7235 GND.n1395 GND 1.27589
R7236 GND.n1403 GND 1.27589
R7237 GND.n1071 GND 1.27589
R7238 GND.n1877 GND 1.27589
R7239 GND.n1743 GND 1.27589
R7240 GND.n2485 GND 1.27589
R7241 GND.n2623 GND 1.27589
R7242 GND.n3039 GND 1.27589
R7243 GND.n3296 GND 1.27589
R7244 GND.n4219 GND 1.27589
R7245 GND.n3582 GND.n225 1.26851
R7246 GND.n3799 GND 1.24694
R7247 GND.n3804 GND 1.15888
R7248 GND.n3472 GND 1.15267
R7249 GND.n3955 GND.n3954 1.14724
R7250 GND.n3433 GND.n3382 1.14724
R7251 GND.n2897 GND.n2896 1.14724
R7252 GND.n2832 GND.n2827 1.14724
R7253 GND.n2255 GND.n2254 1.14724
R7254 GND.n2065 GND.n766 1.14724
R7255 GND.n2131 GND.n670 1.14724
R7256 GND.n261 GND.n260 1.1418
R7257 GND.n3598 GND.n3597 1.1418
R7258 GND.n3578 GND.n3577 1.1418
R7259 GND.n3559 GND.n3558 1.1418
R7260 GND.n3537 GND.n3536 1.1418
R7261 GND.n3496 GND.n3495 1.1418
R7262 GND.n3877 GND.n197 1.1418
R7263 GND.n3809 GND 1.07082
R7264 GND.n246 GND.n244 1.06843
R7265 GND.n3605 GND.n3604 1.06843
R7266 GND.n3586 GND.n3585 1.06843
R7267 GND.n3566 GND.n3565 1.06843
R7268 GND.n3525 GND.n3524 1.06843
R7269 GND.n3503 GND.n3502 1.06843
R7270 GND.n4087 GND 1.01137
R7271 GND.n4060 GND 1.01137
R7272 GND.n4076 GND 1.01137
R7273 GND.n4073 GND 1.01137
R7274 GND.n4038 GND 1.01137
R7275 GND.n4030 GND 1.01137
R7276 GND.n3316 GND 1.01137
R7277 GND.n3326 GND 1.01137
R7278 GND GND.n391 1.01137
R7279 GND GND.n401 1.01137
R7280 GND GND.n425 1.01137
R7281 GND.n430 GND 1.01137
R7282 GND.n3165 GND 1.01137
R7283 GND.n3138 GND 1.01137
R7284 GND.n3154 GND 1.01137
R7285 GND.n3151 GND 1.01137
R7286 GND.n3116 GND 1.01137
R7287 GND.n3108 GND 1.01137
R7288 GND.n2612 GND 1.01137
R7289 GND.n2585 GND 1.01137
R7290 GND.n2601 GND 1.01137
R7291 GND.n2598 GND 1.01137
R7292 GND.n2563 GND 1.01137
R7293 GND.n2555 GND 1.01137
R7294 GND.n1867 GND 1.01137
R7295 GND.n1840 GND 1.01137
R7296 GND.n1856 GND 1.01137
R7297 GND.n1853 GND 1.01137
R7298 GND.n1818 GND 1.01137
R7299 GND.n1810 GND 1.01137
R7300 GND.n1610 GND 1.01137
R7301 GND.n1583 GND 1.01137
R7302 GND.n1599 GND 1.01137
R7303 GND.n1596 GND 1.01137
R7304 GND.n1561 GND 1.01137
R7305 GND.n1553 GND 1.01137
R7306 GND.n1262 GND 1.01137
R7307 GND.n1235 GND 1.01137
R7308 GND.n1251 GND 1.01137
R7309 GND.n1248 GND 1.01137
R7310 GND.n1213 GND 1.01137
R7311 GND.n1205 GND 1.01137
R7312 GND.n1392 GND 1.01137
R7313 GND.n1365 GND 1.01137
R7314 GND.n1381 GND 1.01137
R7315 GND.n1378 GND 1.01137
R7316 GND.n1343 GND 1.01137
R7317 GND.n1335 GND 1.01137
R7318 GND.n1515 GND 1.01137
R7319 GND.n1508 GND 1.01137
R7320 GND.n1501 GND 1.01137
R7321 GND.n1498 GND 1.01137
R7322 GND.n1483 GND 1.01137
R7323 GND.n1475 GND 1.01137
R7324 GND.n1068 GND 1.01137
R7325 GND GND.n1028 1.01137
R7326 GND.n1058 GND 1.01137
R7327 GND.n1046 GND 1.01137
R7328 GND.n1038 GND 1.01137
R7329 GND.n3597 GND 1.01137
R7330 GND.n3577 GND 1.01137
R7331 GND.n3558 GND 1.01137
R7332 GND.n3536 GND 1.01137
R7333 GND.n3514 GND 1.01137
R7334 GND.n3495 GND 1.01137
R7335 GND.n3877 GND 1.01137
R7336 GND.n3942 GND 1.01137
R7337 GND.n3932 GND 1.01137
R7338 GND GND.n3930 1.01137
R7339 GND.n3918 GND 1.01137
R7340 GND.n3422 GND 1.01137
R7341 GND.n3412 GND 1.01137
R7342 GND GND.n3410 1.01137
R7343 GND.n3887 GND 1.01137
R7344 GND GND.n313 1.01137
R7345 GND GND.n3464 1.01137
R7346 GND.n3455 GND 1.01137
R7347 GND.n3444 GND 1.01137
R7348 GND GND.n511 1.01137
R7349 GND.n2854 GND 1.01137
R7350 GND.n2863 GND 1.01137
R7351 GND.n2875 GND 1.01137
R7352 GND.n2242 GND 1.01137
R7353 GND.n2232 GND 1.01137
R7354 GND GND.n2230 1.01137
R7355 GND.n2218 GND 1.01137
R7356 GND.n754 GND 1.01137
R7357 GND.n744 GND 1.01137
R7358 GND.n2107 GND 1.01137
R7359 GND.n2119 GND 1.01137
R7360 GND GND.n661 1.01137
R7361 GND.n2153 GND 1.01137
R7362 GND.n2162 GND 1.01137
R7363 GND.n2174 GND 1.01137
R7364 GND GND.n2092 1.01137
R7365 GND.n2079 GND 1.01137
R7366 GND GND.n2077 1.01137
R7367 GND GND.n2071 1.01137
R7368 GND.n1989 GND 1.01137
R7369 GND.n1982 GND 1.01137
R7370 GND.n1975 GND 1.01137
R7371 GND.n1972 GND 1.01137
R7372 GND.n1957 GND 1.01137
R7373 GND.n1949 GND 1.01137
R7374 GND.n1740 GND 1.01137
R7375 GND.n1713 GND 1.01137
R7376 GND.n1729 GND 1.01137
R7377 GND.n1726 GND 1.01137
R7378 GND.n1691 GND 1.01137
R7379 GND.n1683 GND 1.01137
R7380 GND.n2482 GND 1.01137
R7381 GND.n2455 GND 1.01137
R7382 GND.n2471 GND 1.01137
R7383 GND.n2468 GND 1.01137
R7384 GND.n2433 GND 1.01137
R7385 GND.n2425 GND 1.01137
R7386 GND.n2735 GND 1.01137
R7387 GND.n2728 GND 1.01137
R7388 GND.n2721 GND 1.01137
R7389 GND.n2718 GND 1.01137
R7390 GND.n2703 GND 1.01137
R7391 GND.n2695 GND 1.01137
R7392 GND.n3036 GND 1.01137
R7393 GND.n3009 GND 1.01137
R7394 GND.n3025 GND 1.01137
R7395 GND.n3022 GND 1.01137
R7396 GND.n2987 GND 1.01137
R7397 GND.n2979 GND 1.01137
R7398 GND.n3293 GND 1.01137
R7399 GND.n3266 GND 1.01137
R7400 GND.n3282 GND 1.01137
R7401 GND.n3279 GND 1.01137
R7402 GND.n3244 GND 1.01137
R7403 GND.n3236 GND 1.01137
R7404 GND.n4216 GND 1.01137
R7405 GND.n4189 GND 1.01137
R7406 GND.n4205 GND 1.01137
R7407 GND.n4202 GND 1.01137
R7408 GND.n4167 GND 1.01137
R7409 GND.n4159 GND 1.01137
R7410 GND.n4271 GND 1.01137
R7411 GND GND.n4267 1.01137
R7412 GND GND.n4255 1.01137
R7413 GND GND.n4246 1.01137
R7414 GND.n4282 GND 1.01137
R7415 GND.n3544 GND.n3543 0.995065
R7416 GND.n3814 GND 0.982757
R7417 GND.n3504 GND.n307 0.935283
R7418 GND.n3819 GND 0.894695
R7419 GND.n3515 GND 0.84425
R7420 GND.n1108 GND 0.821929
R7421 GND GND.n2043 0.821929
R7422 GND GND.n2002 0.821929
R7423 GND.n2325 GND 0.821929
R7424 GND GND.n2805 0.821929
R7425 GND GND.n2929 0.821929
R7426 GND GND.n3978 0.821929
R7427 GND GND.n4310 0.821929
R7428 GND.n3824 GND 0.806633
R7429 GND.n3518 GND.n3517 0.804848
R7430 GND.n3484 GND.n3483 0.791261
R7431 GND.n3829 GND 0.718572
R7432 GND.n3663 GND.n3662 0.682785
R7433 GND.n3757 GND.n3756 0.679084
R7434 GND.n3476 GND.n3475 0.645183
R7435 GND.n3498 GND.n3497 0.645183
R7436 GND.n3520 GND.n3519 0.645183
R7437 GND.n3539 GND.n3538 0.645183
R7438 GND.n3561 GND.n3560 0.645183
R7439 GND.n3580 GND.n3579 0.645183
R7440 GND.n3600 GND.n3599 0.645183
R7441 GND.n257 GND.n256 0.645183
R7442 GND.n1020 GND 0.643357
R7443 GND.n1030 GND 0.643357
R7444 GND.n1044 GND 0.643357
R7445 GND.n4269 GND 0.643357
R7446 GND.n4280 GND 0.643357
R7447 GND.n4225 GND 0.643357
R7448 GND.n262 GND 0.630935
R7449 GND.n3834 GND 0.63051
R7450 GND.n3685 GND.n3684 0.61867
R7451 GND.n3688 GND.n3687 0.61867
R7452 GND.n3691 GND.n3690 0.61867
R7453 GND.n3694 GND.n3693 0.61867
R7454 GND.n3697 GND.n3696 0.61867
R7455 GND.n3700 GND.n3699 0.61867
R7456 GND.n3703 GND.n3702 0.61867
R7457 GND.n3706 GND.n3705 0.61867
R7458 GND.n3709 GND.n3708 0.61867
R7459 GND.n3712 GND.n3711 0.61867
R7460 GND.n3715 GND.n3714 0.61867
R7461 GND.n3718 GND.n3717 0.61867
R7462 GND.n3721 GND.n3720 0.61867
R7463 GND.n3724 GND.n3723 0.61867
R7464 GND.n3727 GND.n3726 0.61867
R7465 GND.n1084 GND.n1083 0.609627
R7466 GND.n1083 GND.n1082 0.609627
R7467 GND.n1108 GND.n976 0.609627
R7468 GND.n1119 GND.n976 0.609627
R7469 GND.n2063 GND.n768 0.609627
R7470 GND.n787 GND.n768 0.609627
R7471 GND.n2043 GND.n797 0.609627
R7472 GND.n840 GND.n797 0.609627
R7473 GND.n867 GND.n865 0.609627
R7474 GND.n868 GND.n867 0.609627
R7475 GND.n2002 GND.n878 0.609627
R7476 GND.n881 GND.n878 0.609627
R7477 GND.n645 GND.n617 0.609627
R7478 GND.n2302 GND.n617 0.609627
R7479 GND.n2326 GND.n2325 0.609627
R7480 GND.n2388 GND.n2326 0.609627
R7481 GND.n2825 GND.n521 0.609627
R7482 GND.n540 GND.n521 0.609627
R7483 GND.n2805 GND.n550 0.609627
R7484 GND.n2758 GND.n550 0.609627
R7485 GND.n2900 GND.n2899 0.609627
R7486 GND.n2942 GND.n2900 0.609627
R7487 GND.n2929 GND.n2928 0.609627
R7488 GND.n2928 GND.n2926 0.609627
R7489 GND.n3380 GND.n99 0.609627
R7490 GND.n3991 GND.n99 0.609627
R7491 GND.n3978 GND.n123 0.609627
R7492 GND.n152 GND.n123 0.609627
R7493 GND.n182 GND.n181 0.609627
R7494 GND.n181 GND.n179 0.609627
R7495 GND.n4310 GND.n4309 0.609627
R7496 GND.n4309 GND.n4307 0.609627
R7497 GND.n3901 GND.n3900 0.606478
R7498 GND.n3941 GND.n3902 0.606478
R7499 GND.n3932 GND.n3931 0.606478
R7500 GND.n3917 GND.n3916 0.606478
R7501 GND.n4368 GND.n4367 0.606478
R7502 GND.n3431 GND.n3383 0.606478
R7503 GND.n3421 GND.n3388 0.606478
R7504 GND.n3412 GND.n3411 0.606478
R7505 GND.n3397 GND.n3396 0.606478
R7506 GND.n3890 GND.n3889 0.606478
R7507 GND.n495 GND.n494 0.606478
R7508 GND.n3466 GND.n3465 0.606478
R7509 GND.n3464 GND.n314 0.606478
R7510 GND.n3453 GND.n324 0.606478
R7511 GND.n3442 GND.n329 0.606478
R7512 GND.n2835 GND.n2834 0.606478
R7513 GND.n2852 GND.n2851 0.606478
R7514 GND.n2854 GND.n2853 0.606478
R7515 GND.n2866 GND.n2865 0.606478
R7516 GND.n2878 GND.n2877 0.606478
R7517 GND.n2190 GND.n2189 0.606478
R7518 GND.n2241 GND.n2191 0.606478
R7519 GND.n2232 GND.n2231 0.606478
R7520 GND.n2210 GND.n2209 0.606478
R7521 GND.n2216 GND.n2211 0.606478
R7522 GND.n735 GND.n734 0.606478
R7523 GND.n753 GND.n736 0.606478
R7524 GND.n744 GND.n743 0.606478
R7525 GND.n2110 GND.n2109 0.606478
R7526 GND.n2122 GND.n2121 0.606478
R7527 GND.n2134 GND.n2133 0.606478
R7528 GND.n2151 GND.n2150 0.606478
R7529 GND.n2153 GND.n2152 0.606478
R7530 GND.n2165 GND.n2164 0.606478
R7531 GND.n2177 GND.n2176 0.606478
R7532 GND.n2094 GND.n2093 0.606478
R7533 GND.n701 GND.n690 0.606478
R7534 GND.n2079 GND.n2078 0.606478
R7535 GND.n2073 GND.n2072 0.606478
R7536 GND.n2067 GND.n2066 0.606478
R7537 GND.n3619 GND.n244 0.601043
R7538 GND.n3606 GND.n3605 0.601043
R7539 GND.n3587 GND.n3586 0.601043
R7540 GND.n3567 GND.n3566 0.601043
R7541 GND.n3526 GND.n3525 0.601043
R7542 GND.n3504 GND.n3503 0.601043
R7543 GND.n3485 GND.n3484 0.601043
R7544 GND.n3475 GND 0.590136
R7545 GND.n3497 GND 0.590136
R7546 GND.n3519 GND 0.590136
R7547 GND.n3538 GND 0.590136
R7548 GND.n3560 GND 0.590136
R7549 GND.n3579 GND 0.590136
R7550 GND.n3599 GND 0.590136
R7551 GND.n256 GND 0.590136
R7552 GND.n4088 GND.n4087 0.543978
R7553 GND.n4054 GND.n4053 0.543978
R7554 GND.n4058 GND.n4057 0.543978
R7555 GND.n4074 GND.n4073 0.543978
R7556 GND.n4017 GND.n4006 0.543978
R7557 GND.n4036 GND.n4035 0.543978
R7558 GND.n3316 GND.n3305 0.543978
R7559 GND.n3314 GND.n3313 0.543978
R7560 GND.n3324 GND.n3323 0.543978
R7561 GND.n401 GND.n393 0.543978
R7562 GND.n404 GND.n403 0.543978
R7563 GND.n428 GND.n427 0.543978
R7564 GND.n3166 GND.n3165 0.543978
R7565 GND.n3132 GND.n3131 0.543978
R7566 GND.n3136 GND.n3135 0.543978
R7567 GND.n3152 GND.n3151 0.543978
R7568 GND.n3095 GND.n3084 0.543978
R7569 GND.n3114 GND.n3113 0.543978
R7570 GND.n2613 GND.n2612 0.543978
R7571 GND.n2579 GND.n2578 0.543978
R7572 GND.n2583 GND.n2582 0.543978
R7573 GND.n2599 GND.n2598 0.543978
R7574 GND.n2542 GND.n2531 0.543978
R7575 GND.n2561 GND.n2560 0.543978
R7576 GND.n1868 GND.n1867 0.543978
R7577 GND.n1834 GND.n1833 0.543978
R7578 GND.n1838 GND.n1837 0.543978
R7579 GND.n1854 GND.n1853 0.543978
R7580 GND.n1797 GND.n1786 0.543978
R7581 GND.n1816 GND.n1815 0.543978
R7582 GND.n1611 GND.n1610 0.543978
R7583 GND.n1577 GND.n1576 0.543978
R7584 GND.n1581 GND.n1580 0.543978
R7585 GND.n1597 GND.n1596 0.543978
R7586 GND.n1540 GND.n1529 0.543978
R7587 GND.n1559 GND.n1558 0.543978
R7588 GND.n1263 GND.n1262 0.543978
R7589 GND.n1229 GND.n1228 0.543978
R7590 GND.n1233 GND.n1232 0.543978
R7591 GND.n1249 GND.n1248 0.543978
R7592 GND.n1192 GND.n1181 0.543978
R7593 GND.n1211 GND.n1210 0.543978
R7594 GND.n1393 GND.n1392 0.543978
R7595 GND.n1359 GND.n1358 0.543978
R7596 GND.n1363 GND.n1362 0.543978
R7597 GND.n1379 GND.n1378 0.543978
R7598 GND.n1322 GND.n1311 0.543978
R7599 GND.n1341 GND.n1340 0.543978
R7600 GND.n1515 GND.n1405 0.543978
R7601 GND.n1513 GND.n1512 0.543978
R7602 GND.n1506 GND.n1505 0.543978
R7603 GND.n1499 GND.n1498 0.543978
R7604 GND.n1435 GND.n1434 0.543978
R7605 GND.n1481 GND.n1480 0.543978
R7606 GND.n1069 GND.n1068 0.543978
R7607 GND.n1021 GND.n1020 0.543978
R7608 GND.n1031 GND.n1030 0.543978
R7609 GND.n1056 GND.n1055 0.543978
R7610 GND.n1044 GND.n1043 0.543978
R7611 GND.n1989 GND.n1879 0.543978
R7612 GND.n1987 GND.n1986 0.543978
R7613 GND.n1980 GND.n1979 0.543978
R7614 GND.n1973 GND.n1972 0.543978
R7615 GND.n1909 GND.n1908 0.543978
R7616 GND.n1955 GND.n1954 0.543978
R7617 GND.n1741 GND.n1740 0.543978
R7618 GND.n1707 GND.n1706 0.543978
R7619 GND.n1711 GND.n1710 0.543978
R7620 GND.n1727 GND.n1726 0.543978
R7621 GND.n1670 GND.n1659 0.543978
R7622 GND.n1689 GND.n1688 0.543978
R7623 GND.n2483 GND.n2482 0.543978
R7624 GND.n2449 GND.n2448 0.543978
R7625 GND.n2453 GND.n2452 0.543978
R7626 GND.n2469 GND.n2468 0.543978
R7627 GND.n2412 GND.n2401 0.543978
R7628 GND.n2431 GND.n2430 0.543978
R7629 GND.n2735 GND.n2625 0.543978
R7630 GND.n2733 GND.n2732 0.543978
R7631 GND.n2726 GND.n2725 0.543978
R7632 GND.n2719 GND.n2718 0.543978
R7633 GND.n2655 GND.n2654 0.543978
R7634 GND.n2701 GND.n2700 0.543978
R7635 GND.n3037 GND.n3036 0.543978
R7636 GND.n3003 GND.n3002 0.543978
R7637 GND.n3007 GND.n3006 0.543978
R7638 GND.n3023 GND.n3022 0.543978
R7639 GND.n2966 GND.n2955 0.543978
R7640 GND.n2985 GND.n2984 0.543978
R7641 GND.n3294 GND.n3293 0.543978
R7642 GND.n3260 GND.n3259 0.543978
R7643 GND.n3264 GND.n3263 0.543978
R7644 GND.n3280 GND.n3279 0.543978
R7645 GND.n3223 GND.n3212 0.543978
R7646 GND.n3242 GND.n3241 0.543978
R7647 GND.n4217 GND.n4216 0.543978
R7648 GND.n4183 GND.n4182 0.543978
R7649 GND.n4187 GND.n4186 0.543978
R7650 GND.n4203 GND.n4202 0.543978
R7651 GND.n4146 GND.n4135 0.543978
R7652 GND.n4165 GND.n4164 0.543978
R7653 GND.n4270 GND.n4269 0.543978
R7654 GND.n4258 GND.n4257 0.543978
R7655 GND.n4255 GND.n4248 0.543978
R7656 GND.n4280 GND.n4279 0.543978
R7657 GND.n4227 GND.n4225 0.543978
R7658 GND.n3839 GND 0.542448
R7659 GND.n3649 GND.n3648 0.537085
R7660 GND.n3651 GND.n3650 0.537085
R7661 GND.n3653 GND.n3652 0.537085
R7662 GND.n3655 GND.n3654 0.537085
R7663 GND.n3657 GND.n3656 0.537085
R7664 GND.n3659 GND.n3658 0.537085
R7665 GND.n3661 GND.n3660 0.537085
R7666 GND.n3665 GND.n3664 0.537085
R7667 GND.n3667 GND.n3666 0.537085
R7668 GND.n3669 GND.n3668 0.537085
R7669 GND.n3671 GND.n3670 0.537085
R7670 GND.n3673 GND.n3672 0.537085
R7671 GND.n3675 GND.n3674 0.537085
R7672 GND.n3677 GND.n3676 0.537085
R7673 GND.n3736 GND.n3735 0.533384
R7674 GND.n3739 GND.n3738 0.533384
R7675 GND.n3742 GND.n3741 0.533384
R7676 GND.n3745 GND.n3744 0.533384
R7677 GND.n3748 GND.n3747 0.533384
R7678 GND.n3751 GND.n3750 0.533384
R7679 GND.n3754 GND.n3753 0.533384
R7680 GND.n3760 GND.n3759 0.533384
R7681 GND.n3763 GND.n3762 0.533384
R7682 GND.n3766 GND.n3765 0.533384
R7683 GND.n3769 GND.n3768 0.533384
R7684 GND.n3772 GND.n3771 0.533384
R7685 GND.n3775 GND.n3774 0.533384
R7686 GND.n3778 GND.n3777 0.533384
R7687 GND.n3548 GND.n3547 0.5005
R7688 GND.n3730 GND.n3729 0.485508
R7689 GND.n3682 GND.n3681 0.481462
R7690 GND GND.n264 0.457022
R7691 GND.n3844 GND 0.454387
R7692 GND.n1056 GND 0.424071
R7693 GND.n4257 GND 0.424071
R7694 GND.n3679 GND.n3678 0.420684
R7695 GND.n3582 GND.n3581 0.419583
R7696 GND.n3647 GND.n1 0.417701
R7697 GND.n3782 GND.n3780 0.417343
R7698 GND.n3733 GND.n3732 0.417341
R7699 GND GND.n3901 0.405391
R7700 GND GND.n3902 0.405391
R7701 GND.n3931 GND 0.405391
R7702 GND GND.n3917 0.405391
R7703 GND GND.n4368 0.405391
R7704 GND GND.n3383 0.405391
R7705 GND GND.n3388 0.405391
R7706 GND.n3411 GND 0.405391
R7707 GND.n3396 GND 0.405391
R7708 GND.n3889 GND 0.405391
R7709 GND.n494 GND 0.405391
R7710 GND.n3465 GND 0.405391
R7711 GND GND.n314 0.405391
R7712 GND GND.n324 0.405391
R7713 GND GND.n329 0.405391
R7714 GND.n2834 GND 0.405391
R7715 GND GND.n2852 0.405391
R7716 GND.n2853 GND 0.405391
R7717 GND.n2865 GND 0.405391
R7718 GND.n2877 GND 0.405391
R7719 GND GND.n2190 0.405391
R7720 GND GND.n2191 0.405391
R7721 GND.n2231 GND 0.405391
R7722 GND GND.n2210 0.405391
R7723 GND.n2211 GND 0.405391
R7724 GND GND.n735 0.405391
R7725 GND GND.n736 0.405391
R7726 GND.n743 GND 0.405391
R7727 GND.n2109 GND 0.405391
R7728 GND.n2121 GND 0.405391
R7729 GND.n2133 GND 0.405391
R7730 GND GND.n2151 0.405391
R7731 GND.n2152 GND 0.405391
R7732 GND.n2164 GND 0.405391
R7733 GND.n2176 GND 0.405391
R7734 GND.n2093 GND 0.405391
R7735 GND GND.n701 0.405391
R7736 GND.n2078 GND 0.405391
R7737 GND.n2072 GND 0.405391
R7738 GND.n2066 GND 0.405391
R7739 GND.n262 GND.n261 0.380935
R7740 GND GND.n1080 0.369548
R7741 GND.n1121 GND 0.369548
R7742 GND GND.n2063 0.369548
R7743 GND.n789 GND 0.369548
R7744 GND.n842 GND 0.369548
R7745 GND.n865 GND 0.369548
R7746 GND.n870 GND 0.369548
R7747 GND GND.n629 0.369548
R7748 GND GND.n645 0.369548
R7749 GND.n2304 GND 0.369548
R7750 GND GND.n2386 0.369548
R7751 GND GND.n2825 0.369548
R7752 GND.n542 GND 0.369548
R7753 GND.n2760 GND 0.369548
R7754 GND.n2899 GND 0.369548
R7755 GND GND.n2940 0.369548
R7756 GND.n3347 GND 0.369548
R7757 GND GND.n3380 0.369548
R7758 GND GND.n3989 0.369548
R7759 GND.n154 GND 0.369548
R7760 GND GND.n182 0.369548
R7761 GND GND.n177 0.369548
R7762 GND.n4329 GND 0.369548
R7763 GND.n3849 GND 0.366325
R7764 GND.n255 GND.n246 0.353761
R7765 GND.n3604 GND.n3603 0.353761
R7766 GND.n3585 GND.n3584 0.353761
R7767 GND.n3565 GND.n3564 0.353761
R7768 GND.n3543 GND.n3542 0.353761
R7769 GND.n3524 GND.n3523 0.353761
R7770 GND.n3502 GND.n3501 0.353761
R7771 GND.n3480 GND.n3479 0.353761
R7772 GND.n1165 GND.n1122 0.350698
R7773 GND.n847 GND.n845 0.350698
R7774 GND.n2288 GND.n630 0.350698
R7775 GND.n2375 GND.n2333 0.350698
R7776 GND.n2765 GND.n2763 0.350698
R7777 GND.n3348 GND.n343 0.350698
R7778 GND.n159 GND.n157 0.350698
R7779 GND.n4330 GND.n18 0.350698
R7780 GND.n3786 GND.n3785 0.3483
R7781 GND.n3791 GND.n3790 0.3483
R7782 GND.n3796 GND.n3795 0.3483
R7783 GND.n3801 GND.n3800 0.3483
R7784 GND.n3806 GND.n3805 0.3483
R7785 GND.n3811 GND.n3810 0.3483
R7786 GND.n3816 GND.n3815 0.3483
R7787 GND.n3821 GND.n3820 0.3483
R7788 GND.n3826 GND.n3825 0.3483
R7789 GND.n3831 GND.n3830 0.3483
R7790 GND.n3836 GND.n3835 0.3483
R7791 GND.n3841 GND.n3840 0.3483
R7792 GND.n3846 GND.n3845 0.3483
R7793 GND.n3851 GND.n3850 0.3483
R7794 GND.n3856 GND.n3855 0.3483
R7795 GND.n3871 GND.n3870 0.3483
R7796 GND.n3866 GND.n3 0.3483
R7797 GND.n4053 GND 0.344537
R7798 GND.n4058 GND 0.344537
R7799 GND.n4036 GND 0.344537
R7800 GND.n3314 GND 0.344537
R7801 GND.n3324 GND 0.344537
R7802 GND.n427 GND 0.344537
R7803 GND.n3131 GND 0.344537
R7804 GND.n3136 GND 0.344537
R7805 GND.n3114 GND 0.344537
R7806 GND.n2578 GND 0.344537
R7807 GND.n2583 GND 0.344537
R7808 GND.n2561 GND 0.344537
R7809 GND.n1833 GND 0.344537
R7810 GND.n1838 GND 0.344537
R7811 GND.n1816 GND 0.344537
R7812 GND.n1576 GND 0.344537
R7813 GND.n1581 GND 0.344537
R7814 GND.n1559 GND 0.344537
R7815 GND.n1228 GND 0.344537
R7816 GND.n1233 GND 0.344537
R7817 GND.n1211 GND 0.344537
R7818 GND.n1358 GND 0.344537
R7819 GND.n1363 GND 0.344537
R7820 GND.n1341 GND 0.344537
R7821 GND.n1513 GND 0.344537
R7822 GND.n1506 GND 0.344537
R7823 GND.n1481 GND 0.344537
R7824 GND.n1987 GND 0.344537
R7825 GND.n1980 GND 0.344537
R7826 GND.n1955 GND 0.344537
R7827 GND.n1706 GND 0.344537
R7828 GND.n1711 GND 0.344537
R7829 GND.n1689 GND 0.344537
R7830 GND.n2448 GND 0.344537
R7831 GND.n2453 GND 0.344537
R7832 GND.n2431 GND 0.344537
R7833 GND.n2733 GND 0.344537
R7834 GND.n2726 GND 0.344537
R7835 GND.n2701 GND 0.344537
R7836 GND.n3002 GND 0.344537
R7837 GND.n3007 GND 0.344537
R7838 GND.n2985 GND 0.344537
R7839 GND.n3259 GND 0.344537
R7840 GND.n3264 GND 0.344537
R7841 GND.n3242 GND 0.344537
R7842 GND.n4182 GND 0.344537
R7843 GND.n4187 GND 0.344537
R7844 GND.n4165 GND 0.344537
R7845 GND.n4052 GND 0.342891
R7846 GND GND.n4059 0.342891
R7847 GND GND.n4075 0.342891
R7848 GND.n4005 GND 0.342891
R7849 GND GND.n4037 0.342891
R7850 GND GND.n3315 0.342891
R7851 GND GND.n3325 0.342891
R7852 GND.n392 GND 0.342891
R7853 GND.n402 GND 0.342891
R7854 GND.n426 GND 0.342891
R7855 GND.n3130 GND 0.342891
R7856 GND GND.n3137 0.342891
R7857 GND GND.n3153 0.342891
R7858 GND.n3083 GND 0.342891
R7859 GND GND.n3115 0.342891
R7860 GND.n2577 GND 0.342891
R7861 GND GND.n2584 0.342891
R7862 GND GND.n2600 0.342891
R7863 GND.n2530 GND 0.342891
R7864 GND GND.n2562 0.342891
R7865 GND.n1832 GND 0.342891
R7866 GND GND.n1839 0.342891
R7867 GND GND.n1855 0.342891
R7868 GND.n1785 GND 0.342891
R7869 GND GND.n1817 0.342891
R7870 GND.n1575 GND 0.342891
R7871 GND GND.n1582 0.342891
R7872 GND GND.n1598 0.342891
R7873 GND.n1528 GND 0.342891
R7874 GND GND.n1560 0.342891
R7875 GND.n1227 GND 0.342891
R7876 GND GND.n1234 0.342891
R7877 GND GND.n1250 0.342891
R7878 GND.n1180 GND 0.342891
R7879 GND GND.n1212 0.342891
R7880 GND.n1357 GND 0.342891
R7881 GND GND.n1364 0.342891
R7882 GND GND.n1380 0.342891
R7883 GND.n1310 GND 0.342891
R7884 GND GND.n1342 0.342891
R7885 GND GND.n1514 0.342891
R7886 GND GND.n1507 0.342891
R7887 GND GND.n1500 0.342891
R7888 GND.n1433 GND 0.342891
R7889 GND GND.n1482 0.342891
R7890 GND.n1019 GND 0.342891
R7891 GND.n1029 GND 0.342891
R7892 GND GND.n1045 0.342891
R7893 GND GND.n1988 0.342891
R7894 GND GND.n1981 0.342891
R7895 GND GND.n1974 0.342891
R7896 GND.n1907 GND 0.342891
R7897 GND GND.n1956 0.342891
R7898 GND.n1705 GND 0.342891
R7899 GND GND.n1712 0.342891
R7900 GND GND.n1728 0.342891
R7901 GND.n1658 GND 0.342891
R7902 GND GND.n1690 0.342891
R7903 GND.n2447 GND 0.342891
R7904 GND GND.n2454 0.342891
R7905 GND GND.n2470 0.342891
R7906 GND.n2400 GND 0.342891
R7907 GND GND.n2432 0.342891
R7908 GND GND.n2734 0.342891
R7909 GND GND.n2727 0.342891
R7910 GND GND.n2720 0.342891
R7911 GND.n2653 GND 0.342891
R7912 GND GND.n2702 0.342891
R7913 GND.n3001 GND 0.342891
R7914 GND GND.n3008 0.342891
R7915 GND GND.n3024 0.342891
R7916 GND.n2954 GND 0.342891
R7917 GND GND.n2986 0.342891
R7918 GND.n3258 GND 0.342891
R7919 GND GND.n3265 0.342891
R7920 GND GND.n3281 0.342891
R7921 GND.n3211 GND 0.342891
R7922 GND GND.n3243 0.342891
R7923 GND.n4181 GND 0.342891
R7924 GND GND.n4188 0.342891
R7925 GND GND.n4204 0.342891
R7926 GND.n4134 GND 0.342891
R7927 GND GND.n4166 0.342891
R7928 GND.n4268 GND 0.342891
R7929 GND.n4256 GND 0.342891
R7930 GND.n4247 GND 0.342891
R7931 GND GND.n4281 0.342891
R7932 GND.n264 GND 0.328625
R7933 GND.n1078 GND.n1075 0.323913
R7934 GND.n795 GND.n794 0.323913
R7935 GND.n876 GND.n875 0.323913
R7936 GND.n2307 GND.n2306 0.323913
R7937 GND.n548 GND.n547 0.323913
R7938 GND.n2923 GND.n2922 0.323913
R7939 GND.n121 GND.n120 0.323913
R7940 GND.n4304 GND.n36 0.323913
R7941 GND.n3681 GND.n3680 0.29425
R7942 GND.n3730 GND.n3629 0.29425
R7943 GND.n3854 GND 0.278263
R7944 GND.n3785 GND.n3784 0.27075
R7945 GND.n3787 GND.n3786 0.27075
R7946 GND.n3790 GND.n3789 0.27075
R7947 GND.n3792 GND.n3791 0.27075
R7948 GND.n3795 GND.n3794 0.27075
R7949 GND.n3797 GND.n3796 0.27075
R7950 GND.n3800 GND.n3799 0.27075
R7951 GND.n3802 GND.n3801 0.27075
R7952 GND.n3805 GND.n3804 0.27075
R7953 GND.n3807 GND.n3806 0.27075
R7954 GND.n3810 GND.n3809 0.27075
R7955 GND.n3812 GND.n3811 0.27075
R7956 GND.n3815 GND.n3814 0.27075
R7957 GND.n3817 GND.n3816 0.27075
R7958 GND.n3820 GND.n3819 0.27075
R7959 GND.n3822 GND.n3821 0.27075
R7960 GND.n3825 GND.n3824 0.27075
R7961 GND.n3827 GND.n3826 0.27075
R7962 GND.n3830 GND.n3829 0.27075
R7963 GND.n3832 GND.n3831 0.27075
R7964 GND.n3835 GND.n3834 0.27075
R7965 GND.n3837 GND.n3836 0.27075
R7966 GND.n3840 GND.n3839 0.27075
R7967 GND.n3842 GND.n3841 0.27075
R7968 GND.n3845 GND.n3844 0.27075
R7969 GND.n3847 GND.n3846 0.27075
R7970 GND.n3850 GND.n3849 0.27075
R7971 GND.n3852 GND.n3851 0.27075
R7972 GND.n3855 GND.n3854 0.27075
R7973 GND.n3857 GND.n3856 0.27075
R7974 GND.n3871 GND.n3858 0.27075
R7975 GND.n3870 GND.n3869 0.27075
R7976 GND.n3866 GND.n3865 0.27075
R7977 GND.n3 GND.n2 0.27075
R7978 GND.n4375 GND.n4374 0.27075
R7979 GND.n289 GND 0.26137
R7980 GND.n1133 GND.n1122 0.259429
R7981 GND.n845 GND.n843 0.259429
R7982 GND.n641 GND.n630 0.259429
R7983 GND.n2375 GND.n2374 0.259429
R7984 GND.n2763 GND.n2761 0.259429
R7985 GND.n3364 GND.n343 0.259429
R7986 GND.n157 GND.n155 0.259429
R7987 GND.n4346 GND.n18 0.259429
R7988 GND.n3732 GND.n3629 0.24725
R7989 GND.n3680 GND.n3679 0.24725
R7990 GND.n3783 GND.n3782 0.24725
R7991 GND.n1 GND.n0 0.24725
R7992 GND.n4006 GND 0.227182
R7993 GND.n403 GND 0.227182
R7994 GND.n3084 GND 0.227182
R7995 GND.n2531 GND 0.227182
R7996 GND.n1786 GND 0.227182
R7997 GND.n1529 GND 0.227182
R7998 GND.n1181 GND 0.227182
R7999 GND.n1311 GND 0.227182
R8000 GND.n1434 GND 0.227182
R8001 GND.n1908 GND 0.227182
R8002 GND.n1659 GND 0.227182
R8003 GND.n2401 GND 0.227182
R8004 GND.n2654 GND 0.227182
R8005 GND.n2955 GND 0.227182
R8006 GND.n3212 GND 0.227182
R8007 GND.n4135 GND 0.227182
R8008 GND.n4372 GND.n4371 0.223445
R8009 GND.n3864 GND.n3859 0.223445
R8010 GND.n3874 GND.n199 0.223445
R8011 GND.n202 GND.n201 0.223445
R8012 GND.n205 GND.n204 0.223445
R8013 GND.n208 GND.n207 0.223445
R8014 GND.n211 GND.n210 0.223445
R8015 GND.n214 GND.n213 0.223445
R8016 GND.n217 GND.n216 0.223445
R8017 GND.n220 GND.n219 0.223445
R8018 GND.n223 GND.n222 0.223445
R8019 GND.n229 GND.n228 0.223445
R8020 GND.n232 GND.n231 0.223445
R8021 GND.n235 GND.n234 0.223445
R8022 GND.n238 GND.n237 0.223445
R8023 GND.n241 GND.n240 0.223445
R8024 GND.n1082 GND.n1081 0.22173
R8025 GND.n1079 GND.n1078 0.22173
R8026 GND.n1075 GND.n985 0.22173
R8027 GND.n1120 GND.n1119 0.22173
R8028 GND.n1167 GND.n1121 0.22173
R8029 GND.n1167 GND.n1166 0.22173
R8030 GND.n1134 GND.n1133 0.22173
R8031 GND.n1150 GND.n767 0.22173
R8032 GND.n788 GND.n787 0.22173
R8033 GND.n794 GND.n790 0.22173
R8034 GND.n796 GND.n795 0.22173
R8035 GND.n841 GND.n840 0.22173
R8036 GND.n849 GND.n842 0.22173
R8037 GND.n849 GND.n848 0.22173
R8038 GND.n843 GND.n830 0.22173
R8039 GND.n863 GND.n862 0.22173
R8040 GND.n869 GND.n868 0.22173
R8041 GND.n875 GND.n871 0.22173
R8042 GND.n877 GND.n876 0.22173
R8043 GND.n881 GND.n880 0.22173
R8044 GND.n2290 GND.n629 0.22173
R8045 GND.n2290 GND.n2289 0.22173
R8046 GND.n642 GND.n641 0.22173
R8047 GND.n2273 GND.n2257 0.22173
R8048 GND.n2303 GND.n2302 0.22173
R8049 GND.n2307 GND.n2305 0.22173
R8050 GND.n2306 GND.n604 0.22173
R8051 GND.n2388 GND.n2387 0.22173
R8052 GND.n2386 GND.n2330 0.22173
R8053 GND.n2332 GND.n2330 0.22173
R8054 GND.n2374 GND.n2373 0.22173
R8055 GND.n2365 GND.n520 0.22173
R8056 GND.n541 GND.n540 0.22173
R8057 GND.n547 GND.n543 0.22173
R8058 GND.n549 GND.n548 0.22173
R8059 GND.n2759 GND.n2758 0.22173
R8060 GND.n2767 GND.n2760 0.22173
R8061 GND.n2767 GND.n2766 0.22173
R8062 GND.n2761 GND.n2747 0.22173
R8063 GND.n2780 GND.n491 0.22173
R8064 GND.n2942 GND.n2941 0.22173
R8065 GND.n2922 GND.n2904 0.22173
R8066 GND.n2924 GND.n2923 0.22173
R8067 GND.n2926 GND.n2925 0.22173
R8068 GND.n3350 GND.n3347 0.22173
R8069 GND.n3350 GND.n3349 0.22173
R8070 GND.n3365 GND.n3364 0.22173
R8071 GND.n3379 GND.n3378 0.22173
R8072 GND.n3991 GND.n3990 0.22173
R8073 GND.n120 GND.n103 0.22173
R8074 GND.n122 GND.n121 0.22173
R8075 GND.n153 GND.n152 0.22173
R8076 GND.n161 GND.n154 0.22173
R8077 GND.n161 GND.n160 0.22173
R8078 GND.n155 GND.n142 0.22173
R8079 GND.n3958 GND.n3957 0.22173
R8080 GND.n179 GND.n178 0.22173
R8081 GND.n174 GND.n36 0.22173
R8082 GND.n4305 GND.n4304 0.22173
R8083 GND.n4307 GND.n4306 0.22173
R8084 GND.n4332 GND.n4329 0.22173
R8085 GND.n4332 GND.n4331 0.22173
R8086 GND.n4347 GND.n4346 0.22173
R8087 GND.n4348 GND.n4 0.22173
R8088 GND.n226 GND.n225 0.217933
R8089 GND.n3606 GND.n267 0.217891
R8090 GND.n3627 GND.n242 0.211695
R8091 GND.n4088 GND 0.204786
R8092 GND.n4074 GND 0.204786
R8093 GND.n3305 GND 0.204786
R8094 GND.n393 GND 0.204786
R8095 GND.n3166 GND 0.204786
R8096 GND.n3152 GND 0.204786
R8097 GND.n2613 GND 0.204786
R8098 GND.n2599 GND 0.204786
R8099 GND.n1868 GND 0.204786
R8100 GND.n1854 GND 0.204786
R8101 GND.n1611 GND 0.204786
R8102 GND.n1597 GND 0.204786
R8103 GND.n1263 GND 0.204786
R8104 GND.n1249 GND 0.204786
R8105 GND.n1393 GND 0.204786
R8106 GND.n1379 GND 0.204786
R8107 GND.n1405 GND 0.204786
R8108 GND.n1499 GND 0.204786
R8109 GND.n1069 GND 0.204786
R8110 GND.n1879 GND 0.204786
R8111 GND.n1973 GND 0.204786
R8112 GND.n1741 GND 0.204786
R8113 GND.n1727 GND 0.204786
R8114 GND.n2483 GND 0.204786
R8115 GND.n2469 GND 0.204786
R8116 GND.n2625 GND 0.204786
R8117 GND.n2719 GND 0.204786
R8118 GND.n3037 GND 0.204786
R8119 GND.n3023 GND 0.204786
R8120 GND.n3294 GND 0.204786
R8121 GND.n3280 GND 0.204786
R8122 GND.n4217 GND 0.204786
R8123 GND.n4203 GND 0.204786
R8124 GND.n4248 GND 0.204786
R8125 GND GND.n1151 0.202881
R8126 GND.n861 GND 0.202881
R8127 GND GND.n2274 0.202881
R8128 GND.n2364 GND 0.202881
R8129 GND.n2779 GND 0.202881
R8130 GND GND.n3366 0.202881
R8131 GND.n173 GND 0.202881
R8132 GND GND.n4349 0.202881
R8133 GND.n3858 GND 0.190202
R8134 GND.n3515 GND.n3514 0.163543
R8135 GND.n3683 GND.n3682 0.151458
R8136 GND.n3686 GND.n3685 0.151458
R8137 GND.n3689 GND.n3688 0.151458
R8138 GND.n3692 GND.n3691 0.151458
R8139 GND.n3695 GND.n3694 0.151458
R8140 GND.n3698 GND.n3697 0.151458
R8141 GND.n3701 GND.n3700 0.151458
R8142 GND.n3704 GND.n3703 0.151458
R8143 GND.n3707 GND.n3706 0.151458
R8144 GND.n3710 GND.n3709 0.151458
R8145 GND.n3713 GND.n3712 0.151458
R8146 GND.n3716 GND.n3715 0.151458
R8147 GND.n3719 GND.n3718 0.151458
R8148 GND.n3722 GND.n3721 0.151458
R8149 GND.n3725 GND.n3724 0.151458
R8150 GND.n3728 GND.n3727 0.151458
R8151 GND.n1081 GND 0.148317
R8152 GND GND.n1120 0.148317
R8153 GND.n1166 GND 0.148317
R8154 GND.n1151 GND 0.148317
R8155 GND GND.n788 0.148317
R8156 GND GND.n841 0.148317
R8157 GND.n848 GND 0.148317
R8158 GND GND.n861 0.148317
R8159 GND GND.n869 0.148317
R8160 GND.n880 GND 0.148317
R8161 GND.n2289 GND 0.148317
R8162 GND.n2274 GND 0.148317
R8163 GND GND.n2303 0.148317
R8164 GND.n2387 GND 0.148317
R8165 GND GND.n2332 0.148317
R8166 GND GND.n2364 0.148317
R8167 GND GND.n541 0.148317
R8168 GND GND.n2759 0.148317
R8169 GND.n2766 GND 0.148317
R8170 GND GND.n2779 0.148317
R8171 GND.n2941 GND 0.148317
R8172 GND.n2925 GND 0.148317
R8173 GND.n3349 GND 0.148317
R8174 GND.n3366 GND 0.148317
R8175 GND.n3990 GND 0.148317
R8176 GND GND.n153 0.148317
R8177 GND.n160 GND 0.148317
R8178 GND GND.n173 0.148317
R8179 GND.n178 GND 0.148317
R8180 GND.n4306 GND 0.148317
R8181 GND.n4331 GND 0.148317
R8182 GND.n4349 GND 0.148317
R8183 GND.n3729 GND.n3728 0.14768
R8184 GND.n3726 GND.n3725 0.14768
R8185 GND.n3723 GND.n3722 0.14768
R8186 GND.n3720 GND.n3719 0.14768
R8187 GND.n3717 GND.n3716 0.14768
R8188 GND.n3714 GND.n3713 0.14768
R8189 GND.n3711 GND.n3710 0.14768
R8190 GND.n3708 GND.n3707 0.14768
R8191 GND.n3705 GND.n3704 0.14768
R8192 GND.n3702 GND.n3701 0.14768
R8193 GND.n3699 GND.n3698 0.14768
R8194 GND.n3696 GND.n3695 0.14768
R8195 GND.n3693 GND.n3692 0.14768
R8196 GND.n3690 GND.n3689 0.14768
R8197 GND.n3687 GND.n3686 0.14768
R8198 GND.n3684 GND.n3683 0.14768
R8199 GND.n1152 GND.n1134 0.129468
R8200 GND.n860 GND.n830 0.129468
R8201 GND.n2275 GND.n642 0.129468
R8202 GND.n2373 GND.n2372 0.129468
R8203 GND.n2778 GND.n2747 0.129468
R8204 GND.n3367 GND.n3365 0.129468
R8205 GND.n172 GND.n142 0.129468
R8206 GND.n4350 GND.n4347 0.129468
R8207 GND.n3734 GND.n3733 0.124897
R8208 GND.n3737 GND.n3736 0.124897
R8209 GND.n3740 GND.n3739 0.124897
R8210 GND.n3743 GND.n3742 0.124897
R8211 GND.n3746 GND.n3745 0.124897
R8212 GND.n3749 GND.n3748 0.124897
R8213 GND.n3752 GND.n3751 0.124897
R8214 GND.n3755 GND.n3754 0.124897
R8215 GND.n3758 GND.n3757 0.124897
R8216 GND.n3761 GND.n3760 0.124897
R8217 GND.n3764 GND.n3763 0.124897
R8218 GND.n3767 GND.n3766 0.124897
R8219 GND.n3770 GND.n3769 0.124897
R8220 GND.n3773 GND.n3772 0.124897
R8221 GND.n3776 GND.n3775 0.124897
R8222 GND.n3779 GND.n3778 0.124897
R8223 GND.n3735 GND.n3734 0.124897
R8224 GND.n3738 GND.n3737 0.124897
R8225 GND.n3741 GND.n3740 0.124897
R8226 GND.n3744 GND.n3743 0.124897
R8227 GND.n3747 GND.n3746 0.124897
R8228 GND.n3750 GND.n3749 0.124897
R8229 GND.n3753 GND.n3752 0.124897
R8230 GND.n3756 GND.n3755 0.124897
R8231 GND.n3759 GND.n3758 0.124897
R8232 GND.n3762 GND.n3761 0.124897
R8233 GND.n3765 GND.n3764 0.124897
R8234 GND.n3768 GND.n3767 0.124897
R8235 GND.n3771 GND.n3770 0.124897
R8236 GND.n3774 GND.n3773 0.124897
R8237 GND.n3777 GND.n3776 0.124897
R8238 GND.n3780 GND.n3779 0.124897
R8239 GND.n3647 GND.n3646 0.124539
R8240 GND.n3649 GND.n3645 0.124539
R8241 GND.n3651 GND.n3644 0.124539
R8242 GND.n3653 GND.n3643 0.124539
R8243 GND.n3655 GND.n3642 0.124539
R8244 GND.n3657 GND.n3641 0.124539
R8245 GND.n3659 GND.n3640 0.124539
R8246 GND.n3661 GND.n3639 0.124539
R8247 GND.n3663 GND.n3638 0.124539
R8248 GND.n3665 GND.n3637 0.124539
R8249 GND.n3667 GND.n3636 0.124539
R8250 GND.n3669 GND.n3635 0.124539
R8251 GND.n3671 GND.n3634 0.124539
R8252 GND.n3673 GND.n3633 0.124539
R8253 GND.n3675 GND.n3632 0.124539
R8254 GND.n3677 GND.n3631 0.124539
R8255 GND.n3678 GND.n3631 0.121365
R8256 GND.n3676 GND.n3632 0.121365
R8257 GND.n3674 GND.n3633 0.121365
R8258 GND.n3672 GND.n3634 0.121365
R8259 GND.n3670 GND.n3635 0.121365
R8260 GND.n3668 GND.n3636 0.121365
R8261 GND.n3666 GND.n3637 0.121365
R8262 GND.n3664 GND.n3638 0.121365
R8263 GND.n3662 GND.n3639 0.121365
R8264 GND.n3660 GND.n3640 0.121365
R8265 GND.n3658 GND.n3641 0.121365
R8266 GND.n3656 GND.n3642 0.121365
R8267 GND.n3654 GND.n3643 0.121365
R8268 GND.n3652 GND.n3644 0.121365
R8269 GND.n3650 GND.n3645 0.121365
R8270 GND.n3648 GND.n3646 0.121365
R8271 GND.n3481 GND.n3480 0.103761
R8272 GND.n3865 GND 0.10214
R8273 GND.n4090 GND.n4089 0.0956087
R8274 GND.n3304 GND.n3303 0.0956087
R8275 GND.n3168 GND.n3167 0.0956087
R8276 GND.n2615 GND.n2614 0.0956087
R8277 GND.n1870 GND.n1869 0.0956087
R8278 GND.n1613 GND.n1612 0.0956087
R8279 GND.n1265 GND.n1264 0.0956087
R8280 GND.n1395 GND.n1394 0.0956087
R8281 GND.n1404 GND.n1403 0.0956087
R8282 GND.n1071 GND.n1070 0.0956087
R8283 GND.n1878 GND.n1877 0.0956087
R8284 GND.n1743 GND.n1742 0.0956087
R8285 GND.n2485 GND.n2484 0.0956087
R8286 GND.n2624 GND.n2623 0.0956087
R8287 GND.n3039 GND.n3038 0.0956087
R8288 GND.n3296 GND.n3295 0.0956087
R8289 GND.n4219 GND.n4218 0.0956087
R8290 GND.n2064 GND.n767 0.0897857
R8291 GND.n864 GND.n863 0.0897857
R8292 GND.n2257 GND.n2256 0.0897857
R8293 GND.n2826 GND.n520 0.0897857
R8294 GND.n2898 GND.n491 0.0897857
R8295 GND.n3381 GND.n3379 0.0897857
R8296 GND.n3957 GND.n3956 0.0897857
R8297 GND.n4369 GND.n4 0.0897857
R8298 GND GND.n1107 0.0838333
R8299 GND.n2044 GND 0.0838333
R8300 GND.n2003 GND 0.0838333
R8301 GND GND.n2324 0.0838333
R8302 GND.n2806 GND 0.0838333
R8303 GND.n2930 GND 0.0838333
R8304 GND.n3979 GND 0.0838333
R8305 GND.n4311 GND 0.0838333
R8306 GND.n1080 GND.n1079 0.0649841
R8307 GND.n1107 GND.n985 0.0649841
R8308 GND.n790 GND.n789 0.0649841
R8309 GND.n2044 GND.n796 0.0649841
R8310 GND.n871 GND.n870 0.0649841
R8311 GND.n2003 GND.n877 0.0649841
R8312 GND.n2305 GND.n2304 0.0649841
R8313 GND.n2324 GND.n604 0.0649841
R8314 GND.n543 GND.n542 0.0649841
R8315 GND.n2806 GND.n549 0.0649841
R8316 GND.n2940 GND.n2904 0.0649841
R8317 GND.n2930 GND.n2924 0.0649841
R8318 GND.n3989 GND.n103 0.0649841
R8319 GND.n3979 GND.n122 0.0649841
R8320 GND.n177 GND.n174 0.0649841
R8321 GND.n4311 GND.n4305 0.0649841
R8322 GND.n4091 GND.n4090 0.063
R8323 GND.n3303 GND.n3302 0.063
R8324 GND.n3169 GND.n3168 0.063
R8325 GND.n2616 GND.n2615 0.063
R8326 GND.n1871 GND.n1870 0.063
R8327 GND.n1614 GND.n1613 0.063
R8328 GND.n1266 GND.n1265 0.063
R8329 GND.n1396 GND.n1395 0.063
R8330 GND.n1403 GND.n1402 0.063
R8331 GND.n1072 GND.n1071 0.063
R8332 GND.n3625 GND.n3624 0.063
R8333 GND.n3624 GND.n3623 0.063
R8334 GND.n3622 GND.n3621 0.063
R8335 GND.n3621 GND.n3620 0.063
R8336 GND.n259 GND.n255 0.063
R8337 GND.n260 GND.n259 0.063
R8338 GND.n263 GND.n262 0.063
R8339 GND.n264 GND.n263 0.063
R8340 GND.n266 GND.n265 0.063
R8341 GND.n267 GND.n266 0.063
R8342 GND.n3603 GND.n3602 0.063
R8343 GND.n3602 GND.n3598 0.063
R8344 GND.n274 GND.n273 0.063
R8345 GND.n275 GND.n274 0.063
R8346 GND.n3584 GND.n3583 0.063
R8347 GND.n3583 GND.n3578 0.063
R8348 GND.n282 GND.n281 0.063
R8349 GND.n283 GND.n282 0.063
R8350 GND.n3564 GND.n3563 0.063
R8351 GND.n3563 GND.n3559 0.063
R8352 GND.n290 GND.n289 0.063
R8353 GND.n291 GND.n290 0.063
R8354 GND.n3547 GND.n3546 0.063
R8355 GND.n3542 GND.n3541 0.063
R8356 GND.n3541 GND.n3537 0.063
R8357 GND.n298 GND.n297 0.063
R8358 GND.n299 GND.n298 0.063
R8359 GND.n3523 GND.n3522 0.063
R8360 GND.n3522 GND.n3518 0.063
R8361 GND.n3517 GND.n3516 0.063
R8362 GND.n3516 GND.n3515 0.063
R8363 GND.n306 GND.n305 0.063
R8364 GND.n307 GND.n306 0.063
R8365 GND.n3501 GND.n3500 0.063
R8366 GND.n3500 GND.n3496 0.063
R8367 GND.n3473 GND.n3472 0.063
R8368 GND.n3474 GND.n3473 0.063
R8369 GND.n3483 GND.n3482 0.063
R8370 GND.n3482 GND.n3481 0.063
R8371 GND.n3479 GND.n3478 0.063
R8372 GND.n3478 GND.n197 0.063
R8373 GND.n3876 GND.n3875 0.063
R8374 GND.n3875 GND.n198 0.063
R8375 GND.n3863 GND.n3860 0.063
R8376 GND.n3863 GND.n3862 0.063
R8377 GND.n1877 GND.n1876 0.063
R8378 GND.n1744 GND.n1743 0.063
R8379 GND.n2486 GND.n2485 0.063
R8380 GND.n2623 GND.n2622 0.063
R8381 GND.n3040 GND.n3039 0.063
R8382 GND.n3297 GND.n3296 0.063
R8383 GND.n4220 GND.n4219 0.063
R8384 GND.n2064 GND 0.0590317
R8385 GND GND.n864 0.0590317
R8386 GND.n2256 GND 0.0590317
R8387 GND.n2826 GND 0.0590317
R8388 GND GND.n2898 0.0590317
R8389 GND.n3381 GND 0.0590317
R8390 GND.n3956 GND 0.0590317
R8391 GND GND.n4369 0.0590317
R8392 GND.n3545 GND.n3544 0.0532344
R8393 GND.n4370 GND 0.0512812
R8394 GND.n4221 GND.n4094 0.024
R8395 GND.n4222 GND.n4221 0.024
R8396 GND.n4092 GND.n58 0.024
R8397 GND.n4093 GND.n4092 0.024
R8398 GND.n3299 GND.n3298 0.024
R8399 GND.n3298 GND.n3173 0.024
R8400 GND.n3301 GND.n3172 0.024
R8401 GND.n3301 GND.n3300 0.024
R8402 GND.n3170 GND.n3043 0.024
R8403 GND.n3171 GND.n3170 0.024
R8404 GND.n3041 GND.n452 0.024
R8405 GND.n3042 GND.n3041 0.024
R8406 GND.n2621 GND.n2619 0.024
R8407 GND.n2621 GND.n2620 0.024
R8408 GND.n2617 GND.n2489 0.024
R8409 GND.n2618 GND.n2617 0.024
R8410 GND.n2487 GND.n565 0.024
R8411 GND.n2488 GND.n2487 0.024
R8412 GND.n1746 GND.n1745 0.024
R8413 GND.n1745 GND.n1618 0.024
R8414 GND.n1873 GND.n1872 0.024
R8415 GND.n1872 GND.n1747 0.024
R8416 GND.n1875 GND.n1617 0.024
R8417 GND.n1875 GND.n1874 0.024
R8418 GND.n1615 GND.n894 0.024
R8419 GND.n1616 GND.n1615 0.024
R8420 GND.n1401 GND.n1399 0.024
R8421 GND.n1401 GND.n1400 0.024
R8422 GND.n1397 GND.n1269 0.024
R8423 GND.n1398 GND.n1397 0.024
R8424 GND.n1267 GND.n937 0.024
R8425 GND.n1268 GND.n1267 0.024
R8426 GND.n1073 GND.n1000 0.024
R8427 GND.n3783 GND.n3628 0.024
R8428 GND.n3784 GND.n3783 0.024
R8429 GND.n3788 GND.n3787 0.024
R8430 GND.n3789 GND.n3788 0.024
R8431 GND.n3793 GND.n3792 0.024
R8432 GND.n3794 GND.n3793 0.024
R8433 GND.n3798 GND.n3797 0.024
R8434 GND.n3799 GND.n3798 0.024
R8435 GND.n3803 GND.n3802 0.024
R8436 GND.n3804 GND.n3803 0.024
R8437 GND.n3808 GND.n3807 0.024
R8438 GND.n3809 GND.n3808 0.024
R8439 GND.n3813 GND.n3812 0.024
R8440 GND.n3814 GND.n3813 0.024
R8441 GND.n3818 GND.n3817 0.024
R8442 GND.n3819 GND.n3818 0.024
R8443 GND.n3823 GND.n3822 0.024
R8444 GND.n3824 GND.n3823 0.024
R8445 GND.n3828 GND.n3827 0.024
R8446 GND.n3829 GND.n3828 0.024
R8447 GND.n3833 GND.n3832 0.024
R8448 GND.n3834 GND.n3833 0.024
R8449 GND.n3838 GND.n3837 0.024
R8450 GND.n3839 GND.n3838 0.024
R8451 GND.n3843 GND.n3842 0.024
R8452 GND.n3844 GND.n3843 0.024
R8453 GND.n3848 GND.n3847 0.024
R8454 GND.n3849 GND.n3848 0.024
R8455 GND.n3853 GND.n3852 0.024
R8456 GND.n3854 GND.n3853 0.024
R8457 GND.n3873 GND.n3857 0.024
R8458 GND.n3873 GND.n3858 0.024
R8459 GND.n3869 GND.n3868 0.024
R8460 GND.n3868 GND.n3865 0.024
R8461 GND.n2 GND.n0 0.024
R8462 GND.n4375 GND.n0 0.024
R8463 GND.n4374 GND 0.024
R8464 GND.n3477 GND 0.0204394
R8465 GND.n3499 GND 0.0204394
R8466 GND.n3521 GND 0.0204394
R8467 GND.n3540 GND 0.0204394
R8468 GND.n3562 GND 0.0204394
R8469 GND.n3581 GND 0.0204394
R8470 GND.n3601 GND 0.0204394
R8471 GND.n258 GND 0.0204394
R8472 GND GND.n1165 0.0193492
R8473 GND.n1152 GND 0.0193492
R8474 GND GND.n1150 0.0193492
R8475 GND GND.n847 0.0193492
R8476 GND GND.n860 0.0193492
R8477 GND.n862 GND 0.0193492
R8478 GND GND.n2288 0.0193492
R8479 GND.n2275 GND 0.0193492
R8480 GND GND.n2273 0.0193492
R8481 GND.n2333 GND 0.0193492
R8482 GND.n2372 GND 0.0193492
R8483 GND.n2365 GND 0.0193492
R8484 GND GND.n2765 0.0193492
R8485 GND GND.n2778 0.0193492
R8486 GND.n2780 GND 0.0193492
R8487 GND GND.n3348 0.0193492
R8488 GND.n3367 GND 0.0193492
R8489 GND.n3378 GND 0.0193492
R8490 GND GND.n159 0.0193492
R8491 GND GND.n172 0.0193492
R8492 GND.n3958 GND 0.0193492
R8493 GND GND.n4330 0.0193492
R8494 GND.n4350 GND 0.0193492
R8495 GND GND.n4348 0.0193492
R8496 GND.n3631 GND.t434 0.0180781
R8497 GND.n3632 GND.t406 0.0180781
R8498 GND.n3633 GND.t442 0.0180781
R8499 GND.n3634 GND.t404 0.0180781
R8500 GND.n3635 GND.t436 0.0180781
R8501 GND.n3636 GND.t484 0.0180781
R8502 GND.n3637 GND.t456 0.0180781
R8503 GND.n3638 GND.t490 0.0180781
R8504 GND.n3639 GND.t410 0.0180781
R8505 GND.n3640 GND.t444 0.0180781
R8506 GND.n3641 GND.t454 0.0180781
R8507 GND.n3642 GND.t488 0.0180781
R8508 GND.n3643 GND.t476 0.0180781
R8509 GND.n3644 GND.t376 0.0180781
R8510 GND.n3645 GND.t480 0.0180781
R8511 GND.n3646 GND.t420 0.0180781
R8512 GND.n3680 GND.t486 0.0180781
R8513 GND.n3683 GND.t426 0.0180781
R8514 GND.n3686 GND.t496 0.0180781
R8515 GND.n3689 GND.t396 0.0180781
R8516 GND.n3692 GND.t494 0.0180781
R8517 GND.n3695 GND.t392 0.0180781
R8518 GND.n3698 GND.t498 0.0180781
R8519 GND.n3701 GND.t398 0.0180781
R8520 GND.n3704 GND.t450 0.0180781
R8521 GND.n3707 GND.t428 0.0180781
R8522 GND.n3710 GND.t462 0.0180781
R8523 GND.n3713 GND.t402 0.0180781
R8524 GND.n3716 GND.t482 0.0180781
R8525 GND.n3719 GND.t382 0.0180781
R8526 GND.n3722 GND.t418 0.0180781
R8527 GND.n3725 GND.t390 0.0180781
R8528 GND.n3728 GND.t468 0.0180781
R8529 GND.n3629 GND.t374 0.0180781
R8530 GND.n3734 GND.t422 0.0180781
R8531 GND.n3737 GND.t384 0.0180781
R8532 GND.n3740 GND.t430 0.0180781
R8533 GND.n3743 GND.t460 0.0180781
R8534 GND.n3746 GND.t492 0.0180781
R8535 GND.n3749 GND.t408 0.0180781
R8536 GND.n3752 GND.t372 0.0180781
R8537 GND.n3755 GND.t416 0.0180781
R8538 GND.n3758 GND.t464 0.0180781
R8539 GND.n3761 GND.t368 0.0180781
R8540 GND.n3764 GND.t370 0.0180781
R8541 GND.n3767 GND.t414 0.0180781
R8542 GND.n3770 GND.t388 0.0180781
R8543 GND.n3773 GND.t432 0.0180781
R8544 GND.n3776 GND.t400 0.0180781
R8545 GND.n3779 GND.t478 0.0180781
R8546 GND.n3783 GND.t386 0.0180781
R8547 GND.n3788 GND.t470 0.0180781
R8548 GND.n3793 GND.t412 0.0180781
R8549 GND.n3798 GND.t474 0.0180781
R8550 GND.n3803 GND.t466 0.0180781
R8551 GND.n3808 GND.t448 0.0180781
R8552 GND.n3813 GND.t380 0.0180781
R8553 GND.n3818 GND.t458 0.0180781
R8554 GND.n3823 GND.t452 0.0180781
R8555 GND.n3828 GND.t378 0.0180781
R8556 GND.n3833 GND.t440 0.0180781
R8557 GND.n3838 GND.t438 0.0180781
R8558 GND.n3843 GND.t502 0.0180781
R8559 GND.n3848 GND.t500 0.0180781
R8560 GND.n3853 GND.t424 0.0180781
R8561 GND.n3873 GND.t446 0.0180781
R8562 GND.n3868 GND.t394 0.0180781
R8563 GND.n0 GND.t472 0.0180781
R8564 GND.n4089 GND.n4088 0.0169286
R8565 GND.n4075 GND.n4074 0.0169286
R8566 GND.n3305 GND.n3304 0.0169286
R8567 GND.n393 GND.n392 0.0169286
R8568 GND.n3167 GND.n3166 0.0169286
R8569 GND.n3153 GND.n3152 0.0169286
R8570 GND.n2614 GND.n2613 0.0169286
R8571 GND.n2600 GND.n2599 0.0169286
R8572 GND.n1869 GND.n1868 0.0169286
R8573 GND.n1855 GND.n1854 0.0169286
R8574 GND.n1612 GND.n1611 0.0169286
R8575 GND.n1598 GND.n1597 0.0169286
R8576 GND.n1264 GND.n1263 0.0169286
R8577 GND.n1250 GND.n1249 0.0169286
R8578 GND.n1394 GND.n1393 0.0169286
R8579 GND.n1380 GND.n1379 0.0169286
R8580 GND.n1405 GND.n1404 0.0169286
R8581 GND.n1500 GND.n1499 0.0169286
R8582 GND.n1070 GND.n1069 0.0169286
R8583 GND.n1020 GND.n1019 0.0169286
R8584 GND.n1030 GND.n1029 0.0169286
R8585 GND.n1057 GND.n1056 0.0169286
R8586 GND.n1045 GND.n1044 0.0169286
R8587 GND.n1879 GND.n1878 0.0169286
R8588 GND.n1974 GND.n1973 0.0169286
R8589 GND.n1742 GND.n1741 0.0169286
R8590 GND.n1728 GND.n1727 0.0169286
R8591 GND.n2484 GND.n2483 0.0169286
R8592 GND.n2470 GND.n2469 0.0169286
R8593 GND.n2625 GND.n2624 0.0169286
R8594 GND.n2720 GND.n2719 0.0169286
R8595 GND.n3038 GND.n3037 0.0169286
R8596 GND.n3024 GND.n3023 0.0169286
R8597 GND.n3295 GND.n3294 0.0169286
R8598 GND.n3281 GND.n3280 0.0169286
R8599 GND.n4218 GND.n4217 0.0169286
R8600 GND.n4204 GND.n4203 0.0169286
R8601 GND.n4269 GND.n4268 0.0169286
R8602 GND.n4257 GND.n4256 0.0169286
R8603 GND.n4248 GND.n4247 0.0169286
R8604 GND.n4281 GND.n4280 0.0169286
R8605 GND.n4225 GND.n4224 0.0169286
R8606 GND.n3861 GND 0.0168043
R8607 GND GND.n4375 0.0140786
R8608 GND.t487 GND.n3630 0.01225
R8609 GND.n3731 GND.t375 0.01225
R8610 GND.t473 GND.n4372 0.01225
R8611 GND.t395 GND.n3859 0.01225
R8612 GND.t447 GND.n199 0.01225
R8613 GND.n202 GND.t425 0.01225
R8614 GND.n205 GND.t501 0.01225
R8615 GND.n208 GND.t503 0.01225
R8616 GND.n211 GND.t439 0.01225
R8617 GND.n214 GND.t441 0.01225
R8618 GND.n217 GND.t379 0.01225
R8619 GND.n220 GND.t453 0.01225
R8620 GND.n223 GND.t459 0.01225
R8621 GND.n226 GND.t381 0.01225
R8622 GND.n229 GND.t449 0.01225
R8623 GND.n232 GND.t467 0.01225
R8624 GND.n235 GND.t475 0.01225
R8625 GND.n238 GND.t413 0.01225
R8626 GND.n241 GND.t471 0.01225
R8627 GND.n3781 GND.t387 0.01225
R8628 GND.t387 GND.n242 0.01225
R8629 GND.n3861 GND 0.0122188
R8630 GND.n3546 GND.n3545 0.0102656
R8631 GND.n4053 GND.n4052 0.00929205
R8632 GND.n4059 GND.n4058 0.00929205
R8633 GND.n4006 GND.n4005 0.00929205
R8634 GND.n4037 GND.n4036 0.00929205
R8635 GND.n3315 GND.n3314 0.00929205
R8636 GND.n3325 GND.n3324 0.00929205
R8637 GND.n403 GND.n402 0.00929205
R8638 GND.n427 GND.n426 0.00929205
R8639 GND.n3131 GND.n3130 0.00929205
R8640 GND.n3137 GND.n3136 0.00929205
R8641 GND.n3084 GND.n3083 0.00929205
R8642 GND.n3115 GND.n3114 0.00929205
R8643 GND.n2578 GND.n2577 0.00929205
R8644 GND.n2584 GND.n2583 0.00929205
R8645 GND.n2531 GND.n2530 0.00929205
R8646 GND.n2562 GND.n2561 0.00929205
R8647 GND.n1833 GND.n1832 0.00929205
R8648 GND.n1839 GND.n1838 0.00929205
R8649 GND.n1786 GND.n1785 0.00929205
R8650 GND.n1817 GND.n1816 0.00929205
R8651 GND.n1576 GND.n1575 0.00929205
R8652 GND.n1582 GND.n1581 0.00929205
R8653 GND.n1529 GND.n1528 0.00929205
R8654 GND.n1560 GND.n1559 0.00929205
R8655 GND.n1228 GND.n1227 0.00929205
R8656 GND.n1234 GND.n1233 0.00929205
R8657 GND.n1181 GND.n1180 0.00929205
R8658 GND.n1212 GND.n1211 0.00929205
R8659 GND.n1358 GND.n1357 0.00929205
R8660 GND.n1364 GND.n1363 0.00929205
R8661 GND.n1311 GND.n1310 0.00929205
R8662 GND.n1342 GND.n1341 0.00929205
R8663 GND.n1514 GND.n1513 0.00929205
R8664 GND.n1507 GND.n1506 0.00929205
R8665 GND.n1434 GND.n1433 0.00929205
R8666 GND.n1482 GND.n1481 0.00929205
R8667 GND.n1988 GND.n1987 0.00929205
R8668 GND.n1981 GND.n1980 0.00929205
R8669 GND.n1908 GND.n1907 0.00929205
R8670 GND.n1956 GND.n1955 0.00929205
R8671 GND.n1706 GND.n1705 0.00929205
R8672 GND.n1712 GND.n1711 0.00929205
R8673 GND.n1659 GND.n1658 0.00929205
R8674 GND.n1690 GND.n1689 0.00929205
R8675 GND.n2448 GND.n2447 0.00929205
R8676 GND.n2454 GND.n2453 0.00929205
R8677 GND.n2401 GND.n2400 0.00929205
R8678 GND.n2432 GND.n2431 0.00929205
R8679 GND.n2734 GND.n2733 0.00929205
R8680 GND.n2727 GND.n2726 0.00929205
R8681 GND.n2654 GND.n2653 0.00929205
R8682 GND.n2702 GND.n2701 0.00929205
R8683 GND.n3002 GND.n3001 0.00929205
R8684 GND.n3008 GND.n3007 0.00929205
R8685 GND.n2955 GND.n2954 0.00929205
R8686 GND.n2986 GND.n2985 0.00929205
R8687 GND.n3259 GND.n3258 0.00929205
R8688 GND.n3265 GND.n3264 0.00929205
R8689 GND.n3212 GND.n3211 0.00929205
R8690 GND.n3243 GND.n3242 0.00929205
R8691 GND.n4182 GND.n4181 0.00929205
R8692 GND.n4188 GND.n4187 0.00929205
R8693 GND.n4135 GND.n4134 0.00929205
R8694 GND.n4166 GND.n4165 0.00929205
R8695 GND.t471 GND.n239 0.00476905
R8696 GND.t413 GND.n236 0.00476905
R8697 GND.t475 GND.n233 0.00476905
R8698 GND.t467 GND.n230 0.00476905
R8699 GND.t449 GND.n227 0.00476905
R8700 GND.t381 GND.n224 0.00476905
R8701 GND.t459 GND.n221 0.00476905
R8702 GND.t453 GND.n218 0.00476905
R8703 GND.t379 GND.n215 0.00476905
R8704 GND.t441 GND.n212 0.00476905
R8705 GND.t439 GND.n209 0.00476905
R8706 GND.t503 GND.n206 0.00476905
R8707 GND.t501 GND.n203 0.00476905
R8708 GND.t425 GND.n200 0.00476905
R8709 GND.n3872 GND.t447 0.00476905
R8710 GND.n3867 GND.t395 0.00476905
R8711 GND.n4373 GND.t473 0.00476905
R8712 GND.n3476 GND 0.00441667
R8713 GND.n3498 GND 0.00441667
R8714 GND.n3520 GND 0.00441667
R8715 GND.n3539 GND 0.00441667
R8716 GND.n3561 GND 0.00441667
R8717 GND.n3580 GND 0.00441667
R8718 GND.n3600 GND 0.00441667
R8719 GND.n257 GND 0.00441667
R8720 GND.n4223 GND 0.00441667
R8721 GND GND.n3476 0.00406061
R8722 GND GND.n3498 0.00406061
R8723 GND GND.n3520 0.00406061
R8724 GND GND.n3539 0.00406061
R8725 GND GND.n3561 0.00406061
R8726 GND GND.n3580 0.00406061
R8727 GND GND.n3600 0.00406061
R8728 GND GND.n257 0.00406061
R8729 GND GND.n4223 0.00406061
R8730 EN.t5 EN.t10 322.06
R8731 EN.n24 EN.t87 158.988
R8732 EN.n10 EN.t28 158.988
R8733 EN.n284 EN.t44 158.56
R8734 EN.n268 EN.t34 158.56
R8735 EN.n252 EN.t103 158.56
R8736 EN.n236 EN.t74 158.56
R8737 EN.n220 EN.t82 158.56
R8738 EN.n204 EN.t46 158.56
R8739 EN.n188 EN.t55 158.56
R8740 EN.n172 EN.t61 158.56
R8741 EN.n156 EN.t62 158.56
R8742 EN.n140 EN.t69 158.56
R8743 EN.n124 EN.t57 158.56
R8744 EN.n108 EN.t78 158.56
R8745 EN.n92 EN.t86 158.56
R8746 EN.n76 EN.t43 158.56
R8747 EN.n60 EN.t93 158.56
R8748 EN.n44 EN.t80 158.56
R8749 EN.t44 EN.n283 151.594
R8750 EN.t34 EN.n267 151.594
R8751 EN.t103 EN.n251 151.594
R8752 EN.t74 EN.n235 151.594
R8753 EN.t82 EN.n219 151.594
R8754 EN.t46 EN.n203 151.594
R8755 EN.t55 EN.n187 151.594
R8756 EN.t61 EN.n171 151.594
R8757 EN.t62 EN.n155 151.594
R8758 EN.t69 EN.n139 151.594
R8759 EN.t57 EN.n123 151.594
R8760 EN.t78 EN.n107 151.594
R8761 EN.t86 EN.n91 151.594
R8762 EN.t43 EN.n75 151.594
R8763 EN.t93 EN.n59 151.594
R8764 EN.t80 EN.n43 151.594
R8765 EN.n34 EN.t89 150.56
R8766 EN.n30 EN.t5 150.56
R8767 EN.n15 EN.t23 150.293
R8768 EN.t10 EN.n29 150.293
R8769 EN.n276 EN.t26 150.273
R8770 EN.n272 EN.t40 150.273
R8771 EN.n260 EN.t33 150.273
R8772 EN.n256 EN.t45 150.273
R8773 EN.n244 EN.t13 150.273
R8774 EN.n240 EN.t31 150.273
R8775 EN.n228 EN.t56 150.273
R8776 EN.n224 EN.t81 150.273
R8777 EN.n212 EN.t63 150.273
R8778 EN.n208 EN.t88 150.273
R8779 EN.n196 EN.t105 150.273
R8780 EN.n192 EN.t19 150.273
R8781 EN.n180 EN.t49 150.273
R8782 EN.n176 EN.t60 150.273
R8783 EN.n164 EN.t51 150.273
R8784 EN.n160 EN.t68 150.273
R8785 EN.n148 EN.t95 150.273
R8786 EN.n144 EN.t12 150.273
R8787 EN.n132 EN.t54 150.273
R8788 EN.n128 EN.t77 150.273
R8789 EN.n116 EN.t75 150.273
R8790 EN.n112 EN.t106 150.273
R8791 EN.n100 EN.t59 150.273
R8792 EN.n96 EN.t85 150.273
R8793 EN.n84 EN.t83 150.273
R8794 EN.n80 EN.t3 150.273
R8795 EN.n68 EN.t7 150.273
R8796 EN.n64 EN.t30 150.273
R8797 EN.n52 EN.t72 150.273
R8798 EN.n48 EN.t102 150.273
R8799 EN.t87 EN.n23 150.273
R8800 EN.t28 EN.n9 150.273
R8801 EN.n5 EN.t99 150.273
R8802 EN.n1 EN.t17 150.273
R8803 EN.n9 EN.t36 74.951
R8804 EN.n275 EN.t64 74.4891
R8805 EN.n271 EN.t90 74.4891
R8806 EN.n259 EN.t50 74.4891
R8807 EN.n255 EN.t67 74.4891
R8808 EN.n243 EN.t24 74.4891
R8809 EN.n239 EN.t39 74.4891
R8810 EN.n227 EN.t70 74.4891
R8811 EN.n223 EN.t97 74.4891
R8812 EN.n211 EN.t79 74.4891
R8813 EN.n207 EN.t0 74.4891
R8814 EN.n195 EN.t94 74.4891
R8815 EN.n191 EN.t11 74.4891
R8816 EN.n179 EN.t53 74.4891
R8817 EN.n175 EN.t76 74.4891
R8818 EN.n163 EN.t14 74.4891
R8819 EN.n159 EN.t32 74.4891
R8820 EN.n147 EN.t58 74.4891
R8821 EN.n143 EN.t84 74.4891
R8822 EN.n131 EN.t65 74.4891
R8823 EN.n127 EN.t91 74.4891
R8824 EN.n115 EN.t6 74.4891
R8825 EN.n111 EN.t29 74.4891
R8826 EN.n99 EN.t71 74.4891
R8827 EN.n95 EN.t101 74.4891
R8828 EN.n83 EN.t98 74.4891
R8829 EN.n79 EN.t16 74.4891
R8830 EN.n67 EN.t21 74.4891
R8831 EN.n63 EN.t38 74.4891
R8832 EN.n51 EN.t1 74.4891
R8833 EN.n47 EN.t20 74.4891
R8834 EN.n4 EN.t73 74.4891
R8835 EN.n0 EN.t104 74.4891
R8836 EN.n21 EN.t42 73.6406
R8837 EN.n283 EN.t35 73.6304
R8838 EN.n267 EN.t41 73.6304
R8839 EN.n251 EN.t52 73.6304
R8840 EN.n235 EN.t25 73.6304
R8841 EN.n219 EN.t15 73.6304
R8842 EN.n203 EN.t2 73.6304
R8843 EN.n187 EN.t96 73.6304
R8844 EN.n171 EN.t107 73.6304
R8845 EN.n155 EN.t27 73.6304
R8846 EN.n139 EN.t4 73.6304
R8847 EN.n123 EN.t9 73.6304
R8848 EN.n107 EN.t8 73.6304
R8849 EN.n91 EN.t18 73.6304
R8850 EN.n75 EN.t100 73.6304
R8851 EN.n59 EN.t22 73.6304
R8852 EN.n43 EN.t37 73.6304
R8853 EN.n35 EN.t66 73.6304
R8854 EN.n31 EN.t92 73.6304
R8855 EN.n17 EN.t48 73.6304
R8856 EN.n12 EN.t47 73.6304
R8857 EN.n46 EN 39.9701
R8858 EN.n45 EN 38.0684
R8859 EN.n62 EN 37.1783
R8860 EN.n61 EN 35.5304
R8861 EN.n78 EN 34.3865
R8862 EN.n77 EN 32.9924
R8863 EN.n94 EN 31.5947
R8864 EN.n93 EN 30.4544
R8865 EN.n110 EN 28.8029
R8866 EN.n109 EN 27.9164
R8867 EN.n126 EN 26.0111
R8868 EN.n125 EN 25.3784
R8869 EN.n142 EN 23.2193
R8870 EN.n141 EN 22.8404
R8871 EN.n158 EN 20.4275
R8872 EN.n157 EN 20.3024
R8873 EN.n173 EN 17.7644
R8874 EN.n174 EN 17.6357
R8875 EN.n279 EN.n274 15.5222
R8876 EN.n263 EN.n258 15.5222
R8877 EN.n247 EN.n242 15.5222
R8878 EN.n231 EN.n226 15.5222
R8879 EN.n215 EN.n210 15.5222
R8880 EN.n199 EN.n194 15.5222
R8881 EN.n183 EN.n178 15.5222
R8882 EN.n167 EN.n162 15.5222
R8883 EN.n151 EN.n146 15.5222
R8884 EN.n135 EN.n130 15.5222
R8885 EN.n119 EN.n114 15.5222
R8886 EN.n103 EN.n98 15.5222
R8887 EN.n87 EN.n82 15.5222
R8888 EN.n71 EN.n66 15.5222
R8889 EN.n55 EN.n50 15.5222
R8890 EN.n26 EN.n20 15.5222
R8891 EN.n38 EN.n33 15.5222
R8892 EN.n8 EN.n3 15.5222
R8893 EN.n189 EN 15.2264
R8894 EN.n190 EN 14.8439
R8895 EN.n205 EN 12.6884
R8896 EN.n206 EN 12.0521
R8897 EN.n221 EN 10.1504
R8898 EN.n222 EN 9.26028
R8899 EN.n280 EN.n279 8.24202
R8900 EN.n264 EN.n263 8.24202
R8901 EN.n248 EN.n247 8.24202
R8902 EN.n232 EN.n231 8.24202
R8903 EN.n216 EN.n215 8.24202
R8904 EN.n200 EN.n199 8.24202
R8905 EN.n184 EN.n183 8.24202
R8906 EN.n168 EN.n167 8.24202
R8907 EN.n152 EN.n151 8.24202
R8908 EN.n136 EN.n135 8.24202
R8909 EN.n120 EN.n119 8.24202
R8910 EN.n104 EN.n103 8.24202
R8911 EN.n88 EN.n87 8.24202
R8912 EN.n72 EN.n71 8.24202
R8913 EN.n56 EN.n55 8.24202
R8914 EN.n26 EN 7.85707
R8915 EN.n39 EN.n38 7.83713
R8916 EN.n237 EN 7.61236
R8917 EN.n238 EN 6.46848
R8918 EN.n253 EN 5.07436
R8919 EN.n40 EN.n39 4.9286
R8920 EN.n279 EN.n278 4.5005
R8921 EN.n263 EN.n262 4.5005
R8922 EN.n247 EN.n246 4.5005
R8923 EN.n231 EN.n230 4.5005
R8924 EN.n215 EN.n214 4.5005
R8925 EN.n199 EN.n198 4.5005
R8926 EN.n183 EN.n182 4.5005
R8927 EN.n167 EN.n166 4.5005
R8928 EN.n151 EN.n150 4.5005
R8929 EN.n135 EN.n134 4.5005
R8930 EN.n119 EN.n118 4.5005
R8931 EN.n103 EN.n102 4.5005
R8932 EN.n87 EN.n86 4.5005
R8933 EN.n71 EN.n70 4.5005
R8934 EN.n55 EN.n54 4.5005
R8935 EN.n27 EN.n26 4.5005
R8936 EN.n38 EN.n37 4.5005
R8937 EN.n8 EN.n7 4.5005
R8938 EN.n40 EN.n8 4.42713
R8939 EN.n41 EN.n40 3.7628
R8940 EN.n254 EN 3.67668
R8941 EN.n269 EN 2.53636
R8942 EN.n46 EN.n45 1.90557
R8943 EN.n62 EN.n61 1.90557
R8944 EN.n78 EN.n77 1.90557
R8945 EN.n94 EN.n93 1.90557
R8946 EN.n110 EN.n109 1.90557
R8947 EN.n126 EN.n125 1.90557
R8948 EN.n142 EN.n141 1.90557
R8949 EN.n158 EN.n157 1.90557
R8950 EN.n174 EN.n173 1.90557
R8951 EN.n190 EN.n189 1.90557
R8952 EN.n206 EN.n205 1.90557
R8953 EN.n222 EN.n221 1.90557
R8954 EN.n238 EN.n237 1.90557
R8955 EN.n254 EN.n253 1.90557
R8956 EN.n270 EN.n269 1.90557
R8957 EN.n22 EN.n21 1.19615
R8958 EN.n34 EN 1.09561
R8959 EN.n16 EN 1.09561
R8960 EN.n28 EN 1.09561
R8961 EN.n30 EN 1.09561
R8962 EN.n270 EN 0.884883
R8963 EN.n36 EN.n35 0.859196
R8964 EN.n32 EN.n31 0.859196
R8965 EN.n19 EN.n18 0.796696
R8966 EN.n14 EN.n13 0.796696
R8967 EN.n25 EN.n24 0.783833
R8968 EN.n11 EN.n10 0.783833
R8969 EN.n42 EN.n41 0.783833
R8970 EN.n58 EN.n57 0.783833
R8971 EN.n74 EN.n73 0.783833
R8972 EN.n90 EN.n89 0.783833
R8973 EN.n106 EN.n105 0.783833
R8974 EN.n122 EN.n121 0.783833
R8975 EN.n138 EN.n137 0.783833
R8976 EN.n154 EN.n153 0.783833
R8977 EN.n170 EN.n169 0.783833
R8978 EN.n186 EN.n185 0.783833
R8979 EN.n202 EN.n201 0.783833
R8980 EN.n218 EN.n217 0.783833
R8981 EN.n234 EN.n233 0.783833
R8982 EN.n250 EN.n249 0.783833
R8983 EN.n266 EN.n265 0.783833
R8984 EN.n282 EN.n281 0.783833
R8985 EN.n24 EN 0.716182
R8986 EN.n10 EN 0.716182
R8987 EN.n41 EN 0.716182
R8988 EN.n57 EN 0.716182
R8989 EN.n73 EN 0.716182
R8990 EN.n89 EN 0.716182
R8991 EN.n105 EN 0.716182
R8992 EN.n121 EN 0.716182
R8993 EN.n137 EN 0.716182
R8994 EN.n153 EN 0.716182
R8995 EN.n169 EN 0.716182
R8996 EN.n185 EN 0.716182
R8997 EN.n201 EN 0.716182
R8998 EN.n217 EN 0.716182
R8999 EN.n233 EN 0.716182
R9000 EN.n249 EN 0.716182
R9001 EN.n265 EN 0.716182
R9002 EN.n281 EN 0.716182
R9003 EN.n36 EN 0.662609
R9004 EN.n19 EN 0.662609
R9005 EN.n14 EN 0.662609
R9006 EN.n32 EN 0.662609
R9007 EN.n275 EN 0.524957
R9008 EN.n271 EN 0.524957
R9009 EN.n259 EN 0.524957
R9010 EN.n255 EN 0.524957
R9011 EN.n243 EN 0.524957
R9012 EN.n239 EN 0.524957
R9013 EN.n227 EN 0.524957
R9014 EN.n223 EN 0.524957
R9015 EN.n211 EN 0.524957
R9016 EN.n207 EN 0.524957
R9017 EN.n195 EN 0.524957
R9018 EN.n191 EN 0.524957
R9019 EN.n179 EN 0.524957
R9020 EN.n175 EN 0.524957
R9021 EN.n163 EN 0.524957
R9022 EN.n159 EN 0.524957
R9023 EN.n147 EN 0.524957
R9024 EN.n143 EN 0.524957
R9025 EN.n131 EN 0.524957
R9026 EN.n127 EN 0.524957
R9027 EN.n115 EN 0.524957
R9028 EN.n111 EN 0.524957
R9029 EN.n99 EN 0.524957
R9030 EN.n95 EN 0.524957
R9031 EN.n83 EN 0.524957
R9032 EN.n79 EN 0.524957
R9033 EN.n67 EN 0.524957
R9034 EN.n63 EN 0.524957
R9035 EN.n51 EN 0.524957
R9036 EN.n47 EN 0.524957
R9037 EN.n4 EN 0.524957
R9038 EN.n0 EN 0.524957
R9039 EN.n15 EN 0.447191
R9040 EN.n29 EN 0.447191
R9041 EN.n277 EN.n276 0.288543
R9042 EN.n273 EN.n272 0.288543
R9043 EN.n261 EN.n260 0.288543
R9044 EN.n257 EN.n256 0.288543
R9045 EN.n245 EN.n244 0.288543
R9046 EN.n241 EN.n240 0.288543
R9047 EN.n229 EN.n228 0.288543
R9048 EN.n225 EN.n224 0.288543
R9049 EN.n213 EN.n212 0.288543
R9050 EN.n209 EN.n208 0.288543
R9051 EN.n197 EN.n196 0.288543
R9052 EN.n193 EN.n192 0.288543
R9053 EN.n181 EN.n180 0.288543
R9054 EN.n177 EN.n176 0.288543
R9055 EN.n165 EN.n164 0.288543
R9056 EN.n161 EN.n160 0.288543
R9057 EN.n149 EN.n148 0.288543
R9058 EN.n145 EN.n144 0.288543
R9059 EN.n133 EN.n132 0.288543
R9060 EN.n129 EN.n128 0.288543
R9061 EN.n117 EN.n116 0.288543
R9062 EN.n113 EN.n112 0.288543
R9063 EN.n101 EN.n100 0.288543
R9064 EN.n97 EN.n96 0.288543
R9065 EN.n85 EN.n84 0.288543
R9066 EN.n81 EN.n80 0.288543
R9067 EN.n69 EN.n68 0.288543
R9068 EN.n65 EN.n64 0.288543
R9069 EN.n53 EN.n52 0.288543
R9070 EN.n49 EN.n48 0.288543
R9071 EN.n6 EN.n5 0.288543
R9072 EN.n2 EN.n1 0.288543
R9073 EN.n277 EN 0.252453
R9074 EN.n273 EN 0.252453
R9075 EN.n261 EN 0.252453
R9076 EN.n257 EN 0.252453
R9077 EN.n245 EN 0.252453
R9078 EN.n241 EN 0.252453
R9079 EN.n229 EN 0.252453
R9080 EN.n225 EN 0.252453
R9081 EN.n213 EN 0.252453
R9082 EN.n209 EN 0.252453
R9083 EN.n197 EN 0.252453
R9084 EN.n193 EN 0.252453
R9085 EN.n181 EN 0.252453
R9086 EN.n177 EN 0.252453
R9087 EN.n165 EN 0.252453
R9088 EN.n161 EN 0.252453
R9089 EN.n149 EN 0.252453
R9090 EN.n145 EN 0.252453
R9091 EN.n133 EN 0.252453
R9092 EN.n129 EN 0.252453
R9093 EN.n117 EN 0.252453
R9094 EN.n113 EN 0.252453
R9095 EN.n101 EN 0.252453
R9096 EN.n97 EN 0.252453
R9097 EN.n85 EN 0.252453
R9098 EN.n81 EN 0.252453
R9099 EN.n69 EN 0.252453
R9100 EN.n65 EN 0.252453
R9101 EN.n53 EN 0.252453
R9102 EN.n49 EN 0.252453
R9103 EN.n6 EN 0.252453
R9104 EN.n2 EN 0.252453
R9105 EN.n16 EN.n15 0.226043
R9106 EN.n29 EN.n28 0.226043
R9107 EN.n21 EN 0.217464
R9108 EN.n22 EN 0.1255
R9109 EN.n18 EN 0.1255
R9110 EN.n13 EN 0.1255
R9111 EN.n283 EN 0.063
R9112 EN.n276 EN 0.063
R9113 EN.n278 EN.n275 0.063
R9114 EN.n278 EN.n277 0.063
R9115 EN.n272 EN 0.063
R9116 EN.n274 EN.n271 0.063
R9117 EN.n274 EN.n273 0.063
R9118 EN.n267 EN 0.063
R9119 EN.n260 EN 0.063
R9120 EN.n262 EN.n259 0.063
R9121 EN.n262 EN.n261 0.063
R9122 EN.n256 EN 0.063
R9123 EN.n258 EN.n255 0.063
R9124 EN.n258 EN.n257 0.063
R9125 EN.n251 EN 0.063
R9126 EN.n244 EN 0.063
R9127 EN.n246 EN.n243 0.063
R9128 EN.n246 EN.n245 0.063
R9129 EN.n240 EN 0.063
R9130 EN.n242 EN.n239 0.063
R9131 EN.n242 EN.n241 0.063
R9132 EN.n235 EN 0.063
R9133 EN.n228 EN 0.063
R9134 EN.n230 EN.n227 0.063
R9135 EN.n230 EN.n229 0.063
R9136 EN.n224 EN 0.063
R9137 EN.n226 EN.n223 0.063
R9138 EN.n226 EN.n225 0.063
R9139 EN.n219 EN 0.063
R9140 EN.n212 EN 0.063
R9141 EN.n214 EN.n211 0.063
R9142 EN.n214 EN.n213 0.063
R9143 EN.n208 EN 0.063
R9144 EN.n210 EN.n207 0.063
R9145 EN.n210 EN.n209 0.063
R9146 EN.n203 EN 0.063
R9147 EN.n196 EN 0.063
R9148 EN.n198 EN.n195 0.063
R9149 EN.n198 EN.n197 0.063
R9150 EN.n192 EN 0.063
R9151 EN.n194 EN.n191 0.063
R9152 EN.n194 EN.n193 0.063
R9153 EN.n187 EN 0.063
R9154 EN.n180 EN 0.063
R9155 EN.n182 EN.n179 0.063
R9156 EN.n182 EN.n181 0.063
R9157 EN.n176 EN 0.063
R9158 EN.n178 EN.n175 0.063
R9159 EN.n178 EN.n177 0.063
R9160 EN.n171 EN 0.063
R9161 EN.n164 EN 0.063
R9162 EN.n166 EN.n163 0.063
R9163 EN.n166 EN.n165 0.063
R9164 EN.n160 EN 0.063
R9165 EN.n162 EN.n159 0.063
R9166 EN.n162 EN.n161 0.063
R9167 EN.n155 EN 0.063
R9168 EN.n148 EN 0.063
R9169 EN.n150 EN.n147 0.063
R9170 EN.n150 EN.n149 0.063
R9171 EN.n144 EN 0.063
R9172 EN.n146 EN.n143 0.063
R9173 EN.n146 EN.n145 0.063
R9174 EN.n139 EN 0.063
R9175 EN.n132 EN 0.063
R9176 EN.n134 EN.n131 0.063
R9177 EN.n134 EN.n133 0.063
R9178 EN.n128 EN 0.063
R9179 EN.n130 EN.n127 0.063
R9180 EN.n130 EN.n129 0.063
R9181 EN.n123 EN 0.063
R9182 EN.n116 EN 0.063
R9183 EN.n118 EN.n115 0.063
R9184 EN.n118 EN.n117 0.063
R9185 EN.n112 EN 0.063
R9186 EN.n114 EN.n111 0.063
R9187 EN.n114 EN.n113 0.063
R9188 EN.n107 EN 0.063
R9189 EN.n100 EN 0.063
R9190 EN.n102 EN.n99 0.063
R9191 EN.n102 EN.n101 0.063
R9192 EN.n96 EN 0.063
R9193 EN.n98 EN.n95 0.063
R9194 EN.n98 EN.n97 0.063
R9195 EN.n91 EN 0.063
R9196 EN.n84 EN 0.063
R9197 EN.n86 EN.n83 0.063
R9198 EN.n86 EN.n85 0.063
R9199 EN.n80 EN 0.063
R9200 EN.n82 EN.n79 0.063
R9201 EN.n82 EN.n81 0.063
R9202 EN.n75 EN 0.063
R9203 EN.n68 EN 0.063
R9204 EN.n70 EN.n67 0.063
R9205 EN.n70 EN.n69 0.063
R9206 EN.n64 EN 0.063
R9207 EN.n66 EN.n63 0.063
R9208 EN.n66 EN.n65 0.063
R9209 EN.n59 EN 0.063
R9210 EN.n52 EN 0.063
R9211 EN.n54 EN.n51 0.063
R9212 EN.n54 EN.n53 0.063
R9213 EN.n48 EN 0.063
R9214 EN.n50 EN.n47 0.063
R9215 EN.n50 EN.n49 0.063
R9216 EN.n43 EN 0.063
R9217 EN.n35 EN 0.063
R9218 EN.n37 EN.n34 0.063
R9219 EN.n37 EN.n36 0.063
R9220 EN.n31 EN 0.063
R9221 EN.n20 EN.n16 0.063
R9222 EN.n20 EN.n19 0.063
R9223 EN.n28 EN.n27 0.063
R9224 EN.n27 EN.n14 0.063
R9225 EN.n33 EN.n30 0.063
R9226 EN.n33 EN.n32 0.063
R9227 EN.n9 EN 0.063
R9228 EN.n5 EN 0.063
R9229 EN.n7 EN.n4 0.063
R9230 EN.n7 EN.n6 0.063
R9231 EN.n1 EN 0.063
R9232 EN.n3 EN.n0 0.063
R9233 EN.n3 EN.n2 0.063
R9234 EN.n45 EN.n44 0.024
R9235 EN.n56 EN.n46 0.024
R9236 EN.n57 EN.n56 0.024
R9237 EN.n61 EN.n60 0.024
R9238 EN.n72 EN.n62 0.024
R9239 EN.n73 EN.n72 0.024
R9240 EN.n77 EN.n76 0.024
R9241 EN.n88 EN.n78 0.024
R9242 EN.n89 EN.n88 0.024
R9243 EN.n93 EN.n92 0.024
R9244 EN.n104 EN.n94 0.024
R9245 EN.n105 EN.n104 0.024
R9246 EN.n109 EN.n108 0.024
R9247 EN.n120 EN.n110 0.024
R9248 EN.n121 EN.n120 0.024
R9249 EN.n125 EN.n124 0.024
R9250 EN.n136 EN.n126 0.024
R9251 EN.n137 EN.n136 0.024
R9252 EN.n141 EN.n140 0.024
R9253 EN.n152 EN.n142 0.024
R9254 EN.n153 EN.n152 0.024
R9255 EN.n157 EN.n156 0.024
R9256 EN.n168 EN.n158 0.024
R9257 EN.n169 EN.n168 0.024
R9258 EN.n173 EN.n172 0.024
R9259 EN.n184 EN.n174 0.024
R9260 EN.n185 EN.n184 0.024
R9261 EN.n189 EN.n188 0.024
R9262 EN.n200 EN.n190 0.024
R9263 EN.n201 EN.n200 0.024
R9264 EN.n205 EN.n204 0.024
R9265 EN.n216 EN.n206 0.024
R9266 EN.n217 EN.n216 0.024
R9267 EN.n221 EN.n220 0.024
R9268 EN.n232 EN.n222 0.024
R9269 EN.n233 EN.n232 0.024
R9270 EN.n237 EN.n236 0.024
R9271 EN.n248 EN.n238 0.024
R9272 EN.n249 EN.n248 0.024
R9273 EN.n253 EN.n252 0.024
R9274 EN.n264 EN.n254 0.024
R9275 EN.n265 EN.n264 0.024
R9276 EN.n269 EN.n268 0.024
R9277 EN.n280 EN.n270 0.024
R9278 EN.n281 EN.n280 0.024
R9279 EN EN.n284 0.0218636
R9280 EN.n23 EN.n22 0.0216397
R9281 EN.n23 EN 0.0216397
R9282 EN.n39 EN 0.0204394
R9283 EN.n44 EN 0.0204394
R9284 EN.n60 EN 0.0204394
R9285 EN.n76 EN 0.0204394
R9286 EN.n92 EN 0.0204394
R9287 EN.n108 EN 0.0204394
R9288 EN.n124 EN 0.0204394
R9289 EN.n140 EN 0.0204394
R9290 EN.n156 EN 0.0204394
R9291 EN.n172 EN 0.0204394
R9292 EN.n188 EN 0.0204394
R9293 EN.n204 EN 0.0204394
R9294 EN.n220 EN 0.0204394
R9295 EN.n236 EN 0.0204394
R9296 EN.n252 EN 0.0204394
R9297 EN.n268 EN 0.0204394
R9298 EN.n284 EN 0.0204394
R9299 EN.n18 EN.n17 0.0107679
R9300 EN.n17 EN 0.0107679
R9301 EN.n13 EN.n12 0.0107679
R9302 EN.n12 EN 0.0107679
R9303 EN.n25 EN 0.00441667
R9304 EN.n11 EN 0.00441667
R9305 EN.n42 EN 0.00441667
R9306 EN.n58 EN 0.00441667
R9307 EN.n74 EN 0.00441667
R9308 EN.n90 EN 0.00441667
R9309 EN.n106 EN 0.00441667
R9310 EN.n122 EN 0.00441667
R9311 EN.n138 EN 0.00441667
R9312 EN.n154 EN 0.00441667
R9313 EN.n170 EN 0.00441667
R9314 EN.n186 EN 0.00441667
R9315 EN.n202 EN 0.00441667
R9316 EN.n218 EN 0.00441667
R9317 EN.n234 EN 0.00441667
R9318 EN.n250 EN 0.00441667
R9319 EN.n266 EN 0.00441667
R9320 EN.n282 EN 0.00441667
R9321 EN EN.n25 0.00406061
R9322 EN EN.n11 0.00406061
R9323 EN EN.n42 0.00406061
R9324 EN EN.n58 0.00406061
R9325 EN EN.n74 0.00406061
R9326 EN EN.n90 0.00406061
R9327 EN EN.n106 0.00406061
R9328 EN EN.n122 0.00406061
R9329 EN EN.n138 0.00406061
R9330 EN EN.n154 0.00406061
R9331 EN EN.n170 0.00406061
R9332 EN EN.n186 0.00406061
R9333 EN EN.n202 0.00406061
R9334 EN EN.n218 0.00406061
R9335 EN EN.n234 0.00406061
R9336 EN EN.n250 0.00406061
R9337 EN EN.n266 0.00406061
R9338 EN EN.n282 0.00406061
R9339 Q0.n8 Q0.t3 169.46
R9340 Q0.n10 Q0.t0 167.809
R9341 Q0.n8 Q0.t2 167.809
R9342 Q0.n16 Q0.t8 158.565
R9343 Q0.n2 Q0.t4 150.543
R9344 Q0.n0 Q0.t7 150.543
R9345 Q0.t8 Q0.n15 150.293
R9346 Q0.n2 Q0.t6 74.4613
R9347 Q0.n0 Q0.t9 74.4613
R9348 Q0.n13 Q0.t5 73.6304
R9349 Q0.n6 Q0.t1 60.3809
R9350 Q0.n5 Q0.n4 12.0647
R9351 Q0.n9 Q0.n8 11.4489
R9352 Q0.n17 Q0.n5 10.1791
R9353 Q0.n5 Q0 9.25452
R9354 Q0.n11 Q0.n10 8.21389
R9355 Q0 Q0.n16 5.41669
R9356 Q0.n7 Q0.n6 1.64452
R9357 Q0.n15 Q0.n14 1.19615
R9358 Q0.n1 Q0 0.984196
R9359 Q0.n6 Q0 0.848156
R9360 Q0.n3 Q0.n2 0.747783
R9361 Q0.n1 Q0.n0 0.747783
R9362 Q0.n3 Q0 0.582531
R9363 Q0.n15 Q0 0.447191
R9364 Q0.n12 Q0.n11 0.425067
R9365 Q0.n11 Q0 0.39003
R9366 Q0.n10 Q0.n9 0.280391
R9367 Q0.n9 Q0 0.200143
R9368 Q0.n14 Q0 0.1255
R9369 Q0.n7 Q0 0.1255
R9370 Q0 Q0.n7 0.063
R9371 Q0.n2 Q0 0.063
R9372 Q0.n4 Q0.n1 0.063
R9373 Q0.n4 Q0.n3 0.063
R9374 Q0.n16 Q0 0.0204394
R9375 Q0.n14 Q0.n13 0.0107679
R9376 Q0.n13 Q0 0.0107679
R9377 Q0.n12 Q0 0.00441667
R9378 Q0 Q0.n12 0.00406061
R9379 Q0.n17 Q0 0.00128333
R9380 Q0.n17 Q0 0.00121212
R9381 CDAC_v3_0.switch_8.Z.n0 CDAC_v3_0.switch_8.Z.t4 168.075
R9382 CDAC_v3_0.switch_8.Z.n0 CDAC_v3_0.switch_8.Z.t1 168.075
R9383 CDAC_v3_0.switch_8.Z.n3 CDAC_v3_0.switch_8.Z.t2 65.4994
R9384 CDAC_v3_0.switch_8.Z.n5 CDAC_v3_0.switch_8.Z.t0 60.6851
R9385 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_8.Z.t3 60.6226
R9386 CDAC_v3_0.switch_8.Z.n2 CDAC_v3_0.switch_8.Z.n1 1.34289
R9387 CDAC_v3_0.switch_8.Z.n2 CDAC_v3_0.switch_8.Z 0.42713
R9388 CDAC_v3_0.switch_8.Z.n4 CDAC_v3_0.switch_8.Z 0.182141
R9389 CDAC_v3_0.switch_8.Z.n1 CDAC_v3_0.switch_8.Z 0.178175
R9390 CDAC_v3_0.switch_8.Z.n5 CDAC_v3_0.switch_8.Z.n4 0.128217
R9391 CDAC_v3_0.switch_8.Z.n5 CDAC_v3_0.switch_8.Z 0.1255
R9392 CDAC_v3_0.switch_8.Z.n3 CDAC_v3_0.switch_8.Z.n2 0.063
R9393 CDAC_v3_0.switch_8.Z.n4 CDAC_v3_0.switch_8.Z.n3 0.063
R9394 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_8.Z.n5 0.063
R9395 CDAC_v3_0.switch_8.Z.n1 CDAC_v3_0.switch_8.Z.n0 0.0130546
R9396 VDD.n7318 VDD.n7317 55259.3
R9397 VDD.n7318 VDD.n7316 49126.7
R9398 VDD.n7324 VDD.n7317 32898.4
R9399 VDD.n7325 VDD.n7324 29988.1
R9400 VDD.n7326 VDD.n7325 29374.8
R9401 VDD.n7320 VDD.n7319 27016.6
R9402 VDD.n7326 VDD.n7316 25484.7
R9403 VDD.n7319 VDD.n7313 24146.4
R9404 VDD.n7323 VDD.n7320 16939.4
R9405 VDD.n7323 VDD.n7315 15719.7
R9406 VDD.n7327 VDD.n7315 15072.6
R9407 VDD.n7327 VDD.n7313 13411.9
R9408 VDD.n7293 VDD.n7284 12650.1
R9409 VDD.n7293 VDD.n7285 12650.1
R9410 VDD.n7289 VDD.n7284 12650.1
R9411 VDD.n7302 VDD.n7299 10684.6
R9412 VDD.n7307 VDD.n7282 10684.6
R9413 VDD.n7306 VDD.n7282 10684.6
R9414 VDD.n7296 VDD.n7281 10167.6
R9415 VDD.n7297 VDD.n7296 10167.6
R9416 VDD.n7321 VDD.n7312 6073.28
R9417 VDD.n7329 VDD.n7312 5168.82
R9418 VDD.n7322 VDD.n7321 4059.29
R9419 VDD.n7322 VDD.n7314 3849.04
R9420 VDD.n7328 VDD.n7314 3690.92
R9421 VDD.n7329 VDD.n7328 2993.95
R9422 VDD.n7291 VDD.n7290 2427.48
R9423 VDD.n7292 VDD.n7291 2427.48
R9424 VDD.n7290 VDD.n7287 2349.78
R9425 VDD.n7292 VDD.n7287 2349.78
R9426 VDD.n7288 VDD.n7285 2128.85
R9427 VDD.n7305 VDD.n7280 2051.01
R9428 VDD.n7303 VDD.n7298 2051.01
R9429 VDD.n7308 VDD.n7280 1973.31
R9430 VDD.n7298 VDD.n7279 1973.31
R9431 VDD.n7309 VDD.n7278 1952
R9432 VDD.n7304 VDD.n7278 1952
R9433 VDD.n402 VDD.n187 1084.97
R9434 VDD.n402 VDD.n188 1084.97
R9435 VDD.n377 VDD.n188 1084.97
R9436 VDD.n377 VDD.n187 1084.97
R9437 VDD.n195 VDD.n194 1084.97
R9438 VDD.n394 VDD.n195 1084.97
R9439 VDD.n395 VDD.n394 1084.97
R9440 VDD.n395 VDD.n194 1084.97
R9441 VDD.n239 VDD.n176 1084.97
R9442 VDD.n240 VDD.n176 1084.97
R9443 VDD.n244 VDD.n240 1084.97
R9444 VDD.n244 VDD.n239 1084.97
R9445 VDD.n222 VDD.n199 1084.97
R9446 VDD.n222 VDD.n200 1084.97
R9447 VDD.n200 VDD.n172 1084.97
R9448 VDD.n199 VDD.n172 1084.97
R9449 VDD.n404 VDD.n174 1084.97
R9450 VDD.n404 VDD.n175 1084.97
R9451 VDD.n375 VDD.n175 1084.97
R9452 VDD.n375 VDD.n174 1084.97
R9453 VDD.n282 VDD.n201 1084.97
R9454 VDD.n282 VDD.n202 1084.97
R9455 VDD.n280 VDD.n202 1084.97
R9456 VDD.n280 VDD.n201 1084.97
R9457 VDD.n285 VDD.n177 1084.97
R9458 VDD.n288 VDD.n177 1084.97
R9459 VDD.n288 VDD.n245 1084.97
R9460 VDD.n285 VDD.n245 1084.97
R9461 VDD.n273 VDD.n203 1084.97
R9462 VDD.n273 VDD.n204 1084.97
R9463 VDD.n277 VDD.n204 1084.97
R9464 VDD.n277 VDD.n203 1084.97
R9465 VDD.n269 VDD.n186 1084.97
R9466 VDD.n270 VDD.n186 1084.97
R9467 VDD.n371 VDD.n270 1084.97
R9468 VDD.n371 VDD.n269 1084.97
R9469 VDD.n355 VDD.n205 1084.97
R9470 VDD.n355 VDD.n206 1084.97
R9471 VDD.n353 VDD.n206 1084.97
R9472 VDD.n353 VDD.n205 1084.97
R9473 VDD.n358 VDD.n178 1084.97
R9474 VDD.n361 VDD.n178 1084.97
R9475 VDD.n361 VDD.n246 1084.97
R9476 VDD.n358 VDD.n246 1084.97
R9477 VDD.n339 VDD.n207 1084.97
R9478 VDD.n339 VDD.n208 1084.97
R9479 VDD.n337 VDD.n208 1084.97
R9480 VDD.n337 VDD.n207 1084.97
R9481 VDD.n342 VDD.n185 1084.97
R9482 VDD.n345 VDD.n185 1084.97
R9483 VDD.n345 VDD.n268 1084.97
R9484 VDD.n342 VDD.n268 1084.97
R9485 VDD.n329 VDD.n209 1084.97
R9486 VDD.n329 VDD.n210 1084.97
R9487 VDD.n328 VDD.n210 1084.97
R9488 VDD.n328 VDD.n209 1084.97
R9489 VDD.n316 VDD.n211 1084.97
R9490 VDD.n316 VDD.n212 1084.97
R9491 VDD.n314 VDD.n212 1084.97
R9492 VDD.n314 VDD.n211 1084.97
R9493 VDD.n319 VDD.n179 1084.97
R9494 VDD.n322 VDD.n179 1084.97
R9495 VDD.n322 VDD.n247 1084.97
R9496 VDD.n319 VDD.n247 1084.97
R9497 VDD.n300 VDD.n213 1084.97
R9498 VDD.n300 VDD.n214 1084.97
R9499 VDD.n298 VDD.n214 1084.97
R9500 VDD.n298 VDD.n213 1084.97
R9501 VDD.n303 VDD.n184 1084.97
R9502 VDD.n306 VDD.n184 1084.97
R9503 VDD.n306 VDD.n267 1084.97
R9504 VDD.n303 VDD.n267 1084.97
R9505 VDD.n252 VDD.n215 1084.97
R9506 VDD.n252 VDD.n216 1084.97
R9507 VDD.n256 VDD.n216 1084.97
R9508 VDD.n256 VDD.n215 1084.97
R9509 VDD.n248 VDD.n180 1084.97
R9510 VDD.n249 VDD.n180 1084.97
R9511 VDD.n261 VDD.n249 1084.97
R9512 VDD.n261 VDD.n248 1084.97
R9513 VDD.n233 VDD.n217 1084.97
R9514 VDD.n233 VDD.n218 1084.97
R9515 VDD.n231 VDD.n218 1084.97
R9516 VDD.n231 VDD.n217 1084.97
R9517 VDD.n238 VDD.n183 1084.97
R9518 VDD.n380 VDD.n183 1084.97
R9519 VDD.n380 VDD.n379 1084.97
R9520 VDD.n379 VDD.n238 1084.97
R9521 VDD.n262 VDD.n181 1084.97
R9522 VDD.n263 VDD.n181 1084.97
R9523 VDD.n266 VDD.n263 1084.97
R9524 VDD.n266 VDD.n262 1084.97
R9525 VDD.n393 VDD.n226 1084.97
R9526 VDD.n226 VDD.n224 1084.97
R9527 VDD.n225 VDD.n224 1084.97
R9528 VDD.n393 VDD.n225 1084.97
R9529 VDD.n650 VDD.n435 1084.97
R9530 VDD.n650 VDD.n436 1084.97
R9531 VDD.n625 VDD.n436 1084.97
R9532 VDD.n625 VDD.n435 1084.97
R9533 VDD.n443 VDD.n442 1084.97
R9534 VDD.n642 VDD.n443 1084.97
R9535 VDD.n643 VDD.n642 1084.97
R9536 VDD.n643 VDD.n442 1084.97
R9537 VDD.n487 VDD.n424 1084.97
R9538 VDD.n488 VDD.n424 1084.97
R9539 VDD.n492 VDD.n488 1084.97
R9540 VDD.n492 VDD.n487 1084.97
R9541 VDD.n470 VDD.n447 1084.97
R9542 VDD.n470 VDD.n448 1084.97
R9543 VDD.n448 VDD.n420 1084.97
R9544 VDD.n447 VDD.n420 1084.97
R9545 VDD.n652 VDD.n422 1084.97
R9546 VDD.n652 VDD.n423 1084.97
R9547 VDD.n623 VDD.n423 1084.97
R9548 VDD.n623 VDD.n422 1084.97
R9549 VDD.n530 VDD.n449 1084.97
R9550 VDD.n530 VDD.n450 1084.97
R9551 VDD.n528 VDD.n450 1084.97
R9552 VDD.n528 VDD.n449 1084.97
R9553 VDD.n533 VDD.n425 1084.97
R9554 VDD.n536 VDD.n425 1084.97
R9555 VDD.n536 VDD.n493 1084.97
R9556 VDD.n533 VDD.n493 1084.97
R9557 VDD.n521 VDD.n451 1084.97
R9558 VDD.n521 VDD.n452 1084.97
R9559 VDD.n525 VDD.n452 1084.97
R9560 VDD.n525 VDD.n451 1084.97
R9561 VDD.n517 VDD.n434 1084.97
R9562 VDD.n518 VDD.n434 1084.97
R9563 VDD.n619 VDD.n518 1084.97
R9564 VDD.n619 VDD.n517 1084.97
R9565 VDD.n603 VDD.n453 1084.97
R9566 VDD.n603 VDD.n454 1084.97
R9567 VDD.n601 VDD.n454 1084.97
R9568 VDD.n601 VDD.n453 1084.97
R9569 VDD.n606 VDD.n426 1084.97
R9570 VDD.n609 VDD.n426 1084.97
R9571 VDD.n609 VDD.n494 1084.97
R9572 VDD.n606 VDD.n494 1084.97
R9573 VDD.n587 VDD.n455 1084.97
R9574 VDD.n587 VDD.n456 1084.97
R9575 VDD.n585 VDD.n456 1084.97
R9576 VDD.n585 VDD.n455 1084.97
R9577 VDD.n590 VDD.n433 1084.97
R9578 VDD.n593 VDD.n433 1084.97
R9579 VDD.n593 VDD.n516 1084.97
R9580 VDD.n590 VDD.n516 1084.97
R9581 VDD.n577 VDD.n457 1084.97
R9582 VDD.n577 VDD.n458 1084.97
R9583 VDD.n576 VDD.n458 1084.97
R9584 VDD.n576 VDD.n457 1084.97
R9585 VDD.n564 VDD.n459 1084.97
R9586 VDD.n564 VDD.n460 1084.97
R9587 VDD.n562 VDD.n460 1084.97
R9588 VDD.n562 VDD.n459 1084.97
R9589 VDD.n567 VDD.n427 1084.97
R9590 VDD.n570 VDD.n427 1084.97
R9591 VDD.n570 VDD.n495 1084.97
R9592 VDD.n567 VDD.n495 1084.97
R9593 VDD.n548 VDD.n461 1084.97
R9594 VDD.n548 VDD.n462 1084.97
R9595 VDD.n546 VDD.n462 1084.97
R9596 VDD.n546 VDD.n461 1084.97
R9597 VDD.n551 VDD.n432 1084.97
R9598 VDD.n554 VDD.n432 1084.97
R9599 VDD.n554 VDD.n515 1084.97
R9600 VDD.n551 VDD.n515 1084.97
R9601 VDD.n500 VDD.n463 1084.97
R9602 VDD.n500 VDD.n464 1084.97
R9603 VDD.n504 VDD.n464 1084.97
R9604 VDD.n504 VDD.n463 1084.97
R9605 VDD.n496 VDD.n428 1084.97
R9606 VDD.n497 VDD.n428 1084.97
R9607 VDD.n509 VDD.n497 1084.97
R9608 VDD.n509 VDD.n496 1084.97
R9609 VDD.n481 VDD.n465 1084.97
R9610 VDD.n481 VDD.n466 1084.97
R9611 VDD.n479 VDD.n466 1084.97
R9612 VDD.n479 VDD.n465 1084.97
R9613 VDD.n486 VDD.n431 1084.97
R9614 VDD.n628 VDD.n431 1084.97
R9615 VDD.n628 VDD.n627 1084.97
R9616 VDD.n627 VDD.n486 1084.97
R9617 VDD.n510 VDD.n429 1084.97
R9618 VDD.n511 VDD.n429 1084.97
R9619 VDD.n514 VDD.n511 1084.97
R9620 VDD.n514 VDD.n510 1084.97
R9621 VDD.n641 VDD.n474 1084.97
R9622 VDD.n474 VDD.n472 1084.97
R9623 VDD.n473 VDD.n472 1084.97
R9624 VDD.n641 VDD.n473 1084.97
R9625 VDD.n909 VDD.n694 1084.97
R9626 VDD.n909 VDD.n695 1084.97
R9627 VDD.n884 VDD.n695 1084.97
R9628 VDD.n884 VDD.n694 1084.97
R9629 VDD.n702 VDD.n701 1084.97
R9630 VDD.n901 VDD.n702 1084.97
R9631 VDD.n902 VDD.n901 1084.97
R9632 VDD.n902 VDD.n701 1084.97
R9633 VDD.n746 VDD.n683 1084.97
R9634 VDD.n747 VDD.n683 1084.97
R9635 VDD.n751 VDD.n747 1084.97
R9636 VDD.n751 VDD.n746 1084.97
R9637 VDD.n729 VDD.n706 1084.97
R9638 VDD.n729 VDD.n707 1084.97
R9639 VDD.n707 VDD.n679 1084.97
R9640 VDD.n706 VDD.n679 1084.97
R9641 VDD.n911 VDD.n681 1084.97
R9642 VDD.n911 VDD.n682 1084.97
R9643 VDD.n882 VDD.n682 1084.97
R9644 VDD.n882 VDD.n681 1084.97
R9645 VDD.n789 VDD.n708 1084.97
R9646 VDD.n789 VDD.n709 1084.97
R9647 VDD.n787 VDD.n709 1084.97
R9648 VDD.n787 VDD.n708 1084.97
R9649 VDD.n792 VDD.n684 1084.97
R9650 VDD.n795 VDD.n684 1084.97
R9651 VDD.n795 VDD.n752 1084.97
R9652 VDD.n792 VDD.n752 1084.97
R9653 VDD.n780 VDD.n710 1084.97
R9654 VDD.n780 VDD.n711 1084.97
R9655 VDD.n784 VDD.n711 1084.97
R9656 VDD.n784 VDD.n710 1084.97
R9657 VDD.n776 VDD.n693 1084.97
R9658 VDD.n777 VDD.n693 1084.97
R9659 VDD.n878 VDD.n777 1084.97
R9660 VDD.n878 VDD.n776 1084.97
R9661 VDD.n862 VDD.n712 1084.97
R9662 VDD.n862 VDD.n713 1084.97
R9663 VDD.n860 VDD.n713 1084.97
R9664 VDD.n860 VDD.n712 1084.97
R9665 VDD.n865 VDD.n685 1084.97
R9666 VDD.n868 VDD.n685 1084.97
R9667 VDD.n868 VDD.n753 1084.97
R9668 VDD.n865 VDD.n753 1084.97
R9669 VDD.n846 VDD.n714 1084.97
R9670 VDD.n846 VDD.n715 1084.97
R9671 VDD.n844 VDD.n715 1084.97
R9672 VDD.n844 VDD.n714 1084.97
R9673 VDD.n849 VDD.n692 1084.97
R9674 VDD.n852 VDD.n692 1084.97
R9675 VDD.n852 VDD.n775 1084.97
R9676 VDD.n849 VDD.n775 1084.97
R9677 VDD.n836 VDD.n716 1084.97
R9678 VDD.n836 VDD.n717 1084.97
R9679 VDD.n835 VDD.n717 1084.97
R9680 VDD.n835 VDD.n716 1084.97
R9681 VDD.n823 VDD.n718 1084.97
R9682 VDD.n823 VDD.n719 1084.97
R9683 VDD.n821 VDD.n719 1084.97
R9684 VDD.n821 VDD.n718 1084.97
R9685 VDD.n826 VDD.n686 1084.97
R9686 VDD.n829 VDD.n686 1084.97
R9687 VDD.n829 VDD.n754 1084.97
R9688 VDD.n826 VDD.n754 1084.97
R9689 VDD.n807 VDD.n720 1084.97
R9690 VDD.n807 VDD.n721 1084.97
R9691 VDD.n805 VDD.n721 1084.97
R9692 VDD.n805 VDD.n720 1084.97
R9693 VDD.n810 VDD.n691 1084.97
R9694 VDD.n813 VDD.n691 1084.97
R9695 VDD.n813 VDD.n774 1084.97
R9696 VDD.n810 VDD.n774 1084.97
R9697 VDD.n759 VDD.n722 1084.97
R9698 VDD.n759 VDD.n723 1084.97
R9699 VDD.n763 VDD.n723 1084.97
R9700 VDD.n763 VDD.n722 1084.97
R9701 VDD.n755 VDD.n687 1084.97
R9702 VDD.n756 VDD.n687 1084.97
R9703 VDD.n768 VDD.n756 1084.97
R9704 VDD.n768 VDD.n755 1084.97
R9705 VDD.n740 VDD.n724 1084.97
R9706 VDD.n740 VDD.n725 1084.97
R9707 VDD.n738 VDD.n725 1084.97
R9708 VDD.n738 VDD.n724 1084.97
R9709 VDD.n745 VDD.n690 1084.97
R9710 VDD.n887 VDD.n690 1084.97
R9711 VDD.n887 VDD.n886 1084.97
R9712 VDD.n886 VDD.n745 1084.97
R9713 VDD.n769 VDD.n688 1084.97
R9714 VDD.n770 VDD.n688 1084.97
R9715 VDD.n773 VDD.n770 1084.97
R9716 VDD.n773 VDD.n769 1084.97
R9717 VDD.n900 VDD.n733 1084.97
R9718 VDD.n733 VDD.n731 1084.97
R9719 VDD.n732 VDD.n731 1084.97
R9720 VDD.n900 VDD.n732 1084.97
R9721 VDD.n1168 VDD.n953 1084.97
R9722 VDD.n1168 VDD.n954 1084.97
R9723 VDD.n1143 VDD.n954 1084.97
R9724 VDD.n1143 VDD.n953 1084.97
R9725 VDD.n961 VDD.n960 1084.97
R9726 VDD.n1160 VDD.n961 1084.97
R9727 VDD.n1161 VDD.n1160 1084.97
R9728 VDD.n1161 VDD.n960 1084.97
R9729 VDD.n1005 VDD.n942 1084.97
R9730 VDD.n1006 VDD.n942 1084.97
R9731 VDD.n1010 VDD.n1006 1084.97
R9732 VDD.n1010 VDD.n1005 1084.97
R9733 VDD.n988 VDD.n965 1084.97
R9734 VDD.n988 VDD.n966 1084.97
R9735 VDD.n966 VDD.n938 1084.97
R9736 VDD.n965 VDD.n938 1084.97
R9737 VDD.n1170 VDD.n940 1084.97
R9738 VDD.n1170 VDD.n941 1084.97
R9739 VDD.n1141 VDD.n941 1084.97
R9740 VDD.n1141 VDD.n940 1084.97
R9741 VDD.n1048 VDD.n967 1084.97
R9742 VDD.n1048 VDD.n968 1084.97
R9743 VDD.n1046 VDD.n968 1084.97
R9744 VDD.n1046 VDD.n967 1084.97
R9745 VDD.n1051 VDD.n943 1084.97
R9746 VDD.n1054 VDD.n943 1084.97
R9747 VDD.n1054 VDD.n1011 1084.97
R9748 VDD.n1051 VDD.n1011 1084.97
R9749 VDD.n1039 VDD.n969 1084.97
R9750 VDD.n1039 VDD.n970 1084.97
R9751 VDD.n1043 VDD.n970 1084.97
R9752 VDD.n1043 VDD.n969 1084.97
R9753 VDD.n1035 VDD.n952 1084.97
R9754 VDD.n1036 VDD.n952 1084.97
R9755 VDD.n1137 VDD.n1036 1084.97
R9756 VDD.n1137 VDD.n1035 1084.97
R9757 VDD.n1121 VDD.n971 1084.97
R9758 VDD.n1121 VDD.n972 1084.97
R9759 VDD.n1119 VDD.n972 1084.97
R9760 VDD.n1119 VDD.n971 1084.97
R9761 VDD.n1124 VDD.n944 1084.97
R9762 VDD.n1127 VDD.n944 1084.97
R9763 VDD.n1127 VDD.n1012 1084.97
R9764 VDD.n1124 VDD.n1012 1084.97
R9765 VDD.n1105 VDD.n973 1084.97
R9766 VDD.n1105 VDD.n974 1084.97
R9767 VDD.n1103 VDD.n974 1084.97
R9768 VDD.n1103 VDD.n973 1084.97
R9769 VDD.n1108 VDD.n951 1084.97
R9770 VDD.n1111 VDD.n951 1084.97
R9771 VDD.n1111 VDD.n1034 1084.97
R9772 VDD.n1108 VDD.n1034 1084.97
R9773 VDD.n1095 VDD.n975 1084.97
R9774 VDD.n1095 VDD.n976 1084.97
R9775 VDD.n1094 VDD.n976 1084.97
R9776 VDD.n1094 VDD.n975 1084.97
R9777 VDD.n1082 VDD.n977 1084.97
R9778 VDD.n1082 VDD.n978 1084.97
R9779 VDD.n1080 VDD.n978 1084.97
R9780 VDD.n1080 VDD.n977 1084.97
R9781 VDD.n1085 VDD.n945 1084.97
R9782 VDD.n1088 VDD.n945 1084.97
R9783 VDD.n1088 VDD.n1013 1084.97
R9784 VDD.n1085 VDD.n1013 1084.97
R9785 VDD.n1066 VDD.n979 1084.97
R9786 VDD.n1066 VDD.n980 1084.97
R9787 VDD.n1064 VDD.n980 1084.97
R9788 VDD.n1064 VDD.n979 1084.97
R9789 VDD.n1069 VDD.n950 1084.97
R9790 VDD.n1072 VDD.n950 1084.97
R9791 VDD.n1072 VDD.n1033 1084.97
R9792 VDD.n1069 VDD.n1033 1084.97
R9793 VDD.n1018 VDD.n981 1084.97
R9794 VDD.n1018 VDD.n982 1084.97
R9795 VDD.n1022 VDD.n982 1084.97
R9796 VDD.n1022 VDD.n981 1084.97
R9797 VDD.n1014 VDD.n946 1084.97
R9798 VDD.n1015 VDD.n946 1084.97
R9799 VDD.n1027 VDD.n1015 1084.97
R9800 VDD.n1027 VDD.n1014 1084.97
R9801 VDD.n999 VDD.n983 1084.97
R9802 VDD.n999 VDD.n984 1084.97
R9803 VDD.n997 VDD.n984 1084.97
R9804 VDD.n997 VDD.n983 1084.97
R9805 VDD.n1004 VDD.n949 1084.97
R9806 VDD.n1146 VDD.n949 1084.97
R9807 VDD.n1146 VDD.n1145 1084.97
R9808 VDD.n1145 VDD.n1004 1084.97
R9809 VDD.n1028 VDD.n947 1084.97
R9810 VDD.n1029 VDD.n947 1084.97
R9811 VDD.n1032 VDD.n1029 1084.97
R9812 VDD.n1032 VDD.n1028 1084.97
R9813 VDD.n1159 VDD.n992 1084.97
R9814 VDD.n992 VDD.n990 1084.97
R9815 VDD.n991 VDD.n990 1084.97
R9816 VDD.n1159 VDD.n991 1084.97
R9817 VDD.n1427 VDD.n1212 1084.97
R9818 VDD.n1427 VDD.n1213 1084.97
R9819 VDD.n1402 VDD.n1213 1084.97
R9820 VDD.n1402 VDD.n1212 1084.97
R9821 VDD.n1220 VDD.n1219 1084.97
R9822 VDD.n1419 VDD.n1220 1084.97
R9823 VDD.n1420 VDD.n1419 1084.97
R9824 VDD.n1420 VDD.n1219 1084.97
R9825 VDD.n1264 VDD.n1201 1084.97
R9826 VDD.n1265 VDD.n1201 1084.97
R9827 VDD.n1269 VDD.n1265 1084.97
R9828 VDD.n1269 VDD.n1264 1084.97
R9829 VDD.n1247 VDD.n1224 1084.97
R9830 VDD.n1247 VDD.n1225 1084.97
R9831 VDD.n1225 VDD.n1197 1084.97
R9832 VDD.n1224 VDD.n1197 1084.97
R9833 VDD.n1429 VDD.n1199 1084.97
R9834 VDD.n1429 VDD.n1200 1084.97
R9835 VDD.n1400 VDD.n1200 1084.97
R9836 VDD.n1400 VDD.n1199 1084.97
R9837 VDD.n1307 VDD.n1226 1084.97
R9838 VDD.n1307 VDD.n1227 1084.97
R9839 VDD.n1305 VDD.n1227 1084.97
R9840 VDD.n1305 VDD.n1226 1084.97
R9841 VDD.n1310 VDD.n1202 1084.97
R9842 VDD.n1313 VDD.n1202 1084.97
R9843 VDD.n1313 VDD.n1270 1084.97
R9844 VDD.n1310 VDD.n1270 1084.97
R9845 VDD.n1298 VDD.n1228 1084.97
R9846 VDD.n1298 VDD.n1229 1084.97
R9847 VDD.n1302 VDD.n1229 1084.97
R9848 VDD.n1302 VDD.n1228 1084.97
R9849 VDD.n1294 VDD.n1211 1084.97
R9850 VDD.n1295 VDD.n1211 1084.97
R9851 VDD.n1396 VDD.n1295 1084.97
R9852 VDD.n1396 VDD.n1294 1084.97
R9853 VDD.n1380 VDD.n1230 1084.97
R9854 VDD.n1380 VDD.n1231 1084.97
R9855 VDD.n1378 VDD.n1231 1084.97
R9856 VDD.n1378 VDD.n1230 1084.97
R9857 VDD.n1383 VDD.n1203 1084.97
R9858 VDD.n1386 VDD.n1203 1084.97
R9859 VDD.n1386 VDD.n1271 1084.97
R9860 VDD.n1383 VDD.n1271 1084.97
R9861 VDD.n1364 VDD.n1232 1084.97
R9862 VDD.n1364 VDD.n1233 1084.97
R9863 VDD.n1362 VDD.n1233 1084.97
R9864 VDD.n1362 VDD.n1232 1084.97
R9865 VDD.n1367 VDD.n1210 1084.97
R9866 VDD.n1370 VDD.n1210 1084.97
R9867 VDD.n1370 VDD.n1293 1084.97
R9868 VDD.n1367 VDD.n1293 1084.97
R9869 VDD.n1354 VDD.n1234 1084.97
R9870 VDD.n1354 VDD.n1235 1084.97
R9871 VDD.n1353 VDD.n1235 1084.97
R9872 VDD.n1353 VDD.n1234 1084.97
R9873 VDD.n1341 VDD.n1236 1084.97
R9874 VDD.n1341 VDD.n1237 1084.97
R9875 VDD.n1339 VDD.n1237 1084.97
R9876 VDD.n1339 VDD.n1236 1084.97
R9877 VDD.n1344 VDD.n1204 1084.97
R9878 VDD.n1347 VDD.n1204 1084.97
R9879 VDD.n1347 VDD.n1272 1084.97
R9880 VDD.n1344 VDD.n1272 1084.97
R9881 VDD.n1325 VDD.n1238 1084.97
R9882 VDD.n1325 VDD.n1239 1084.97
R9883 VDD.n1323 VDD.n1239 1084.97
R9884 VDD.n1323 VDD.n1238 1084.97
R9885 VDD.n1328 VDD.n1209 1084.97
R9886 VDD.n1331 VDD.n1209 1084.97
R9887 VDD.n1331 VDD.n1292 1084.97
R9888 VDD.n1328 VDD.n1292 1084.97
R9889 VDD.n1277 VDD.n1240 1084.97
R9890 VDD.n1277 VDD.n1241 1084.97
R9891 VDD.n1281 VDD.n1241 1084.97
R9892 VDD.n1281 VDD.n1240 1084.97
R9893 VDD.n1273 VDD.n1205 1084.97
R9894 VDD.n1274 VDD.n1205 1084.97
R9895 VDD.n1286 VDD.n1274 1084.97
R9896 VDD.n1286 VDD.n1273 1084.97
R9897 VDD.n1258 VDD.n1242 1084.97
R9898 VDD.n1258 VDD.n1243 1084.97
R9899 VDD.n1256 VDD.n1243 1084.97
R9900 VDD.n1256 VDD.n1242 1084.97
R9901 VDD.n1263 VDD.n1208 1084.97
R9902 VDD.n1405 VDD.n1208 1084.97
R9903 VDD.n1405 VDD.n1404 1084.97
R9904 VDD.n1404 VDD.n1263 1084.97
R9905 VDD.n1287 VDD.n1206 1084.97
R9906 VDD.n1288 VDD.n1206 1084.97
R9907 VDD.n1291 VDD.n1288 1084.97
R9908 VDD.n1291 VDD.n1287 1084.97
R9909 VDD.n1418 VDD.n1251 1084.97
R9910 VDD.n1251 VDD.n1249 1084.97
R9911 VDD.n1250 VDD.n1249 1084.97
R9912 VDD.n1418 VDD.n1250 1084.97
R9913 VDD.n1686 VDD.n1471 1084.97
R9914 VDD.n1686 VDD.n1472 1084.97
R9915 VDD.n1661 VDD.n1472 1084.97
R9916 VDD.n1661 VDD.n1471 1084.97
R9917 VDD.n1479 VDD.n1478 1084.97
R9918 VDD.n1678 VDD.n1479 1084.97
R9919 VDD.n1679 VDD.n1678 1084.97
R9920 VDD.n1679 VDD.n1478 1084.97
R9921 VDD.n1523 VDD.n1460 1084.97
R9922 VDD.n1524 VDD.n1460 1084.97
R9923 VDD.n1528 VDD.n1524 1084.97
R9924 VDD.n1528 VDD.n1523 1084.97
R9925 VDD.n1506 VDD.n1483 1084.97
R9926 VDD.n1506 VDD.n1484 1084.97
R9927 VDD.n1484 VDD.n1456 1084.97
R9928 VDD.n1483 VDD.n1456 1084.97
R9929 VDD.n1688 VDD.n1458 1084.97
R9930 VDD.n1688 VDD.n1459 1084.97
R9931 VDD.n1659 VDD.n1459 1084.97
R9932 VDD.n1659 VDD.n1458 1084.97
R9933 VDD.n1566 VDD.n1485 1084.97
R9934 VDD.n1566 VDD.n1486 1084.97
R9935 VDD.n1564 VDD.n1486 1084.97
R9936 VDD.n1564 VDD.n1485 1084.97
R9937 VDD.n1569 VDD.n1461 1084.97
R9938 VDD.n1572 VDD.n1461 1084.97
R9939 VDD.n1572 VDD.n1529 1084.97
R9940 VDD.n1569 VDD.n1529 1084.97
R9941 VDD.n1557 VDD.n1487 1084.97
R9942 VDD.n1557 VDD.n1488 1084.97
R9943 VDD.n1561 VDD.n1488 1084.97
R9944 VDD.n1561 VDD.n1487 1084.97
R9945 VDD.n1553 VDD.n1470 1084.97
R9946 VDD.n1554 VDD.n1470 1084.97
R9947 VDD.n1655 VDD.n1554 1084.97
R9948 VDD.n1655 VDD.n1553 1084.97
R9949 VDD.n1639 VDD.n1489 1084.97
R9950 VDD.n1639 VDD.n1490 1084.97
R9951 VDD.n1637 VDD.n1490 1084.97
R9952 VDD.n1637 VDD.n1489 1084.97
R9953 VDD.n1642 VDD.n1462 1084.97
R9954 VDD.n1645 VDD.n1462 1084.97
R9955 VDD.n1645 VDD.n1530 1084.97
R9956 VDD.n1642 VDD.n1530 1084.97
R9957 VDD.n1623 VDD.n1491 1084.97
R9958 VDD.n1623 VDD.n1492 1084.97
R9959 VDD.n1621 VDD.n1492 1084.97
R9960 VDD.n1621 VDD.n1491 1084.97
R9961 VDD.n1626 VDD.n1469 1084.97
R9962 VDD.n1629 VDD.n1469 1084.97
R9963 VDD.n1629 VDD.n1552 1084.97
R9964 VDD.n1626 VDD.n1552 1084.97
R9965 VDD.n1613 VDD.n1493 1084.97
R9966 VDD.n1613 VDD.n1494 1084.97
R9967 VDD.n1612 VDD.n1494 1084.97
R9968 VDD.n1612 VDD.n1493 1084.97
R9969 VDD.n1600 VDD.n1495 1084.97
R9970 VDD.n1600 VDD.n1496 1084.97
R9971 VDD.n1598 VDD.n1496 1084.97
R9972 VDD.n1598 VDD.n1495 1084.97
R9973 VDD.n1603 VDD.n1463 1084.97
R9974 VDD.n1606 VDD.n1463 1084.97
R9975 VDD.n1606 VDD.n1531 1084.97
R9976 VDD.n1603 VDD.n1531 1084.97
R9977 VDD.n1584 VDD.n1497 1084.97
R9978 VDD.n1584 VDD.n1498 1084.97
R9979 VDD.n1582 VDD.n1498 1084.97
R9980 VDD.n1582 VDD.n1497 1084.97
R9981 VDD.n1587 VDD.n1468 1084.97
R9982 VDD.n1590 VDD.n1468 1084.97
R9983 VDD.n1590 VDD.n1551 1084.97
R9984 VDD.n1587 VDD.n1551 1084.97
R9985 VDD.n1536 VDD.n1499 1084.97
R9986 VDD.n1536 VDD.n1500 1084.97
R9987 VDD.n1540 VDD.n1500 1084.97
R9988 VDD.n1540 VDD.n1499 1084.97
R9989 VDD.n1532 VDD.n1464 1084.97
R9990 VDD.n1533 VDD.n1464 1084.97
R9991 VDD.n1545 VDD.n1533 1084.97
R9992 VDD.n1545 VDD.n1532 1084.97
R9993 VDD.n1517 VDD.n1501 1084.97
R9994 VDD.n1517 VDD.n1502 1084.97
R9995 VDD.n1515 VDD.n1502 1084.97
R9996 VDD.n1515 VDD.n1501 1084.97
R9997 VDD.n1522 VDD.n1467 1084.97
R9998 VDD.n1664 VDD.n1467 1084.97
R9999 VDD.n1664 VDD.n1663 1084.97
R10000 VDD.n1663 VDD.n1522 1084.97
R10001 VDD.n1546 VDD.n1465 1084.97
R10002 VDD.n1547 VDD.n1465 1084.97
R10003 VDD.n1550 VDD.n1547 1084.97
R10004 VDD.n1550 VDD.n1546 1084.97
R10005 VDD.n1677 VDD.n1510 1084.97
R10006 VDD.n1510 VDD.n1508 1084.97
R10007 VDD.n1509 VDD.n1508 1084.97
R10008 VDD.n1677 VDD.n1509 1084.97
R10009 VDD.n1945 VDD.n1730 1084.97
R10010 VDD.n1945 VDD.n1731 1084.97
R10011 VDD.n1920 VDD.n1731 1084.97
R10012 VDD.n1920 VDD.n1730 1084.97
R10013 VDD.n1738 VDD.n1737 1084.97
R10014 VDD.n1937 VDD.n1738 1084.97
R10015 VDD.n1938 VDD.n1937 1084.97
R10016 VDD.n1938 VDD.n1737 1084.97
R10017 VDD.n1782 VDD.n1719 1084.97
R10018 VDD.n1783 VDD.n1719 1084.97
R10019 VDD.n1787 VDD.n1783 1084.97
R10020 VDD.n1787 VDD.n1782 1084.97
R10021 VDD.n1765 VDD.n1742 1084.97
R10022 VDD.n1765 VDD.n1743 1084.97
R10023 VDD.n1743 VDD.n1715 1084.97
R10024 VDD.n1742 VDD.n1715 1084.97
R10025 VDD.n1947 VDD.n1717 1084.97
R10026 VDD.n1947 VDD.n1718 1084.97
R10027 VDD.n1918 VDD.n1718 1084.97
R10028 VDD.n1918 VDD.n1717 1084.97
R10029 VDD.n1825 VDD.n1744 1084.97
R10030 VDD.n1825 VDD.n1745 1084.97
R10031 VDD.n1823 VDD.n1745 1084.97
R10032 VDD.n1823 VDD.n1744 1084.97
R10033 VDD.n1828 VDD.n1720 1084.97
R10034 VDD.n1831 VDD.n1720 1084.97
R10035 VDD.n1831 VDD.n1788 1084.97
R10036 VDD.n1828 VDD.n1788 1084.97
R10037 VDD.n1816 VDD.n1746 1084.97
R10038 VDD.n1816 VDD.n1747 1084.97
R10039 VDD.n1820 VDD.n1747 1084.97
R10040 VDD.n1820 VDD.n1746 1084.97
R10041 VDD.n1812 VDD.n1729 1084.97
R10042 VDD.n1813 VDD.n1729 1084.97
R10043 VDD.n1914 VDD.n1813 1084.97
R10044 VDD.n1914 VDD.n1812 1084.97
R10045 VDD.n1898 VDD.n1748 1084.97
R10046 VDD.n1898 VDD.n1749 1084.97
R10047 VDD.n1896 VDD.n1749 1084.97
R10048 VDD.n1896 VDD.n1748 1084.97
R10049 VDD.n1901 VDD.n1721 1084.97
R10050 VDD.n1904 VDD.n1721 1084.97
R10051 VDD.n1904 VDD.n1789 1084.97
R10052 VDD.n1901 VDD.n1789 1084.97
R10053 VDD.n1882 VDD.n1750 1084.97
R10054 VDD.n1882 VDD.n1751 1084.97
R10055 VDD.n1880 VDD.n1751 1084.97
R10056 VDD.n1880 VDD.n1750 1084.97
R10057 VDD.n1885 VDD.n1728 1084.97
R10058 VDD.n1888 VDD.n1728 1084.97
R10059 VDD.n1888 VDD.n1811 1084.97
R10060 VDD.n1885 VDD.n1811 1084.97
R10061 VDD.n1872 VDD.n1752 1084.97
R10062 VDD.n1872 VDD.n1753 1084.97
R10063 VDD.n1871 VDD.n1753 1084.97
R10064 VDD.n1871 VDD.n1752 1084.97
R10065 VDD.n1859 VDD.n1754 1084.97
R10066 VDD.n1859 VDD.n1755 1084.97
R10067 VDD.n1857 VDD.n1755 1084.97
R10068 VDD.n1857 VDD.n1754 1084.97
R10069 VDD.n1862 VDD.n1722 1084.97
R10070 VDD.n1865 VDD.n1722 1084.97
R10071 VDD.n1865 VDD.n1790 1084.97
R10072 VDD.n1862 VDD.n1790 1084.97
R10073 VDD.n1843 VDD.n1756 1084.97
R10074 VDD.n1843 VDD.n1757 1084.97
R10075 VDD.n1841 VDD.n1757 1084.97
R10076 VDD.n1841 VDD.n1756 1084.97
R10077 VDD.n1846 VDD.n1727 1084.97
R10078 VDD.n1849 VDD.n1727 1084.97
R10079 VDD.n1849 VDD.n1810 1084.97
R10080 VDD.n1846 VDD.n1810 1084.97
R10081 VDD.n1795 VDD.n1758 1084.97
R10082 VDD.n1795 VDD.n1759 1084.97
R10083 VDD.n1799 VDD.n1759 1084.97
R10084 VDD.n1799 VDD.n1758 1084.97
R10085 VDD.n1791 VDD.n1723 1084.97
R10086 VDD.n1792 VDD.n1723 1084.97
R10087 VDD.n1804 VDD.n1792 1084.97
R10088 VDD.n1804 VDD.n1791 1084.97
R10089 VDD.n1776 VDD.n1760 1084.97
R10090 VDD.n1776 VDD.n1761 1084.97
R10091 VDD.n1774 VDD.n1761 1084.97
R10092 VDD.n1774 VDD.n1760 1084.97
R10093 VDD.n1781 VDD.n1726 1084.97
R10094 VDD.n1923 VDD.n1726 1084.97
R10095 VDD.n1923 VDD.n1922 1084.97
R10096 VDD.n1922 VDD.n1781 1084.97
R10097 VDD.n1805 VDD.n1724 1084.97
R10098 VDD.n1806 VDD.n1724 1084.97
R10099 VDD.n1809 VDD.n1806 1084.97
R10100 VDD.n1809 VDD.n1805 1084.97
R10101 VDD.n1936 VDD.n1769 1084.97
R10102 VDD.n1769 VDD.n1767 1084.97
R10103 VDD.n1768 VDD.n1767 1084.97
R10104 VDD.n1936 VDD.n1768 1084.97
R10105 VDD.n2204 VDD.n1989 1084.97
R10106 VDD.n2204 VDD.n1990 1084.97
R10107 VDD.n2179 VDD.n1990 1084.97
R10108 VDD.n2179 VDD.n1989 1084.97
R10109 VDD.n1997 VDD.n1996 1084.97
R10110 VDD.n2196 VDD.n1997 1084.97
R10111 VDD.n2197 VDD.n2196 1084.97
R10112 VDD.n2197 VDD.n1996 1084.97
R10113 VDD.n2041 VDD.n1978 1084.97
R10114 VDD.n2042 VDD.n1978 1084.97
R10115 VDD.n2046 VDD.n2042 1084.97
R10116 VDD.n2046 VDD.n2041 1084.97
R10117 VDD.n2024 VDD.n2001 1084.97
R10118 VDD.n2024 VDD.n2002 1084.97
R10119 VDD.n2002 VDD.n1974 1084.97
R10120 VDD.n2001 VDD.n1974 1084.97
R10121 VDD.n2206 VDD.n1976 1084.97
R10122 VDD.n2206 VDD.n1977 1084.97
R10123 VDD.n2177 VDD.n1977 1084.97
R10124 VDD.n2177 VDD.n1976 1084.97
R10125 VDD.n2084 VDD.n2003 1084.97
R10126 VDD.n2084 VDD.n2004 1084.97
R10127 VDD.n2082 VDD.n2004 1084.97
R10128 VDD.n2082 VDD.n2003 1084.97
R10129 VDD.n2087 VDD.n1979 1084.97
R10130 VDD.n2090 VDD.n1979 1084.97
R10131 VDD.n2090 VDD.n2047 1084.97
R10132 VDD.n2087 VDD.n2047 1084.97
R10133 VDD.n2075 VDD.n2005 1084.97
R10134 VDD.n2075 VDD.n2006 1084.97
R10135 VDD.n2079 VDD.n2006 1084.97
R10136 VDD.n2079 VDD.n2005 1084.97
R10137 VDD.n2071 VDD.n1988 1084.97
R10138 VDD.n2072 VDD.n1988 1084.97
R10139 VDD.n2173 VDD.n2072 1084.97
R10140 VDD.n2173 VDD.n2071 1084.97
R10141 VDD.n2157 VDD.n2007 1084.97
R10142 VDD.n2157 VDD.n2008 1084.97
R10143 VDD.n2155 VDD.n2008 1084.97
R10144 VDD.n2155 VDD.n2007 1084.97
R10145 VDD.n2160 VDD.n1980 1084.97
R10146 VDD.n2163 VDD.n1980 1084.97
R10147 VDD.n2163 VDD.n2048 1084.97
R10148 VDD.n2160 VDD.n2048 1084.97
R10149 VDD.n2141 VDD.n2009 1084.97
R10150 VDD.n2141 VDD.n2010 1084.97
R10151 VDD.n2139 VDD.n2010 1084.97
R10152 VDD.n2139 VDD.n2009 1084.97
R10153 VDD.n2144 VDD.n1987 1084.97
R10154 VDD.n2147 VDD.n1987 1084.97
R10155 VDD.n2147 VDD.n2070 1084.97
R10156 VDD.n2144 VDD.n2070 1084.97
R10157 VDD.n2131 VDD.n2011 1084.97
R10158 VDD.n2131 VDD.n2012 1084.97
R10159 VDD.n2130 VDD.n2012 1084.97
R10160 VDD.n2130 VDD.n2011 1084.97
R10161 VDD.n2118 VDD.n2013 1084.97
R10162 VDD.n2118 VDD.n2014 1084.97
R10163 VDD.n2116 VDD.n2014 1084.97
R10164 VDD.n2116 VDD.n2013 1084.97
R10165 VDD.n2121 VDD.n1981 1084.97
R10166 VDD.n2124 VDD.n1981 1084.97
R10167 VDD.n2124 VDD.n2049 1084.97
R10168 VDD.n2121 VDD.n2049 1084.97
R10169 VDD.n2102 VDD.n2015 1084.97
R10170 VDD.n2102 VDD.n2016 1084.97
R10171 VDD.n2100 VDD.n2016 1084.97
R10172 VDD.n2100 VDD.n2015 1084.97
R10173 VDD.n2105 VDD.n1986 1084.97
R10174 VDD.n2108 VDD.n1986 1084.97
R10175 VDD.n2108 VDD.n2069 1084.97
R10176 VDD.n2105 VDD.n2069 1084.97
R10177 VDD.n2054 VDD.n2017 1084.97
R10178 VDD.n2054 VDD.n2018 1084.97
R10179 VDD.n2058 VDD.n2018 1084.97
R10180 VDD.n2058 VDD.n2017 1084.97
R10181 VDD.n2050 VDD.n1982 1084.97
R10182 VDD.n2051 VDD.n1982 1084.97
R10183 VDD.n2063 VDD.n2051 1084.97
R10184 VDD.n2063 VDD.n2050 1084.97
R10185 VDD.n2035 VDD.n2019 1084.97
R10186 VDD.n2035 VDD.n2020 1084.97
R10187 VDD.n2033 VDD.n2020 1084.97
R10188 VDD.n2033 VDD.n2019 1084.97
R10189 VDD.n2040 VDD.n1985 1084.97
R10190 VDD.n2182 VDD.n1985 1084.97
R10191 VDD.n2182 VDD.n2181 1084.97
R10192 VDD.n2181 VDD.n2040 1084.97
R10193 VDD.n2064 VDD.n1983 1084.97
R10194 VDD.n2065 VDD.n1983 1084.97
R10195 VDD.n2068 VDD.n2065 1084.97
R10196 VDD.n2068 VDD.n2064 1084.97
R10197 VDD.n2195 VDD.n2028 1084.97
R10198 VDD.n2028 VDD.n2026 1084.97
R10199 VDD.n2027 VDD.n2026 1084.97
R10200 VDD.n2195 VDD.n2027 1084.97
R10201 VDD.n2463 VDD.n2248 1084.97
R10202 VDD.n2463 VDD.n2249 1084.97
R10203 VDD.n2438 VDD.n2249 1084.97
R10204 VDD.n2438 VDD.n2248 1084.97
R10205 VDD.n2256 VDD.n2255 1084.97
R10206 VDD.n2455 VDD.n2256 1084.97
R10207 VDD.n2456 VDD.n2455 1084.97
R10208 VDD.n2456 VDD.n2255 1084.97
R10209 VDD.n2300 VDD.n2237 1084.97
R10210 VDD.n2301 VDD.n2237 1084.97
R10211 VDD.n2305 VDD.n2301 1084.97
R10212 VDD.n2305 VDD.n2300 1084.97
R10213 VDD.n2283 VDD.n2260 1084.97
R10214 VDD.n2283 VDD.n2261 1084.97
R10215 VDD.n2261 VDD.n2233 1084.97
R10216 VDD.n2260 VDD.n2233 1084.97
R10217 VDD.n2465 VDD.n2235 1084.97
R10218 VDD.n2465 VDD.n2236 1084.97
R10219 VDD.n2436 VDD.n2236 1084.97
R10220 VDD.n2436 VDD.n2235 1084.97
R10221 VDD.n2343 VDD.n2262 1084.97
R10222 VDD.n2343 VDD.n2263 1084.97
R10223 VDD.n2341 VDD.n2263 1084.97
R10224 VDD.n2341 VDD.n2262 1084.97
R10225 VDD.n2346 VDD.n2238 1084.97
R10226 VDD.n2349 VDD.n2238 1084.97
R10227 VDD.n2349 VDD.n2306 1084.97
R10228 VDD.n2346 VDD.n2306 1084.97
R10229 VDD.n2334 VDD.n2264 1084.97
R10230 VDD.n2334 VDD.n2265 1084.97
R10231 VDD.n2338 VDD.n2265 1084.97
R10232 VDD.n2338 VDD.n2264 1084.97
R10233 VDD.n2330 VDD.n2247 1084.97
R10234 VDD.n2331 VDD.n2247 1084.97
R10235 VDD.n2432 VDD.n2331 1084.97
R10236 VDD.n2432 VDD.n2330 1084.97
R10237 VDD.n2416 VDD.n2266 1084.97
R10238 VDD.n2416 VDD.n2267 1084.97
R10239 VDD.n2414 VDD.n2267 1084.97
R10240 VDD.n2414 VDD.n2266 1084.97
R10241 VDD.n2419 VDD.n2239 1084.97
R10242 VDD.n2422 VDD.n2239 1084.97
R10243 VDD.n2422 VDD.n2307 1084.97
R10244 VDD.n2419 VDD.n2307 1084.97
R10245 VDD.n2400 VDD.n2268 1084.97
R10246 VDD.n2400 VDD.n2269 1084.97
R10247 VDD.n2398 VDD.n2269 1084.97
R10248 VDD.n2398 VDD.n2268 1084.97
R10249 VDD.n2403 VDD.n2246 1084.97
R10250 VDD.n2406 VDD.n2246 1084.97
R10251 VDD.n2406 VDD.n2329 1084.97
R10252 VDD.n2403 VDD.n2329 1084.97
R10253 VDD.n2390 VDD.n2270 1084.97
R10254 VDD.n2390 VDD.n2271 1084.97
R10255 VDD.n2389 VDD.n2271 1084.97
R10256 VDD.n2389 VDD.n2270 1084.97
R10257 VDD.n2377 VDD.n2272 1084.97
R10258 VDD.n2377 VDD.n2273 1084.97
R10259 VDD.n2375 VDD.n2273 1084.97
R10260 VDD.n2375 VDD.n2272 1084.97
R10261 VDD.n2380 VDD.n2240 1084.97
R10262 VDD.n2383 VDD.n2240 1084.97
R10263 VDD.n2383 VDD.n2308 1084.97
R10264 VDD.n2380 VDD.n2308 1084.97
R10265 VDD.n2361 VDD.n2274 1084.97
R10266 VDD.n2361 VDD.n2275 1084.97
R10267 VDD.n2359 VDD.n2275 1084.97
R10268 VDD.n2359 VDD.n2274 1084.97
R10269 VDD.n2364 VDD.n2245 1084.97
R10270 VDD.n2367 VDD.n2245 1084.97
R10271 VDD.n2367 VDD.n2328 1084.97
R10272 VDD.n2364 VDD.n2328 1084.97
R10273 VDD.n2313 VDD.n2276 1084.97
R10274 VDD.n2313 VDD.n2277 1084.97
R10275 VDD.n2317 VDD.n2277 1084.97
R10276 VDD.n2317 VDD.n2276 1084.97
R10277 VDD.n2309 VDD.n2241 1084.97
R10278 VDD.n2310 VDD.n2241 1084.97
R10279 VDD.n2322 VDD.n2310 1084.97
R10280 VDD.n2322 VDD.n2309 1084.97
R10281 VDD.n2294 VDD.n2278 1084.97
R10282 VDD.n2294 VDD.n2279 1084.97
R10283 VDD.n2292 VDD.n2279 1084.97
R10284 VDD.n2292 VDD.n2278 1084.97
R10285 VDD.n2299 VDD.n2244 1084.97
R10286 VDD.n2441 VDD.n2244 1084.97
R10287 VDD.n2441 VDD.n2440 1084.97
R10288 VDD.n2440 VDD.n2299 1084.97
R10289 VDD.n2323 VDD.n2242 1084.97
R10290 VDD.n2324 VDD.n2242 1084.97
R10291 VDD.n2327 VDD.n2324 1084.97
R10292 VDD.n2327 VDD.n2323 1084.97
R10293 VDD.n2454 VDD.n2287 1084.97
R10294 VDD.n2287 VDD.n2285 1084.97
R10295 VDD.n2286 VDD.n2285 1084.97
R10296 VDD.n2454 VDD.n2286 1084.97
R10297 VDD.n2722 VDD.n2507 1084.97
R10298 VDD.n2722 VDD.n2508 1084.97
R10299 VDD.n2697 VDD.n2508 1084.97
R10300 VDD.n2697 VDD.n2507 1084.97
R10301 VDD.n2515 VDD.n2514 1084.97
R10302 VDD.n2714 VDD.n2515 1084.97
R10303 VDD.n2715 VDD.n2714 1084.97
R10304 VDD.n2715 VDD.n2514 1084.97
R10305 VDD.n2559 VDD.n2496 1084.97
R10306 VDD.n2560 VDD.n2496 1084.97
R10307 VDD.n2564 VDD.n2560 1084.97
R10308 VDD.n2564 VDD.n2559 1084.97
R10309 VDD.n2542 VDD.n2519 1084.97
R10310 VDD.n2542 VDD.n2520 1084.97
R10311 VDD.n2520 VDD.n2492 1084.97
R10312 VDD.n2519 VDD.n2492 1084.97
R10313 VDD.n2724 VDD.n2494 1084.97
R10314 VDD.n2724 VDD.n2495 1084.97
R10315 VDD.n2695 VDD.n2495 1084.97
R10316 VDD.n2695 VDD.n2494 1084.97
R10317 VDD.n2602 VDD.n2521 1084.97
R10318 VDD.n2602 VDD.n2522 1084.97
R10319 VDD.n2600 VDD.n2522 1084.97
R10320 VDD.n2600 VDD.n2521 1084.97
R10321 VDD.n2605 VDD.n2497 1084.97
R10322 VDD.n2608 VDD.n2497 1084.97
R10323 VDD.n2608 VDD.n2565 1084.97
R10324 VDD.n2605 VDD.n2565 1084.97
R10325 VDD.n2593 VDD.n2523 1084.97
R10326 VDD.n2593 VDD.n2524 1084.97
R10327 VDD.n2597 VDD.n2524 1084.97
R10328 VDD.n2597 VDD.n2523 1084.97
R10329 VDD.n2589 VDD.n2506 1084.97
R10330 VDD.n2590 VDD.n2506 1084.97
R10331 VDD.n2691 VDD.n2590 1084.97
R10332 VDD.n2691 VDD.n2589 1084.97
R10333 VDD.n2675 VDD.n2525 1084.97
R10334 VDD.n2675 VDD.n2526 1084.97
R10335 VDD.n2673 VDD.n2526 1084.97
R10336 VDD.n2673 VDD.n2525 1084.97
R10337 VDD.n2678 VDD.n2498 1084.97
R10338 VDD.n2681 VDD.n2498 1084.97
R10339 VDD.n2681 VDD.n2566 1084.97
R10340 VDD.n2678 VDD.n2566 1084.97
R10341 VDD.n2659 VDD.n2527 1084.97
R10342 VDD.n2659 VDD.n2528 1084.97
R10343 VDD.n2657 VDD.n2528 1084.97
R10344 VDD.n2657 VDD.n2527 1084.97
R10345 VDD.n2662 VDD.n2505 1084.97
R10346 VDD.n2665 VDD.n2505 1084.97
R10347 VDD.n2665 VDD.n2588 1084.97
R10348 VDD.n2662 VDD.n2588 1084.97
R10349 VDD.n2649 VDD.n2529 1084.97
R10350 VDD.n2649 VDD.n2530 1084.97
R10351 VDD.n2648 VDD.n2530 1084.97
R10352 VDD.n2648 VDD.n2529 1084.97
R10353 VDD.n2636 VDD.n2531 1084.97
R10354 VDD.n2636 VDD.n2532 1084.97
R10355 VDD.n2634 VDD.n2532 1084.97
R10356 VDD.n2634 VDD.n2531 1084.97
R10357 VDD.n2639 VDD.n2499 1084.97
R10358 VDD.n2642 VDD.n2499 1084.97
R10359 VDD.n2642 VDD.n2567 1084.97
R10360 VDD.n2639 VDD.n2567 1084.97
R10361 VDD.n2620 VDD.n2533 1084.97
R10362 VDD.n2620 VDD.n2534 1084.97
R10363 VDD.n2618 VDD.n2534 1084.97
R10364 VDD.n2618 VDD.n2533 1084.97
R10365 VDD.n2623 VDD.n2504 1084.97
R10366 VDD.n2626 VDD.n2504 1084.97
R10367 VDD.n2626 VDD.n2587 1084.97
R10368 VDD.n2623 VDD.n2587 1084.97
R10369 VDD.n2572 VDD.n2535 1084.97
R10370 VDD.n2572 VDD.n2536 1084.97
R10371 VDD.n2576 VDD.n2536 1084.97
R10372 VDD.n2576 VDD.n2535 1084.97
R10373 VDD.n2568 VDD.n2500 1084.97
R10374 VDD.n2569 VDD.n2500 1084.97
R10375 VDD.n2581 VDD.n2569 1084.97
R10376 VDD.n2581 VDD.n2568 1084.97
R10377 VDD.n2553 VDD.n2537 1084.97
R10378 VDD.n2553 VDD.n2538 1084.97
R10379 VDD.n2551 VDD.n2538 1084.97
R10380 VDD.n2551 VDD.n2537 1084.97
R10381 VDD.n2558 VDD.n2503 1084.97
R10382 VDD.n2700 VDD.n2503 1084.97
R10383 VDD.n2700 VDD.n2699 1084.97
R10384 VDD.n2699 VDD.n2558 1084.97
R10385 VDD.n2582 VDD.n2501 1084.97
R10386 VDD.n2583 VDD.n2501 1084.97
R10387 VDD.n2586 VDD.n2583 1084.97
R10388 VDD.n2586 VDD.n2582 1084.97
R10389 VDD.n2713 VDD.n2546 1084.97
R10390 VDD.n2546 VDD.n2544 1084.97
R10391 VDD.n2545 VDD.n2544 1084.97
R10392 VDD.n2713 VDD.n2545 1084.97
R10393 VDD.n2981 VDD.n2766 1084.97
R10394 VDD.n2981 VDD.n2767 1084.97
R10395 VDD.n2956 VDD.n2767 1084.97
R10396 VDD.n2956 VDD.n2766 1084.97
R10397 VDD.n2774 VDD.n2773 1084.97
R10398 VDD.n2973 VDD.n2774 1084.97
R10399 VDD.n2974 VDD.n2973 1084.97
R10400 VDD.n2974 VDD.n2773 1084.97
R10401 VDD.n2818 VDD.n2755 1084.97
R10402 VDD.n2819 VDD.n2755 1084.97
R10403 VDD.n2823 VDD.n2819 1084.97
R10404 VDD.n2823 VDD.n2818 1084.97
R10405 VDD.n2801 VDD.n2778 1084.97
R10406 VDD.n2801 VDD.n2779 1084.97
R10407 VDD.n2779 VDD.n2751 1084.97
R10408 VDD.n2778 VDD.n2751 1084.97
R10409 VDD.n2983 VDD.n2753 1084.97
R10410 VDD.n2983 VDD.n2754 1084.97
R10411 VDD.n2954 VDD.n2754 1084.97
R10412 VDD.n2954 VDD.n2753 1084.97
R10413 VDD.n2861 VDD.n2780 1084.97
R10414 VDD.n2861 VDD.n2781 1084.97
R10415 VDD.n2859 VDD.n2781 1084.97
R10416 VDD.n2859 VDD.n2780 1084.97
R10417 VDD.n2864 VDD.n2756 1084.97
R10418 VDD.n2867 VDD.n2756 1084.97
R10419 VDD.n2867 VDD.n2824 1084.97
R10420 VDD.n2864 VDD.n2824 1084.97
R10421 VDD.n2852 VDD.n2782 1084.97
R10422 VDD.n2852 VDD.n2783 1084.97
R10423 VDD.n2856 VDD.n2783 1084.97
R10424 VDD.n2856 VDD.n2782 1084.97
R10425 VDD.n2848 VDD.n2765 1084.97
R10426 VDD.n2849 VDD.n2765 1084.97
R10427 VDD.n2950 VDD.n2849 1084.97
R10428 VDD.n2950 VDD.n2848 1084.97
R10429 VDD.n2934 VDD.n2784 1084.97
R10430 VDD.n2934 VDD.n2785 1084.97
R10431 VDD.n2932 VDD.n2785 1084.97
R10432 VDD.n2932 VDD.n2784 1084.97
R10433 VDD.n2937 VDD.n2757 1084.97
R10434 VDD.n2940 VDD.n2757 1084.97
R10435 VDD.n2940 VDD.n2825 1084.97
R10436 VDD.n2937 VDD.n2825 1084.97
R10437 VDD.n2918 VDD.n2786 1084.97
R10438 VDD.n2918 VDD.n2787 1084.97
R10439 VDD.n2916 VDD.n2787 1084.97
R10440 VDD.n2916 VDD.n2786 1084.97
R10441 VDD.n2921 VDD.n2764 1084.97
R10442 VDD.n2924 VDD.n2764 1084.97
R10443 VDD.n2924 VDD.n2847 1084.97
R10444 VDD.n2921 VDD.n2847 1084.97
R10445 VDD.n2908 VDD.n2788 1084.97
R10446 VDD.n2908 VDD.n2789 1084.97
R10447 VDD.n2907 VDD.n2789 1084.97
R10448 VDD.n2907 VDD.n2788 1084.97
R10449 VDD.n2895 VDD.n2790 1084.97
R10450 VDD.n2895 VDD.n2791 1084.97
R10451 VDD.n2893 VDD.n2791 1084.97
R10452 VDD.n2893 VDD.n2790 1084.97
R10453 VDD.n2898 VDD.n2758 1084.97
R10454 VDD.n2901 VDD.n2758 1084.97
R10455 VDD.n2901 VDD.n2826 1084.97
R10456 VDD.n2898 VDD.n2826 1084.97
R10457 VDD.n2879 VDD.n2792 1084.97
R10458 VDD.n2879 VDD.n2793 1084.97
R10459 VDD.n2877 VDD.n2793 1084.97
R10460 VDD.n2877 VDD.n2792 1084.97
R10461 VDD.n2882 VDD.n2763 1084.97
R10462 VDD.n2885 VDD.n2763 1084.97
R10463 VDD.n2885 VDD.n2846 1084.97
R10464 VDD.n2882 VDD.n2846 1084.97
R10465 VDD.n2831 VDD.n2794 1084.97
R10466 VDD.n2831 VDD.n2795 1084.97
R10467 VDD.n2835 VDD.n2795 1084.97
R10468 VDD.n2835 VDD.n2794 1084.97
R10469 VDD.n2827 VDD.n2759 1084.97
R10470 VDD.n2828 VDD.n2759 1084.97
R10471 VDD.n2840 VDD.n2828 1084.97
R10472 VDD.n2840 VDD.n2827 1084.97
R10473 VDD.n2812 VDD.n2796 1084.97
R10474 VDD.n2812 VDD.n2797 1084.97
R10475 VDD.n2810 VDD.n2797 1084.97
R10476 VDD.n2810 VDD.n2796 1084.97
R10477 VDD.n2817 VDD.n2762 1084.97
R10478 VDD.n2959 VDD.n2762 1084.97
R10479 VDD.n2959 VDD.n2958 1084.97
R10480 VDD.n2958 VDD.n2817 1084.97
R10481 VDD.n2841 VDD.n2760 1084.97
R10482 VDD.n2842 VDD.n2760 1084.97
R10483 VDD.n2845 VDD.n2842 1084.97
R10484 VDD.n2845 VDD.n2841 1084.97
R10485 VDD.n2972 VDD.n2805 1084.97
R10486 VDD.n2805 VDD.n2803 1084.97
R10487 VDD.n2804 VDD.n2803 1084.97
R10488 VDD.n2972 VDD.n2804 1084.97
R10489 VDD.n3240 VDD.n3025 1084.97
R10490 VDD.n3240 VDD.n3026 1084.97
R10491 VDD.n3215 VDD.n3026 1084.97
R10492 VDD.n3215 VDD.n3025 1084.97
R10493 VDD.n3033 VDD.n3032 1084.97
R10494 VDD.n3232 VDD.n3033 1084.97
R10495 VDD.n3233 VDD.n3232 1084.97
R10496 VDD.n3233 VDD.n3032 1084.97
R10497 VDD.n3077 VDD.n3014 1084.97
R10498 VDD.n3078 VDD.n3014 1084.97
R10499 VDD.n3082 VDD.n3078 1084.97
R10500 VDD.n3082 VDD.n3077 1084.97
R10501 VDD.n3060 VDD.n3037 1084.97
R10502 VDD.n3060 VDD.n3038 1084.97
R10503 VDD.n3038 VDD.n3010 1084.97
R10504 VDD.n3037 VDD.n3010 1084.97
R10505 VDD.n3242 VDD.n3012 1084.97
R10506 VDD.n3242 VDD.n3013 1084.97
R10507 VDD.n3213 VDD.n3013 1084.97
R10508 VDD.n3213 VDD.n3012 1084.97
R10509 VDD.n3120 VDD.n3039 1084.97
R10510 VDD.n3120 VDD.n3040 1084.97
R10511 VDD.n3118 VDD.n3040 1084.97
R10512 VDD.n3118 VDD.n3039 1084.97
R10513 VDD.n3123 VDD.n3015 1084.97
R10514 VDD.n3126 VDD.n3015 1084.97
R10515 VDD.n3126 VDD.n3083 1084.97
R10516 VDD.n3123 VDD.n3083 1084.97
R10517 VDD.n3111 VDD.n3041 1084.97
R10518 VDD.n3111 VDD.n3042 1084.97
R10519 VDD.n3115 VDD.n3042 1084.97
R10520 VDD.n3115 VDD.n3041 1084.97
R10521 VDD.n3107 VDD.n3024 1084.97
R10522 VDD.n3108 VDD.n3024 1084.97
R10523 VDD.n3209 VDD.n3108 1084.97
R10524 VDD.n3209 VDD.n3107 1084.97
R10525 VDD.n3193 VDD.n3043 1084.97
R10526 VDD.n3193 VDD.n3044 1084.97
R10527 VDD.n3191 VDD.n3044 1084.97
R10528 VDD.n3191 VDD.n3043 1084.97
R10529 VDD.n3196 VDD.n3016 1084.97
R10530 VDD.n3199 VDD.n3016 1084.97
R10531 VDD.n3199 VDD.n3084 1084.97
R10532 VDD.n3196 VDD.n3084 1084.97
R10533 VDD.n3177 VDD.n3045 1084.97
R10534 VDD.n3177 VDD.n3046 1084.97
R10535 VDD.n3175 VDD.n3046 1084.97
R10536 VDD.n3175 VDD.n3045 1084.97
R10537 VDD.n3180 VDD.n3023 1084.97
R10538 VDD.n3183 VDD.n3023 1084.97
R10539 VDD.n3183 VDD.n3106 1084.97
R10540 VDD.n3180 VDD.n3106 1084.97
R10541 VDD.n3167 VDD.n3047 1084.97
R10542 VDD.n3167 VDD.n3048 1084.97
R10543 VDD.n3166 VDD.n3048 1084.97
R10544 VDD.n3166 VDD.n3047 1084.97
R10545 VDD.n3154 VDD.n3049 1084.97
R10546 VDD.n3154 VDD.n3050 1084.97
R10547 VDD.n3152 VDD.n3050 1084.97
R10548 VDD.n3152 VDD.n3049 1084.97
R10549 VDD.n3157 VDD.n3017 1084.97
R10550 VDD.n3160 VDD.n3017 1084.97
R10551 VDD.n3160 VDD.n3085 1084.97
R10552 VDD.n3157 VDD.n3085 1084.97
R10553 VDD.n3138 VDD.n3051 1084.97
R10554 VDD.n3138 VDD.n3052 1084.97
R10555 VDD.n3136 VDD.n3052 1084.97
R10556 VDD.n3136 VDD.n3051 1084.97
R10557 VDD.n3141 VDD.n3022 1084.97
R10558 VDD.n3144 VDD.n3022 1084.97
R10559 VDD.n3144 VDD.n3105 1084.97
R10560 VDD.n3141 VDD.n3105 1084.97
R10561 VDD.n3090 VDD.n3053 1084.97
R10562 VDD.n3090 VDD.n3054 1084.97
R10563 VDD.n3094 VDD.n3054 1084.97
R10564 VDD.n3094 VDD.n3053 1084.97
R10565 VDD.n3086 VDD.n3018 1084.97
R10566 VDD.n3087 VDD.n3018 1084.97
R10567 VDD.n3099 VDD.n3087 1084.97
R10568 VDD.n3099 VDD.n3086 1084.97
R10569 VDD.n3071 VDD.n3055 1084.97
R10570 VDD.n3071 VDD.n3056 1084.97
R10571 VDD.n3069 VDD.n3056 1084.97
R10572 VDD.n3069 VDD.n3055 1084.97
R10573 VDD.n3076 VDD.n3021 1084.97
R10574 VDD.n3218 VDD.n3021 1084.97
R10575 VDD.n3218 VDD.n3217 1084.97
R10576 VDD.n3217 VDD.n3076 1084.97
R10577 VDD.n3100 VDD.n3019 1084.97
R10578 VDD.n3101 VDD.n3019 1084.97
R10579 VDD.n3104 VDD.n3101 1084.97
R10580 VDD.n3104 VDD.n3100 1084.97
R10581 VDD.n3231 VDD.n3064 1084.97
R10582 VDD.n3064 VDD.n3062 1084.97
R10583 VDD.n3063 VDD.n3062 1084.97
R10584 VDD.n3231 VDD.n3063 1084.97
R10585 VDD.n3499 VDD.n3284 1084.97
R10586 VDD.n3499 VDD.n3285 1084.97
R10587 VDD.n3474 VDD.n3285 1084.97
R10588 VDD.n3474 VDD.n3284 1084.97
R10589 VDD.n3292 VDD.n3291 1084.97
R10590 VDD.n3491 VDD.n3292 1084.97
R10591 VDD.n3492 VDD.n3491 1084.97
R10592 VDD.n3492 VDD.n3291 1084.97
R10593 VDD.n3336 VDD.n3273 1084.97
R10594 VDD.n3337 VDD.n3273 1084.97
R10595 VDD.n3341 VDD.n3337 1084.97
R10596 VDD.n3341 VDD.n3336 1084.97
R10597 VDD.n3319 VDD.n3296 1084.97
R10598 VDD.n3319 VDD.n3297 1084.97
R10599 VDD.n3297 VDD.n3269 1084.97
R10600 VDD.n3296 VDD.n3269 1084.97
R10601 VDD.n3501 VDD.n3271 1084.97
R10602 VDD.n3501 VDD.n3272 1084.97
R10603 VDD.n3472 VDD.n3272 1084.97
R10604 VDD.n3472 VDD.n3271 1084.97
R10605 VDD.n3379 VDD.n3298 1084.97
R10606 VDD.n3379 VDD.n3299 1084.97
R10607 VDD.n3377 VDD.n3299 1084.97
R10608 VDD.n3377 VDD.n3298 1084.97
R10609 VDD.n3382 VDD.n3274 1084.97
R10610 VDD.n3385 VDD.n3274 1084.97
R10611 VDD.n3385 VDD.n3342 1084.97
R10612 VDD.n3382 VDD.n3342 1084.97
R10613 VDD.n3370 VDD.n3300 1084.97
R10614 VDD.n3370 VDD.n3301 1084.97
R10615 VDD.n3374 VDD.n3301 1084.97
R10616 VDD.n3374 VDD.n3300 1084.97
R10617 VDD.n3366 VDD.n3283 1084.97
R10618 VDD.n3367 VDD.n3283 1084.97
R10619 VDD.n3468 VDD.n3367 1084.97
R10620 VDD.n3468 VDD.n3366 1084.97
R10621 VDD.n3452 VDD.n3302 1084.97
R10622 VDD.n3452 VDD.n3303 1084.97
R10623 VDD.n3450 VDD.n3303 1084.97
R10624 VDD.n3450 VDD.n3302 1084.97
R10625 VDD.n3455 VDD.n3275 1084.97
R10626 VDD.n3458 VDD.n3275 1084.97
R10627 VDD.n3458 VDD.n3343 1084.97
R10628 VDD.n3455 VDD.n3343 1084.97
R10629 VDD.n3436 VDD.n3304 1084.97
R10630 VDD.n3436 VDD.n3305 1084.97
R10631 VDD.n3434 VDD.n3305 1084.97
R10632 VDD.n3434 VDD.n3304 1084.97
R10633 VDD.n3439 VDD.n3282 1084.97
R10634 VDD.n3442 VDD.n3282 1084.97
R10635 VDD.n3442 VDD.n3365 1084.97
R10636 VDD.n3439 VDD.n3365 1084.97
R10637 VDD.n3426 VDD.n3306 1084.97
R10638 VDD.n3426 VDD.n3307 1084.97
R10639 VDD.n3425 VDD.n3307 1084.97
R10640 VDD.n3425 VDD.n3306 1084.97
R10641 VDD.n3413 VDD.n3308 1084.97
R10642 VDD.n3413 VDD.n3309 1084.97
R10643 VDD.n3411 VDD.n3309 1084.97
R10644 VDD.n3411 VDD.n3308 1084.97
R10645 VDD.n3416 VDD.n3276 1084.97
R10646 VDD.n3419 VDD.n3276 1084.97
R10647 VDD.n3419 VDD.n3344 1084.97
R10648 VDD.n3416 VDD.n3344 1084.97
R10649 VDD.n3397 VDD.n3310 1084.97
R10650 VDD.n3397 VDD.n3311 1084.97
R10651 VDD.n3395 VDD.n3311 1084.97
R10652 VDD.n3395 VDD.n3310 1084.97
R10653 VDD.n3400 VDD.n3281 1084.97
R10654 VDD.n3403 VDD.n3281 1084.97
R10655 VDD.n3403 VDD.n3364 1084.97
R10656 VDD.n3400 VDD.n3364 1084.97
R10657 VDD.n3349 VDD.n3312 1084.97
R10658 VDD.n3349 VDD.n3313 1084.97
R10659 VDD.n3353 VDD.n3313 1084.97
R10660 VDD.n3353 VDD.n3312 1084.97
R10661 VDD.n3345 VDD.n3277 1084.97
R10662 VDD.n3346 VDD.n3277 1084.97
R10663 VDD.n3358 VDD.n3346 1084.97
R10664 VDD.n3358 VDD.n3345 1084.97
R10665 VDD.n3330 VDD.n3314 1084.97
R10666 VDD.n3330 VDD.n3315 1084.97
R10667 VDD.n3328 VDD.n3315 1084.97
R10668 VDD.n3328 VDD.n3314 1084.97
R10669 VDD.n3335 VDD.n3280 1084.97
R10670 VDD.n3477 VDD.n3280 1084.97
R10671 VDD.n3477 VDD.n3476 1084.97
R10672 VDD.n3476 VDD.n3335 1084.97
R10673 VDD.n3359 VDD.n3278 1084.97
R10674 VDD.n3360 VDD.n3278 1084.97
R10675 VDD.n3363 VDD.n3360 1084.97
R10676 VDD.n3363 VDD.n3359 1084.97
R10677 VDD.n3490 VDD.n3323 1084.97
R10678 VDD.n3323 VDD.n3321 1084.97
R10679 VDD.n3322 VDD.n3321 1084.97
R10680 VDD.n3490 VDD.n3322 1084.97
R10681 VDD.n3758 VDD.n3543 1084.97
R10682 VDD.n3758 VDD.n3544 1084.97
R10683 VDD.n3733 VDD.n3544 1084.97
R10684 VDD.n3733 VDD.n3543 1084.97
R10685 VDD.n3551 VDD.n3550 1084.97
R10686 VDD.n3750 VDD.n3551 1084.97
R10687 VDD.n3751 VDD.n3750 1084.97
R10688 VDD.n3751 VDD.n3550 1084.97
R10689 VDD.n3595 VDD.n3532 1084.97
R10690 VDD.n3596 VDD.n3532 1084.97
R10691 VDD.n3600 VDD.n3596 1084.97
R10692 VDD.n3600 VDD.n3595 1084.97
R10693 VDD.n3578 VDD.n3555 1084.97
R10694 VDD.n3578 VDD.n3556 1084.97
R10695 VDD.n3556 VDD.n3528 1084.97
R10696 VDD.n3555 VDD.n3528 1084.97
R10697 VDD.n3760 VDD.n3530 1084.97
R10698 VDD.n3760 VDD.n3531 1084.97
R10699 VDD.n3731 VDD.n3531 1084.97
R10700 VDD.n3731 VDD.n3530 1084.97
R10701 VDD.n3638 VDD.n3557 1084.97
R10702 VDD.n3638 VDD.n3558 1084.97
R10703 VDD.n3636 VDD.n3558 1084.97
R10704 VDD.n3636 VDD.n3557 1084.97
R10705 VDD.n3641 VDD.n3533 1084.97
R10706 VDD.n3644 VDD.n3533 1084.97
R10707 VDD.n3644 VDD.n3601 1084.97
R10708 VDD.n3641 VDD.n3601 1084.97
R10709 VDD.n3629 VDD.n3559 1084.97
R10710 VDD.n3629 VDD.n3560 1084.97
R10711 VDD.n3633 VDD.n3560 1084.97
R10712 VDD.n3633 VDD.n3559 1084.97
R10713 VDD.n3625 VDD.n3542 1084.97
R10714 VDD.n3626 VDD.n3542 1084.97
R10715 VDD.n3727 VDD.n3626 1084.97
R10716 VDD.n3727 VDD.n3625 1084.97
R10717 VDD.n3711 VDD.n3561 1084.97
R10718 VDD.n3711 VDD.n3562 1084.97
R10719 VDD.n3709 VDD.n3562 1084.97
R10720 VDD.n3709 VDD.n3561 1084.97
R10721 VDD.n3714 VDD.n3534 1084.97
R10722 VDD.n3717 VDD.n3534 1084.97
R10723 VDD.n3717 VDD.n3602 1084.97
R10724 VDD.n3714 VDD.n3602 1084.97
R10725 VDD.n3695 VDD.n3563 1084.97
R10726 VDD.n3695 VDD.n3564 1084.97
R10727 VDD.n3693 VDD.n3564 1084.97
R10728 VDD.n3693 VDD.n3563 1084.97
R10729 VDD.n3698 VDD.n3541 1084.97
R10730 VDD.n3701 VDD.n3541 1084.97
R10731 VDD.n3701 VDD.n3624 1084.97
R10732 VDD.n3698 VDD.n3624 1084.97
R10733 VDD.n3685 VDD.n3565 1084.97
R10734 VDD.n3685 VDD.n3566 1084.97
R10735 VDD.n3684 VDD.n3566 1084.97
R10736 VDD.n3684 VDD.n3565 1084.97
R10737 VDD.n3672 VDD.n3567 1084.97
R10738 VDD.n3672 VDD.n3568 1084.97
R10739 VDD.n3670 VDD.n3568 1084.97
R10740 VDD.n3670 VDD.n3567 1084.97
R10741 VDD.n3675 VDD.n3535 1084.97
R10742 VDD.n3678 VDD.n3535 1084.97
R10743 VDD.n3678 VDD.n3603 1084.97
R10744 VDD.n3675 VDD.n3603 1084.97
R10745 VDD.n3656 VDD.n3569 1084.97
R10746 VDD.n3656 VDD.n3570 1084.97
R10747 VDD.n3654 VDD.n3570 1084.97
R10748 VDD.n3654 VDD.n3569 1084.97
R10749 VDD.n3659 VDD.n3540 1084.97
R10750 VDD.n3662 VDD.n3540 1084.97
R10751 VDD.n3662 VDD.n3623 1084.97
R10752 VDD.n3659 VDD.n3623 1084.97
R10753 VDD.n3608 VDD.n3571 1084.97
R10754 VDD.n3608 VDD.n3572 1084.97
R10755 VDD.n3612 VDD.n3572 1084.97
R10756 VDD.n3612 VDD.n3571 1084.97
R10757 VDD.n3604 VDD.n3536 1084.97
R10758 VDD.n3605 VDD.n3536 1084.97
R10759 VDD.n3617 VDD.n3605 1084.97
R10760 VDD.n3617 VDD.n3604 1084.97
R10761 VDD.n3589 VDD.n3573 1084.97
R10762 VDD.n3589 VDD.n3574 1084.97
R10763 VDD.n3587 VDD.n3574 1084.97
R10764 VDD.n3587 VDD.n3573 1084.97
R10765 VDD.n3594 VDD.n3539 1084.97
R10766 VDD.n3736 VDD.n3539 1084.97
R10767 VDD.n3736 VDD.n3735 1084.97
R10768 VDD.n3735 VDD.n3594 1084.97
R10769 VDD.n3618 VDD.n3537 1084.97
R10770 VDD.n3619 VDD.n3537 1084.97
R10771 VDD.n3622 VDD.n3619 1084.97
R10772 VDD.n3622 VDD.n3618 1084.97
R10773 VDD.n3749 VDD.n3582 1084.97
R10774 VDD.n3582 VDD.n3580 1084.97
R10775 VDD.n3581 VDD.n3580 1084.97
R10776 VDD.n3749 VDD.n3581 1084.97
R10777 VDD.n4017 VDD.n3802 1084.97
R10778 VDD.n4017 VDD.n3803 1084.97
R10779 VDD.n3992 VDD.n3803 1084.97
R10780 VDD.n3992 VDD.n3802 1084.97
R10781 VDD.n3810 VDD.n3809 1084.97
R10782 VDD.n4009 VDD.n3810 1084.97
R10783 VDD.n4010 VDD.n4009 1084.97
R10784 VDD.n4010 VDD.n3809 1084.97
R10785 VDD.n3854 VDD.n3791 1084.97
R10786 VDD.n3855 VDD.n3791 1084.97
R10787 VDD.n3859 VDD.n3855 1084.97
R10788 VDD.n3859 VDD.n3854 1084.97
R10789 VDD.n3837 VDD.n3814 1084.97
R10790 VDD.n3837 VDD.n3815 1084.97
R10791 VDD.n3815 VDD.n3787 1084.97
R10792 VDD.n3814 VDD.n3787 1084.97
R10793 VDD.n4019 VDD.n3789 1084.97
R10794 VDD.n4019 VDD.n3790 1084.97
R10795 VDD.n3990 VDD.n3790 1084.97
R10796 VDD.n3990 VDD.n3789 1084.97
R10797 VDD.n3897 VDD.n3816 1084.97
R10798 VDD.n3897 VDD.n3817 1084.97
R10799 VDD.n3895 VDD.n3817 1084.97
R10800 VDD.n3895 VDD.n3816 1084.97
R10801 VDD.n3900 VDD.n3792 1084.97
R10802 VDD.n3903 VDD.n3792 1084.97
R10803 VDD.n3903 VDD.n3860 1084.97
R10804 VDD.n3900 VDD.n3860 1084.97
R10805 VDD.n3888 VDD.n3818 1084.97
R10806 VDD.n3888 VDD.n3819 1084.97
R10807 VDD.n3892 VDD.n3819 1084.97
R10808 VDD.n3892 VDD.n3818 1084.97
R10809 VDD.n3884 VDD.n3801 1084.97
R10810 VDD.n3885 VDD.n3801 1084.97
R10811 VDD.n3986 VDD.n3885 1084.97
R10812 VDD.n3986 VDD.n3884 1084.97
R10813 VDD.n3970 VDD.n3820 1084.97
R10814 VDD.n3970 VDD.n3821 1084.97
R10815 VDD.n3968 VDD.n3821 1084.97
R10816 VDD.n3968 VDD.n3820 1084.97
R10817 VDD.n3973 VDD.n3793 1084.97
R10818 VDD.n3976 VDD.n3793 1084.97
R10819 VDD.n3976 VDD.n3861 1084.97
R10820 VDD.n3973 VDD.n3861 1084.97
R10821 VDD.n3954 VDD.n3822 1084.97
R10822 VDD.n3954 VDD.n3823 1084.97
R10823 VDD.n3952 VDD.n3823 1084.97
R10824 VDD.n3952 VDD.n3822 1084.97
R10825 VDD.n3957 VDD.n3800 1084.97
R10826 VDD.n3960 VDD.n3800 1084.97
R10827 VDD.n3960 VDD.n3883 1084.97
R10828 VDD.n3957 VDD.n3883 1084.97
R10829 VDD.n3944 VDD.n3824 1084.97
R10830 VDD.n3944 VDD.n3825 1084.97
R10831 VDD.n3943 VDD.n3825 1084.97
R10832 VDD.n3943 VDD.n3824 1084.97
R10833 VDD.n3931 VDD.n3826 1084.97
R10834 VDD.n3931 VDD.n3827 1084.97
R10835 VDD.n3929 VDD.n3827 1084.97
R10836 VDD.n3929 VDD.n3826 1084.97
R10837 VDD.n3934 VDD.n3794 1084.97
R10838 VDD.n3937 VDD.n3794 1084.97
R10839 VDD.n3937 VDD.n3862 1084.97
R10840 VDD.n3934 VDD.n3862 1084.97
R10841 VDD.n3915 VDD.n3828 1084.97
R10842 VDD.n3915 VDD.n3829 1084.97
R10843 VDD.n3913 VDD.n3829 1084.97
R10844 VDD.n3913 VDD.n3828 1084.97
R10845 VDD.n3918 VDD.n3799 1084.97
R10846 VDD.n3921 VDD.n3799 1084.97
R10847 VDD.n3921 VDD.n3882 1084.97
R10848 VDD.n3918 VDD.n3882 1084.97
R10849 VDD.n3867 VDD.n3830 1084.97
R10850 VDD.n3867 VDD.n3831 1084.97
R10851 VDD.n3871 VDD.n3831 1084.97
R10852 VDD.n3871 VDD.n3830 1084.97
R10853 VDD.n3863 VDD.n3795 1084.97
R10854 VDD.n3864 VDD.n3795 1084.97
R10855 VDD.n3876 VDD.n3864 1084.97
R10856 VDD.n3876 VDD.n3863 1084.97
R10857 VDD.n3848 VDD.n3832 1084.97
R10858 VDD.n3848 VDD.n3833 1084.97
R10859 VDD.n3846 VDD.n3833 1084.97
R10860 VDD.n3846 VDD.n3832 1084.97
R10861 VDD.n3853 VDD.n3798 1084.97
R10862 VDD.n3995 VDD.n3798 1084.97
R10863 VDD.n3995 VDD.n3994 1084.97
R10864 VDD.n3994 VDD.n3853 1084.97
R10865 VDD.n3877 VDD.n3796 1084.97
R10866 VDD.n3878 VDD.n3796 1084.97
R10867 VDD.n3881 VDD.n3878 1084.97
R10868 VDD.n3881 VDD.n3877 1084.97
R10869 VDD.n4008 VDD.n3841 1084.97
R10870 VDD.n3841 VDD.n3839 1084.97
R10871 VDD.n3840 VDD.n3839 1084.97
R10872 VDD.n4008 VDD.n3840 1084.97
R10873 VDD.n4276 VDD.n4061 1084.97
R10874 VDD.n4276 VDD.n4062 1084.97
R10875 VDD.n4251 VDD.n4062 1084.97
R10876 VDD.n4251 VDD.n4061 1084.97
R10877 VDD.n4069 VDD.n4068 1084.97
R10878 VDD.n4268 VDD.n4069 1084.97
R10879 VDD.n4269 VDD.n4268 1084.97
R10880 VDD.n4269 VDD.n4068 1084.97
R10881 VDD.n4113 VDD.n4050 1084.97
R10882 VDD.n4114 VDD.n4050 1084.97
R10883 VDD.n4118 VDD.n4114 1084.97
R10884 VDD.n4118 VDD.n4113 1084.97
R10885 VDD.n4096 VDD.n4073 1084.97
R10886 VDD.n4096 VDD.n4074 1084.97
R10887 VDD.n4074 VDD.n4046 1084.97
R10888 VDD.n4073 VDD.n4046 1084.97
R10889 VDD.n4278 VDD.n4048 1084.97
R10890 VDD.n4278 VDD.n4049 1084.97
R10891 VDD.n4249 VDD.n4049 1084.97
R10892 VDD.n4249 VDD.n4048 1084.97
R10893 VDD.n4156 VDD.n4075 1084.97
R10894 VDD.n4156 VDD.n4076 1084.97
R10895 VDD.n4154 VDD.n4076 1084.97
R10896 VDD.n4154 VDD.n4075 1084.97
R10897 VDD.n4159 VDD.n4051 1084.97
R10898 VDD.n4162 VDD.n4051 1084.97
R10899 VDD.n4162 VDD.n4119 1084.97
R10900 VDD.n4159 VDD.n4119 1084.97
R10901 VDD.n4147 VDD.n4077 1084.97
R10902 VDD.n4147 VDD.n4078 1084.97
R10903 VDD.n4151 VDD.n4078 1084.97
R10904 VDD.n4151 VDD.n4077 1084.97
R10905 VDD.n4143 VDD.n4060 1084.97
R10906 VDD.n4144 VDD.n4060 1084.97
R10907 VDD.n4245 VDD.n4144 1084.97
R10908 VDD.n4245 VDD.n4143 1084.97
R10909 VDD.n4229 VDD.n4079 1084.97
R10910 VDD.n4229 VDD.n4080 1084.97
R10911 VDD.n4227 VDD.n4080 1084.97
R10912 VDD.n4227 VDD.n4079 1084.97
R10913 VDD.n4232 VDD.n4052 1084.97
R10914 VDD.n4235 VDD.n4052 1084.97
R10915 VDD.n4235 VDD.n4120 1084.97
R10916 VDD.n4232 VDD.n4120 1084.97
R10917 VDD.n4213 VDD.n4081 1084.97
R10918 VDD.n4213 VDD.n4082 1084.97
R10919 VDD.n4211 VDD.n4082 1084.97
R10920 VDD.n4211 VDD.n4081 1084.97
R10921 VDD.n4216 VDD.n4059 1084.97
R10922 VDD.n4219 VDD.n4059 1084.97
R10923 VDD.n4219 VDD.n4142 1084.97
R10924 VDD.n4216 VDD.n4142 1084.97
R10925 VDD.n4203 VDD.n4083 1084.97
R10926 VDD.n4203 VDD.n4084 1084.97
R10927 VDD.n4202 VDD.n4084 1084.97
R10928 VDD.n4202 VDD.n4083 1084.97
R10929 VDD.n4190 VDD.n4085 1084.97
R10930 VDD.n4190 VDD.n4086 1084.97
R10931 VDD.n4188 VDD.n4086 1084.97
R10932 VDD.n4188 VDD.n4085 1084.97
R10933 VDD.n4193 VDD.n4053 1084.97
R10934 VDD.n4196 VDD.n4053 1084.97
R10935 VDD.n4196 VDD.n4121 1084.97
R10936 VDD.n4193 VDD.n4121 1084.97
R10937 VDD.n4174 VDD.n4087 1084.97
R10938 VDD.n4174 VDD.n4088 1084.97
R10939 VDD.n4172 VDD.n4088 1084.97
R10940 VDD.n4172 VDD.n4087 1084.97
R10941 VDD.n4177 VDD.n4058 1084.97
R10942 VDD.n4180 VDD.n4058 1084.97
R10943 VDD.n4180 VDD.n4141 1084.97
R10944 VDD.n4177 VDD.n4141 1084.97
R10945 VDD.n4126 VDD.n4089 1084.97
R10946 VDD.n4126 VDD.n4090 1084.97
R10947 VDD.n4130 VDD.n4090 1084.97
R10948 VDD.n4130 VDD.n4089 1084.97
R10949 VDD.n4122 VDD.n4054 1084.97
R10950 VDD.n4123 VDD.n4054 1084.97
R10951 VDD.n4135 VDD.n4123 1084.97
R10952 VDD.n4135 VDD.n4122 1084.97
R10953 VDD.n4107 VDD.n4091 1084.97
R10954 VDD.n4107 VDD.n4092 1084.97
R10955 VDD.n4105 VDD.n4092 1084.97
R10956 VDD.n4105 VDD.n4091 1084.97
R10957 VDD.n4112 VDD.n4057 1084.97
R10958 VDD.n4254 VDD.n4057 1084.97
R10959 VDD.n4254 VDD.n4253 1084.97
R10960 VDD.n4253 VDD.n4112 1084.97
R10961 VDD.n4136 VDD.n4055 1084.97
R10962 VDD.n4137 VDD.n4055 1084.97
R10963 VDD.n4140 VDD.n4137 1084.97
R10964 VDD.n4140 VDD.n4136 1084.97
R10965 VDD.n4267 VDD.n4100 1084.97
R10966 VDD.n4100 VDD.n4098 1084.97
R10967 VDD.n4099 VDD.n4098 1084.97
R10968 VDD.n4267 VDD.n4099 1084.97
R10969 VDD.n4510 VDD.n4320 1084.97
R10970 VDD.n4535 VDD.n4320 1084.97
R10971 VDD.n4535 VDD.n4321 1084.97
R10972 VDD.n4510 VDD.n4321 1084.97
R10973 VDD.n4328 VDD.n4327 1084.97
R10974 VDD.n4527 VDD.n4328 1084.97
R10975 VDD.n4528 VDD.n4527 1084.97
R10976 VDD.n4528 VDD.n4327 1084.97
R10977 VDD.n4372 VDD.n4309 1084.97
R10978 VDD.n4373 VDD.n4309 1084.97
R10979 VDD.n4377 VDD.n4373 1084.97
R10980 VDD.n4377 VDD.n4372 1084.97
R10981 VDD.n4355 VDD.n4332 1084.97
R10982 VDD.n4355 VDD.n4333 1084.97
R10983 VDD.n4333 VDD.n4305 1084.97
R10984 VDD.n4332 VDD.n4305 1084.97
R10985 VDD.n4537 VDD.n4307 1084.97
R10986 VDD.n4537 VDD.n4308 1084.97
R10987 VDD.n4508 VDD.n4308 1084.97
R10988 VDD.n4508 VDD.n4307 1084.97
R10989 VDD.n4415 VDD.n4334 1084.97
R10990 VDD.n4415 VDD.n4335 1084.97
R10991 VDD.n4413 VDD.n4335 1084.97
R10992 VDD.n4413 VDD.n4334 1084.97
R10993 VDD.n4418 VDD.n4310 1084.97
R10994 VDD.n4421 VDD.n4310 1084.97
R10995 VDD.n4421 VDD.n4378 1084.97
R10996 VDD.n4418 VDD.n4378 1084.97
R10997 VDD.n4406 VDD.n4336 1084.97
R10998 VDD.n4406 VDD.n4337 1084.97
R10999 VDD.n4410 VDD.n4337 1084.97
R11000 VDD.n4410 VDD.n4336 1084.97
R11001 VDD.n4402 VDD.n4319 1084.97
R11002 VDD.n4403 VDD.n4319 1084.97
R11003 VDD.n4504 VDD.n4403 1084.97
R11004 VDD.n4504 VDD.n4402 1084.97
R11005 VDD.n4488 VDD.n4338 1084.97
R11006 VDD.n4488 VDD.n4339 1084.97
R11007 VDD.n4486 VDD.n4339 1084.97
R11008 VDD.n4486 VDD.n4338 1084.97
R11009 VDD.n4491 VDD.n4311 1084.97
R11010 VDD.n4494 VDD.n4311 1084.97
R11011 VDD.n4494 VDD.n4379 1084.97
R11012 VDD.n4491 VDD.n4379 1084.97
R11013 VDD.n4472 VDD.n4340 1084.97
R11014 VDD.n4472 VDD.n4341 1084.97
R11015 VDD.n4470 VDD.n4341 1084.97
R11016 VDD.n4470 VDD.n4340 1084.97
R11017 VDD.n4475 VDD.n4318 1084.97
R11018 VDD.n4478 VDD.n4318 1084.97
R11019 VDD.n4478 VDD.n4401 1084.97
R11020 VDD.n4475 VDD.n4401 1084.97
R11021 VDD.n4462 VDD.n4342 1084.97
R11022 VDD.n4462 VDD.n4343 1084.97
R11023 VDD.n4461 VDD.n4343 1084.97
R11024 VDD.n4461 VDD.n4342 1084.97
R11025 VDD.n4449 VDD.n4344 1084.97
R11026 VDD.n4449 VDD.n4345 1084.97
R11027 VDD.n4447 VDD.n4345 1084.97
R11028 VDD.n4447 VDD.n4344 1084.97
R11029 VDD.n4452 VDD.n4312 1084.97
R11030 VDD.n4455 VDD.n4312 1084.97
R11031 VDD.n4455 VDD.n4380 1084.97
R11032 VDD.n4452 VDD.n4380 1084.97
R11033 VDD.n4433 VDD.n4346 1084.97
R11034 VDD.n4433 VDD.n4347 1084.97
R11035 VDD.n4431 VDD.n4347 1084.97
R11036 VDD.n4431 VDD.n4346 1084.97
R11037 VDD.n4436 VDD.n4317 1084.97
R11038 VDD.n4439 VDD.n4317 1084.97
R11039 VDD.n4439 VDD.n4400 1084.97
R11040 VDD.n4436 VDD.n4400 1084.97
R11041 VDD.n4385 VDD.n4348 1084.97
R11042 VDD.n4385 VDD.n4349 1084.97
R11043 VDD.n4389 VDD.n4349 1084.97
R11044 VDD.n4389 VDD.n4348 1084.97
R11045 VDD.n4381 VDD.n4313 1084.97
R11046 VDD.n4382 VDD.n4313 1084.97
R11047 VDD.n4394 VDD.n4382 1084.97
R11048 VDD.n4394 VDD.n4381 1084.97
R11049 VDD.n4366 VDD.n4350 1084.97
R11050 VDD.n4366 VDD.n4351 1084.97
R11051 VDD.n4364 VDD.n4351 1084.97
R11052 VDD.n4364 VDD.n4350 1084.97
R11053 VDD.n4371 VDD.n4316 1084.97
R11054 VDD.n4513 VDD.n4316 1084.97
R11055 VDD.n4513 VDD.n4512 1084.97
R11056 VDD.n4512 VDD.n4371 1084.97
R11057 VDD.n4395 VDD.n4314 1084.97
R11058 VDD.n4396 VDD.n4314 1084.97
R11059 VDD.n4399 VDD.n4396 1084.97
R11060 VDD.n4399 VDD.n4395 1084.97
R11061 VDD.n4526 VDD.n4359 1084.97
R11062 VDD.n4359 VDD.n4357 1084.97
R11063 VDD.n4358 VDD.n4357 1084.97
R11064 VDD.n4526 VDD.n4358 1084.97
R11065 VDD.n5031 VDD.n4560 1084.97
R11066 VDD.n5029 VDD.n4559 1084.97
R11067 VDD.n5031 VDD.n4559 1084.97
R11068 VDD.n5025 VDD.n4561 1084.97
R11069 VDD.n5025 VDD.n4562 1084.97
R11070 VDD.n5021 VDD.n4562 1084.97
R11071 VDD.n5021 VDD.n4561 1084.97
R11072 VDD.n5018 VDD.n4564 1084.97
R11073 VDD.n5014 VDD.n4565 1084.97
R11074 VDD.n5018 VDD.n4565 1084.97
R11075 VDD.n5006 VDD.n4571 1084.97
R11076 VDD.n5004 VDD.n4570 1084.97
R11077 VDD.n5006 VDD.n4570 1084.97
R11078 VDD.n5000 VDD.n4572 1084.97
R11079 VDD.n4996 VDD.n4573 1084.97
R11080 VDD.n5000 VDD.n4573 1084.97
R11081 VDD.n4990 VDD.n4579 1084.97
R11082 VDD.n4988 VDD.n4578 1084.97
R11083 VDD.n4990 VDD.n4578 1084.97
R11084 VDD.n4984 VDD.n4580 1084.97
R11085 VDD.n4984 VDD.n4581 1084.97
R11086 VDD.n4980 VDD.n4581 1084.97
R11087 VDD.n4980 VDD.n4580 1084.97
R11088 VDD.n4977 VDD.n4583 1084.97
R11089 VDD.n4973 VDD.n4584 1084.97
R11090 VDD.n4977 VDD.n4584 1084.97
R11091 VDD.n4965 VDD.n4590 1084.97
R11092 VDD.n4963 VDD.n4589 1084.97
R11093 VDD.n4965 VDD.n4589 1084.97
R11094 VDD.n4959 VDD.n4591 1084.97
R11095 VDD.n4955 VDD.n4592 1084.97
R11096 VDD.n4959 VDD.n4592 1084.97
R11097 VDD.n4949 VDD.n4598 1084.97
R11098 VDD.n4947 VDD.n4597 1084.97
R11099 VDD.n4949 VDD.n4597 1084.97
R11100 VDD.n4943 VDD.n4599 1084.97
R11101 VDD.n4943 VDD.n4600 1084.97
R11102 VDD.n4939 VDD.n4600 1084.97
R11103 VDD.n4939 VDD.n4599 1084.97
R11104 VDD.n4936 VDD.n4602 1084.97
R11105 VDD.n4932 VDD.n4603 1084.97
R11106 VDD.n4936 VDD.n4603 1084.97
R11107 VDD.n4924 VDD.n4609 1084.97
R11108 VDD.n4922 VDD.n4608 1084.97
R11109 VDD.n4924 VDD.n4608 1084.97
R11110 VDD.n4918 VDD.n4610 1084.97
R11111 VDD.n4914 VDD.n4611 1084.97
R11112 VDD.n4918 VDD.n4611 1084.97
R11113 VDD.n4908 VDD.n4617 1084.97
R11114 VDD.n4906 VDD.n4616 1084.97
R11115 VDD.n4908 VDD.n4616 1084.97
R11116 VDD.n4902 VDD.n4618 1084.97
R11117 VDD.n4902 VDD.n4619 1084.97
R11118 VDD.n4898 VDD.n4619 1084.97
R11119 VDD.n4898 VDD.n4618 1084.97
R11120 VDD.n4895 VDD.n4621 1084.97
R11121 VDD.n4891 VDD.n4622 1084.97
R11122 VDD.n4895 VDD.n4622 1084.97
R11123 VDD.n4883 VDD.n4628 1084.97
R11124 VDD.n4881 VDD.n4627 1084.97
R11125 VDD.n4883 VDD.n4627 1084.97
R11126 VDD.n4877 VDD.n4629 1084.97
R11127 VDD.n4873 VDD.n4630 1084.97
R11128 VDD.n4877 VDD.n4630 1084.97
R11129 VDD.n4867 VDD.n4636 1084.97
R11130 VDD.n4865 VDD.n4635 1084.97
R11131 VDD.n4867 VDD.n4635 1084.97
R11132 VDD.n4861 VDD.n4637 1084.97
R11133 VDD.n4861 VDD.n4638 1084.97
R11134 VDD.n4857 VDD.n4638 1084.97
R11135 VDD.n4857 VDD.n4637 1084.97
R11136 VDD.n4854 VDD.n4640 1084.97
R11137 VDD.n4850 VDD.n4641 1084.97
R11138 VDD.n4854 VDD.n4641 1084.97
R11139 VDD.n4842 VDD.n4647 1084.97
R11140 VDD.n4840 VDD.n4646 1084.97
R11141 VDD.n4842 VDD.n4646 1084.97
R11142 VDD.n4836 VDD.n4648 1084.97
R11143 VDD.n4832 VDD.n4649 1084.97
R11144 VDD.n4836 VDD.n4649 1084.97
R11145 VDD.n4826 VDD.n4655 1084.97
R11146 VDD.n4824 VDD.n4654 1084.97
R11147 VDD.n4826 VDD.n4654 1084.97
R11148 VDD.n4820 VDD.n4656 1084.97
R11149 VDD.n4820 VDD.n4657 1084.97
R11150 VDD.n4816 VDD.n4657 1084.97
R11151 VDD.n4816 VDD.n4656 1084.97
R11152 VDD.n4813 VDD.n4659 1084.97
R11153 VDD.n4809 VDD.n4660 1084.97
R11154 VDD.n4813 VDD.n4660 1084.97
R11155 VDD.n4801 VDD.n4666 1084.97
R11156 VDD.n4799 VDD.n4665 1084.97
R11157 VDD.n4801 VDD.n4665 1084.97
R11158 VDD.n4795 VDD.n4667 1084.97
R11159 VDD.n4791 VDD.n4668 1084.97
R11160 VDD.n4795 VDD.n4668 1084.97
R11161 VDD.n4785 VDD.n4674 1084.97
R11162 VDD.n4783 VDD.n4673 1084.97
R11163 VDD.n4785 VDD.n4673 1084.97
R11164 VDD.n4779 VDD.n4675 1084.97
R11165 VDD.n4779 VDD.n4676 1084.97
R11166 VDD.n4775 VDD.n4676 1084.97
R11167 VDD.n4775 VDD.n4675 1084.97
R11168 VDD.n4772 VDD.n4678 1084.97
R11169 VDD.n4768 VDD.n4679 1084.97
R11170 VDD.n4772 VDD.n4679 1084.97
R11171 VDD.n4760 VDD.n4685 1084.97
R11172 VDD.n4758 VDD.n4684 1084.97
R11173 VDD.n4760 VDD.n4684 1084.97
R11174 VDD.n4754 VDD.n4686 1084.97
R11175 VDD.n4750 VDD.n4687 1084.97
R11176 VDD.n4754 VDD.n4687 1084.97
R11177 VDD.n4744 VDD.n4693 1084.97
R11178 VDD.n4742 VDD.n4692 1084.97
R11179 VDD.n4744 VDD.n4692 1084.97
R11180 VDD.n4738 VDD.n4694 1084.97
R11181 VDD.n4738 VDD.n4695 1084.97
R11182 VDD.n4734 VDD.n4695 1084.97
R11183 VDD.n4734 VDD.n4694 1084.97
R11184 VDD.n4731 VDD.n4697 1084.97
R11185 VDD.n4727 VDD.n4698 1084.97
R11186 VDD.n4731 VDD.n4698 1084.97
R11187 VDD.n4719 VDD.n4704 1084.97
R11188 VDD.n4717 VDD.n4703 1084.97
R11189 VDD.n4719 VDD.n4703 1084.97
R11190 VDD.n4713 VDD.n4705 1084.97
R11191 VDD.n4709 VDD.n4706 1084.97
R11192 VDD.n4713 VDD.n4706 1084.97
R11193 VDD.n7101 VDD.n5038 1084.97
R11194 VDD.n7098 VDD.n5036 1084.97
R11195 VDD.n7098 VDD.n5038 1084.97
R11196 VDD.n7096 VDD.n5040 1084.97
R11197 VDD.n7096 VDD.n5041 1084.97
R11198 VDD.n7089 VDD.n5041 1084.97
R11199 VDD.n7089 VDD.n5040 1084.97
R11200 VDD.n7086 VDD.n5051 1084.97
R11201 VDD.n7086 VDD.n5052 1084.97
R11202 VDD.n7079 VDD.n5052 1084.97
R11203 VDD.n7079 VDD.n5051 1084.97
R11204 VDD.n7076 VDD.n5061 1084.97
R11205 VDD.n7076 VDD.n5062 1084.97
R11206 VDD.n7069 VDD.n5062 1084.97
R11207 VDD.n7069 VDD.n5061 1084.97
R11208 VDD.n7066 VDD.n5074 1084.97
R11209 VDD.n7066 VDD.n5075 1084.97
R11210 VDD.n7059 VDD.n5075 1084.97
R11211 VDD.n7059 VDD.n5074 1084.97
R11212 VDD.n7056 VDD.n5085 1084.97
R11213 VDD.n7056 VDD.n5086 1084.97
R11214 VDD.n7049 VDD.n5086 1084.97
R11215 VDD.n7049 VDD.n5085 1084.97
R11216 VDD.n7046 VDD.n5095 1084.97
R11217 VDD.n7046 VDD.n5096 1084.97
R11218 VDD.n7039 VDD.n5096 1084.97
R11219 VDD.n7039 VDD.n5095 1084.97
R11220 VDD.n7029 VDD.n5111 1084.97
R11221 VDD.n7029 VDD.n5112 1084.97
R11222 VDD.n7022 VDD.n5112 1084.97
R11223 VDD.n7022 VDD.n5111 1084.97
R11224 VDD.n7019 VDD.n5123 1084.97
R11225 VDD.n7019 VDD.n5124 1084.97
R11226 VDD.n7012 VDD.n5124 1084.97
R11227 VDD.n7012 VDD.n5123 1084.97
R11228 VDD.n7009 VDD.n5136 1084.97
R11229 VDD.n7009 VDD.n5137 1084.97
R11230 VDD.n7002 VDD.n5137 1084.97
R11231 VDD.n7002 VDD.n5136 1084.97
R11232 VDD.n6999 VDD.n5147 1084.97
R11233 VDD.n6999 VDD.n5148 1084.97
R11234 VDD.n6992 VDD.n5148 1084.97
R11235 VDD.n6992 VDD.n5147 1084.97
R11236 VDD.n6989 VDD.n5157 1084.97
R11237 VDD.n6989 VDD.n5158 1084.97
R11238 VDD.n6982 VDD.n5158 1084.97
R11239 VDD.n6982 VDD.n5157 1084.97
R11240 VDD.n6979 VDD.n5169 1084.97
R11241 VDD.n6979 VDD.n5170 1084.97
R11242 VDD.n6962 VDD.n5170 1084.97
R11243 VDD.n6962 VDD.n5169 1084.97
R11244 VDD.n6970 VDD.n6966 1084.97
R11245 VDD.n6966 VDD.n5175 1084.97
R11246 VDD.n6965 VDD.n5175 1084.97
R11247 VDD.n6970 VDD.n6965 1084.97
R11248 VDD.n6955 VDD.n5180 1084.97
R11249 VDD.n6955 VDD.n5181 1084.97
R11250 VDD.n6948 VDD.n5181 1084.97
R11251 VDD.n6948 VDD.n5180 1084.97
R11252 VDD.n6945 VDD.n5189 1084.97
R11253 VDD.n6945 VDD.n5190 1084.97
R11254 VDD.n6938 VDD.n5190 1084.97
R11255 VDD.n6938 VDD.n5189 1084.97
R11256 VDD.n6935 VDD.n5202 1084.97
R11257 VDD.n6935 VDD.n5203 1084.97
R11258 VDD.n6928 VDD.n5203 1084.97
R11259 VDD.n6928 VDD.n5202 1084.97
R11260 VDD.n6925 VDD.n5213 1084.97
R11261 VDD.n6925 VDD.n5214 1084.97
R11262 VDD.n6918 VDD.n5214 1084.97
R11263 VDD.n6918 VDD.n5213 1084.97
R11264 VDD.n6915 VDD.n5223 1084.97
R11265 VDD.n6915 VDD.n5224 1084.97
R11266 VDD.n6908 VDD.n5224 1084.97
R11267 VDD.n6908 VDD.n5223 1084.97
R11268 VDD.n6898 VDD.n5239 1084.97
R11269 VDD.n6898 VDD.n5240 1084.97
R11270 VDD.n6891 VDD.n5240 1084.97
R11271 VDD.n6891 VDD.n5239 1084.97
R11272 VDD.n6888 VDD.n5251 1084.97
R11273 VDD.n6888 VDD.n5252 1084.97
R11274 VDD.n6881 VDD.n5252 1084.97
R11275 VDD.n6881 VDD.n5251 1084.97
R11276 VDD.n6878 VDD.n5264 1084.97
R11277 VDD.n6878 VDD.n5265 1084.97
R11278 VDD.n6871 VDD.n5265 1084.97
R11279 VDD.n6871 VDD.n5264 1084.97
R11280 VDD.n6868 VDD.n5275 1084.97
R11281 VDD.n6868 VDD.n5276 1084.97
R11282 VDD.n6861 VDD.n5276 1084.97
R11283 VDD.n6861 VDD.n5275 1084.97
R11284 VDD.n6858 VDD.n5285 1084.97
R11285 VDD.n6858 VDD.n5286 1084.97
R11286 VDD.n6851 VDD.n5286 1084.97
R11287 VDD.n6851 VDD.n5285 1084.97
R11288 VDD.n6848 VDD.n5297 1084.97
R11289 VDD.n6848 VDD.n5298 1084.97
R11290 VDD.n6831 VDD.n5298 1084.97
R11291 VDD.n6831 VDD.n5297 1084.97
R11292 VDD.n6839 VDD.n6835 1084.97
R11293 VDD.n6835 VDD.n5303 1084.97
R11294 VDD.n6834 VDD.n5303 1084.97
R11295 VDD.n6839 VDD.n6834 1084.97
R11296 VDD.n6824 VDD.n5308 1084.97
R11297 VDD.n6824 VDD.n5309 1084.97
R11298 VDD.n6817 VDD.n5309 1084.97
R11299 VDD.n6817 VDD.n5308 1084.97
R11300 VDD.n6814 VDD.n5317 1084.97
R11301 VDD.n6814 VDD.n5318 1084.97
R11302 VDD.n6807 VDD.n5318 1084.97
R11303 VDD.n6807 VDD.n5317 1084.97
R11304 VDD.n6804 VDD.n5330 1084.97
R11305 VDD.n6804 VDD.n5331 1084.97
R11306 VDD.n6797 VDD.n5331 1084.97
R11307 VDD.n6797 VDD.n5330 1084.97
R11308 VDD.n6794 VDD.n5341 1084.97
R11309 VDD.n6794 VDD.n5342 1084.97
R11310 VDD.n6787 VDD.n5342 1084.97
R11311 VDD.n6787 VDD.n5341 1084.97
R11312 VDD.n6784 VDD.n5351 1084.97
R11313 VDD.n6784 VDD.n5352 1084.97
R11314 VDD.n6777 VDD.n5352 1084.97
R11315 VDD.n6777 VDD.n5351 1084.97
R11316 VDD.n6767 VDD.n5367 1084.97
R11317 VDD.n6767 VDD.n5368 1084.97
R11318 VDD.n6760 VDD.n5368 1084.97
R11319 VDD.n6760 VDD.n5367 1084.97
R11320 VDD.n6757 VDD.n5379 1084.97
R11321 VDD.n6757 VDD.n5380 1084.97
R11322 VDD.n6750 VDD.n5380 1084.97
R11323 VDD.n6750 VDD.n5379 1084.97
R11324 VDD.n6747 VDD.n5392 1084.97
R11325 VDD.n6747 VDD.n5393 1084.97
R11326 VDD.n6740 VDD.n5393 1084.97
R11327 VDD.n6740 VDD.n5392 1084.97
R11328 VDD.n6737 VDD.n5403 1084.97
R11329 VDD.n6737 VDD.n5404 1084.97
R11330 VDD.n6730 VDD.n5404 1084.97
R11331 VDD.n6730 VDD.n5403 1084.97
R11332 VDD.n6727 VDD.n5413 1084.97
R11333 VDD.n6727 VDD.n5414 1084.97
R11334 VDD.n6720 VDD.n5414 1084.97
R11335 VDD.n6720 VDD.n5413 1084.97
R11336 VDD.n6717 VDD.n5425 1084.97
R11337 VDD.n6717 VDD.n5426 1084.97
R11338 VDD.n6700 VDD.n5426 1084.97
R11339 VDD.n6700 VDD.n5425 1084.97
R11340 VDD.n6708 VDD.n6704 1084.97
R11341 VDD.n6704 VDD.n5431 1084.97
R11342 VDD.n6703 VDD.n5431 1084.97
R11343 VDD.n6708 VDD.n6703 1084.97
R11344 VDD.n6693 VDD.n5436 1084.97
R11345 VDD.n6693 VDD.n5437 1084.97
R11346 VDD.n6686 VDD.n5437 1084.97
R11347 VDD.n6686 VDD.n5436 1084.97
R11348 VDD.n6683 VDD.n5445 1084.97
R11349 VDD.n6683 VDD.n5446 1084.97
R11350 VDD.n6676 VDD.n5446 1084.97
R11351 VDD.n6676 VDD.n5445 1084.97
R11352 VDD.n6673 VDD.n5458 1084.97
R11353 VDD.n6673 VDD.n5459 1084.97
R11354 VDD.n6666 VDD.n5459 1084.97
R11355 VDD.n6666 VDD.n5458 1084.97
R11356 VDD.n6663 VDD.n5469 1084.97
R11357 VDD.n6663 VDD.n5470 1084.97
R11358 VDD.n6656 VDD.n5470 1084.97
R11359 VDD.n6656 VDD.n5469 1084.97
R11360 VDD.n6653 VDD.n5479 1084.97
R11361 VDD.n6653 VDD.n5480 1084.97
R11362 VDD.n6646 VDD.n5480 1084.97
R11363 VDD.n6646 VDD.n5479 1084.97
R11364 VDD.n6636 VDD.n5495 1084.97
R11365 VDD.n6636 VDD.n5496 1084.97
R11366 VDD.n6629 VDD.n5496 1084.97
R11367 VDD.n6629 VDD.n5495 1084.97
R11368 VDD.n6626 VDD.n5507 1084.97
R11369 VDD.n6626 VDD.n5508 1084.97
R11370 VDD.n6619 VDD.n5508 1084.97
R11371 VDD.n6619 VDD.n5507 1084.97
R11372 VDD.n6616 VDD.n5520 1084.97
R11373 VDD.n6616 VDD.n5521 1084.97
R11374 VDD.n6609 VDD.n5521 1084.97
R11375 VDD.n6609 VDD.n5520 1084.97
R11376 VDD.n6606 VDD.n5531 1084.97
R11377 VDD.n6606 VDD.n5532 1084.97
R11378 VDD.n6599 VDD.n5532 1084.97
R11379 VDD.n6599 VDD.n5531 1084.97
R11380 VDD.n6596 VDD.n5541 1084.97
R11381 VDD.n6596 VDD.n5542 1084.97
R11382 VDD.n6589 VDD.n5542 1084.97
R11383 VDD.n6589 VDD.n5541 1084.97
R11384 VDD.n6586 VDD.n5553 1084.97
R11385 VDD.n6586 VDD.n5554 1084.97
R11386 VDD.n6569 VDD.n5554 1084.97
R11387 VDD.n6569 VDD.n5553 1084.97
R11388 VDD.n6577 VDD.n6573 1084.97
R11389 VDD.n6573 VDD.n5559 1084.97
R11390 VDD.n6572 VDD.n5559 1084.97
R11391 VDD.n6577 VDD.n6572 1084.97
R11392 VDD.n6562 VDD.n5564 1084.97
R11393 VDD.n6562 VDD.n5565 1084.97
R11394 VDD.n6555 VDD.n5565 1084.97
R11395 VDD.n6555 VDD.n5564 1084.97
R11396 VDD.n6552 VDD.n5573 1084.97
R11397 VDD.n6552 VDD.n5574 1084.97
R11398 VDD.n6545 VDD.n5574 1084.97
R11399 VDD.n6545 VDD.n5573 1084.97
R11400 VDD.n6542 VDD.n5586 1084.97
R11401 VDD.n6542 VDD.n5587 1084.97
R11402 VDD.n6535 VDD.n5587 1084.97
R11403 VDD.n6535 VDD.n5586 1084.97
R11404 VDD.n6532 VDD.n5597 1084.97
R11405 VDD.n6532 VDD.n5598 1084.97
R11406 VDD.n6525 VDD.n5598 1084.97
R11407 VDD.n6525 VDD.n5597 1084.97
R11408 VDD.n6522 VDD.n5607 1084.97
R11409 VDD.n6522 VDD.n5608 1084.97
R11410 VDD.n6515 VDD.n5608 1084.97
R11411 VDD.n6515 VDD.n5607 1084.97
R11412 VDD.n6505 VDD.n5623 1084.97
R11413 VDD.n6505 VDD.n5624 1084.97
R11414 VDD.n6498 VDD.n5624 1084.97
R11415 VDD.n6498 VDD.n5623 1084.97
R11416 VDD.n6495 VDD.n5635 1084.97
R11417 VDD.n6495 VDD.n5636 1084.97
R11418 VDD.n6488 VDD.n5636 1084.97
R11419 VDD.n6488 VDD.n5635 1084.97
R11420 VDD.n6485 VDD.n5648 1084.97
R11421 VDD.n6485 VDD.n5649 1084.97
R11422 VDD.n6478 VDD.n5649 1084.97
R11423 VDD.n6478 VDD.n5648 1084.97
R11424 VDD.n6475 VDD.n5659 1084.97
R11425 VDD.n6475 VDD.n5660 1084.97
R11426 VDD.n6468 VDD.n5660 1084.97
R11427 VDD.n6468 VDD.n5659 1084.97
R11428 VDD.n6465 VDD.n5669 1084.97
R11429 VDD.n6465 VDD.n5670 1084.97
R11430 VDD.n6458 VDD.n5670 1084.97
R11431 VDD.n6458 VDD.n5669 1084.97
R11432 VDD.n6455 VDD.n5681 1084.97
R11433 VDD.n6455 VDD.n5682 1084.97
R11434 VDD.n6438 VDD.n5682 1084.97
R11435 VDD.n6438 VDD.n5681 1084.97
R11436 VDD.n6446 VDD.n6442 1084.97
R11437 VDD.n6442 VDD.n5687 1084.97
R11438 VDD.n6441 VDD.n5687 1084.97
R11439 VDD.n6446 VDD.n6441 1084.97
R11440 VDD.n6431 VDD.n5692 1084.97
R11441 VDD.n6431 VDD.n5693 1084.97
R11442 VDD.n6424 VDD.n5693 1084.97
R11443 VDD.n6424 VDD.n5692 1084.97
R11444 VDD.n6421 VDD.n5701 1084.97
R11445 VDD.n6421 VDD.n5702 1084.97
R11446 VDD.n6414 VDD.n5702 1084.97
R11447 VDD.n6414 VDD.n5701 1084.97
R11448 VDD.n6411 VDD.n5714 1084.97
R11449 VDD.n6411 VDD.n5715 1084.97
R11450 VDD.n6404 VDD.n5715 1084.97
R11451 VDD.n6404 VDD.n5714 1084.97
R11452 VDD.n6401 VDD.n5725 1084.97
R11453 VDD.n6401 VDD.n5726 1084.97
R11454 VDD.n6394 VDD.n5726 1084.97
R11455 VDD.n6394 VDD.n5725 1084.97
R11456 VDD.n6391 VDD.n5735 1084.97
R11457 VDD.n6391 VDD.n5736 1084.97
R11458 VDD.n6384 VDD.n5736 1084.97
R11459 VDD.n6384 VDD.n5735 1084.97
R11460 VDD.n6374 VDD.n5751 1084.97
R11461 VDD.n6374 VDD.n5752 1084.97
R11462 VDD.n6367 VDD.n5752 1084.97
R11463 VDD.n6367 VDD.n5751 1084.97
R11464 VDD.n6364 VDD.n5763 1084.97
R11465 VDD.n6364 VDD.n5764 1084.97
R11466 VDD.n6357 VDD.n5764 1084.97
R11467 VDD.n6357 VDD.n5763 1084.97
R11468 VDD.n6354 VDD.n5776 1084.97
R11469 VDD.n6354 VDD.n5777 1084.97
R11470 VDD.n6347 VDD.n5777 1084.97
R11471 VDD.n6347 VDD.n5776 1084.97
R11472 VDD.n6344 VDD.n5787 1084.97
R11473 VDD.n6344 VDD.n5788 1084.97
R11474 VDD.n6337 VDD.n5788 1084.97
R11475 VDD.n6337 VDD.n5787 1084.97
R11476 VDD.n6334 VDD.n5797 1084.97
R11477 VDD.n6334 VDD.n5798 1084.97
R11478 VDD.n6327 VDD.n5798 1084.97
R11479 VDD.n6327 VDD.n5797 1084.97
R11480 VDD.n6324 VDD.n5809 1084.97
R11481 VDD.n6324 VDD.n5810 1084.97
R11482 VDD.n6307 VDD.n5810 1084.97
R11483 VDD.n6307 VDD.n5809 1084.97
R11484 VDD.n6315 VDD.n6311 1084.97
R11485 VDD.n6311 VDD.n5815 1084.97
R11486 VDD.n6310 VDD.n5815 1084.97
R11487 VDD.n6315 VDD.n6310 1084.97
R11488 VDD.n6300 VDD.n5820 1084.97
R11489 VDD.n6300 VDD.n5821 1084.97
R11490 VDD.n6293 VDD.n5821 1084.97
R11491 VDD.n6293 VDD.n5820 1084.97
R11492 VDD.n6290 VDD.n5829 1084.97
R11493 VDD.n6290 VDD.n5830 1084.97
R11494 VDD.n6283 VDD.n5830 1084.97
R11495 VDD.n6283 VDD.n5829 1084.97
R11496 VDD.n6280 VDD.n5842 1084.97
R11497 VDD.n6280 VDD.n5843 1084.97
R11498 VDD.n6273 VDD.n5843 1084.97
R11499 VDD.n6273 VDD.n5842 1084.97
R11500 VDD.n6270 VDD.n5853 1084.97
R11501 VDD.n6270 VDD.n5854 1084.97
R11502 VDD.n6263 VDD.n5854 1084.97
R11503 VDD.n6263 VDD.n5853 1084.97
R11504 VDD.n6260 VDD.n5863 1084.97
R11505 VDD.n6260 VDD.n5864 1084.97
R11506 VDD.n6253 VDD.n5864 1084.97
R11507 VDD.n6253 VDD.n5863 1084.97
R11508 VDD.n6243 VDD.n5879 1084.97
R11509 VDD.n6243 VDD.n5880 1084.97
R11510 VDD.n6236 VDD.n5880 1084.97
R11511 VDD.n6236 VDD.n5879 1084.97
R11512 VDD.n6233 VDD.n5891 1084.97
R11513 VDD.n6233 VDD.n5892 1084.97
R11514 VDD.n6226 VDD.n5892 1084.97
R11515 VDD.n6226 VDD.n5891 1084.97
R11516 VDD.n6223 VDD.n5904 1084.97
R11517 VDD.n6223 VDD.n5905 1084.97
R11518 VDD.n6216 VDD.n5905 1084.97
R11519 VDD.n6216 VDD.n5904 1084.97
R11520 VDD.n6213 VDD.n5915 1084.97
R11521 VDD.n6213 VDD.n5916 1084.97
R11522 VDD.n6206 VDD.n5916 1084.97
R11523 VDD.n6206 VDD.n5915 1084.97
R11524 VDD.n6203 VDD.n5925 1084.97
R11525 VDD.n6203 VDD.n5926 1084.97
R11526 VDD.n6196 VDD.n5926 1084.97
R11527 VDD.n6196 VDD.n5925 1084.97
R11528 VDD.n6193 VDD.n5937 1084.97
R11529 VDD.n6193 VDD.n5938 1084.97
R11530 VDD.n6176 VDD.n5938 1084.97
R11531 VDD.n6176 VDD.n5937 1084.97
R11532 VDD.n6184 VDD.n6180 1084.97
R11533 VDD.n6180 VDD.n5943 1084.97
R11534 VDD.n6179 VDD.n5943 1084.97
R11535 VDD.n6184 VDD.n6179 1084.97
R11536 VDD.n6169 VDD.n5948 1084.97
R11537 VDD.n6169 VDD.n5949 1084.97
R11538 VDD.n6162 VDD.n5949 1084.97
R11539 VDD.n6162 VDD.n5948 1084.97
R11540 VDD.n6159 VDD.n5957 1084.97
R11541 VDD.n6159 VDD.n5958 1084.97
R11542 VDD.n6152 VDD.n5958 1084.97
R11543 VDD.n6152 VDD.n5957 1084.97
R11544 VDD.n6149 VDD.n5970 1084.97
R11545 VDD.n6149 VDD.n5971 1084.97
R11546 VDD.n6142 VDD.n5971 1084.97
R11547 VDD.n6142 VDD.n5970 1084.97
R11548 VDD.n6139 VDD.n5981 1084.97
R11549 VDD.n6139 VDD.n5982 1084.97
R11550 VDD.n6132 VDD.n5982 1084.97
R11551 VDD.n6132 VDD.n5981 1084.97
R11552 VDD.n6129 VDD.n5991 1084.97
R11553 VDD.n6129 VDD.n5992 1084.97
R11554 VDD.n6122 VDD.n5992 1084.97
R11555 VDD.n6122 VDD.n5991 1084.97
R11556 VDD.n6112 VDD.n6007 1084.97
R11557 VDD.n6112 VDD.n6008 1084.97
R11558 VDD.n6105 VDD.n6008 1084.97
R11559 VDD.n6105 VDD.n6007 1084.97
R11560 VDD.n6102 VDD.n6019 1084.97
R11561 VDD.n6102 VDD.n6020 1084.97
R11562 VDD.n6095 VDD.n6020 1084.97
R11563 VDD.n6095 VDD.n6019 1084.97
R11564 VDD.n6092 VDD.n6032 1084.97
R11565 VDD.n6092 VDD.n6033 1084.97
R11566 VDD.n6085 VDD.n6033 1084.97
R11567 VDD.n6085 VDD.n6032 1084.97
R11568 VDD.n6082 VDD.n6043 1084.97
R11569 VDD.n6082 VDD.n6044 1084.97
R11570 VDD.n6075 VDD.n6044 1084.97
R11571 VDD.n6075 VDD.n6043 1084.97
R11572 VDD.n7092 VDD.n5039 1084.97
R11573 VDD.n5047 VDD.n5039 1084.97
R11574 VDD.n7091 VDD.n5047 1084.97
R11575 VDD.n7092 VDD.n7091 1084.97
R11576 VDD.n7082 VDD.n5050 1084.97
R11577 VDD.n5057 VDD.n5050 1084.97
R11578 VDD.n7081 VDD.n5057 1084.97
R11579 VDD.n7082 VDD.n7081 1084.97
R11580 VDD.n7072 VDD.n5060 1084.97
R11581 VDD.n5070 VDD.n5060 1084.97
R11582 VDD.n7071 VDD.n5070 1084.97
R11583 VDD.n7072 VDD.n7071 1084.97
R11584 VDD.n7062 VDD.n5073 1084.97
R11585 VDD.n5081 VDD.n5073 1084.97
R11586 VDD.n7061 VDD.n5081 1084.97
R11587 VDD.n7062 VDD.n7061 1084.97
R11588 VDD.n7052 VDD.n5084 1084.97
R11589 VDD.n5091 VDD.n5084 1084.97
R11590 VDD.n7051 VDD.n5091 1084.97
R11591 VDD.n7052 VDD.n7051 1084.97
R11592 VDD.n7042 VDD.n5094 1084.97
R11593 VDD.n5104 VDD.n5094 1084.97
R11594 VDD.n7041 VDD.n5104 1084.97
R11595 VDD.n7042 VDD.n7041 1084.97
R11596 VDD.n7036 VDD.n5107 1084.97
R11597 VDD.n7036 VDD.n5108 1084.97
R11598 VDD.n7032 VDD.n5108 1084.97
R11599 VDD.n7032 VDD.n5107 1084.97
R11600 VDD.n7025 VDD.n5110 1084.97
R11601 VDD.n5119 VDD.n5110 1084.97
R11602 VDD.n7024 VDD.n5119 1084.97
R11603 VDD.n7025 VDD.n7024 1084.97
R11604 VDD.n7015 VDD.n5122 1084.97
R11605 VDD.n5132 VDD.n5122 1084.97
R11606 VDD.n7014 VDD.n5132 1084.97
R11607 VDD.n7015 VDD.n7014 1084.97
R11608 VDD.n7005 VDD.n5135 1084.97
R11609 VDD.n5143 VDD.n5135 1084.97
R11610 VDD.n7004 VDD.n5143 1084.97
R11611 VDD.n7005 VDD.n7004 1084.97
R11612 VDD.n6995 VDD.n5146 1084.97
R11613 VDD.n5153 VDD.n5146 1084.97
R11614 VDD.n6994 VDD.n5153 1084.97
R11615 VDD.n6995 VDD.n6994 1084.97
R11616 VDD.n6985 VDD.n5156 1084.97
R11617 VDD.n5166 VDD.n5156 1084.97
R11618 VDD.n6984 VDD.n5166 1084.97
R11619 VDD.n6985 VDD.n6984 1084.97
R11620 VDD.n6971 VDD.n5178 1084.97
R11621 VDD.n6961 VDD.n5178 1084.97
R11622 VDD.n6961 VDD.n5177 1084.97
R11623 VDD.n6971 VDD.n5177 1084.97
R11624 VDD.n6951 VDD.n5179 1084.97
R11625 VDD.n5185 VDD.n5179 1084.97
R11626 VDD.n6950 VDD.n5185 1084.97
R11627 VDD.n6951 VDD.n6950 1084.97
R11628 VDD.n6941 VDD.n5188 1084.97
R11629 VDD.n5198 VDD.n5188 1084.97
R11630 VDD.n6940 VDD.n5198 1084.97
R11631 VDD.n6941 VDD.n6940 1084.97
R11632 VDD.n6931 VDD.n5201 1084.97
R11633 VDD.n5209 VDD.n5201 1084.97
R11634 VDD.n6930 VDD.n5209 1084.97
R11635 VDD.n6931 VDD.n6930 1084.97
R11636 VDD.n6921 VDD.n5212 1084.97
R11637 VDD.n5219 VDD.n5212 1084.97
R11638 VDD.n6920 VDD.n5219 1084.97
R11639 VDD.n6921 VDD.n6920 1084.97
R11640 VDD.n6911 VDD.n5222 1084.97
R11641 VDD.n5232 VDD.n5222 1084.97
R11642 VDD.n6910 VDD.n5232 1084.97
R11643 VDD.n6911 VDD.n6910 1084.97
R11644 VDD.n6905 VDD.n5235 1084.97
R11645 VDD.n6905 VDD.n5236 1084.97
R11646 VDD.n6901 VDD.n5236 1084.97
R11647 VDD.n6901 VDD.n5235 1084.97
R11648 VDD.n6894 VDD.n5238 1084.97
R11649 VDD.n5247 VDD.n5238 1084.97
R11650 VDD.n6893 VDD.n5247 1084.97
R11651 VDD.n6894 VDD.n6893 1084.97
R11652 VDD.n6884 VDD.n5250 1084.97
R11653 VDD.n5260 VDD.n5250 1084.97
R11654 VDD.n6883 VDD.n5260 1084.97
R11655 VDD.n6884 VDD.n6883 1084.97
R11656 VDD.n6874 VDD.n5263 1084.97
R11657 VDD.n5271 VDD.n5263 1084.97
R11658 VDD.n6873 VDD.n5271 1084.97
R11659 VDD.n6874 VDD.n6873 1084.97
R11660 VDD.n6864 VDD.n5274 1084.97
R11661 VDD.n5281 VDD.n5274 1084.97
R11662 VDD.n6863 VDD.n5281 1084.97
R11663 VDD.n6864 VDD.n6863 1084.97
R11664 VDD.n6854 VDD.n5284 1084.97
R11665 VDD.n5294 VDD.n5284 1084.97
R11666 VDD.n6853 VDD.n5294 1084.97
R11667 VDD.n6854 VDD.n6853 1084.97
R11668 VDD.n6840 VDD.n5306 1084.97
R11669 VDD.n6830 VDD.n5306 1084.97
R11670 VDD.n6830 VDD.n5305 1084.97
R11671 VDD.n6840 VDD.n5305 1084.97
R11672 VDD.n6820 VDD.n5307 1084.97
R11673 VDD.n5313 VDD.n5307 1084.97
R11674 VDD.n6819 VDD.n5313 1084.97
R11675 VDD.n6820 VDD.n6819 1084.97
R11676 VDD.n6810 VDD.n5316 1084.97
R11677 VDD.n5326 VDD.n5316 1084.97
R11678 VDD.n6809 VDD.n5326 1084.97
R11679 VDD.n6810 VDD.n6809 1084.97
R11680 VDD.n6800 VDD.n5329 1084.97
R11681 VDD.n5337 VDD.n5329 1084.97
R11682 VDD.n6799 VDD.n5337 1084.97
R11683 VDD.n6800 VDD.n6799 1084.97
R11684 VDD.n6790 VDD.n5340 1084.97
R11685 VDD.n5347 VDD.n5340 1084.97
R11686 VDD.n6789 VDD.n5347 1084.97
R11687 VDD.n6790 VDD.n6789 1084.97
R11688 VDD.n6780 VDD.n5350 1084.97
R11689 VDD.n5360 VDD.n5350 1084.97
R11690 VDD.n6779 VDD.n5360 1084.97
R11691 VDD.n6780 VDD.n6779 1084.97
R11692 VDD.n6774 VDD.n5363 1084.97
R11693 VDD.n6774 VDD.n5364 1084.97
R11694 VDD.n6770 VDD.n5364 1084.97
R11695 VDD.n6770 VDD.n5363 1084.97
R11696 VDD.n6763 VDD.n5366 1084.97
R11697 VDD.n5375 VDD.n5366 1084.97
R11698 VDD.n6762 VDD.n5375 1084.97
R11699 VDD.n6763 VDD.n6762 1084.97
R11700 VDD.n6753 VDD.n5378 1084.97
R11701 VDD.n5388 VDD.n5378 1084.97
R11702 VDD.n6752 VDD.n5388 1084.97
R11703 VDD.n6753 VDD.n6752 1084.97
R11704 VDD.n6743 VDD.n5391 1084.97
R11705 VDD.n5399 VDD.n5391 1084.97
R11706 VDD.n6742 VDD.n5399 1084.97
R11707 VDD.n6743 VDD.n6742 1084.97
R11708 VDD.n6733 VDD.n5402 1084.97
R11709 VDD.n5409 VDD.n5402 1084.97
R11710 VDD.n6732 VDD.n5409 1084.97
R11711 VDD.n6733 VDD.n6732 1084.97
R11712 VDD.n6723 VDD.n5412 1084.97
R11713 VDD.n5422 VDD.n5412 1084.97
R11714 VDD.n6722 VDD.n5422 1084.97
R11715 VDD.n6723 VDD.n6722 1084.97
R11716 VDD.n6709 VDD.n5434 1084.97
R11717 VDD.n6699 VDD.n5434 1084.97
R11718 VDD.n6699 VDD.n5433 1084.97
R11719 VDD.n6709 VDD.n5433 1084.97
R11720 VDD.n6689 VDD.n5435 1084.97
R11721 VDD.n5441 VDD.n5435 1084.97
R11722 VDD.n6688 VDD.n5441 1084.97
R11723 VDD.n6689 VDD.n6688 1084.97
R11724 VDD.n6679 VDD.n5444 1084.97
R11725 VDD.n5454 VDD.n5444 1084.97
R11726 VDD.n6678 VDD.n5454 1084.97
R11727 VDD.n6679 VDD.n6678 1084.97
R11728 VDD.n6669 VDD.n5457 1084.97
R11729 VDD.n5465 VDD.n5457 1084.97
R11730 VDD.n6668 VDD.n5465 1084.97
R11731 VDD.n6669 VDD.n6668 1084.97
R11732 VDD.n6659 VDD.n5468 1084.97
R11733 VDD.n5475 VDD.n5468 1084.97
R11734 VDD.n6658 VDD.n5475 1084.97
R11735 VDD.n6659 VDD.n6658 1084.97
R11736 VDD.n6649 VDD.n5478 1084.97
R11737 VDD.n5488 VDD.n5478 1084.97
R11738 VDD.n6648 VDD.n5488 1084.97
R11739 VDD.n6649 VDD.n6648 1084.97
R11740 VDD.n6643 VDD.n5491 1084.97
R11741 VDD.n6643 VDD.n5492 1084.97
R11742 VDD.n6639 VDD.n5492 1084.97
R11743 VDD.n6639 VDD.n5491 1084.97
R11744 VDD.n6632 VDD.n5494 1084.97
R11745 VDD.n5503 VDD.n5494 1084.97
R11746 VDD.n6631 VDD.n5503 1084.97
R11747 VDD.n6632 VDD.n6631 1084.97
R11748 VDD.n6622 VDD.n5506 1084.97
R11749 VDD.n5516 VDD.n5506 1084.97
R11750 VDD.n6621 VDD.n5516 1084.97
R11751 VDD.n6622 VDD.n6621 1084.97
R11752 VDD.n6612 VDD.n5519 1084.97
R11753 VDD.n5527 VDD.n5519 1084.97
R11754 VDD.n6611 VDD.n5527 1084.97
R11755 VDD.n6612 VDD.n6611 1084.97
R11756 VDD.n6602 VDD.n5530 1084.97
R11757 VDD.n5537 VDD.n5530 1084.97
R11758 VDD.n6601 VDD.n5537 1084.97
R11759 VDD.n6602 VDD.n6601 1084.97
R11760 VDD.n6592 VDD.n5540 1084.97
R11761 VDD.n5550 VDD.n5540 1084.97
R11762 VDD.n6591 VDD.n5550 1084.97
R11763 VDD.n6592 VDD.n6591 1084.97
R11764 VDD.n6578 VDD.n5562 1084.97
R11765 VDD.n6568 VDD.n5562 1084.97
R11766 VDD.n6568 VDD.n5561 1084.97
R11767 VDD.n6578 VDD.n5561 1084.97
R11768 VDD.n6558 VDD.n5563 1084.97
R11769 VDD.n5569 VDD.n5563 1084.97
R11770 VDD.n6557 VDD.n5569 1084.97
R11771 VDD.n6558 VDD.n6557 1084.97
R11772 VDD.n6548 VDD.n5572 1084.97
R11773 VDD.n5582 VDD.n5572 1084.97
R11774 VDD.n6547 VDD.n5582 1084.97
R11775 VDD.n6548 VDD.n6547 1084.97
R11776 VDD.n6538 VDD.n5585 1084.97
R11777 VDD.n5593 VDD.n5585 1084.97
R11778 VDD.n6537 VDD.n5593 1084.97
R11779 VDD.n6538 VDD.n6537 1084.97
R11780 VDD.n6528 VDD.n5596 1084.97
R11781 VDD.n5603 VDD.n5596 1084.97
R11782 VDD.n6527 VDD.n5603 1084.97
R11783 VDD.n6528 VDD.n6527 1084.97
R11784 VDD.n6518 VDD.n5606 1084.97
R11785 VDD.n5616 VDD.n5606 1084.97
R11786 VDD.n6517 VDD.n5616 1084.97
R11787 VDD.n6518 VDD.n6517 1084.97
R11788 VDD.n6512 VDD.n5619 1084.97
R11789 VDD.n6512 VDD.n5620 1084.97
R11790 VDD.n6508 VDD.n5620 1084.97
R11791 VDD.n6508 VDD.n5619 1084.97
R11792 VDD.n6501 VDD.n5622 1084.97
R11793 VDD.n5631 VDD.n5622 1084.97
R11794 VDD.n6500 VDD.n5631 1084.97
R11795 VDD.n6501 VDD.n6500 1084.97
R11796 VDD.n6491 VDD.n5634 1084.97
R11797 VDD.n5644 VDD.n5634 1084.97
R11798 VDD.n6490 VDD.n5644 1084.97
R11799 VDD.n6491 VDD.n6490 1084.97
R11800 VDD.n6481 VDD.n5647 1084.97
R11801 VDD.n5655 VDD.n5647 1084.97
R11802 VDD.n6480 VDD.n5655 1084.97
R11803 VDD.n6481 VDD.n6480 1084.97
R11804 VDD.n6471 VDD.n5658 1084.97
R11805 VDD.n5665 VDD.n5658 1084.97
R11806 VDD.n6470 VDD.n5665 1084.97
R11807 VDD.n6471 VDD.n6470 1084.97
R11808 VDD.n6461 VDD.n5668 1084.97
R11809 VDD.n5678 VDD.n5668 1084.97
R11810 VDD.n6460 VDD.n5678 1084.97
R11811 VDD.n6461 VDD.n6460 1084.97
R11812 VDD.n6447 VDD.n5690 1084.97
R11813 VDD.n6437 VDD.n5690 1084.97
R11814 VDD.n6437 VDD.n5689 1084.97
R11815 VDD.n6447 VDD.n5689 1084.97
R11816 VDD.n6427 VDD.n5691 1084.97
R11817 VDD.n5697 VDD.n5691 1084.97
R11818 VDD.n6426 VDD.n5697 1084.97
R11819 VDD.n6427 VDD.n6426 1084.97
R11820 VDD.n6417 VDD.n5700 1084.97
R11821 VDD.n5710 VDD.n5700 1084.97
R11822 VDD.n6416 VDD.n5710 1084.97
R11823 VDD.n6417 VDD.n6416 1084.97
R11824 VDD.n6407 VDD.n5713 1084.97
R11825 VDD.n5721 VDD.n5713 1084.97
R11826 VDD.n6406 VDD.n5721 1084.97
R11827 VDD.n6407 VDD.n6406 1084.97
R11828 VDD.n6397 VDD.n5724 1084.97
R11829 VDD.n5731 VDD.n5724 1084.97
R11830 VDD.n6396 VDD.n5731 1084.97
R11831 VDD.n6397 VDD.n6396 1084.97
R11832 VDD.n6387 VDD.n5734 1084.97
R11833 VDD.n5744 VDD.n5734 1084.97
R11834 VDD.n6386 VDD.n5744 1084.97
R11835 VDD.n6387 VDD.n6386 1084.97
R11836 VDD.n6381 VDD.n5747 1084.97
R11837 VDD.n6381 VDD.n5748 1084.97
R11838 VDD.n6377 VDD.n5748 1084.97
R11839 VDD.n6377 VDD.n5747 1084.97
R11840 VDD.n6370 VDD.n5750 1084.97
R11841 VDD.n5759 VDD.n5750 1084.97
R11842 VDD.n6369 VDD.n5759 1084.97
R11843 VDD.n6370 VDD.n6369 1084.97
R11844 VDD.n6360 VDD.n5762 1084.97
R11845 VDD.n5772 VDD.n5762 1084.97
R11846 VDD.n6359 VDD.n5772 1084.97
R11847 VDD.n6360 VDD.n6359 1084.97
R11848 VDD.n6350 VDD.n5775 1084.97
R11849 VDD.n5783 VDD.n5775 1084.97
R11850 VDD.n6349 VDD.n5783 1084.97
R11851 VDD.n6350 VDD.n6349 1084.97
R11852 VDD.n6340 VDD.n5786 1084.97
R11853 VDD.n5793 VDD.n5786 1084.97
R11854 VDD.n6339 VDD.n5793 1084.97
R11855 VDD.n6340 VDD.n6339 1084.97
R11856 VDD.n6330 VDD.n5796 1084.97
R11857 VDD.n5806 VDD.n5796 1084.97
R11858 VDD.n6329 VDD.n5806 1084.97
R11859 VDD.n6330 VDD.n6329 1084.97
R11860 VDD.n6316 VDD.n5818 1084.97
R11861 VDD.n6306 VDD.n5818 1084.97
R11862 VDD.n6306 VDD.n5817 1084.97
R11863 VDD.n6316 VDD.n5817 1084.97
R11864 VDD.n6296 VDD.n5819 1084.97
R11865 VDD.n5825 VDD.n5819 1084.97
R11866 VDD.n6295 VDD.n5825 1084.97
R11867 VDD.n6296 VDD.n6295 1084.97
R11868 VDD.n6286 VDD.n5828 1084.97
R11869 VDD.n5838 VDD.n5828 1084.97
R11870 VDD.n6285 VDD.n5838 1084.97
R11871 VDD.n6286 VDD.n6285 1084.97
R11872 VDD.n6276 VDD.n5841 1084.97
R11873 VDD.n5849 VDD.n5841 1084.97
R11874 VDD.n6275 VDD.n5849 1084.97
R11875 VDD.n6276 VDD.n6275 1084.97
R11876 VDD.n6266 VDD.n5852 1084.97
R11877 VDD.n5859 VDD.n5852 1084.97
R11878 VDD.n6265 VDD.n5859 1084.97
R11879 VDD.n6266 VDD.n6265 1084.97
R11880 VDD.n6256 VDD.n5862 1084.97
R11881 VDD.n5872 VDD.n5862 1084.97
R11882 VDD.n6255 VDD.n5872 1084.97
R11883 VDD.n6256 VDD.n6255 1084.97
R11884 VDD.n6250 VDD.n5875 1084.97
R11885 VDD.n6250 VDD.n5876 1084.97
R11886 VDD.n6246 VDD.n5876 1084.97
R11887 VDD.n6246 VDD.n5875 1084.97
R11888 VDD.n6239 VDD.n5878 1084.97
R11889 VDD.n5887 VDD.n5878 1084.97
R11890 VDD.n6238 VDD.n5887 1084.97
R11891 VDD.n6239 VDD.n6238 1084.97
R11892 VDD.n6229 VDD.n5890 1084.97
R11893 VDD.n5900 VDD.n5890 1084.97
R11894 VDD.n6228 VDD.n5900 1084.97
R11895 VDD.n6229 VDD.n6228 1084.97
R11896 VDD.n6219 VDD.n5903 1084.97
R11897 VDD.n5911 VDD.n5903 1084.97
R11898 VDD.n6218 VDD.n5911 1084.97
R11899 VDD.n6219 VDD.n6218 1084.97
R11900 VDD.n6209 VDD.n5914 1084.97
R11901 VDD.n5921 VDD.n5914 1084.97
R11902 VDD.n6208 VDD.n5921 1084.97
R11903 VDD.n6209 VDD.n6208 1084.97
R11904 VDD.n6199 VDD.n5924 1084.97
R11905 VDD.n5934 VDD.n5924 1084.97
R11906 VDD.n6198 VDD.n5934 1084.97
R11907 VDD.n6199 VDD.n6198 1084.97
R11908 VDD.n6185 VDD.n5946 1084.97
R11909 VDD.n6175 VDD.n5946 1084.97
R11910 VDD.n6175 VDD.n5945 1084.97
R11911 VDD.n6185 VDD.n5945 1084.97
R11912 VDD.n6165 VDD.n5947 1084.97
R11913 VDD.n5953 VDD.n5947 1084.97
R11914 VDD.n6164 VDD.n5953 1084.97
R11915 VDD.n6165 VDD.n6164 1084.97
R11916 VDD.n6155 VDD.n5956 1084.97
R11917 VDD.n5966 VDD.n5956 1084.97
R11918 VDD.n6154 VDD.n5966 1084.97
R11919 VDD.n6155 VDD.n6154 1084.97
R11920 VDD.n6145 VDD.n5969 1084.97
R11921 VDD.n5977 VDD.n5969 1084.97
R11922 VDD.n6144 VDD.n5977 1084.97
R11923 VDD.n6145 VDD.n6144 1084.97
R11924 VDD.n6135 VDD.n5980 1084.97
R11925 VDD.n5987 VDD.n5980 1084.97
R11926 VDD.n6134 VDD.n5987 1084.97
R11927 VDD.n6135 VDD.n6134 1084.97
R11928 VDD.n6125 VDD.n5990 1084.97
R11929 VDD.n6000 VDD.n5990 1084.97
R11930 VDD.n6124 VDD.n6000 1084.97
R11931 VDD.n6125 VDD.n6124 1084.97
R11932 VDD.n6119 VDD.n6003 1084.97
R11933 VDD.n6119 VDD.n6004 1084.97
R11934 VDD.n6115 VDD.n6004 1084.97
R11935 VDD.n6115 VDD.n6003 1084.97
R11936 VDD.n6108 VDD.n6006 1084.97
R11937 VDD.n6015 VDD.n6006 1084.97
R11938 VDD.n6107 VDD.n6015 1084.97
R11939 VDD.n6108 VDD.n6107 1084.97
R11940 VDD.n6098 VDD.n6018 1084.97
R11941 VDD.n6028 VDD.n6018 1084.97
R11942 VDD.n6097 VDD.n6028 1084.97
R11943 VDD.n6098 VDD.n6097 1084.97
R11944 VDD.n6088 VDD.n6031 1084.97
R11945 VDD.n6039 VDD.n6031 1084.97
R11946 VDD.n6087 VDD.n6039 1084.97
R11947 VDD.n6088 VDD.n6087 1084.97
R11948 VDD.n6078 VDD.n6042 1084.97
R11949 VDD.n6049 VDD.n6042 1084.97
R11950 VDD.n6077 VDD.n6049 1084.97
R11951 VDD.n6078 VDD.n6077 1084.97
R11952 VDD.n6065 VDD.n6064 1084.97
R11953 VDD.n6065 VDD.n6052 1084.97
R11954 VDD.n6058 VDD.n6052 1084.97
R11955 VDD.n6064 VDD.n6058 1084.97
R11956 VDD.n6062 VDD.n6053 1084.97
R11957 VDD.n6072 VDD.n6053 1084.97
R11958 VDD.n6062 VDD.n6054 1084.97
R11959 VDD.n6072 VDD.n6054 1084.97
R11960 VDD.n7110 VDD.n144 1084.97
R11961 VDD.n7114 VDD.n145 1084.97
R11962 VDD.n7114 VDD.n144 1084.97
R11963 VDD.n7117 VDD.n141 1084.97
R11964 VDD.n7117 VDD.n142 1084.97
R11965 VDD.n7121 VDD.n142 1084.97
R11966 VDD.n7121 VDD.n141 1084.97
R11967 VDD.n7124 VDD.n136 1084.97
R11968 VDD.n139 VDD.n138 1084.97
R11969 VDD.n7124 VDD.n138 1084.97
R11970 VDD.n7131 VDD.n125 1084.97
R11971 VDD.n7135 VDD.n126 1084.97
R11972 VDD.n7135 VDD.n125 1084.97
R11973 VDD.n7138 VDD.n122 1084.97
R11974 VDD.n7138 VDD.n123 1084.97
R11975 VDD.n7142 VDD.n123 1084.97
R11976 VDD.n7142 VDD.n122 1084.97
R11977 VDD.n7145 VDD.n117 1084.97
R11978 VDD.n120 VDD.n119 1084.97
R11979 VDD.n7145 VDD.n119 1084.97
R11980 VDD.n7152 VDD.n106 1084.97
R11981 VDD.n7156 VDD.n107 1084.97
R11982 VDD.n7156 VDD.n106 1084.97
R11983 VDD.n7159 VDD.n103 1084.97
R11984 VDD.n7159 VDD.n104 1084.97
R11985 VDD.n7163 VDD.n104 1084.97
R11986 VDD.n7163 VDD.n103 1084.97
R11987 VDD.n7166 VDD.n98 1084.97
R11988 VDD.n101 VDD.n100 1084.97
R11989 VDD.n7166 VDD.n100 1084.97
R11990 VDD.n7173 VDD.n87 1084.97
R11991 VDD.n7177 VDD.n88 1084.97
R11992 VDD.n7177 VDD.n87 1084.97
R11993 VDD.n7180 VDD.n84 1084.97
R11994 VDD.n7180 VDD.n85 1084.97
R11995 VDD.n7184 VDD.n85 1084.97
R11996 VDD.n7184 VDD.n84 1084.97
R11997 VDD.n7187 VDD.n79 1084.97
R11998 VDD.n82 VDD.n81 1084.97
R11999 VDD.n7187 VDD.n81 1084.97
R12000 VDD.n7194 VDD.n68 1084.97
R12001 VDD.n7198 VDD.n69 1084.97
R12002 VDD.n7198 VDD.n68 1084.97
R12003 VDD.n7201 VDD.n65 1084.97
R12004 VDD.n7201 VDD.n66 1084.97
R12005 VDD.n7205 VDD.n66 1084.97
R12006 VDD.n7205 VDD.n65 1084.97
R12007 VDD.n7208 VDD.n60 1084.97
R12008 VDD.n63 VDD.n62 1084.97
R12009 VDD.n7208 VDD.n62 1084.97
R12010 VDD.n7215 VDD.n49 1084.97
R12011 VDD.n7219 VDD.n50 1084.97
R12012 VDD.n7219 VDD.n49 1084.97
R12013 VDD.n7222 VDD.n46 1084.97
R12014 VDD.n7222 VDD.n47 1084.97
R12015 VDD.n7226 VDD.n47 1084.97
R12016 VDD.n7226 VDD.n46 1084.97
R12017 VDD.n7229 VDD.n41 1084.97
R12018 VDD.n44 VDD.n43 1084.97
R12019 VDD.n7229 VDD.n43 1084.97
R12020 VDD.n7236 VDD.n30 1084.97
R12021 VDD.n7240 VDD.n31 1084.97
R12022 VDD.n7240 VDD.n30 1084.97
R12023 VDD.n7243 VDD.n27 1084.97
R12024 VDD.n7243 VDD.n28 1084.97
R12025 VDD.n7247 VDD.n28 1084.97
R12026 VDD.n7247 VDD.n27 1084.97
R12027 VDD.n7250 VDD.n22 1084.97
R12028 VDD.n25 VDD.n24 1084.97
R12029 VDD.n7250 VDD.n24 1084.97
R12030 VDD.n7257 VDD.n11 1084.97
R12031 VDD.n7261 VDD.n12 1084.97
R12032 VDD.n7261 VDD.n11 1084.97
R12033 VDD.n7264 VDD.n8 1084.97
R12034 VDD.n7264 VDD.n9 1084.97
R12035 VDD.n7268 VDD.n9 1084.97
R12036 VDD.n7268 VDD.n8 1084.97
R12037 VDD.n7271 VDD.n3 1084.97
R12038 VDD.n6 VDD.n5 1084.97
R12039 VDD.n7271 VDD.n5 1084.97
R12040 VDD.n7300 VDD.n7281 516.932
R12041 VDD.n7307 VDD.n7281 516.932
R12042 VDD.n7302 VDD.n7297 516.932
R12043 VDD.n7306 VDD.n7297 516.932
R12044 VDD.n5020 VDD.n5019 295.125
R12045 VDD.n4979 VDD.n4978 295.125
R12046 VDD.n4938 VDD.n4937 295.125
R12047 VDD.n4897 VDD.n4896 295.125
R12048 VDD.n4856 VDD.n4855 295.125
R12049 VDD.n4815 VDD.n4814 295.125
R12050 VDD.n4774 VDD.n4773 295.125
R12051 VDD.n4733 VDD.n4732 295.125
R12052 VDD.n5019 VDD.t332 253.119
R12053 VDD.n5020 VDD.t819 253.119
R12054 VDD.n5026 VDD.t819 253.119
R12055 VDD.t796 VDD.n5027 253.119
R12056 VDD.n5001 VDD.t468 253.119
R12057 VDD.t269 VDD.n5002 253.119
R12058 VDD.n4978 VDD.t585 253.119
R12059 VDD.n4979 VDD.t252 253.119
R12060 VDD.n4985 VDD.t252 253.119
R12061 VDD.t583 VDD.n4986 253.119
R12062 VDD.n4960 VDD.t888 253.119
R12063 VDD.t703 VDD.n4961 253.119
R12064 VDD.n4937 VDD.t549 253.119
R12065 VDD.n4938 VDD.t292 253.119
R12066 VDD.n4944 VDD.t292 253.119
R12067 VDD.t598 VDD.n4945 253.119
R12068 VDD.n4919 VDD.t31 253.119
R12069 VDD.t732 VDD.n4920 253.119
R12070 VDD.n4896 VDD.t526 253.119
R12071 VDD.n4897 VDD.t828 253.119
R12072 VDD.n4903 VDD.t828 253.119
R12073 VDD.t891 VDD.n4904 253.119
R12074 VDD.n4878 VDD.t59 253.119
R12075 VDD.t454 VDD.n4879 253.119
R12076 VDD.n4855 VDD.t596 253.119
R12077 VDD.n4856 VDD.t744 253.119
R12078 VDD.n4862 VDD.t744 253.119
R12079 VDD.t594 VDD.n4863 253.119
R12080 VDD.n4837 VDD.t553 253.119
R12081 VDD.t368 VDD.n4838 253.119
R12082 VDD.n4814 VDD.t645 253.119
R12083 VDD.n4815 VDD.t822 253.119
R12084 VDD.n4821 VDD.t822 253.119
R12085 VDD.t296 VDD.n4822 253.119
R12086 VDD.n4796 VDD.t87 253.119
R12087 VDD.t794 VDD.n4797 253.119
R12088 VDD.n4773 VDD.t725 253.119
R12089 VDD.n4774 VDD.t224 253.119
R12090 VDD.n4780 VDD.t224 253.119
R12091 VDD.t422 VDD.n4781 253.119
R12092 VDD.n4755 VDD.t747 253.119
R12093 VDD.t878 VDD.n4756 253.119
R12094 VDD.n4732 VDD.t869 253.119
R12095 VDD.n4733 VDD.t812 253.119
R12096 VDD.n4739 VDD.t812 253.119
R12097 VDD.t842 VDD.n4740 253.119
R12098 VDD.n4714 VDD.t340 253.119
R12099 VDD.t571 VDD.n4715 253.119
R12100 VDD.n7123 VDD.t773 253.119
R12101 VDD.n7122 VDD.t776 253.119
R12102 VDD.n7116 VDD.t776 253.119
R12103 VDD.n7115 VDD.t915 253.119
R12104 VDD.n7144 VDD.t903 253.119
R12105 VDD.n7143 VDD.t905 253.119
R12106 VDD.n7137 VDD.t905 253.119
R12107 VDD.n7136 VDD.t880 253.119
R12108 VDD.n7165 VDD.t855 253.119
R12109 VDD.n7164 VDD.t866 253.119
R12110 VDD.n7158 VDD.t866 253.119
R12111 VDD.n7157 VDD.t544 253.119
R12112 VDD.n7186 VDD.t298 253.119
R12113 VDD.n7185 VDD.t790 253.119
R12114 VDD.n7179 VDD.t790 253.119
R12115 VDD.n7178 VDD.t96 253.119
R12116 VDD.n7207 VDD.t714 253.119
R12117 VDD.n7206 VDD.t713 253.119
R12118 VDD.n7200 VDD.t713 253.119
R12119 VDD.n7199 VDD.t402 253.119
R12120 VDD.n7228 VDD.t383 253.119
R12121 VDD.n7227 VDD.t427 253.119
R12122 VDD.n7221 VDD.t427 253.119
R12123 VDD.n7220 VDD.t630 253.119
R12124 VDD.n7249 VDD.t895 253.119
R12125 VDD.n7248 VDD.t894 253.119
R12126 VDD.n7242 VDD.t894 253.119
R12127 VDD.n7241 VDD.t301 253.119
R12128 VDD.n7270 VDD.t509 253.119
R12129 VDD.n7269 VDD.t911 253.119
R12130 VDD.n7263 VDD.t911 253.119
R12131 VDD.n7262 VDD.t314 253.119
R12132 VDD.n5030 VDD.n4560 214.357
R12133 VDD.n5014 VDD.n5013 214.357
R12134 VDD.n5005 VDD.n4571 214.357
R12135 VDD.n4996 VDD.n4995 214.357
R12136 VDD.n4989 VDD.n4579 214.357
R12137 VDD.n4973 VDD.n4972 214.357
R12138 VDD.n4964 VDD.n4590 214.357
R12139 VDD.n4955 VDD.n4954 214.357
R12140 VDD.n4948 VDD.n4598 214.357
R12141 VDD.n4932 VDD.n4931 214.357
R12142 VDD.n4923 VDD.n4609 214.357
R12143 VDD.n4914 VDD.n4913 214.357
R12144 VDD.n4907 VDD.n4617 214.357
R12145 VDD.n4891 VDD.n4890 214.357
R12146 VDD.n4882 VDD.n4628 214.357
R12147 VDD.n4873 VDD.n4872 214.357
R12148 VDD.n4866 VDD.n4636 214.357
R12149 VDD.n4850 VDD.n4849 214.357
R12150 VDD.n4841 VDD.n4647 214.357
R12151 VDD.n4832 VDD.n4831 214.357
R12152 VDD.n4825 VDD.n4655 214.357
R12153 VDD.n4809 VDD.n4808 214.357
R12154 VDD.n4800 VDD.n4666 214.357
R12155 VDD.n4791 VDD.n4790 214.357
R12156 VDD.n4784 VDD.n4674 214.357
R12157 VDD.n4768 VDD.n4767 214.357
R12158 VDD.n4759 VDD.n4685 214.357
R12159 VDD.n4750 VDD.n4749 214.357
R12160 VDD.n4743 VDD.n4693 214.357
R12161 VDD.n4727 VDD.n4726 214.357
R12162 VDD.n4718 VDD.n4704 214.357
R12163 VDD.n4709 VDD.n4708 214.357
R12164 VDD.n7110 VDD.n7109 214.357
R12165 VDD.n140 VDD.n139 214.357
R12166 VDD.n7131 VDD.n7130 214.357
R12167 VDD.n121 VDD.n120 214.357
R12168 VDD.n7152 VDD.n7151 214.357
R12169 VDD.n102 VDD.n101 214.357
R12170 VDD.n7173 VDD.n7172 214.357
R12171 VDD.n83 VDD.n82 214.357
R12172 VDD.n7194 VDD.n7193 214.357
R12173 VDD.n64 VDD.n63 214.357
R12174 VDD.n7215 VDD.n7214 214.357
R12175 VDD.n45 VDD.n44 214.357
R12176 VDD.n7236 VDD.n7235 214.357
R12177 VDD.n26 VDD.n25 214.357
R12178 VDD.n7257 VDD.n7256 214.357
R12179 VDD.n7 VDD.n6 214.357
R12180 VDD.n376 VDD.n189 212.329
R12181 VDD.n376 VDD.n190 212.329
R12182 VDD.n198 VDD.n197 212.329
R12183 VDD.n197 VDD.n196 212.329
R12184 VDD.n243 VDD.n242 212.329
R12185 VDD.n243 VDD.n241 212.329
R12186 VDD.n221 VDD.n220 212.329
R12187 VDD.n221 VDD.n219 212.329
R12188 VDD.n374 VDD.n373 212.329
R12189 VDD.n374 VDD.n372 212.329
R12190 VDD.n284 VDD.n283 212.329
R12191 VDD.n283 VDD.n281 212.329
R12192 VDD.n289 VDD.n287 212.329
R12193 VDD.n287 VDD.n286 212.329
R12194 VDD.n274 VDD.n272 212.329
R12195 VDD.n275 VDD.n274 212.329
R12196 VDD.n370 VDD.n369 212.329
R12197 VDD.n370 VDD.n271 212.329
R12198 VDD.n357 VDD.n356 212.329
R12199 VDD.n356 VDD.n354 212.329
R12200 VDD.n362 VDD.n360 212.329
R12201 VDD.n360 VDD.n359 212.329
R12202 VDD.n341 VDD.n340 212.329
R12203 VDD.n340 VDD.n338 212.329
R12204 VDD.n346 VDD.n344 212.329
R12205 VDD.n344 VDD.n343 212.329
R12206 VDD.n330 VDD.n327 212.329
R12207 VDD.n331 VDD.n330 212.329
R12208 VDD.n318 VDD.n317 212.329
R12209 VDD.n317 VDD.n315 212.329
R12210 VDD.n323 VDD.n321 212.329
R12211 VDD.n321 VDD.n320 212.329
R12212 VDD.n302 VDD.n301 212.329
R12213 VDD.n301 VDD.n299 212.329
R12214 VDD.n307 VDD.n305 212.329
R12215 VDD.n305 VDD.n304 212.329
R12216 VDD.n253 VDD.n251 212.329
R12217 VDD.n254 VDD.n253 212.329
R12218 VDD.n260 VDD.n259 212.329
R12219 VDD.n260 VDD.n250 212.329
R12220 VDD.n235 VDD.n234 212.329
R12221 VDD.n234 VDD.n232 212.329
R12222 VDD.n381 VDD.n236 212.329
R12223 VDD.n237 VDD.n236 212.329
R12224 VDD.n265 VDD.n228 212.329
R12225 VDD.n265 VDD.n264 212.329
R12226 VDD.n392 VDD.n391 212.329
R12227 VDD.n391 VDD.n390 212.329
R12228 VDD.n624 VDD.n437 212.329
R12229 VDD.n624 VDD.n438 212.329
R12230 VDD.n446 VDD.n445 212.329
R12231 VDD.n445 VDD.n444 212.329
R12232 VDD.n491 VDD.n490 212.329
R12233 VDD.n491 VDD.n489 212.329
R12234 VDD.n469 VDD.n468 212.329
R12235 VDD.n469 VDD.n467 212.329
R12236 VDD.n622 VDD.n621 212.329
R12237 VDD.n622 VDD.n620 212.329
R12238 VDD.n532 VDD.n531 212.329
R12239 VDD.n531 VDD.n529 212.329
R12240 VDD.n537 VDD.n535 212.329
R12241 VDD.n535 VDD.n534 212.329
R12242 VDD.n522 VDD.n520 212.329
R12243 VDD.n523 VDD.n522 212.329
R12244 VDD.n618 VDD.n617 212.329
R12245 VDD.n618 VDD.n519 212.329
R12246 VDD.n605 VDD.n604 212.329
R12247 VDD.n604 VDD.n602 212.329
R12248 VDD.n610 VDD.n608 212.329
R12249 VDD.n608 VDD.n607 212.329
R12250 VDD.n589 VDD.n588 212.329
R12251 VDD.n588 VDD.n586 212.329
R12252 VDD.n594 VDD.n592 212.329
R12253 VDD.n592 VDD.n591 212.329
R12254 VDD.n578 VDD.n575 212.329
R12255 VDD.n579 VDD.n578 212.329
R12256 VDD.n566 VDD.n565 212.329
R12257 VDD.n565 VDD.n563 212.329
R12258 VDD.n571 VDD.n569 212.329
R12259 VDD.n569 VDD.n568 212.329
R12260 VDD.n550 VDD.n549 212.329
R12261 VDD.n549 VDD.n547 212.329
R12262 VDD.n555 VDD.n553 212.329
R12263 VDD.n553 VDD.n552 212.329
R12264 VDD.n501 VDD.n499 212.329
R12265 VDD.n502 VDD.n501 212.329
R12266 VDD.n508 VDD.n507 212.329
R12267 VDD.n508 VDD.n498 212.329
R12268 VDD.n483 VDD.n482 212.329
R12269 VDD.n482 VDD.n480 212.329
R12270 VDD.n629 VDD.n484 212.329
R12271 VDD.n485 VDD.n484 212.329
R12272 VDD.n513 VDD.n476 212.329
R12273 VDD.n513 VDD.n512 212.329
R12274 VDD.n640 VDD.n639 212.329
R12275 VDD.n639 VDD.n638 212.329
R12276 VDD.n883 VDD.n696 212.329
R12277 VDD.n883 VDD.n697 212.329
R12278 VDD.n705 VDD.n704 212.329
R12279 VDD.n704 VDD.n703 212.329
R12280 VDD.n750 VDD.n749 212.329
R12281 VDD.n750 VDD.n748 212.329
R12282 VDD.n728 VDD.n727 212.329
R12283 VDD.n728 VDD.n726 212.329
R12284 VDD.n881 VDD.n880 212.329
R12285 VDD.n881 VDD.n879 212.329
R12286 VDD.n791 VDD.n790 212.329
R12287 VDD.n790 VDD.n788 212.329
R12288 VDD.n796 VDD.n794 212.329
R12289 VDD.n794 VDD.n793 212.329
R12290 VDD.n781 VDD.n779 212.329
R12291 VDD.n782 VDD.n781 212.329
R12292 VDD.n877 VDD.n876 212.329
R12293 VDD.n877 VDD.n778 212.329
R12294 VDD.n864 VDD.n863 212.329
R12295 VDD.n863 VDD.n861 212.329
R12296 VDD.n869 VDD.n867 212.329
R12297 VDD.n867 VDD.n866 212.329
R12298 VDD.n848 VDD.n847 212.329
R12299 VDD.n847 VDD.n845 212.329
R12300 VDD.n853 VDD.n851 212.329
R12301 VDD.n851 VDD.n850 212.329
R12302 VDD.n837 VDD.n834 212.329
R12303 VDD.n838 VDD.n837 212.329
R12304 VDD.n825 VDD.n824 212.329
R12305 VDD.n824 VDD.n822 212.329
R12306 VDD.n830 VDD.n828 212.329
R12307 VDD.n828 VDD.n827 212.329
R12308 VDD.n809 VDD.n808 212.329
R12309 VDD.n808 VDD.n806 212.329
R12310 VDD.n814 VDD.n812 212.329
R12311 VDD.n812 VDD.n811 212.329
R12312 VDD.n760 VDD.n758 212.329
R12313 VDD.n761 VDD.n760 212.329
R12314 VDD.n767 VDD.n766 212.329
R12315 VDD.n767 VDD.n757 212.329
R12316 VDD.n742 VDD.n741 212.329
R12317 VDD.n741 VDD.n739 212.329
R12318 VDD.n888 VDD.n743 212.329
R12319 VDD.n744 VDD.n743 212.329
R12320 VDD.n772 VDD.n735 212.329
R12321 VDD.n772 VDD.n771 212.329
R12322 VDD.n899 VDD.n898 212.329
R12323 VDD.n898 VDD.n897 212.329
R12324 VDD.n1142 VDD.n955 212.329
R12325 VDD.n1142 VDD.n956 212.329
R12326 VDD.n964 VDD.n963 212.329
R12327 VDD.n963 VDD.n962 212.329
R12328 VDD.n1009 VDD.n1008 212.329
R12329 VDD.n1009 VDD.n1007 212.329
R12330 VDD.n987 VDD.n986 212.329
R12331 VDD.n987 VDD.n985 212.329
R12332 VDD.n1140 VDD.n1139 212.329
R12333 VDD.n1140 VDD.n1138 212.329
R12334 VDD.n1050 VDD.n1049 212.329
R12335 VDD.n1049 VDD.n1047 212.329
R12336 VDD.n1055 VDD.n1053 212.329
R12337 VDD.n1053 VDD.n1052 212.329
R12338 VDD.n1040 VDD.n1038 212.329
R12339 VDD.n1041 VDD.n1040 212.329
R12340 VDD.n1136 VDD.n1135 212.329
R12341 VDD.n1136 VDD.n1037 212.329
R12342 VDD.n1123 VDD.n1122 212.329
R12343 VDD.n1122 VDD.n1120 212.329
R12344 VDD.n1128 VDD.n1126 212.329
R12345 VDD.n1126 VDD.n1125 212.329
R12346 VDD.n1107 VDD.n1106 212.329
R12347 VDD.n1106 VDD.n1104 212.329
R12348 VDD.n1112 VDD.n1110 212.329
R12349 VDD.n1110 VDD.n1109 212.329
R12350 VDD.n1096 VDD.n1093 212.329
R12351 VDD.n1097 VDD.n1096 212.329
R12352 VDD.n1084 VDD.n1083 212.329
R12353 VDD.n1083 VDD.n1081 212.329
R12354 VDD.n1089 VDD.n1087 212.329
R12355 VDD.n1087 VDD.n1086 212.329
R12356 VDD.n1068 VDD.n1067 212.329
R12357 VDD.n1067 VDD.n1065 212.329
R12358 VDD.n1073 VDD.n1071 212.329
R12359 VDD.n1071 VDD.n1070 212.329
R12360 VDD.n1019 VDD.n1017 212.329
R12361 VDD.n1020 VDD.n1019 212.329
R12362 VDD.n1026 VDD.n1025 212.329
R12363 VDD.n1026 VDD.n1016 212.329
R12364 VDD.n1001 VDD.n1000 212.329
R12365 VDD.n1000 VDD.n998 212.329
R12366 VDD.n1147 VDD.n1002 212.329
R12367 VDD.n1003 VDD.n1002 212.329
R12368 VDD.n1031 VDD.n994 212.329
R12369 VDD.n1031 VDD.n1030 212.329
R12370 VDD.n1158 VDD.n1157 212.329
R12371 VDD.n1157 VDD.n1156 212.329
R12372 VDD.n1401 VDD.n1214 212.329
R12373 VDD.n1401 VDD.n1215 212.329
R12374 VDD.n1223 VDD.n1222 212.329
R12375 VDD.n1222 VDD.n1221 212.329
R12376 VDD.n1268 VDD.n1267 212.329
R12377 VDD.n1268 VDD.n1266 212.329
R12378 VDD.n1246 VDD.n1245 212.329
R12379 VDD.n1246 VDD.n1244 212.329
R12380 VDD.n1399 VDD.n1398 212.329
R12381 VDD.n1399 VDD.n1397 212.329
R12382 VDD.n1309 VDD.n1308 212.329
R12383 VDD.n1308 VDD.n1306 212.329
R12384 VDD.n1314 VDD.n1312 212.329
R12385 VDD.n1312 VDD.n1311 212.329
R12386 VDD.n1299 VDD.n1297 212.329
R12387 VDD.n1300 VDD.n1299 212.329
R12388 VDD.n1395 VDD.n1394 212.329
R12389 VDD.n1395 VDD.n1296 212.329
R12390 VDD.n1382 VDD.n1381 212.329
R12391 VDD.n1381 VDD.n1379 212.329
R12392 VDD.n1387 VDD.n1385 212.329
R12393 VDD.n1385 VDD.n1384 212.329
R12394 VDD.n1366 VDD.n1365 212.329
R12395 VDD.n1365 VDD.n1363 212.329
R12396 VDD.n1371 VDD.n1369 212.329
R12397 VDD.n1369 VDD.n1368 212.329
R12398 VDD.n1355 VDD.n1352 212.329
R12399 VDD.n1356 VDD.n1355 212.329
R12400 VDD.n1343 VDD.n1342 212.329
R12401 VDD.n1342 VDD.n1340 212.329
R12402 VDD.n1348 VDD.n1346 212.329
R12403 VDD.n1346 VDD.n1345 212.329
R12404 VDD.n1327 VDD.n1326 212.329
R12405 VDD.n1326 VDD.n1324 212.329
R12406 VDD.n1332 VDD.n1330 212.329
R12407 VDD.n1330 VDD.n1329 212.329
R12408 VDD.n1278 VDD.n1276 212.329
R12409 VDD.n1279 VDD.n1278 212.329
R12410 VDD.n1285 VDD.n1284 212.329
R12411 VDD.n1285 VDD.n1275 212.329
R12412 VDD.n1260 VDD.n1259 212.329
R12413 VDD.n1259 VDD.n1257 212.329
R12414 VDD.n1406 VDD.n1261 212.329
R12415 VDD.n1262 VDD.n1261 212.329
R12416 VDD.n1290 VDD.n1253 212.329
R12417 VDD.n1290 VDD.n1289 212.329
R12418 VDD.n1417 VDD.n1416 212.329
R12419 VDD.n1416 VDD.n1415 212.329
R12420 VDD.n1660 VDD.n1473 212.329
R12421 VDD.n1660 VDD.n1474 212.329
R12422 VDD.n1482 VDD.n1481 212.329
R12423 VDD.n1481 VDD.n1480 212.329
R12424 VDD.n1527 VDD.n1526 212.329
R12425 VDD.n1527 VDD.n1525 212.329
R12426 VDD.n1505 VDD.n1504 212.329
R12427 VDD.n1505 VDD.n1503 212.329
R12428 VDD.n1658 VDD.n1657 212.329
R12429 VDD.n1658 VDD.n1656 212.329
R12430 VDD.n1568 VDD.n1567 212.329
R12431 VDD.n1567 VDD.n1565 212.329
R12432 VDD.n1573 VDD.n1571 212.329
R12433 VDD.n1571 VDD.n1570 212.329
R12434 VDD.n1558 VDD.n1556 212.329
R12435 VDD.n1559 VDD.n1558 212.329
R12436 VDD.n1654 VDD.n1653 212.329
R12437 VDD.n1654 VDD.n1555 212.329
R12438 VDD.n1641 VDD.n1640 212.329
R12439 VDD.n1640 VDD.n1638 212.329
R12440 VDD.n1646 VDD.n1644 212.329
R12441 VDD.n1644 VDD.n1643 212.329
R12442 VDD.n1625 VDD.n1624 212.329
R12443 VDD.n1624 VDD.n1622 212.329
R12444 VDD.n1630 VDD.n1628 212.329
R12445 VDD.n1628 VDD.n1627 212.329
R12446 VDD.n1614 VDD.n1611 212.329
R12447 VDD.n1615 VDD.n1614 212.329
R12448 VDD.n1602 VDD.n1601 212.329
R12449 VDD.n1601 VDD.n1599 212.329
R12450 VDD.n1607 VDD.n1605 212.329
R12451 VDD.n1605 VDD.n1604 212.329
R12452 VDD.n1586 VDD.n1585 212.329
R12453 VDD.n1585 VDD.n1583 212.329
R12454 VDD.n1591 VDD.n1589 212.329
R12455 VDD.n1589 VDD.n1588 212.329
R12456 VDD.n1537 VDD.n1535 212.329
R12457 VDD.n1538 VDD.n1537 212.329
R12458 VDD.n1544 VDD.n1543 212.329
R12459 VDD.n1544 VDD.n1534 212.329
R12460 VDD.n1519 VDD.n1518 212.329
R12461 VDD.n1518 VDD.n1516 212.329
R12462 VDD.n1665 VDD.n1520 212.329
R12463 VDD.n1521 VDD.n1520 212.329
R12464 VDD.n1549 VDD.n1512 212.329
R12465 VDD.n1549 VDD.n1548 212.329
R12466 VDD.n1676 VDD.n1675 212.329
R12467 VDD.n1675 VDD.n1674 212.329
R12468 VDD.n1919 VDD.n1732 212.329
R12469 VDD.n1919 VDD.n1733 212.329
R12470 VDD.n1741 VDD.n1740 212.329
R12471 VDD.n1740 VDD.n1739 212.329
R12472 VDD.n1786 VDD.n1785 212.329
R12473 VDD.n1786 VDD.n1784 212.329
R12474 VDD.n1764 VDD.n1763 212.329
R12475 VDD.n1764 VDD.n1762 212.329
R12476 VDD.n1917 VDD.n1916 212.329
R12477 VDD.n1917 VDD.n1915 212.329
R12478 VDD.n1827 VDD.n1826 212.329
R12479 VDD.n1826 VDD.n1824 212.329
R12480 VDD.n1832 VDD.n1830 212.329
R12481 VDD.n1830 VDD.n1829 212.329
R12482 VDD.n1817 VDD.n1815 212.329
R12483 VDD.n1818 VDD.n1817 212.329
R12484 VDD.n1913 VDD.n1912 212.329
R12485 VDD.n1913 VDD.n1814 212.329
R12486 VDD.n1900 VDD.n1899 212.329
R12487 VDD.n1899 VDD.n1897 212.329
R12488 VDD.n1905 VDD.n1903 212.329
R12489 VDD.n1903 VDD.n1902 212.329
R12490 VDD.n1884 VDD.n1883 212.329
R12491 VDD.n1883 VDD.n1881 212.329
R12492 VDD.n1889 VDD.n1887 212.329
R12493 VDD.n1887 VDD.n1886 212.329
R12494 VDD.n1873 VDD.n1870 212.329
R12495 VDD.n1874 VDD.n1873 212.329
R12496 VDD.n1861 VDD.n1860 212.329
R12497 VDD.n1860 VDD.n1858 212.329
R12498 VDD.n1866 VDD.n1864 212.329
R12499 VDD.n1864 VDD.n1863 212.329
R12500 VDD.n1845 VDD.n1844 212.329
R12501 VDD.n1844 VDD.n1842 212.329
R12502 VDD.n1850 VDD.n1848 212.329
R12503 VDD.n1848 VDD.n1847 212.329
R12504 VDD.n1796 VDD.n1794 212.329
R12505 VDD.n1797 VDD.n1796 212.329
R12506 VDD.n1803 VDD.n1802 212.329
R12507 VDD.n1803 VDD.n1793 212.329
R12508 VDD.n1778 VDD.n1777 212.329
R12509 VDD.n1777 VDD.n1775 212.329
R12510 VDD.n1924 VDD.n1779 212.329
R12511 VDD.n1780 VDD.n1779 212.329
R12512 VDD.n1808 VDD.n1771 212.329
R12513 VDD.n1808 VDD.n1807 212.329
R12514 VDD.n1935 VDD.n1934 212.329
R12515 VDD.n1934 VDD.n1933 212.329
R12516 VDD.n2178 VDD.n1991 212.329
R12517 VDD.n2178 VDD.n1992 212.329
R12518 VDD.n2000 VDD.n1999 212.329
R12519 VDD.n1999 VDD.n1998 212.329
R12520 VDD.n2045 VDD.n2044 212.329
R12521 VDD.n2045 VDD.n2043 212.329
R12522 VDD.n2023 VDD.n2022 212.329
R12523 VDD.n2023 VDD.n2021 212.329
R12524 VDD.n2176 VDD.n2175 212.329
R12525 VDD.n2176 VDD.n2174 212.329
R12526 VDD.n2086 VDD.n2085 212.329
R12527 VDD.n2085 VDD.n2083 212.329
R12528 VDD.n2091 VDD.n2089 212.329
R12529 VDD.n2089 VDD.n2088 212.329
R12530 VDD.n2076 VDD.n2074 212.329
R12531 VDD.n2077 VDD.n2076 212.329
R12532 VDD.n2172 VDD.n2171 212.329
R12533 VDD.n2172 VDD.n2073 212.329
R12534 VDD.n2159 VDD.n2158 212.329
R12535 VDD.n2158 VDD.n2156 212.329
R12536 VDD.n2164 VDD.n2162 212.329
R12537 VDD.n2162 VDD.n2161 212.329
R12538 VDD.n2143 VDD.n2142 212.329
R12539 VDD.n2142 VDD.n2140 212.329
R12540 VDD.n2148 VDD.n2146 212.329
R12541 VDD.n2146 VDD.n2145 212.329
R12542 VDD.n2132 VDD.n2129 212.329
R12543 VDD.n2133 VDD.n2132 212.329
R12544 VDD.n2120 VDD.n2119 212.329
R12545 VDD.n2119 VDD.n2117 212.329
R12546 VDD.n2125 VDD.n2123 212.329
R12547 VDD.n2123 VDD.n2122 212.329
R12548 VDD.n2104 VDD.n2103 212.329
R12549 VDD.n2103 VDD.n2101 212.329
R12550 VDD.n2109 VDD.n2107 212.329
R12551 VDD.n2107 VDD.n2106 212.329
R12552 VDD.n2055 VDD.n2053 212.329
R12553 VDD.n2056 VDD.n2055 212.329
R12554 VDD.n2062 VDD.n2061 212.329
R12555 VDD.n2062 VDD.n2052 212.329
R12556 VDD.n2037 VDD.n2036 212.329
R12557 VDD.n2036 VDD.n2034 212.329
R12558 VDD.n2183 VDD.n2038 212.329
R12559 VDD.n2039 VDD.n2038 212.329
R12560 VDD.n2067 VDD.n2030 212.329
R12561 VDD.n2067 VDD.n2066 212.329
R12562 VDD.n2194 VDD.n2193 212.329
R12563 VDD.n2193 VDD.n2192 212.329
R12564 VDD.n2437 VDD.n2250 212.329
R12565 VDD.n2437 VDD.n2251 212.329
R12566 VDD.n2259 VDD.n2258 212.329
R12567 VDD.n2258 VDD.n2257 212.329
R12568 VDD.n2304 VDD.n2303 212.329
R12569 VDD.n2304 VDD.n2302 212.329
R12570 VDD.n2282 VDD.n2281 212.329
R12571 VDD.n2282 VDD.n2280 212.329
R12572 VDD.n2435 VDD.n2434 212.329
R12573 VDD.n2435 VDD.n2433 212.329
R12574 VDD.n2345 VDD.n2344 212.329
R12575 VDD.n2344 VDD.n2342 212.329
R12576 VDD.n2350 VDD.n2348 212.329
R12577 VDD.n2348 VDD.n2347 212.329
R12578 VDD.n2335 VDD.n2333 212.329
R12579 VDD.n2336 VDD.n2335 212.329
R12580 VDD.n2431 VDD.n2430 212.329
R12581 VDD.n2431 VDD.n2332 212.329
R12582 VDD.n2418 VDD.n2417 212.329
R12583 VDD.n2417 VDD.n2415 212.329
R12584 VDD.n2423 VDD.n2421 212.329
R12585 VDD.n2421 VDD.n2420 212.329
R12586 VDD.n2402 VDD.n2401 212.329
R12587 VDD.n2401 VDD.n2399 212.329
R12588 VDD.n2407 VDD.n2405 212.329
R12589 VDD.n2405 VDD.n2404 212.329
R12590 VDD.n2391 VDD.n2388 212.329
R12591 VDD.n2392 VDD.n2391 212.329
R12592 VDD.n2379 VDD.n2378 212.329
R12593 VDD.n2378 VDD.n2376 212.329
R12594 VDD.n2384 VDD.n2382 212.329
R12595 VDD.n2382 VDD.n2381 212.329
R12596 VDD.n2363 VDD.n2362 212.329
R12597 VDD.n2362 VDD.n2360 212.329
R12598 VDD.n2368 VDD.n2366 212.329
R12599 VDD.n2366 VDD.n2365 212.329
R12600 VDD.n2314 VDD.n2312 212.329
R12601 VDD.n2315 VDD.n2314 212.329
R12602 VDD.n2321 VDD.n2320 212.329
R12603 VDD.n2321 VDD.n2311 212.329
R12604 VDD.n2296 VDD.n2295 212.329
R12605 VDD.n2295 VDD.n2293 212.329
R12606 VDD.n2442 VDD.n2297 212.329
R12607 VDD.n2298 VDD.n2297 212.329
R12608 VDD.n2326 VDD.n2289 212.329
R12609 VDD.n2326 VDD.n2325 212.329
R12610 VDD.n2453 VDD.n2452 212.329
R12611 VDD.n2452 VDD.n2451 212.329
R12612 VDD.n2696 VDD.n2509 212.329
R12613 VDD.n2696 VDD.n2510 212.329
R12614 VDD.n2518 VDD.n2517 212.329
R12615 VDD.n2517 VDD.n2516 212.329
R12616 VDD.n2563 VDD.n2562 212.329
R12617 VDD.n2563 VDD.n2561 212.329
R12618 VDD.n2541 VDD.n2540 212.329
R12619 VDD.n2541 VDD.n2539 212.329
R12620 VDD.n2694 VDD.n2693 212.329
R12621 VDD.n2694 VDD.n2692 212.329
R12622 VDD.n2604 VDD.n2603 212.329
R12623 VDD.n2603 VDD.n2601 212.329
R12624 VDD.n2609 VDD.n2607 212.329
R12625 VDD.n2607 VDD.n2606 212.329
R12626 VDD.n2594 VDD.n2592 212.329
R12627 VDD.n2595 VDD.n2594 212.329
R12628 VDD.n2690 VDD.n2689 212.329
R12629 VDD.n2690 VDD.n2591 212.329
R12630 VDD.n2677 VDD.n2676 212.329
R12631 VDD.n2676 VDD.n2674 212.329
R12632 VDD.n2682 VDD.n2680 212.329
R12633 VDD.n2680 VDD.n2679 212.329
R12634 VDD.n2661 VDD.n2660 212.329
R12635 VDD.n2660 VDD.n2658 212.329
R12636 VDD.n2666 VDD.n2664 212.329
R12637 VDD.n2664 VDD.n2663 212.329
R12638 VDD.n2650 VDD.n2647 212.329
R12639 VDD.n2651 VDD.n2650 212.329
R12640 VDD.n2638 VDD.n2637 212.329
R12641 VDD.n2637 VDD.n2635 212.329
R12642 VDD.n2643 VDD.n2641 212.329
R12643 VDD.n2641 VDD.n2640 212.329
R12644 VDD.n2622 VDD.n2621 212.329
R12645 VDD.n2621 VDD.n2619 212.329
R12646 VDD.n2627 VDD.n2625 212.329
R12647 VDD.n2625 VDD.n2624 212.329
R12648 VDD.n2573 VDD.n2571 212.329
R12649 VDD.n2574 VDD.n2573 212.329
R12650 VDD.n2580 VDD.n2579 212.329
R12651 VDD.n2580 VDD.n2570 212.329
R12652 VDD.n2555 VDD.n2554 212.329
R12653 VDD.n2554 VDD.n2552 212.329
R12654 VDD.n2701 VDD.n2556 212.329
R12655 VDD.n2557 VDD.n2556 212.329
R12656 VDD.n2585 VDD.n2548 212.329
R12657 VDD.n2585 VDD.n2584 212.329
R12658 VDD.n2712 VDD.n2711 212.329
R12659 VDD.n2711 VDD.n2710 212.329
R12660 VDD.n2955 VDD.n2768 212.329
R12661 VDD.n2955 VDD.n2769 212.329
R12662 VDD.n2777 VDD.n2776 212.329
R12663 VDD.n2776 VDD.n2775 212.329
R12664 VDD.n2822 VDD.n2821 212.329
R12665 VDD.n2822 VDD.n2820 212.329
R12666 VDD.n2800 VDD.n2799 212.329
R12667 VDD.n2800 VDD.n2798 212.329
R12668 VDD.n2953 VDD.n2952 212.329
R12669 VDD.n2953 VDD.n2951 212.329
R12670 VDD.n2863 VDD.n2862 212.329
R12671 VDD.n2862 VDD.n2860 212.329
R12672 VDD.n2868 VDD.n2866 212.329
R12673 VDD.n2866 VDD.n2865 212.329
R12674 VDD.n2853 VDD.n2851 212.329
R12675 VDD.n2854 VDD.n2853 212.329
R12676 VDD.n2949 VDD.n2948 212.329
R12677 VDD.n2949 VDD.n2850 212.329
R12678 VDD.n2936 VDD.n2935 212.329
R12679 VDD.n2935 VDD.n2933 212.329
R12680 VDD.n2941 VDD.n2939 212.329
R12681 VDD.n2939 VDD.n2938 212.329
R12682 VDD.n2920 VDD.n2919 212.329
R12683 VDD.n2919 VDD.n2917 212.329
R12684 VDD.n2925 VDD.n2923 212.329
R12685 VDD.n2923 VDD.n2922 212.329
R12686 VDD.n2909 VDD.n2906 212.329
R12687 VDD.n2910 VDD.n2909 212.329
R12688 VDD.n2897 VDD.n2896 212.329
R12689 VDD.n2896 VDD.n2894 212.329
R12690 VDD.n2902 VDD.n2900 212.329
R12691 VDD.n2900 VDD.n2899 212.329
R12692 VDD.n2881 VDD.n2880 212.329
R12693 VDD.n2880 VDD.n2878 212.329
R12694 VDD.n2886 VDD.n2884 212.329
R12695 VDD.n2884 VDD.n2883 212.329
R12696 VDD.n2832 VDD.n2830 212.329
R12697 VDD.n2833 VDD.n2832 212.329
R12698 VDD.n2839 VDD.n2838 212.329
R12699 VDD.n2839 VDD.n2829 212.329
R12700 VDD.n2814 VDD.n2813 212.329
R12701 VDD.n2813 VDD.n2811 212.329
R12702 VDD.n2960 VDD.n2815 212.329
R12703 VDD.n2816 VDD.n2815 212.329
R12704 VDD.n2844 VDD.n2807 212.329
R12705 VDD.n2844 VDD.n2843 212.329
R12706 VDD.n2971 VDD.n2970 212.329
R12707 VDD.n2970 VDD.n2969 212.329
R12708 VDD.n3214 VDD.n3027 212.329
R12709 VDD.n3214 VDD.n3028 212.329
R12710 VDD.n3036 VDD.n3035 212.329
R12711 VDD.n3035 VDD.n3034 212.329
R12712 VDD.n3081 VDD.n3080 212.329
R12713 VDD.n3081 VDD.n3079 212.329
R12714 VDD.n3059 VDD.n3058 212.329
R12715 VDD.n3059 VDD.n3057 212.329
R12716 VDD.n3212 VDD.n3211 212.329
R12717 VDD.n3212 VDD.n3210 212.329
R12718 VDD.n3122 VDD.n3121 212.329
R12719 VDD.n3121 VDD.n3119 212.329
R12720 VDD.n3127 VDD.n3125 212.329
R12721 VDD.n3125 VDD.n3124 212.329
R12722 VDD.n3112 VDD.n3110 212.329
R12723 VDD.n3113 VDD.n3112 212.329
R12724 VDD.n3208 VDD.n3207 212.329
R12725 VDD.n3208 VDD.n3109 212.329
R12726 VDD.n3195 VDD.n3194 212.329
R12727 VDD.n3194 VDD.n3192 212.329
R12728 VDD.n3200 VDD.n3198 212.329
R12729 VDD.n3198 VDD.n3197 212.329
R12730 VDD.n3179 VDD.n3178 212.329
R12731 VDD.n3178 VDD.n3176 212.329
R12732 VDD.n3184 VDD.n3182 212.329
R12733 VDD.n3182 VDD.n3181 212.329
R12734 VDD.n3168 VDD.n3165 212.329
R12735 VDD.n3169 VDD.n3168 212.329
R12736 VDD.n3156 VDD.n3155 212.329
R12737 VDD.n3155 VDD.n3153 212.329
R12738 VDD.n3161 VDD.n3159 212.329
R12739 VDD.n3159 VDD.n3158 212.329
R12740 VDD.n3140 VDD.n3139 212.329
R12741 VDD.n3139 VDD.n3137 212.329
R12742 VDD.n3145 VDD.n3143 212.329
R12743 VDD.n3143 VDD.n3142 212.329
R12744 VDD.n3091 VDD.n3089 212.329
R12745 VDD.n3092 VDD.n3091 212.329
R12746 VDD.n3098 VDD.n3097 212.329
R12747 VDD.n3098 VDD.n3088 212.329
R12748 VDD.n3073 VDD.n3072 212.329
R12749 VDD.n3072 VDD.n3070 212.329
R12750 VDD.n3219 VDD.n3074 212.329
R12751 VDD.n3075 VDD.n3074 212.329
R12752 VDD.n3103 VDD.n3066 212.329
R12753 VDD.n3103 VDD.n3102 212.329
R12754 VDD.n3230 VDD.n3229 212.329
R12755 VDD.n3229 VDD.n3228 212.329
R12756 VDD.n3473 VDD.n3286 212.329
R12757 VDD.n3473 VDD.n3287 212.329
R12758 VDD.n3295 VDD.n3294 212.329
R12759 VDD.n3294 VDD.n3293 212.329
R12760 VDD.n3340 VDD.n3339 212.329
R12761 VDD.n3340 VDD.n3338 212.329
R12762 VDD.n3318 VDD.n3317 212.329
R12763 VDD.n3318 VDD.n3316 212.329
R12764 VDD.n3471 VDD.n3470 212.329
R12765 VDD.n3471 VDD.n3469 212.329
R12766 VDD.n3381 VDD.n3380 212.329
R12767 VDD.n3380 VDD.n3378 212.329
R12768 VDD.n3386 VDD.n3384 212.329
R12769 VDD.n3384 VDD.n3383 212.329
R12770 VDD.n3371 VDD.n3369 212.329
R12771 VDD.n3372 VDD.n3371 212.329
R12772 VDD.n3467 VDD.n3466 212.329
R12773 VDD.n3467 VDD.n3368 212.329
R12774 VDD.n3454 VDD.n3453 212.329
R12775 VDD.n3453 VDD.n3451 212.329
R12776 VDD.n3459 VDD.n3457 212.329
R12777 VDD.n3457 VDD.n3456 212.329
R12778 VDD.n3438 VDD.n3437 212.329
R12779 VDD.n3437 VDD.n3435 212.329
R12780 VDD.n3443 VDD.n3441 212.329
R12781 VDD.n3441 VDD.n3440 212.329
R12782 VDD.n3427 VDD.n3424 212.329
R12783 VDD.n3428 VDD.n3427 212.329
R12784 VDD.n3415 VDD.n3414 212.329
R12785 VDD.n3414 VDD.n3412 212.329
R12786 VDD.n3420 VDD.n3418 212.329
R12787 VDD.n3418 VDD.n3417 212.329
R12788 VDD.n3399 VDD.n3398 212.329
R12789 VDD.n3398 VDD.n3396 212.329
R12790 VDD.n3404 VDD.n3402 212.329
R12791 VDD.n3402 VDD.n3401 212.329
R12792 VDD.n3350 VDD.n3348 212.329
R12793 VDD.n3351 VDD.n3350 212.329
R12794 VDD.n3357 VDD.n3356 212.329
R12795 VDD.n3357 VDD.n3347 212.329
R12796 VDD.n3332 VDD.n3331 212.329
R12797 VDD.n3331 VDD.n3329 212.329
R12798 VDD.n3478 VDD.n3333 212.329
R12799 VDD.n3334 VDD.n3333 212.329
R12800 VDD.n3362 VDD.n3325 212.329
R12801 VDD.n3362 VDD.n3361 212.329
R12802 VDD.n3489 VDD.n3488 212.329
R12803 VDD.n3488 VDD.n3487 212.329
R12804 VDD.n3732 VDD.n3545 212.329
R12805 VDD.n3732 VDD.n3546 212.329
R12806 VDD.n3554 VDD.n3553 212.329
R12807 VDD.n3553 VDD.n3552 212.329
R12808 VDD.n3599 VDD.n3598 212.329
R12809 VDD.n3599 VDD.n3597 212.329
R12810 VDD.n3577 VDD.n3576 212.329
R12811 VDD.n3577 VDD.n3575 212.329
R12812 VDD.n3730 VDD.n3729 212.329
R12813 VDD.n3730 VDD.n3728 212.329
R12814 VDD.n3640 VDD.n3639 212.329
R12815 VDD.n3639 VDD.n3637 212.329
R12816 VDD.n3645 VDD.n3643 212.329
R12817 VDD.n3643 VDD.n3642 212.329
R12818 VDD.n3630 VDD.n3628 212.329
R12819 VDD.n3631 VDD.n3630 212.329
R12820 VDD.n3726 VDD.n3725 212.329
R12821 VDD.n3726 VDD.n3627 212.329
R12822 VDD.n3713 VDD.n3712 212.329
R12823 VDD.n3712 VDD.n3710 212.329
R12824 VDD.n3718 VDD.n3716 212.329
R12825 VDD.n3716 VDD.n3715 212.329
R12826 VDD.n3697 VDD.n3696 212.329
R12827 VDD.n3696 VDD.n3694 212.329
R12828 VDD.n3702 VDD.n3700 212.329
R12829 VDD.n3700 VDD.n3699 212.329
R12830 VDD.n3686 VDD.n3683 212.329
R12831 VDD.n3687 VDD.n3686 212.329
R12832 VDD.n3674 VDD.n3673 212.329
R12833 VDD.n3673 VDD.n3671 212.329
R12834 VDD.n3679 VDD.n3677 212.329
R12835 VDD.n3677 VDD.n3676 212.329
R12836 VDD.n3658 VDD.n3657 212.329
R12837 VDD.n3657 VDD.n3655 212.329
R12838 VDD.n3663 VDD.n3661 212.329
R12839 VDD.n3661 VDD.n3660 212.329
R12840 VDD.n3609 VDD.n3607 212.329
R12841 VDD.n3610 VDD.n3609 212.329
R12842 VDD.n3616 VDD.n3615 212.329
R12843 VDD.n3616 VDD.n3606 212.329
R12844 VDD.n3591 VDD.n3590 212.329
R12845 VDD.n3590 VDD.n3588 212.329
R12846 VDD.n3737 VDD.n3592 212.329
R12847 VDD.n3593 VDD.n3592 212.329
R12848 VDD.n3621 VDD.n3584 212.329
R12849 VDD.n3621 VDD.n3620 212.329
R12850 VDD.n3748 VDD.n3747 212.329
R12851 VDD.n3747 VDD.n3746 212.329
R12852 VDD.n3991 VDD.n3804 212.329
R12853 VDD.n3991 VDD.n3805 212.329
R12854 VDD.n3813 VDD.n3812 212.329
R12855 VDD.n3812 VDD.n3811 212.329
R12856 VDD.n3858 VDD.n3857 212.329
R12857 VDD.n3858 VDD.n3856 212.329
R12858 VDD.n3836 VDD.n3835 212.329
R12859 VDD.n3836 VDD.n3834 212.329
R12860 VDD.n3989 VDD.n3988 212.329
R12861 VDD.n3989 VDD.n3987 212.329
R12862 VDD.n3899 VDD.n3898 212.329
R12863 VDD.n3898 VDD.n3896 212.329
R12864 VDD.n3904 VDD.n3902 212.329
R12865 VDD.n3902 VDD.n3901 212.329
R12866 VDD.n3889 VDD.n3887 212.329
R12867 VDD.n3890 VDD.n3889 212.329
R12868 VDD.n3985 VDD.n3984 212.329
R12869 VDD.n3985 VDD.n3886 212.329
R12870 VDD.n3972 VDD.n3971 212.329
R12871 VDD.n3971 VDD.n3969 212.329
R12872 VDD.n3977 VDD.n3975 212.329
R12873 VDD.n3975 VDD.n3974 212.329
R12874 VDD.n3956 VDD.n3955 212.329
R12875 VDD.n3955 VDD.n3953 212.329
R12876 VDD.n3961 VDD.n3959 212.329
R12877 VDD.n3959 VDD.n3958 212.329
R12878 VDD.n3945 VDD.n3942 212.329
R12879 VDD.n3946 VDD.n3945 212.329
R12880 VDD.n3933 VDD.n3932 212.329
R12881 VDD.n3932 VDD.n3930 212.329
R12882 VDD.n3938 VDD.n3936 212.329
R12883 VDD.n3936 VDD.n3935 212.329
R12884 VDD.n3917 VDD.n3916 212.329
R12885 VDD.n3916 VDD.n3914 212.329
R12886 VDD.n3922 VDD.n3920 212.329
R12887 VDD.n3920 VDD.n3919 212.329
R12888 VDD.n3868 VDD.n3866 212.329
R12889 VDD.n3869 VDD.n3868 212.329
R12890 VDD.n3875 VDD.n3874 212.329
R12891 VDD.n3875 VDD.n3865 212.329
R12892 VDD.n3850 VDD.n3849 212.329
R12893 VDD.n3849 VDD.n3847 212.329
R12894 VDD.n3996 VDD.n3851 212.329
R12895 VDD.n3852 VDD.n3851 212.329
R12896 VDD.n3880 VDD.n3843 212.329
R12897 VDD.n3880 VDD.n3879 212.329
R12898 VDD.n4007 VDD.n4006 212.329
R12899 VDD.n4006 VDD.n4005 212.329
R12900 VDD.n4250 VDD.n4063 212.329
R12901 VDD.n4250 VDD.n4064 212.329
R12902 VDD.n4072 VDD.n4071 212.329
R12903 VDD.n4071 VDD.n4070 212.329
R12904 VDD.n4117 VDD.n4116 212.329
R12905 VDD.n4117 VDD.n4115 212.329
R12906 VDD.n4095 VDD.n4094 212.329
R12907 VDD.n4095 VDD.n4093 212.329
R12908 VDD.n4248 VDD.n4247 212.329
R12909 VDD.n4248 VDD.n4246 212.329
R12910 VDD.n4158 VDD.n4157 212.329
R12911 VDD.n4157 VDD.n4155 212.329
R12912 VDD.n4163 VDD.n4161 212.329
R12913 VDD.n4161 VDD.n4160 212.329
R12914 VDD.n4148 VDD.n4146 212.329
R12915 VDD.n4149 VDD.n4148 212.329
R12916 VDD.n4244 VDD.n4243 212.329
R12917 VDD.n4244 VDD.n4145 212.329
R12918 VDD.n4231 VDD.n4230 212.329
R12919 VDD.n4230 VDD.n4228 212.329
R12920 VDD.n4236 VDD.n4234 212.329
R12921 VDD.n4234 VDD.n4233 212.329
R12922 VDD.n4215 VDD.n4214 212.329
R12923 VDD.n4214 VDD.n4212 212.329
R12924 VDD.n4220 VDD.n4218 212.329
R12925 VDD.n4218 VDD.n4217 212.329
R12926 VDD.n4204 VDD.n4201 212.329
R12927 VDD.n4205 VDD.n4204 212.329
R12928 VDD.n4192 VDD.n4191 212.329
R12929 VDD.n4191 VDD.n4189 212.329
R12930 VDD.n4197 VDD.n4195 212.329
R12931 VDD.n4195 VDD.n4194 212.329
R12932 VDD.n4176 VDD.n4175 212.329
R12933 VDD.n4175 VDD.n4173 212.329
R12934 VDD.n4181 VDD.n4179 212.329
R12935 VDD.n4179 VDD.n4178 212.329
R12936 VDD.n4127 VDD.n4125 212.329
R12937 VDD.n4128 VDD.n4127 212.329
R12938 VDD.n4134 VDD.n4133 212.329
R12939 VDD.n4134 VDD.n4124 212.329
R12940 VDD.n4109 VDD.n4108 212.329
R12941 VDD.n4108 VDD.n4106 212.329
R12942 VDD.n4255 VDD.n4110 212.329
R12943 VDD.n4111 VDD.n4110 212.329
R12944 VDD.n4139 VDD.n4102 212.329
R12945 VDD.n4139 VDD.n4138 212.329
R12946 VDD.n4266 VDD.n4265 212.329
R12947 VDD.n4265 VDD.n4264 212.329
R12948 VDD.n4509 VDD.n4322 212.329
R12949 VDD.n4509 VDD.n4323 212.329
R12950 VDD.n4331 VDD.n4330 212.329
R12951 VDD.n4330 VDD.n4329 212.329
R12952 VDD.n4376 VDD.n4375 212.329
R12953 VDD.n4376 VDD.n4374 212.329
R12954 VDD.n4354 VDD.n4353 212.329
R12955 VDD.n4354 VDD.n4352 212.329
R12956 VDD.n4507 VDD.n4506 212.329
R12957 VDD.n4507 VDD.n4505 212.329
R12958 VDD.n4417 VDD.n4416 212.329
R12959 VDD.n4416 VDD.n4414 212.329
R12960 VDD.n4422 VDD.n4420 212.329
R12961 VDD.n4420 VDD.n4419 212.329
R12962 VDD.n4407 VDD.n4405 212.329
R12963 VDD.n4408 VDD.n4407 212.329
R12964 VDD.n4503 VDD.n4502 212.329
R12965 VDD.n4503 VDD.n4404 212.329
R12966 VDD.n4490 VDD.n4489 212.329
R12967 VDD.n4489 VDD.n4487 212.329
R12968 VDD.n4495 VDD.n4493 212.329
R12969 VDD.n4493 VDD.n4492 212.329
R12970 VDD.n4474 VDD.n4473 212.329
R12971 VDD.n4473 VDD.n4471 212.329
R12972 VDD.n4479 VDD.n4477 212.329
R12973 VDD.n4477 VDD.n4476 212.329
R12974 VDD.n4463 VDD.n4460 212.329
R12975 VDD.n4464 VDD.n4463 212.329
R12976 VDD.n4451 VDD.n4450 212.329
R12977 VDD.n4450 VDD.n4448 212.329
R12978 VDD.n4456 VDD.n4454 212.329
R12979 VDD.n4454 VDD.n4453 212.329
R12980 VDD.n4435 VDD.n4434 212.329
R12981 VDD.n4434 VDD.n4432 212.329
R12982 VDD.n4440 VDD.n4438 212.329
R12983 VDD.n4438 VDD.n4437 212.329
R12984 VDD.n4386 VDD.n4384 212.329
R12985 VDD.n4387 VDD.n4386 212.329
R12986 VDD.n4393 VDD.n4392 212.329
R12987 VDD.n4393 VDD.n4383 212.329
R12988 VDD.n4368 VDD.n4367 212.329
R12989 VDD.n4367 VDD.n4365 212.329
R12990 VDD.n4514 VDD.n4369 212.329
R12991 VDD.n4370 VDD.n4369 212.329
R12992 VDD.n4398 VDD.n4361 212.329
R12993 VDD.n4398 VDD.n4397 212.329
R12994 VDD.n4525 VDD.n4524 212.329
R12995 VDD.n4524 VDD.n4523 212.329
R12996 VDD.n5028 VDD.n4558 212.329
R12997 VDD.n5028 VDD.n4557 212.329
R12998 VDD.n5024 VDD.n5023 212.329
R12999 VDD.n5023 VDD.n5022 212.329
R13000 VDD.n5017 VDD.n5016 212.329
R13001 VDD.n5016 VDD.n5015 212.329
R13002 VDD.n5003 VDD.n4569 212.329
R13003 VDD.n5003 VDD.n4568 212.329
R13004 VDD.n4999 VDD.n4998 212.329
R13005 VDD.n4998 VDD.n4997 212.329
R13006 VDD.n4987 VDD.n4577 212.329
R13007 VDD.n4987 VDD.n4576 212.329
R13008 VDD.n4983 VDD.n4982 212.329
R13009 VDD.n4982 VDD.n4981 212.329
R13010 VDD.n4976 VDD.n4975 212.329
R13011 VDD.n4975 VDD.n4974 212.329
R13012 VDD.n4962 VDD.n4588 212.329
R13013 VDD.n4962 VDD.n4587 212.329
R13014 VDD.n4958 VDD.n4957 212.329
R13015 VDD.n4957 VDD.n4956 212.329
R13016 VDD.n4946 VDD.n4596 212.329
R13017 VDD.n4946 VDD.n4595 212.329
R13018 VDD.n4942 VDD.n4941 212.329
R13019 VDD.n4941 VDD.n4940 212.329
R13020 VDD.n4935 VDD.n4934 212.329
R13021 VDD.n4934 VDD.n4933 212.329
R13022 VDD.n4921 VDD.n4607 212.329
R13023 VDD.n4921 VDD.n4606 212.329
R13024 VDD.n4917 VDD.n4916 212.329
R13025 VDD.n4916 VDD.n4915 212.329
R13026 VDD.n4905 VDD.n4615 212.329
R13027 VDD.n4905 VDD.n4614 212.329
R13028 VDD.n4901 VDD.n4900 212.329
R13029 VDD.n4900 VDD.n4899 212.329
R13030 VDD.n4894 VDD.n4893 212.329
R13031 VDD.n4893 VDD.n4892 212.329
R13032 VDD.n4880 VDD.n4626 212.329
R13033 VDD.n4880 VDD.n4625 212.329
R13034 VDD.n4876 VDD.n4875 212.329
R13035 VDD.n4875 VDD.n4874 212.329
R13036 VDD.n4864 VDD.n4634 212.329
R13037 VDD.n4864 VDD.n4633 212.329
R13038 VDD.n4860 VDD.n4859 212.329
R13039 VDD.n4859 VDD.n4858 212.329
R13040 VDD.n4853 VDD.n4852 212.329
R13041 VDD.n4852 VDD.n4851 212.329
R13042 VDD.n4839 VDD.n4645 212.329
R13043 VDD.n4839 VDD.n4644 212.329
R13044 VDD.n4835 VDD.n4834 212.329
R13045 VDD.n4834 VDD.n4833 212.329
R13046 VDD.n4823 VDD.n4653 212.329
R13047 VDD.n4823 VDD.n4652 212.329
R13048 VDD.n4819 VDD.n4818 212.329
R13049 VDD.n4818 VDD.n4817 212.329
R13050 VDD.n4812 VDD.n4811 212.329
R13051 VDD.n4811 VDD.n4810 212.329
R13052 VDD.n4798 VDD.n4664 212.329
R13053 VDD.n4798 VDD.n4663 212.329
R13054 VDD.n4794 VDD.n4793 212.329
R13055 VDD.n4793 VDD.n4792 212.329
R13056 VDD.n4782 VDD.n4672 212.329
R13057 VDD.n4782 VDD.n4671 212.329
R13058 VDD.n4778 VDD.n4777 212.329
R13059 VDD.n4777 VDD.n4776 212.329
R13060 VDD.n4771 VDD.n4770 212.329
R13061 VDD.n4770 VDD.n4769 212.329
R13062 VDD.n4757 VDD.n4683 212.329
R13063 VDD.n4757 VDD.n4682 212.329
R13064 VDD.n4753 VDD.n4752 212.329
R13065 VDD.n4752 VDD.n4751 212.329
R13066 VDD.n4741 VDD.n4691 212.329
R13067 VDD.n4741 VDD.n4690 212.329
R13068 VDD.n4737 VDD.n4736 212.329
R13069 VDD.n4736 VDD.n4735 212.329
R13070 VDD.n4730 VDD.n4729 212.329
R13071 VDD.n4729 VDD.n4728 212.329
R13072 VDD.n4716 VDD.n4702 212.329
R13073 VDD.n4716 VDD.n4701 212.329
R13074 VDD.n4712 VDD.n4711 212.329
R13075 VDD.n4711 VDD.n4710 212.329
R13076 VDD.n7102 VDD.n5037 212.329
R13077 VDD.n5037 VDD.n5035 212.329
R13078 VDD.n6978 VDD.n5171 212.329
R13079 VDD.n5172 VDD.n5171 212.329
R13080 VDD.n6847 VDD.n5299 212.329
R13081 VDD.n5300 VDD.n5299 212.329
R13082 VDD.n6716 VDD.n5427 212.329
R13083 VDD.n5428 VDD.n5427 212.329
R13084 VDD.n6585 VDD.n5555 212.329
R13085 VDD.n5556 VDD.n5555 212.329
R13086 VDD.n6454 VDD.n5683 212.329
R13087 VDD.n5684 VDD.n5683 212.329
R13088 VDD.n6323 VDD.n5811 212.329
R13089 VDD.n5812 VDD.n5811 212.329
R13090 VDD.n6192 VDD.n5939 212.329
R13091 VDD.n5940 VDD.n5939 212.329
R13092 VDD.n5048 VDD.n5043 212.329
R13093 VDD.n5049 VDD.n5048 212.329
R13094 VDD.n7095 VDD.n5042 212.329
R13095 VDD.n7088 VDD.n5042 212.329
R13096 VDD.n5058 VDD.n5054 212.329
R13097 VDD.n5059 VDD.n5058 212.329
R13098 VDD.n7085 VDD.n5053 212.329
R13099 VDD.n7078 VDD.n5053 212.329
R13100 VDD.n5071 VDD.n5064 212.329
R13101 VDD.n5072 VDD.n5071 212.329
R13102 VDD.n7075 VDD.n5063 212.329
R13103 VDD.n7068 VDD.n5063 212.329
R13104 VDD.n5082 VDD.n5077 212.329
R13105 VDD.n5083 VDD.n5082 212.329
R13106 VDD.n7065 VDD.n5076 212.329
R13107 VDD.n7058 VDD.n5076 212.329
R13108 VDD.n5092 VDD.n5088 212.329
R13109 VDD.n5093 VDD.n5092 212.329
R13110 VDD.n7055 VDD.n5087 212.329
R13111 VDD.n7048 VDD.n5087 212.329
R13112 VDD.n5105 VDD.n5098 212.329
R13113 VDD.n5106 VDD.n5105 212.329
R13114 VDD.n7045 VDD.n5097 212.329
R13115 VDD.n7038 VDD.n5097 212.329
R13116 VDD.n7035 VDD.n7034 212.329
R13117 VDD.n7034 VDD.n7033 212.329
R13118 VDD.n5120 VDD.n5114 212.329
R13119 VDD.n5121 VDD.n5120 212.329
R13120 VDD.n7028 VDD.n5113 212.329
R13121 VDD.n7021 VDD.n5113 212.329
R13122 VDD.n5133 VDD.n5126 212.329
R13123 VDD.n5134 VDD.n5133 212.329
R13124 VDD.n7018 VDD.n5125 212.329
R13125 VDD.n7011 VDD.n5125 212.329
R13126 VDD.n5144 VDD.n5139 212.329
R13127 VDD.n5145 VDD.n5144 212.329
R13128 VDD.n7008 VDD.n5138 212.329
R13129 VDD.n7001 VDD.n5138 212.329
R13130 VDD.n5154 VDD.n5150 212.329
R13131 VDD.n5155 VDD.n5154 212.329
R13132 VDD.n6998 VDD.n5149 212.329
R13133 VDD.n6991 VDD.n5149 212.329
R13134 VDD.n5167 VDD.n5160 212.329
R13135 VDD.n5168 VDD.n5167 212.329
R13136 VDD.n6988 VDD.n5159 212.329
R13137 VDD.n6981 VDD.n5159 212.329
R13138 VDD.n6960 VDD.n6959 212.329
R13139 VDD.n6960 VDD.n6958 212.329
R13140 VDD.n6969 VDD.n6968 212.329
R13141 VDD.n6969 VDD.n6967 212.329
R13142 VDD.n5186 VDD.n5183 212.329
R13143 VDD.n5187 VDD.n5186 212.329
R13144 VDD.n6954 VDD.n5182 212.329
R13145 VDD.n6947 VDD.n5182 212.329
R13146 VDD.n5199 VDD.n5192 212.329
R13147 VDD.n5200 VDD.n5199 212.329
R13148 VDD.n6944 VDD.n5191 212.329
R13149 VDD.n6937 VDD.n5191 212.329
R13150 VDD.n5210 VDD.n5205 212.329
R13151 VDD.n5211 VDD.n5210 212.329
R13152 VDD.n6934 VDD.n5204 212.329
R13153 VDD.n6927 VDD.n5204 212.329
R13154 VDD.n5220 VDD.n5216 212.329
R13155 VDD.n5221 VDD.n5220 212.329
R13156 VDD.n6924 VDD.n5215 212.329
R13157 VDD.n6917 VDD.n5215 212.329
R13158 VDD.n5233 VDD.n5226 212.329
R13159 VDD.n5234 VDD.n5233 212.329
R13160 VDD.n6914 VDD.n5225 212.329
R13161 VDD.n6907 VDD.n5225 212.329
R13162 VDD.n6904 VDD.n6903 212.329
R13163 VDD.n6903 VDD.n6902 212.329
R13164 VDD.n5248 VDD.n5242 212.329
R13165 VDD.n5249 VDD.n5248 212.329
R13166 VDD.n6897 VDD.n5241 212.329
R13167 VDD.n6890 VDD.n5241 212.329
R13168 VDD.n5261 VDD.n5254 212.329
R13169 VDD.n5262 VDD.n5261 212.329
R13170 VDD.n6887 VDD.n5253 212.329
R13171 VDD.n6880 VDD.n5253 212.329
R13172 VDD.n5272 VDD.n5267 212.329
R13173 VDD.n5273 VDD.n5272 212.329
R13174 VDD.n6877 VDD.n5266 212.329
R13175 VDD.n6870 VDD.n5266 212.329
R13176 VDD.n5282 VDD.n5278 212.329
R13177 VDD.n5283 VDD.n5282 212.329
R13178 VDD.n6867 VDD.n5277 212.329
R13179 VDD.n6860 VDD.n5277 212.329
R13180 VDD.n5295 VDD.n5288 212.329
R13181 VDD.n5296 VDD.n5295 212.329
R13182 VDD.n6857 VDD.n5287 212.329
R13183 VDD.n6850 VDD.n5287 212.329
R13184 VDD.n6829 VDD.n6828 212.329
R13185 VDD.n6829 VDD.n6827 212.329
R13186 VDD.n6838 VDD.n6837 212.329
R13187 VDD.n6838 VDD.n6836 212.329
R13188 VDD.n5314 VDD.n5311 212.329
R13189 VDD.n5315 VDD.n5314 212.329
R13190 VDD.n6823 VDD.n5310 212.329
R13191 VDD.n6816 VDD.n5310 212.329
R13192 VDD.n5327 VDD.n5320 212.329
R13193 VDD.n5328 VDD.n5327 212.329
R13194 VDD.n6813 VDD.n5319 212.329
R13195 VDD.n6806 VDD.n5319 212.329
R13196 VDD.n5338 VDD.n5333 212.329
R13197 VDD.n5339 VDD.n5338 212.329
R13198 VDD.n6803 VDD.n5332 212.329
R13199 VDD.n6796 VDD.n5332 212.329
R13200 VDD.n5348 VDD.n5344 212.329
R13201 VDD.n5349 VDD.n5348 212.329
R13202 VDD.n6793 VDD.n5343 212.329
R13203 VDD.n6786 VDD.n5343 212.329
R13204 VDD.n5361 VDD.n5354 212.329
R13205 VDD.n5362 VDD.n5361 212.329
R13206 VDD.n6783 VDD.n5353 212.329
R13207 VDD.n6776 VDD.n5353 212.329
R13208 VDD.n6773 VDD.n6772 212.329
R13209 VDD.n6772 VDD.n6771 212.329
R13210 VDD.n5376 VDD.n5370 212.329
R13211 VDD.n5377 VDD.n5376 212.329
R13212 VDD.n6766 VDD.n5369 212.329
R13213 VDD.n6759 VDD.n5369 212.329
R13214 VDD.n5389 VDD.n5382 212.329
R13215 VDD.n5390 VDD.n5389 212.329
R13216 VDD.n6756 VDD.n5381 212.329
R13217 VDD.n6749 VDD.n5381 212.329
R13218 VDD.n5400 VDD.n5395 212.329
R13219 VDD.n5401 VDD.n5400 212.329
R13220 VDD.n6746 VDD.n5394 212.329
R13221 VDD.n6739 VDD.n5394 212.329
R13222 VDD.n5410 VDD.n5406 212.329
R13223 VDD.n5411 VDD.n5410 212.329
R13224 VDD.n6736 VDD.n5405 212.329
R13225 VDD.n6729 VDD.n5405 212.329
R13226 VDD.n5423 VDD.n5416 212.329
R13227 VDD.n5424 VDD.n5423 212.329
R13228 VDD.n6726 VDD.n5415 212.329
R13229 VDD.n6719 VDD.n5415 212.329
R13230 VDD.n6698 VDD.n6697 212.329
R13231 VDD.n6698 VDD.n6696 212.329
R13232 VDD.n6707 VDD.n6706 212.329
R13233 VDD.n6707 VDD.n6705 212.329
R13234 VDD.n5442 VDD.n5439 212.329
R13235 VDD.n5443 VDD.n5442 212.329
R13236 VDD.n6692 VDD.n5438 212.329
R13237 VDD.n6685 VDD.n5438 212.329
R13238 VDD.n5455 VDD.n5448 212.329
R13239 VDD.n5456 VDD.n5455 212.329
R13240 VDD.n6682 VDD.n5447 212.329
R13241 VDD.n6675 VDD.n5447 212.329
R13242 VDD.n5466 VDD.n5461 212.329
R13243 VDD.n5467 VDD.n5466 212.329
R13244 VDD.n6672 VDD.n5460 212.329
R13245 VDD.n6665 VDD.n5460 212.329
R13246 VDD.n5476 VDD.n5472 212.329
R13247 VDD.n5477 VDD.n5476 212.329
R13248 VDD.n6662 VDD.n5471 212.329
R13249 VDD.n6655 VDD.n5471 212.329
R13250 VDD.n5489 VDD.n5482 212.329
R13251 VDD.n5490 VDD.n5489 212.329
R13252 VDD.n6652 VDD.n5481 212.329
R13253 VDD.n6645 VDD.n5481 212.329
R13254 VDD.n6642 VDD.n6641 212.329
R13255 VDD.n6641 VDD.n6640 212.329
R13256 VDD.n5504 VDD.n5498 212.329
R13257 VDD.n5505 VDD.n5504 212.329
R13258 VDD.n6635 VDD.n5497 212.329
R13259 VDD.n6628 VDD.n5497 212.329
R13260 VDD.n5517 VDD.n5510 212.329
R13261 VDD.n5518 VDD.n5517 212.329
R13262 VDD.n6625 VDD.n5509 212.329
R13263 VDD.n6618 VDD.n5509 212.329
R13264 VDD.n5528 VDD.n5523 212.329
R13265 VDD.n5529 VDD.n5528 212.329
R13266 VDD.n6615 VDD.n5522 212.329
R13267 VDD.n6608 VDD.n5522 212.329
R13268 VDD.n5538 VDD.n5534 212.329
R13269 VDD.n5539 VDD.n5538 212.329
R13270 VDD.n6605 VDD.n5533 212.329
R13271 VDD.n6598 VDD.n5533 212.329
R13272 VDD.n5551 VDD.n5544 212.329
R13273 VDD.n5552 VDD.n5551 212.329
R13274 VDD.n6595 VDD.n5543 212.329
R13275 VDD.n6588 VDD.n5543 212.329
R13276 VDD.n6567 VDD.n6566 212.329
R13277 VDD.n6567 VDD.n6565 212.329
R13278 VDD.n6576 VDD.n6575 212.329
R13279 VDD.n6576 VDD.n6574 212.329
R13280 VDD.n5570 VDD.n5567 212.329
R13281 VDD.n5571 VDD.n5570 212.329
R13282 VDD.n6561 VDD.n5566 212.329
R13283 VDD.n6554 VDD.n5566 212.329
R13284 VDD.n5583 VDD.n5576 212.329
R13285 VDD.n5584 VDD.n5583 212.329
R13286 VDD.n6551 VDD.n5575 212.329
R13287 VDD.n6544 VDD.n5575 212.329
R13288 VDD.n5594 VDD.n5589 212.329
R13289 VDD.n5595 VDD.n5594 212.329
R13290 VDD.n6541 VDD.n5588 212.329
R13291 VDD.n6534 VDD.n5588 212.329
R13292 VDD.n5604 VDD.n5600 212.329
R13293 VDD.n5605 VDD.n5604 212.329
R13294 VDD.n6531 VDD.n5599 212.329
R13295 VDD.n6524 VDD.n5599 212.329
R13296 VDD.n5617 VDD.n5610 212.329
R13297 VDD.n5618 VDD.n5617 212.329
R13298 VDD.n6521 VDD.n5609 212.329
R13299 VDD.n6514 VDD.n5609 212.329
R13300 VDD.n6511 VDD.n6510 212.329
R13301 VDD.n6510 VDD.n6509 212.329
R13302 VDD.n5632 VDD.n5626 212.329
R13303 VDD.n5633 VDD.n5632 212.329
R13304 VDD.n6504 VDD.n5625 212.329
R13305 VDD.n6497 VDD.n5625 212.329
R13306 VDD.n5645 VDD.n5638 212.329
R13307 VDD.n5646 VDD.n5645 212.329
R13308 VDD.n6494 VDD.n5637 212.329
R13309 VDD.n6487 VDD.n5637 212.329
R13310 VDD.n5656 VDD.n5651 212.329
R13311 VDD.n5657 VDD.n5656 212.329
R13312 VDD.n6484 VDD.n5650 212.329
R13313 VDD.n6477 VDD.n5650 212.329
R13314 VDD.n5666 VDD.n5662 212.329
R13315 VDD.n5667 VDD.n5666 212.329
R13316 VDD.n6474 VDD.n5661 212.329
R13317 VDD.n6467 VDD.n5661 212.329
R13318 VDD.n5679 VDD.n5672 212.329
R13319 VDD.n5680 VDD.n5679 212.329
R13320 VDD.n6464 VDD.n5671 212.329
R13321 VDD.n6457 VDD.n5671 212.329
R13322 VDD.n6436 VDD.n6435 212.329
R13323 VDD.n6436 VDD.n6434 212.329
R13324 VDD.n6445 VDD.n6444 212.329
R13325 VDD.n6445 VDD.n6443 212.329
R13326 VDD.n5698 VDD.n5695 212.329
R13327 VDD.n5699 VDD.n5698 212.329
R13328 VDD.n6430 VDD.n5694 212.329
R13329 VDD.n6423 VDD.n5694 212.329
R13330 VDD.n5711 VDD.n5704 212.329
R13331 VDD.n5712 VDD.n5711 212.329
R13332 VDD.n6420 VDD.n5703 212.329
R13333 VDD.n6413 VDD.n5703 212.329
R13334 VDD.n5722 VDD.n5717 212.329
R13335 VDD.n5723 VDD.n5722 212.329
R13336 VDD.n6410 VDD.n5716 212.329
R13337 VDD.n6403 VDD.n5716 212.329
R13338 VDD.n5732 VDD.n5728 212.329
R13339 VDD.n5733 VDD.n5732 212.329
R13340 VDD.n6400 VDD.n5727 212.329
R13341 VDD.n6393 VDD.n5727 212.329
R13342 VDD.n5745 VDD.n5738 212.329
R13343 VDD.n5746 VDD.n5745 212.329
R13344 VDD.n6390 VDD.n5737 212.329
R13345 VDD.n6383 VDD.n5737 212.329
R13346 VDD.n6380 VDD.n6379 212.329
R13347 VDD.n6379 VDD.n6378 212.329
R13348 VDD.n5760 VDD.n5754 212.329
R13349 VDD.n5761 VDD.n5760 212.329
R13350 VDD.n6373 VDD.n5753 212.329
R13351 VDD.n6366 VDD.n5753 212.329
R13352 VDD.n5773 VDD.n5766 212.329
R13353 VDD.n5774 VDD.n5773 212.329
R13354 VDD.n6363 VDD.n5765 212.329
R13355 VDD.n6356 VDD.n5765 212.329
R13356 VDD.n5784 VDD.n5779 212.329
R13357 VDD.n5785 VDD.n5784 212.329
R13358 VDD.n6353 VDD.n5778 212.329
R13359 VDD.n6346 VDD.n5778 212.329
R13360 VDD.n5794 VDD.n5790 212.329
R13361 VDD.n5795 VDD.n5794 212.329
R13362 VDD.n6343 VDD.n5789 212.329
R13363 VDD.n6336 VDD.n5789 212.329
R13364 VDD.n5807 VDD.n5800 212.329
R13365 VDD.n5808 VDD.n5807 212.329
R13366 VDD.n6333 VDD.n5799 212.329
R13367 VDD.n6326 VDD.n5799 212.329
R13368 VDD.n6305 VDD.n6304 212.329
R13369 VDD.n6305 VDD.n6303 212.329
R13370 VDD.n6314 VDD.n6313 212.329
R13371 VDD.n6314 VDD.n6312 212.329
R13372 VDD.n5826 VDD.n5823 212.329
R13373 VDD.n5827 VDD.n5826 212.329
R13374 VDD.n6299 VDD.n5822 212.329
R13375 VDD.n6292 VDD.n5822 212.329
R13376 VDD.n5839 VDD.n5832 212.329
R13377 VDD.n5840 VDD.n5839 212.329
R13378 VDD.n6289 VDD.n5831 212.329
R13379 VDD.n6282 VDD.n5831 212.329
R13380 VDD.n5850 VDD.n5845 212.329
R13381 VDD.n5851 VDD.n5850 212.329
R13382 VDD.n6279 VDD.n5844 212.329
R13383 VDD.n6272 VDD.n5844 212.329
R13384 VDD.n5860 VDD.n5856 212.329
R13385 VDD.n5861 VDD.n5860 212.329
R13386 VDD.n6269 VDD.n5855 212.329
R13387 VDD.n6262 VDD.n5855 212.329
R13388 VDD.n5873 VDD.n5866 212.329
R13389 VDD.n5874 VDD.n5873 212.329
R13390 VDD.n6259 VDD.n5865 212.329
R13391 VDD.n6252 VDD.n5865 212.329
R13392 VDD.n6249 VDD.n6248 212.329
R13393 VDD.n6248 VDD.n6247 212.329
R13394 VDD.n5888 VDD.n5882 212.329
R13395 VDD.n5889 VDD.n5888 212.329
R13396 VDD.n6242 VDD.n5881 212.329
R13397 VDD.n6235 VDD.n5881 212.329
R13398 VDD.n5901 VDD.n5894 212.329
R13399 VDD.n5902 VDD.n5901 212.329
R13400 VDD.n6232 VDD.n5893 212.329
R13401 VDD.n6225 VDD.n5893 212.329
R13402 VDD.n5912 VDD.n5907 212.329
R13403 VDD.n5913 VDD.n5912 212.329
R13404 VDD.n6222 VDD.n5906 212.329
R13405 VDD.n6215 VDD.n5906 212.329
R13406 VDD.n5922 VDD.n5918 212.329
R13407 VDD.n5923 VDD.n5922 212.329
R13408 VDD.n6212 VDD.n5917 212.329
R13409 VDD.n6205 VDD.n5917 212.329
R13410 VDD.n5935 VDD.n5928 212.329
R13411 VDD.n5936 VDD.n5935 212.329
R13412 VDD.n6202 VDD.n5927 212.329
R13413 VDD.n6195 VDD.n5927 212.329
R13414 VDD.n6174 VDD.n6173 212.329
R13415 VDD.n6174 VDD.n6172 212.329
R13416 VDD.n6183 VDD.n6182 212.329
R13417 VDD.n6183 VDD.n6181 212.329
R13418 VDD.n5954 VDD.n5951 212.329
R13419 VDD.n5955 VDD.n5954 212.329
R13420 VDD.n6168 VDD.n5950 212.329
R13421 VDD.n6161 VDD.n5950 212.329
R13422 VDD.n5967 VDD.n5960 212.329
R13423 VDD.n5968 VDD.n5967 212.329
R13424 VDD.n6158 VDD.n5959 212.329
R13425 VDD.n6151 VDD.n5959 212.329
R13426 VDD.n5978 VDD.n5973 212.329
R13427 VDD.n5979 VDD.n5978 212.329
R13428 VDD.n6148 VDD.n5972 212.329
R13429 VDD.n6141 VDD.n5972 212.329
R13430 VDD.n5988 VDD.n5984 212.329
R13431 VDD.n5989 VDD.n5988 212.329
R13432 VDD.n6138 VDD.n5983 212.329
R13433 VDD.n6131 VDD.n5983 212.329
R13434 VDD.n6001 VDD.n5994 212.329
R13435 VDD.n6002 VDD.n6001 212.329
R13436 VDD.n6128 VDD.n5993 212.329
R13437 VDD.n6121 VDD.n5993 212.329
R13438 VDD.n6118 VDD.n6117 212.329
R13439 VDD.n6117 VDD.n6116 212.329
R13440 VDD.n6016 VDD.n6010 212.329
R13441 VDD.n6017 VDD.n6016 212.329
R13442 VDD.n6111 VDD.n6009 212.329
R13443 VDD.n6104 VDD.n6009 212.329
R13444 VDD.n6029 VDD.n6022 212.329
R13445 VDD.n6030 VDD.n6029 212.329
R13446 VDD.n6101 VDD.n6021 212.329
R13447 VDD.n6094 VDD.n6021 212.329
R13448 VDD.n6040 VDD.n6035 212.329
R13449 VDD.n6041 VDD.n6040 212.329
R13450 VDD.n6091 VDD.n6034 212.329
R13451 VDD.n6084 VDD.n6034 212.329
R13452 VDD.n6050 VDD.n6046 212.329
R13453 VDD.n6051 VDD.n6050 212.329
R13454 VDD.n6081 VDD.n6045 212.329
R13455 VDD.n6074 VDD.n6045 212.329
R13456 VDD.n6059 VDD.n6056 212.329
R13457 VDD.n6060 VDD.n6059 212.329
R13458 VDD.n6071 VDD.n6055 212.329
R13459 VDD.n6061 VDD.n6055 212.329
R13460 VDD.n7112 VDD.n7111 212.329
R13461 VDD.n7113 VDD.n7112 212.329
R13462 VDD.n7119 VDD.n7118 212.329
R13463 VDD.n7120 VDD.n7119 212.329
R13464 VDD.n7125 VDD.n137 212.329
R13465 VDD.n137 VDD.n135 212.329
R13466 VDD.n7133 VDD.n7132 212.329
R13467 VDD.n7134 VDD.n7133 212.329
R13468 VDD.n7140 VDD.n7139 212.329
R13469 VDD.n7141 VDD.n7140 212.329
R13470 VDD.n7146 VDD.n118 212.329
R13471 VDD.n118 VDD.n116 212.329
R13472 VDD.n7154 VDD.n7153 212.329
R13473 VDD.n7155 VDD.n7154 212.329
R13474 VDD.n7161 VDD.n7160 212.329
R13475 VDD.n7162 VDD.n7161 212.329
R13476 VDD.n7167 VDD.n99 212.329
R13477 VDD.n99 VDD.n97 212.329
R13478 VDD.n7175 VDD.n7174 212.329
R13479 VDD.n7176 VDD.n7175 212.329
R13480 VDD.n7182 VDD.n7181 212.329
R13481 VDD.n7183 VDD.n7182 212.329
R13482 VDD.n7188 VDD.n80 212.329
R13483 VDD.n80 VDD.n78 212.329
R13484 VDD.n7196 VDD.n7195 212.329
R13485 VDD.n7197 VDD.n7196 212.329
R13486 VDD.n7203 VDD.n7202 212.329
R13487 VDD.n7204 VDD.n7203 212.329
R13488 VDD.n7209 VDD.n61 212.329
R13489 VDD.n61 VDD.n59 212.329
R13490 VDD.n7217 VDD.n7216 212.329
R13491 VDD.n7218 VDD.n7217 212.329
R13492 VDD.n7224 VDD.n7223 212.329
R13493 VDD.n7225 VDD.n7224 212.329
R13494 VDD.n7230 VDD.n42 212.329
R13495 VDD.n42 VDD.n40 212.329
R13496 VDD.n7238 VDD.n7237 212.329
R13497 VDD.n7239 VDD.n7238 212.329
R13498 VDD.n7245 VDD.n7244 212.329
R13499 VDD.n7246 VDD.n7245 212.329
R13500 VDD.n7251 VDD.n23 212.329
R13501 VDD.n23 VDD.n21 212.329
R13502 VDD.n7259 VDD.n7258 212.329
R13503 VDD.n7260 VDD.n7259 212.329
R13504 VDD.n7266 VDD.n7265 212.329
R13505 VDD.n7267 VDD.n7266 212.329
R13506 VDD.n7272 VDD.n4 212.329
R13507 VDD.n4 VDD.n2 212.329
R13508 VDD.n150 VDD.t916 176.65
R13509 VDD.n131 VDD.t881 176.65
R13510 VDD.n112 VDD.t545 176.65
R13511 VDD.n93 VDD.t97 176.65
R13512 VDD.n74 VDD.t403 176.65
R13513 VDD.n55 VDD.t631 176.65
R13514 VDD.n36 VDD.t302 176.65
R13515 VDD.n17 VDD.t315 176.65
R13516 VDD.n5010 VDD.t333 169.018
R13517 VDD.n4969 VDD.t586 169.018
R13518 VDD.n4928 VDD.t550 169.018
R13519 VDD.n4887 VDD.t527 169.018
R13520 VDD.n4846 VDD.t597 169.018
R13521 VDD.n4805 VDD.t646 169.018
R13522 VDD.n4764 VDD.t726 169.018
R13523 VDD.n4723 VDD.t870 169.018
R13524 VDD.n6037 VDD.t692 169.018
R13525 VDD.n6037 VDD.t357 169.018
R13526 VDD.n5975 VDD.t697 169.018
R13527 VDD.n5975 VDD.t389 169.018
R13528 VDD.n6188 VDD.t475 169.018
R13529 VDD.n6188 VDD.t656 169.018
R13530 VDD.n6189 VDD.t717 169.018
R13531 VDD.n5909 VDD.t559 169.018
R13532 VDD.n5909 VDD.t541 169.018
R13533 VDD.n5847 VDD.t766 169.018
R13534 VDD.n5847 VDD.t539 169.018
R13535 VDD.n6319 VDD.t537 169.018
R13536 VDD.n6319 VDD.t570 169.018
R13537 VDD.n6320 VDD.t721 169.018
R13538 VDD.n5781 VDD.t391 169.018
R13539 VDD.n5781 VDD.t739 169.018
R13540 VDD.n5719 VDD.t562 169.018
R13541 VDD.n5719 VDD.t792 169.018
R13542 VDD.n6450 VDD.t286 169.018
R13543 VDD.n6450 VDD.t765 169.018
R13544 VDD.n6451 VDD.t451 169.018
R13545 VDD.n5653 VDD.t640 169.018
R13546 VDD.n5653 VDD.t753 169.018
R13547 VDD.n5591 VDD.t638 169.018
R13548 VDD.n5591 VDD.t752 169.018
R13549 VDD.n6581 VDD.t754 169.018
R13550 VDD.n6581 VDD.t564 169.018
R13551 VDD.n6582 VDD.t17 169.018
R13552 VDD.n5525 VDD.t636 169.018
R13553 VDD.n5525 VDD.t788 169.018
R13554 VDD.n5463 VDD.t898 169.018
R13555 VDD.n5463 VDD.t353 169.018
R13556 VDD.n6712 VDD.t365 169.018
R13557 VDD.n6712 VDD.t560 169.018
R13558 VDD.n6713 VDD.t719 169.018
R13559 VDD.n5397 VDD.t569 169.018
R13560 VDD.n5397 VDD.t731 169.018
R13561 VDD.n5335 VDD.t359 169.018
R13562 VDD.n5335 VDD.t590 169.018
R13563 VDD.n6843 VDD.t494 169.018
R13564 VDD.n6843 VDD.t565 169.018
R13565 VDD.n6844 VDD.t276 169.018
R13566 VDD.n5269 VDD.t392 169.018
R13567 VDD.n5269 VDD.t91 169.018
R13568 VDD.n5207 VDD.t567 169.018
R13569 VDD.n5207 VDD.t705 169.018
R13570 VDD.n6974 VDD.t479 169.018
R13571 VDD.n6974 VDD.t767 169.018
R13572 VDD.n6975 VDD.t453 169.018
R13573 VDD.n5141 VDD.t764 169.018
R13574 VDD.n5141 VDD.t914 169.018
R13575 VDD.n5079 VDD.t476 169.018
R13576 VDD.n5079 VDD.t409 169.018
R13577 VDD.n5045 VDD.t913 169.018
R13578 VDD.n5045 VDD.t644 169.018
R13579 VDD.n7105 VDD.t756 169.018
R13580 VDD.n5116 VDD.t615 169.018
R13581 VDD.n5244 VDD.t377 169.018
R13582 VDD.n5372 VDD.t486 169.018
R13583 VDD.n5500 VDD.t41 169.018
R13584 VDD.n5628 VDD.t900 169.018
R13585 VDD.n5756 VDD.t736 169.018
R13586 VDD.n5884 VDD.t840 169.018
R13587 VDD.n6012 VDD.t461 169.018
R13588 VDD.n1 VDD.t510 169.012
R13589 VDD.n20 VDD.t896 169.012
R13590 VDD.n39 VDD.t384 169.012
R13591 VDD.n58 VDD.t715 169.012
R13592 VDD.n77 VDD.t299 169.012
R13593 VDD.n96 VDD.t856 169.012
R13594 VDD.n115 VDD.t904 169.012
R13595 VDD.n134 VDD.t774 169.012
R13596 VDD.n4555 VDD.t797 168.635
R13597 VDD.n4555 VDD.t820 168.635
R13598 VDD.n4566 VDD.t270 168.635
R13599 VDD.n4566 VDD.t469 168.635
R13600 VDD.n4574 VDD.t584 168.635
R13601 VDD.n4574 VDD.t253 168.635
R13602 VDD.n4585 VDD.t704 168.635
R13603 VDD.n4585 VDD.t889 168.635
R13604 VDD.n4593 VDD.t599 168.635
R13605 VDD.n4593 VDD.t293 168.635
R13606 VDD.n4604 VDD.t733 168.635
R13607 VDD.n4604 VDD.t32 168.635
R13608 VDD.n4612 VDD.t892 168.635
R13609 VDD.n4612 VDD.t829 168.635
R13610 VDD.n4623 VDD.t455 168.635
R13611 VDD.n4623 VDD.t60 168.635
R13612 VDD.n4631 VDD.t595 168.635
R13613 VDD.n4631 VDD.t745 168.635
R13614 VDD.n4642 VDD.t369 168.635
R13615 VDD.n4642 VDD.t554 168.635
R13616 VDD.n4650 VDD.t297 168.635
R13617 VDD.n4650 VDD.t823 168.635
R13618 VDD.n4661 VDD.t795 168.635
R13619 VDD.n4661 VDD.t88 168.635
R13620 VDD.n4669 VDD.t423 168.635
R13621 VDD.n4669 VDD.t225 168.635
R13622 VDD.n4680 VDD.t879 168.635
R13623 VDD.n4680 VDD.t748 168.635
R13624 VDD.n4688 VDD.t843 168.635
R13625 VDD.n4688 VDD.t813 168.635
R13626 VDD.n4699 VDD.t572 168.635
R13627 VDD.n4699 VDD.t341 168.635
R13628 VDD.n6067 VDD.t372 168.635
R13629 VDD.n6067 VDD.t910 168.635
R13630 VDD.n6066 VDD.t524 168.635
R13631 VDD.n6066 VDD.t873 168.635
R13632 VDD.n6025 VDD.t327 168.635
R13633 VDD.n6025 VDD.t317 168.635
R13634 VDD.n6024 VDD.t318 168.635
R13635 VDD.n6024 VDD.t546 168.635
R13636 VDD.n5997 VDD.t619 168.635
R13637 VDD.n5997 VDD.t5 168.635
R13638 VDD.n5996 VDD.t325 168.635
R13639 VDD.n5996 VDD.t885 168.635
R13640 VDD.n5963 VDD.t289 168.635
R13641 VDD.n5963 VDD.t459 168.635
R13642 VDD.n5962 VDD.t784 168.635
R13643 VDD.n5962 VDD.t21 168.635
R13644 VDD.n5931 VDD.t82 168.635
R13645 VDD.n5931 VDD.t28 168.635
R13646 VDD.n5930 VDD.t477 168.635
R13647 VDD.n5930 VDD.t532 168.635
R13648 VDD.n5897 VDD.t283 168.635
R13649 VDD.n5897 VDD.t396 168.635
R13650 VDD.n5896 VDD.t397 168.635
R13651 VDD.n5896 VDD.t574 168.635
R13652 VDD.n5869 VDD.t573 168.635
R13653 VDD.n5869 VDD.t457 168.635
R13654 VDD.n5868 VDD.t281 168.635
R13655 VDD.n5868 VDD.t548 168.635
R13656 VDD.n5835 VDD.t543 168.635
R13657 VDD.n5835 VDD.t838 168.635
R13658 VDD.n5834 VDD.t837 168.635
R13659 VDD.n5834 VDD.t760 168.635
R13660 VDD.n5803 VDD.t875 168.635
R13661 VDD.n5803 VDD.t386 168.635
R13662 VDD.n5802 VDD.t847 168.635
R13663 VDD.n5802 VDD.t805 168.635
R13664 VDD.n5769 VDD.t534 168.635
R13665 VDD.n5769 VDD.t65 168.635
R13666 VDD.n5768 VDD.t66 168.635
R13667 VDD.n5768 VDD.t1 168.635
R13668 VDD.n5741 VDD.t701 168.635
R13669 VDD.n5741 VDD.t3 168.635
R13670 VDD.n5740 VDD.t535 168.635
R13671 VDD.n5740 VDD.t350 168.635
R13672 VDD.n5707 VDD.t424 168.635
R13673 VDD.n5707 VDD.t864 168.635
R13674 VDD.n5706 VDD.t863 168.635
R13675 VDD.n5706 VDD.t278 168.635
R13676 VDD.n5675 VDD.t577 168.635
R13677 VDD.n5675 VDD.t712 168.635
R13678 VDD.n5674 VDD.t496 168.635
R13679 VDD.n5674 VDD.t348 168.635
R13680 VDD.n5641 VDD.t431 168.635
R13681 VDD.n5641 VDD.t504 168.635
R13682 VDD.n5640 VDD.t505 168.635
R13683 VDD.n5640 VDD.t610 168.635
R13684 VDD.n5613 VDD.t528 168.635
R13685 VDD.n5613 VDD.t432 168.635
R13686 VDD.n5612 VDD.t429 168.635
R13687 VDD.n5612 VDD.t79 168.635
R13688 VDD.n5579 VDD.t576 168.635
R13689 VDD.n5579 VDD.t258 168.635
R13690 VDD.n5578 VDD.t901 168.635
R13691 VDD.n5578 VDD.t19 168.635
R13692 VDD.n5547 VDD.t401 168.635
R13693 VDD.n5547 VDD.t300 168.635
R13694 VDD.n5546 VDD.t71 168.635
R13695 VDD.n5546 VDD.t438 168.635
R13696 VDD.n5513 VDD.t738 168.635
R13697 VDD.n5513 VDD.t626 168.635
R13698 VDD.n5512 VDD.t627 168.635
R13699 VDD.n5512 VDD.t307 168.635
R13700 VDD.n5485 VDD.t466 168.635
R13701 VDD.n5485 VDD.t421 168.635
R13702 VDD.n5484 VDD.t737 168.635
R13703 VDD.n5484 VDD.t922 168.635
R13704 VDD.n5451 VDD.t69 168.635
R13705 VDD.n5451 VDD.t39 168.635
R13706 VDD.n5450 VDD.t38 168.635
R13707 VDD.n5450 VDD.t757 168.635
R13708 VDD.n5419 VDD.t288 168.635
R13709 VDD.n5419 VDD.t854 168.635
R13710 VDD.n5418 VDD.t412 168.635
R13711 VDD.n5418 VDD.t499 168.635
R13712 VDD.n5385 VDD.t827 168.635
R13713 VDD.n5385 VDD.t440 168.635
R13714 VDD.n5384 VDD.t441 168.635
R13715 VDD.n5384 VDD.t216 168.635
R13716 VDD.n5357 VDD.t605 168.635
R13717 VDD.n5357 VDD.t75 168.635
R13718 VDD.n5356 VDD.t826 168.635
R13719 VDD.n5356 VDD.t770 168.635
R13720 VDD.n5323 VDD.t95 168.635
R13721 VDD.n5323 VDD.t484 168.635
R13722 VDD.n5322 VDD.t483 168.635
R13723 VDD.n5322 VDD.t758 168.635
R13724 VDD.n5291 VDD.t419 168.635
R13725 VDD.n5291 VDD.t449 168.635
R13726 VDD.n5290 VDD.t309 168.635
R13727 VDD.n5290 VDD.t902 168.635
R13728 VDD.n5257 VDD.t782 168.635
R13729 VDD.n5257 VDD.t443 168.635
R13730 VDD.n5256 VDD.t444 168.635
R13731 VDD.n5256 VDD.t502 168.635
R13732 VDD.n5229 VDD.t877 168.635
R13733 VDD.n5229 VDD.t262 168.635
R13734 VDD.n5228 VDD.t394 168.635
R13735 VDD.n5228 VDD.t336 168.635
R13736 VDD.n5195 VDD.t488 168.635
R13737 VDD.n5195 VDD.t375 168.635
R13738 VDD.n5194 VDD.t344 168.635
R13739 VDD.n5194 VDD.t722 168.635
R13740 VDD.n5163 VDD.t578 168.635
R13741 VDD.n5163 VDD.t772 168.635
R13742 VDD.n5162 VDD.t426 168.635
R13743 VDD.n5162 VDD.t507 168.635
R13744 VDD.n5129 VDD.t223 168.635
R13745 VDD.n5129 VDD.t531 168.635
R13746 VDD.n5128 VDD.t530 168.635
R13747 VDD.n5128 VDD.t330 168.635
R13748 VDD.n5101 VDD.t558 168.635
R13749 VDD.n5101 VDD.t304 168.635
R13750 VDD.n5100 VDD.t617 168.635
R13751 VDD.n5100 VDD.t63 168.635
R13752 VDD.n5067 VDD.t629 168.635
R13753 VDD.n5067 VDD.t613 168.635
R13754 VDD.n5066 VDD.t612 168.635
R13755 VDD.n5066 VDD.t759 168.635
R13756 VDD.n170 VDD.t219 168.571
R13757 VDD.n170 VDD.t897 168.571
R13758 VDD.n351 VDD.t362 168.571
R13759 VDD.n351 VDD.t771 168.571
R13760 VDD.n312 VDD.t446 168.571
R13761 VDD.n312 VDD.t845 168.571
R13762 VDD.n385 VDD.t607 168.571
R13763 VDD.n385 VDD.t800 168.571
R13764 VDD.n386 VDD.t876 168.571
R13765 VDD.n386 VDD.t641 168.571
R13766 VDD.n311 VDD.t435 168.571
R13767 VDD.n311 VDD.t434 168.571
R13768 VDD.n350 VDD.t844 168.571
R13769 VDD.n350 VDD.t447 168.571
R13770 VDD.n278 VDD.t251 168.571
R13771 VDD.n278 VDD.t815 168.571
R13772 VDD.n418 VDD.t387 168.571
R13773 VDD.n418 VDD.t848 168.571
R13774 VDD.n599 VDD.t313 168.571
R13775 VDD.n599 VDD.t342 168.571
R13776 VDD.n560 VDD.t762 168.571
R13777 VDD.n560 VDD.t708 168.571
R13778 VDD.n633 VDD.t634 168.571
R13779 VDD.n633 VDD.t606 168.571
R13780 VDD.n634 VDD.t886 168.571
R13781 VDD.n634 VDD.t339 168.571
R13782 VDD.n559 VDD.t462 168.571
R13783 VDD.n559 VDD.t620 168.571
R13784 VDD.n598 VDD.t707 168.571
R13785 VDD.n598 VDD.t399 168.571
R13786 VDD.n526 VDD.t818 168.571
R13787 VDD.n526 VDD.t226 168.571
R13788 VDD.n677 VDD.t329 168.571
R13789 VDD.n677 VDD.t709 168.571
R13790 VDD.n858 VDD.t511 168.571
R13791 VDD.n858 VDD.t497 168.571
R13792 VDD.n819 VDD.t328 168.571
R13793 VDD.n819 VDD.t803 168.571
R13794 VDD.n892 VDD.t923 168.571
R13795 VDD.n892 VDD.t345 168.571
R13796 VDD.n893 VDD.t525 168.571
R13797 VDD.n893 VDD.t858 168.571
R13798 VDD.n818 VDD.t273 168.571
R13799 VDD.n818 VDD.t498 168.571
R13800 VDD.n857 VDD.t807 168.571
R13801 VDD.n857 VDD.t602 168.571
R13802 VDD.n785 VDD.t228 168.571
R13803 VDD.n785 VDD.t809 168.571
R13804 VDD.n936 VDD.t857 168.571
R13805 VDD.n936 VDD.t80 168.571
R13806 VDD.n1117 VDD.t603 168.571
R13807 VDD.n1117 VDD.t791 168.571
R13808 VDD.n1078 VDD.t381 168.571
R13809 VDD.n1078 VDD.t355 168.571
R13810 VDD.n1151 VDD.t67 168.571
R13811 VDD.n1151 VDD.t52 168.571
R13812 VDD.n1152 VDD.t50 168.571
R13813 VDD.n1152 VDD.t749 168.571
R13814 VDD.n1077 VDD.t13 168.571
R13815 VDD.n1077 VDD.t556 168.571
R13816 VDD.n1116 VDD.t354 168.571
R13817 VDD.n1116 VDD.t268 168.571
R13818 VDD.n1044 VDD.t832 168.571
R13819 VDD.n1044 VDD.t234 168.571
R13820 VDD.n1195 VDD.t263 168.571
R13821 VDD.n1195 VDD.t290 168.571
R13822 VDD.n1376 VDD.t798 168.571
R13823 VDD.n1376 VDD.t918 168.571
R13824 VDD.n1337 VDD.t320 168.571
R13825 VDD.n1337 VDD.t54 168.571
R13826 VDD.n1410 VDD.t310 168.571
R13827 VDD.n1410 VDD.t702 168.571
R13828 VDD.n1411 VDD.t266 168.571
R13829 VDD.n1411 VDD.t741 168.571
R13830 VDD.n1336 VDD.t516 168.571
R13831 VDD.n1336 VDD.t514 168.571
R13832 VDD.n1375 VDD.t841 168.571
R13833 VDD.n1375 VDD.t593 168.571
R13834 VDD.n1303 VDD.t810 168.571
R13835 VDD.n1303 VDD.t229 168.571
R13836 VDD.n1454 VDD.t793 168.571
R13837 VDD.n1454 VDD.t557 168.571
R13838 VDD.n1635 VDD.t906 168.571
R13839 VDD.n1635 VDD.t849 168.571
R13840 VDD.n1596 VDD.t473 168.571
R13841 VDD.n1596 VDD.t768 168.571
R13842 VDD.n1669 VDD.t398 168.571
R13843 VDD.n1669 VDD.t47 168.571
R13844 VDD.n1670 VDD.t835 168.571
R13845 VDD.n1670 VDD.t85 168.571
R13846 VDD.n1595 VDD.t750 168.571
R13847 VDD.n1595 VDD.t751 168.571
R13848 VDD.n1634 VDD.t769 168.571
R13849 VDD.n1634 VDD.t472 168.571
R13850 VDD.n1562 VDD.t243 168.571
R13851 VDD.n1562 VDD.t247 168.571
R13852 VDD.n1713 VDD.t23 168.571
R13853 VDD.n1713 VDD.t729 168.571
R13854 VDD.n1894 VDD.t921 168.571
R13855 VDD.n1894 VDD.t445 168.571
R13856 VDD.n1855 VDD.t311 168.571
R13857 VDD.n1855 VDD.t433 168.571
R13858 VDD.n1928 VDD.t491 168.571
R13859 VDD.n1928 VDD.t360 168.571
R13860 VDD.n1929 VDD.t907 168.571
R13861 VDD.n1929 VDD.t711 168.571
R13862 VDD.n1854 VDD.t591 168.571
R13863 VDD.n1854 VDD.t274 168.571
R13864 VDD.n1893 VDD.t417 168.571
R13865 VDD.n1893 VDD.t312 168.571
R13866 VDD.n1821 VDD.t230 168.571
R13867 VDD.n1821 VDD.t233 168.571
R13868 VDD.n1972 VDD.t367 168.571
R13869 VDD.n1972 VDD.t217 168.571
R13870 VDD.n2153 VDD.t582 168.571
R13871 VDD.n2153 VDD.t284 168.571
R13872 VDD.n2114 VDD.t515 168.571
R13873 VDD.n2114 VDD.t882 168.571
R13874 VDD.n2187 VDD.t522 168.571
R13875 VDD.n2187 VDD.t366 168.571
R13876 VDD.n2188 VDD.t533 168.571
R13877 VDD.n2188 VDD.t551 168.571
R13878 VDD.n2113 VDD.t264 168.571
R13879 VDD.n2113 VDD.t265 168.571
R13880 VDD.n2152 VDD.t786 168.571
R13881 VDD.n2152 VDD.t36 168.571
R13882 VDD.n2080 VDD.t321 168.571
R13883 VDD.n2080 VDD.t244 168.571
R13884 VDD.n2231 VDD.t909 168.571
R13885 VDD.n2231 VDD.t633 168.571
R13886 VDD.n2412 VDD.t920 168.571
R13887 VDD.n2412 VDD.t616 168.571
R13888 VDD.n2373 VDD.t334 168.571
R13889 VDD.n2373 VDD.t867 168.571
R13890 VDD.n2446 VDD.t785 168.571
R13891 VDD.n2446 VDD.t404 168.571
R13892 VDD.n2447 VDD.t363 168.571
R13893 VDD.n2447 VDD.t787 168.571
R13894 VDD.n2372 VDD.t218 168.571
R13895 VDD.n2372 VDD.t30 168.571
R13896 VDD.n2411 VDD.t868 168.571
R13897 VDD.n2411 VDD.t723 168.571
R13898 VDD.n2339 VDD.t817 168.571
R13899 VDD.n2339 VDD.t322 168.571
R13900 VDD.n2490 VDD.t351 168.571
R13901 VDD.n2490 VDD.t84 168.571
R13902 VDD.n2671 VDD.t806 168.571
R13903 VDD.n2671 VDD.t600 168.571
R13904 VDD.n2632 VDD.t414 168.571
R13905 VDD.n2632 VDD.t393 168.571
R13906 VDD.n2705 VDD.t410 168.571
R13907 VDD.n2705 VDD.t575 168.571
R13908 VDD.n2706 VDD.t73 168.571
R13909 VDD.n2706 VDD.t436 168.571
R13910 VDD.n2631 VDD.t917 168.571
R13911 VDD.n2631 VDD.t489 168.571
R13912 VDD.n2670 VDD.t919 168.571
R13913 VDD.n2670 VDD.t513 168.571
R13914 VDD.n2598 VDD.t231 168.571
R13915 VDD.n2598 VDD.t323 168.571
R13916 VDD.n2749 VDD.t58 168.571
R13917 VDD.n2749 VDD.t490 168.571
R13918 VDD.n2930 VDD.t512 168.571
R13919 VDD.n2930 VDD.t279 168.571
R13920 VDD.n2891 VDD.t374 168.571
R13921 VDD.n2891 VDD.t851 168.571
R13922 VDD.n2964 VDD.t587 168.571
R13923 VDD.n2964 VDD.t11 168.571
R13924 VDD.n2965 VDD.t706 168.571
R13925 VDD.n2965 VDD.t588 168.571
R13926 VDD.n2890 VDD.t621 168.571
R13927 VDD.n2890 VDD.t622 168.571
R13928 VDD.n2929 VDD.t852 168.571
R13929 VDD.n2929 VDD.t337 168.571
R13930 VDD.n2857 VDD.t250 168.571
R13931 VDD.n2857 VDD.t232 168.571
R13932 VDD.n3008 VDD.t589 168.571
R13933 VDD.n3008 VDD.t56 168.571
R13934 VDD.n3189 VDD.t872 168.571
R13935 VDD.n3189 VDD.t373 168.571
R13936 VDD.n3150 VDD.t623 168.571
R13937 VDD.n3150 VDD.t781 168.571
R13938 VDD.n3223 VDD.t49 168.571
R13939 VDD.n3223 VDD.t519 168.571
R13940 VDD.n3224 VDD.t305 168.571
R13941 VDD.n3224 VDD.t406 168.571
R13942 VDD.n3149 VDD.t734 168.571
R13943 VDD.n3149 VDD.t908 168.571
R13944 VDD.n3188 VDD.t780 168.571
R13945 VDD.n3188 VDD.t624 168.571
R13946 VDD.n3116 VDD.t821 168.571
R13947 VDD.n3116 VDD.t743 168.571
R13948 VDD.n3267 VDD.t405 168.571
R13949 VDD.n3267 VDD.t874 168.571
R13950 VDD.n3448 VDD.t608 168.571
R13951 VDD.n3448 VDD.t850 168.571
R13952 VDD.n3409 VDD.t464 168.571
R13953 VDD.n3409 VDD.t860 168.571
R13954 VDD.n3482 VDD.t267 168.571
R13955 VDD.n3482 VDD.t632 168.571
R13956 VDD.n3483 VDD.t500 168.571
R13957 VDD.n3483 VDD.t93 168.571
R13958 VDD.n3408 VDD.t520 168.571
R13959 VDD.n3408 VDD.t521 168.571
R13960 VDD.n3447 VDD.t861 168.571
R13961 VDD.n3447 VDD.t463 168.571
R13962 VDD.n3375 VDD.t245 168.571
R13963 VDD.n3375 VDD.t227 168.571
R13964 VDD.n3526 VDD.t480 168.571
R13965 VDD.n3526 VDD.t801 168.571
R13966 VDD.n3707 VDD.t581 168.571
R13967 VDD.n3707 VDD.t331 168.571
R13968 VDD.n3668 VDD.t592 168.571
R13969 VDD.n3668 VDD.t33 168.571
R13970 VDD.n3741 VDD.t724 168.571
R13971 VDD.n3741 VDD.t727 168.571
R13972 VDD.n3742 VDD.t555 168.571
R13973 VDD.n3742 VDD.t380 168.571
R13974 VDD.n3667 VDD.t25 168.571
R13975 VDD.n3667 VDD.t26 168.571
R13976 VDD.n3706 VDD.t34 168.571
R13977 VDD.n3706 VDD.t15 168.571
R13978 VDD.n3634 VDD.t324 168.571
R13979 VDD.n3634 VDD.t246 168.571
R13980 VDD.n3785 VDD.t887 168.571
R13981 VDD.n3785 VDD.t272 168.571
R13982 VDD.n3966 VDD.t777 168.571
R13983 VDD.n3966 VDD.t730 168.571
R13984 VDD.n3927 VDD.t825 168.571
R13985 VDD.n3927 VDD.t779 168.571
R13986 VDD.n4000 VDD.t609 168.571
R13987 VDD.n4000 VDD.t834 168.571
R13988 VDD.n4001 VDD.t865 168.571
R13989 VDD.n4001 VDD.t271 168.571
R13990 VDD.n3926 VDD.t517 168.571
R13991 VDD.n3926 VDD.t518 168.571
R13992 VDD.n3965 VDD.t778 168.571
R13993 VDD.n3965 VDD.t814 168.571
R13994 VDD.n3893 VDD.t833 168.571
R13995 VDD.n3893 VDD.t816 168.571
R13996 VDD.n4044 VDD.t912 168.571
R13997 VDD.n4044 VDD.t319 168.571
R13998 VDD.n4225 VDD.t580 168.571
R13999 VDD.n4225 VDD.t378 168.571
R14000 VDD.n4186 VDD.t783 168.571
R14001 VDD.n4186 VDD.t416 168.571
R14002 VDD.n4259 VDD.t799 168.571
R14003 VDD.n4259 VDD.t481 168.571
R14004 VDD.n4260 VDD.t601 168.571
R14005 VDD.n4260 VDD.t471 168.571
R14006 VDD.n4185 VDD.t9 168.571
R14007 VDD.n4185 VDD.t7 168.571
R14008 VDD.n4224 VDD.t415 168.571
R14009 VDD.n4224 VDD.t221 168.571
R14010 VDD.n4152 VDD.t242 168.571
R14011 VDD.n4152 VDD.t239 168.571
R14012 VDD.n4303 VDD.t467 168.571
R14013 VDD.n4303 VDD.t437 168.571
R14014 VDD.n4484 VDD.t77 168.571
R14015 VDD.n4484 VDD.t346 168.571
R14016 VDD.n4445 VDD.t260 168.571
R14017 VDD.n4445 VDD.t761 168.571
R14018 VDD.n4518 VDD.t413 168.571
R14019 VDD.n4518 VDD.t846 168.571
R14020 VDD.n4519 VDD.t871 168.571
R14021 VDD.n4519 VDD.t808 168.571
R14022 VDD.n4444 VDD.t379 168.571
R14023 VDD.n4444 VDD.t579 168.571
R14024 VDD.n4483 VDD.t742 168.571
R14025 VDD.n4483 VDD.t259 168.571
R14026 VDD.n4411 VDD.t254 168.571
R14027 VDD.n4411 VDD.t236 168.571
R14028 VDD.n398 VDD.t102 168.148
R14029 VDD.n398 VDD.t690 168.148
R14030 VDD.n191 VDD.t220 168.148
R14031 VDD.n295 VDD.t191 168.148
R14032 VDD.n295 VDD.t699 168.148
R14033 VDD.n334 VDD.t248 168.148
R14034 VDD.n294 VDD.t197 168.148
R14035 VDD.n294 VDD.t654 168.148
R14036 VDD.n646 VDD.t662 168.148
R14037 VDD.n646 VDD.t211 168.148
R14038 VDD.n439 VDD.t642 168.148
R14039 VDD.n543 VDD.t694 168.148
R14040 VDD.n543 VDD.t107 168.148
R14041 VDD.n582 VDD.t235 168.148
R14042 VDD.n542 VDD.t651 168.148
R14043 VDD.n542 VDD.t145 168.148
R14044 VDD.n905 VDD.t653 168.148
R14045 VDD.n905 VDD.t124 168.148
R14046 VDD.n698 VDD.t338 168.148
R14047 VDD.n802 VDD.t650 168.148
R14048 VDD.n802 VDD.t208 168.148
R14049 VDD.n841 VDD.t746 168.148
R14050 VDD.n801 VDD.t667 168.148
R14051 VDD.n801 VDD.t127 168.148
R14052 VDD.n1164 VDD.t684 168.148
R14053 VDD.n1164 VDD.t202 168.148
R14054 VDD.n957 VDD.t859 168.148
R14055 VDD.n1061 VDD.t689 168.148
R14056 VDD.n1061 VDD.t178 168.148
R14057 VDD.n1100 VDD.t824 168.148
R14058 VDD.n1060 VDD.t698 168.148
R14059 VDD.n1060 VDD.t186 168.148
R14060 VDD.n1423 VDD.t657 168.148
R14061 VDD.n1423 VDD.t112 168.148
R14062 VDD.n1216 VDD.t370 168.148
R14063 VDD.n1320 VDD.t700 168.148
R14064 VDD.n1320 VDD.t99 168.148
R14065 VDD.n1359 VDD.t238 168.148
R14066 VDD.n1319 VDD.t659 168.148
R14067 VDD.n1319 VDD.t133 168.148
R14068 VDD.n1682 VDD.t663 168.148
R14069 VDD.n1682 VDD.t148 168.148
R14070 VDD.n1475 VDD.t740 168.148
R14071 VDD.n1579 VDD.t658 168.148
R14072 VDD.n1579 VDD.t109 168.148
R14073 VDD.n1618 VDD.t295 168.148
R14074 VDD.n1578 VDD.t674 168.148
R14075 VDD.n1578 VDD.t150 168.148
R14076 VDD.n1941 VDD.t675 168.148
R14077 VDD.n1941 VDD.t121 168.148
R14078 VDD.n1734 VDD.t86 168.148
R14079 VDD.n1838 VDD.t647 168.148
R14080 VDD.n1838 VDD.t141 168.148
R14081 VDD.n1877 VDD.t256 168.148
R14082 VDD.n1837 VDD.t665 168.148
R14083 VDD.n1837 VDD.t167 168.148
R14084 VDD.n2200 VDD.t668 168.148
R14085 VDD.n2200 VDD.t157 168.148
R14086 VDD.n1993 VDD.t710 168.148
R14087 VDD.n2097 VDD.t664 168.148
R14088 VDD.n2097 VDD.t119 168.148
R14089 VDD.n2136 VDD.t291 168.148
R14090 VDD.n2096 VDD.t678 168.148
R14091 VDD.n2096 VDD.t159 168.148
R14092 VDD.n2459 VDD.t671 168.148
R14093 VDD.n2459 VDD.t214 168.148
R14094 VDD.n2252 VDD.t552 168.148
R14095 VDD.n2356 VDD.t696 168.148
R14096 VDD.n2356 VDD.t131 168.148
R14097 VDD.n2395 VDD.t240 168.148
R14098 VDD.n2355 VDD.t652 168.148
R14099 VDD.n2355 VDD.t165 168.148
R14100 VDD.n2718 VDD.t672 168.148
R14101 VDD.n2718 VDD.t161 168.148
R14102 VDD.n2511 VDD.t456 168.148
R14103 VDD.n2615 VDD.t669 168.148
R14104 VDD.n2615 VDD.t129 168.148
R14105 VDD.n2654 VDD.t241 168.148
R14106 VDD.n2614 VDD.t679 168.148
R14107 VDD.n2614 VDD.t163 168.148
R14108 VDD.n2977 VDD.t677 168.148
R14109 VDD.n2977 VDD.t171 168.148
R14110 VDD.n2770 VDD.t61 168.148
R14111 VDD.n2874 VDD.t673 168.148
R14112 VDD.n2874 VDD.t143 168.148
R14113 VDD.n2913 VDD.t255 168.148
R14114 VDD.n2873 VDD.t680 168.148
R14115 VDD.n2873 VDD.t173 168.148
R14116 VDD.n3236 VDD.t681 168.148
R14117 VDD.n3236 VDD.t206 168.148
R14118 VDD.n3029 VDD.t492 168.148
R14119 VDD.n3133 VDD.t693 168.148
R14120 VDD.n3133 VDD.t169 168.148
R14121 VDD.n3172 VDD.t831 168.148
R14122 VDD.n3132 VDD.t648 168.148
R14123 VDD.n3132 VDD.t180 168.148
R14124 VDD.n3495 VDD.t660 168.148
R14125 VDD.n3495 VDD.t136 168.148
R14126 VDD.n3288 VDD.t802 168.148
R14127 VDD.n3392 VDD.t655 168.148
R14128 VDD.n3392 VDD.t104 168.148
R14129 VDD.n3431 VDD.t237 168.148
R14130 VDD.n3391 VDD.t670 168.148
R14131 VDD.n3391 VDD.t138 168.148
R14132 VDD.n3754 VDD.t666 168.148
R14133 VDD.n3754 VDD.t152 168.148
R14134 VDD.n3547 VDD.t89 168.148
R14135 VDD.n3651 VDD.t661 168.148
R14136 VDD.n3651 VDD.t114 168.148
R14137 VDD.n3690 VDD.t294 168.148
R14138 VDD.n3650 VDD.t676 168.148
R14139 VDD.n3650 VDD.t154 168.148
R14140 VDD.n4013 VDD.t649 168.148
R14141 VDD.n4013 VDD.t200 168.148
R14142 VDD.n3806 VDD.t890 168.148
R14143 VDD.n3910 VDD.t688 168.148
R14144 VDD.n3910 VDD.t204 168.148
R14145 VDD.n3949 VDD.t249 168.148
R14146 VDD.n3909 VDD.t695 168.148
R14147 VDD.n3909 VDD.t117 168.148
R14148 VDD.n4272 VDD.t686 168.148
R14149 VDD.n4272 VDD.t188 168.148
R14150 VDD.n4065 VDD.t407 168.148
R14151 VDD.n4169 VDD.t682 168.148
R14152 VDD.n4169 VDD.t182 168.148
R14153 VDD.n4208 VDD.t811 168.148
R14154 VDD.n4168 VDD.t687 168.148
R14155 VDD.n4168 VDD.t195 168.148
R14156 VDD.n4531 VDD.t683 168.148
R14157 VDD.n4531 VDD.t193 168.148
R14158 VDD.n4324 VDD.t470 168.148
R14159 VDD.n4428 VDD.t685 168.148
R14160 VDD.n4428 VDD.t176 168.148
R14161 VDD.n4467 VDD.t830 168.148
R14162 VDD.n4427 VDD.t691 168.148
R14163 VDD.n4427 VDD.t184 168.148
R14164 VDD.n401 VDD.n189 166.238
R14165 VDD.n401 VDD.n190 166.238
R14166 VDD.n332 VDD.n331 166.238
R14167 VDD.n332 VDD.n327 166.238
R14168 VDD.n649 VDD.n437 166.238
R14169 VDD.n649 VDD.n438 166.238
R14170 VDD.n580 VDD.n579 166.238
R14171 VDD.n580 VDD.n575 166.238
R14172 VDD.n908 VDD.n696 166.238
R14173 VDD.n908 VDD.n697 166.238
R14174 VDD.n839 VDD.n838 166.238
R14175 VDD.n839 VDD.n834 166.238
R14176 VDD.n1167 VDD.n955 166.238
R14177 VDD.n1167 VDD.n956 166.238
R14178 VDD.n1098 VDD.n1097 166.238
R14179 VDD.n1098 VDD.n1093 166.238
R14180 VDD.n1426 VDD.n1214 166.238
R14181 VDD.n1426 VDD.n1215 166.238
R14182 VDD.n1357 VDD.n1356 166.238
R14183 VDD.n1357 VDD.n1352 166.238
R14184 VDD.n1685 VDD.n1473 166.238
R14185 VDD.n1685 VDD.n1474 166.238
R14186 VDD.n1616 VDD.n1615 166.238
R14187 VDD.n1616 VDD.n1611 166.238
R14188 VDD.n1944 VDD.n1732 166.238
R14189 VDD.n1944 VDD.n1733 166.238
R14190 VDD.n1875 VDD.n1874 166.238
R14191 VDD.n1875 VDD.n1870 166.238
R14192 VDD.n2203 VDD.n1991 166.238
R14193 VDD.n2203 VDD.n1992 166.238
R14194 VDD.n2134 VDD.n2133 166.238
R14195 VDD.n2134 VDD.n2129 166.238
R14196 VDD.n2462 VDD.n2250 166.238
R14197 VDD.n2462 VDD.n2251 166.238
R14198 VDD.n2393 VDD.n2392 166.238
R14199 VDD.n2393 VDD.n2388 166.238
R14200 VDD.n2721 VDD.n2509 166.238
R14201 VDD.n2721 VDD.n2510 166.238
R14202 VDD.n2652 VDD.n2651 166.238
R14203 VDD.n2652 VDD.n2647 166.238
R14204 VDD.n2980 VDD.n2768 166.238
R14205 VDD.n2980 VDD.n2769 166.238
R14206 VDD.n2911 VDD.n2910 166.238
R14207 VDD.n2911 VDD.n2906 166.238
R14208 VDD.n3239 VDD.n3027 166.238
R14209 VDD.n3239 VDD.n3028 166.238
R14210 VDD.n3170 VDD.n3169 166.238
R14211 VDD.n3170 VDD.n3165 166.238
R14212 VDD.n3498 VDD.n3286 166.238
R14213 VDD.n3498 VDD.n3287 166.238
R14214 VDD.n3429 VDD.n3428 166.238
R14215 VDD.n3429 VDD.n3424 166.238
R14216 VDD.n3757 VDD.n3545 166.238
R14217 VDD.n3757 VDD.n3546 166.238
R14218 VDD.n3688 VDD.n3687 166.238
R14219 VDD.n3688 VDD.n3683 166.238
R14220 VDD.n4016 VDD.n3804 166.238
R14221 VDD.n4016 VDD.n3805 166.238
R14222 VDD.n3947 VDD.n3946 166.238
R14223 VDD.n3947 VDD.n3942 166.238
R14224 VDD.n4275 VDD.n4063 166.238
R14225 VDD.n4275 VDD.n4064 166.238
R14226 VDD.n4206 VDD.n4205 166.238
R14227 VDD.n4206 VDD.n4201 166.238
R14228 VDD.n4534 VDD.n4322 166.238
R14229 VDD.n4534 VDD.n4323 166.238
R14230 VDD.n4465 VDD.n4464 166.238
R14231 VDD.n4465 VDD.n4460 166.238
R14232 VDD.n5032 VDD.n4558 166.238
R14233 VDD.n5032 VDD.n4557 166.238
R14234 VDD.n5024 VDD.n4563 166.238
R14235 VDD.n5022 VDD.n4563 166.238
R14236 VDD.n5017 VDD.n5012 166.238
R14237 VDD.n5015 VDD.n5012 166.238
R14238 VDD.n5007 VDD.n4569 166.238
R14239 VDD.n5007 VDD.n4568 166.238
R14240 VDD.n4999 VDD.n4994 166.238
R14241 VDD.n4997 VDD.n4994 166.238
R14242 VDD.n4991 VDD.n4577 166.238
R14243 VDD.n4991 VDD.n4576 166.238
R14244 VDD.n4983 VDD.n4582 166.238
R14245 VDD.n4981 VDD.n4582 166.238
R14246 VDD.n4976 VDD.n4971 166.238
R14247 VDD.n4974 VDD.n4971 166.238
R14248 VDD.n4966 VDD.n4588 166.238
R14249 VDD.n4966 VDD.n4587 166.238
R14250 VDD.n4958 VDD.n4953 166.238
R14251 VDD.n4956 VDD.n4953 166.238
R14252 VDD.n4950 VDD.n4596 166.238
R14253 VDD.n4950 VDD.n4595 166.238
R14254 VDD.n4942 VDD.n4601 166.238
R14255 VDD.n4940 VDD.n4601 166.238
R14256 VDD.n4935 VDD.n4930 166.238
R14257 VDD.n4933 VDD.n4930 166.238
R14258 VDD.n4925 VDD.n4607 166.238
R14259 VDD.n4925 VDD.n4606 166.238
R14260 VDD.n4917 VDD.n4912 166.238
R14261 VDD.n4915 VDD.n4912 166.238
R14262 VDD.n4909 VDD.n4615 166.238
R14263 VDD.n4909 VDD.n4614 166.238
R14264 VDD.n4901 VDD.n4620 166.238
R14265 VDD.n4899 VDD.n4620 166.238
R14266 VDD.n4894 VDD.n4889 166.238
R14267 VDD.n4892 VDD.n4889 166.238
R14268 VDD.n4884 VDD.n4626 166.238
R14269 VDD.n4884 VDD.n4625 166.238
R14270 VDD.n4876 VDD.n4871 166.238
R14271 VDD.n4874 VDD.n4871 166.238
R14272 VDD.n4868 VDD.n4634 166.238
R14273 VDD.n4868 VDD.n4633 166.238
R14274 VDD.n4860 VDD.n4639 166.238
R14275 VDD.n4858 VDD.n4639 166.238
R14276 VDD.n4853 VDD.n4848 166.238
R14277 VDD.n4851 VDD.n4848 166.238
R14278 VDD.n4843 VDD.n4645 166.238
R14279 VDD.n4843 VDD.n4644 166.238
R14280 VDD.n4835 VDD.n4830 166.238
R14281 VDD.n4833 VDD.n4830 166.238
R14282 VDD.n4827 VDD.n4653 166.238
R14283 VDD.n4827 VDD.n4652 166.238
R14284 VDD.n4819 VDD.n4658 166.238
R14285 VDD.n4817 VDD.n4658 166.238
R14286 VDD.n4812 VDD.n4807 166.238
R14287 VDD.n4810 VDD.n4807 166.238
R14288 VDD.n4802 VDD.n4664 166.238
R14289 VDD.n4802 VDD.n4663 166.238
R14290 VDD.n4794 VDD.n4789 166.238
R14291 VDD.n4792 VDD.n4789 166.238
R14292 VDD.n4786 VDD.n4672 166.238
R14293 VDD.n4786 VDD.n4671 166.238
R14294 VDD.n4778 VDD.n4677 166.238
R14295 VDD.n4776 VDD.n4677 166.238
R14296 VDD.n4771 VDD.n4766 166.238
R14297 VDD.n4769 VDD.n4766 166.238
R14298 VDD.n4761 VDD.n4683 166.238
R14299 VDD.n4761 VDD.n4682 166.238
R14300 VDD.n4753 VDD.n4748 166.238
R14301 VDD.n4751 VDD.n4748 166.238
R14302 VDD.n4745 VDD.n4691 166.238
R14303 VDD.n4745 VDD.n4690 166.238
R14304 VDD.n4737 VDD.n4696 166.238
R14305 VDD.n4735 VDD.n4696 166.238
R14306 VDD.n4730 VDD.n4725 166.238
R14307 VDD.n4728 VDD.n4725 166.238
R14308 VDD.n4720 VDD.n4702 166.238
R14309 VDD.n4720 VDD.n4701 166.238
R14310 VDD.n4712 VDD.n4707 166.238
R14311 VDD.n4710 VDD.n4707 166.238
R14312 VDD.n7103 VDD.n7102 166.238
R14313 VDD.n7103 VDD.n5035 166.238
R14314 VDD.n6978 VDD.n6977 166.238
R14315 VDD.n6977 VDD.n5172 166.238
R14316 VDD.n6847 VDD.n6846 166.238
R14317 VDD.n6846 VDD.n5300 166.238
R14318 VDD.n6716 VDD.n6715 166.238
R14319 VDD.n6715 VDD.n5428 166.238
R14320 VDD.n6585 VDD.n6584 166.238
R14321 VDD.n6584 VDD.n5556 166.238
R14322 VDD.n6454 VDD.n6453 166.238
R14323 VDD.n6453 VDD.n5684 166.238
R14324 VDD.n6323 VDD.n6322 166.238
R14325 VDD.n6322 VDD.n5812 166.238
R14326 VDD.n6192 VDD.n6191 166.238
R14327 VDD.n6191 VDD.n5940 166.238
R14328 VDD.n7035 VDD.n5109 166.238
R14329 VDD.n7033 VDD.n5109 166.238
R14330 VDD.n6904 VDD.n5237 166.238
R14331 VDD.n6902 VDD.n5237 166.238
R14332 VDD.n6773 VDD.n5365 166.238
R14333 VDD.n6771 VDD.n5365 166.238
R14334 VDD.n6642 VDD.n5493 166.238
R14335 VDD.n6640 VDD.n5493 166.238
R14336 VDD.n6511 VDD.n5621 166.238
R14337 VDD.n6509 VDD.n5621 166.238
R14338 VDD.n6380 VDD.n5749 166.238
R14339 VDD.n6378 VDD.n5749 166.238
R14340 VDD.n6249 VDD.n5877 166.238
R14341 VDD.n6247 VDD.n5877 166.238
R14342 VDD.n6118 VDD.n6005 166.238
R14343 VDD.n6116 VDD.n6005 166.238
R14344 VDD.n7111 VDD.n7108 166.238
R14345 VDD.n7113 VDD.n7108 166.238
R14346 VDD.n7118 VDD.n143 166.238
R14347 VDD.n7120 VDD.n143 166.238
R14348 VDD.n7126 VDD.n7125 166.238
R14349 VDD.n7126 VDD.n135 166.238
R14350 VDD.n7132 VDD.n7129 166.238
R14351 VDD.n7134 VDD.n7129 166.238
R14352 VDD.n7139 VDD.n124 166.238
R14353 VDD.n7141 VDD.n124 166.238
R14354 VDD.n7147 VDD.n7146 166.238
R14355 VDD.n7147 VDD.n116 166.238
R14356 VDD.n7153 VDD.n7150 166.238
R14357 VDD.n7155 VDD.n7150 166.238
R14358 VDD.n7160 VDD.n105 166.238
R14359 VDD.n7162 VDD.n105 166.238
R14360 VDD.n7168 VDD.n7167 166.238
R14361 VDD.n7168 VDD.n97 166.238
R14362 VDD.n7174 VDD.n7171 166.238
R14363 VDD.n7176 VDD.n7171 166.238
R14364 VDD.n7181 VDD.n86 166.238
R14365 VDD.n7183 VDD.n86 166.238
R14366 VDD.n7189 VDD.n7188 166.238
R14367 VDD.n7189 VDD.n78 166.238
R14368 VDD.n7195 VDD.n7192 166.238
R14369 VDD.n7197 VDD.n7192 166.238
R14370 VDD.n7202 VDD.n67 166.238
R14371 VDD.n7204 VDD.n67 166.238
R14372 VDD.n7210 VDD.n7209 166.238
R14373 VDD.n7210 VDD.n59 166.238
R14374 VDD.n7216 VDD.n7213 166.238
R14375 VDD.n7218 VDD.n7213 166.238
R14376 VDD.n7223 VDD.n48 166.238
R14377 VDD.n7225 VDD.n48 166.238
R14378 VDD.n7231 VDD.n7230 166.238
R14379 VDD.n7231 VDD.n40 166.238
R14380 VDD.n7237 VDD.n7234 166.238
R14381 VDD.n7239 VDD.n7234 166.238
R14382 VDD.n7244 VDD.n29 166.238
R14383 VDD.n7246 VDD.n29 166.238
R14384 VDD.n7252 VDD.n7251 166.238
R14385 VDD.n7252 VDD.n21 166.238
R14386 VDD.n7258 VDD.n7255 166.238
R14387 VDD.n7260 VDD.n7255 166.238
R14388 VDD.n7265 VDD.n10 166.238
R14389 VDD.n7267 VDD.n10 166.238
R14390 VDD.n7273 VDD.n7272 166.238
R14391 VDD.n7273 VDD.n2 166.238
R14392 VDD.n673 VDD.t122 158.965
R14393 VDD.n932 VDD.t201 158.965
R14394 VDD.n1191 VDD.t110 158.965
R14395 VDD.n1450 VDD.t146 158.965
R14396 VDD.n1709 VDD.t120 158.965
R14397 VDD.n1968 VDD.t155 158.965
R14398 VDD.n2227 VDD.t212 158.965
R14399 VDD.n2486 VDD.t160 158.965
R14400 VDD.n2745 VDD.t170 158.965
R14401 VDD.n3004 VDD.t205 158.965
R14402 VDD.n3263 VDD.t134 158.965
R14403 VDD.n3522 VDD.t151 158.965
R14404 VDD.n3781 VDD.t198 158.965
R14405 VDD.n4040 VDD.t187 158.965
R14406 VDD.n4299 VDD.t192 158.965
R14407 VDD.n5027 VDD.n5026 155.102
R14408 VDD.n5002 VDD.n5001 155.102
R14409 VDD.n4986 VDD.n4985 155.102
R14410 VDD.n4961 VDD.n4960 155.102
R14411 VDD.n4945 VDD.n4944 155.102
R14412 VDD.n4920 VDD.n4919 155.102
R14413 VDD.n4904 VDD.n4903 155.102
R14414 VDD.n4879 VDD.n4878 155.102
R14415 VDD.n4863 VDD.n4862 155.102
R14416 VDD.n4838 VDD.n4837 155.102
R14417 VDD.n4822 VDD.n4821 155.102
R14418 VDD.n4797 VDD.n4796 155.102
R14419 VDD.n4781 VDD.n4780 155.102
R14420 VDD.n4756 VDD.n4755 155.102
R14421 VDD.n4740 VDD.n4739 155.102
R14422 VDD.n4715 VDD.n4714 155.102
R14423 VDD.n7123 VDD.n7122 155.102
R14424 VDD.n7116 VDD.n7115 155.102
R14425 VDD.n7144 VDD.n7143 155.102
R14426 VDD.n7137 VDD.n7136 155.102
R14427 VDD.n7165 VDD.n7164 155.102
R14428 VDD.n7158 VDD.n7157 155.102
R14429 VDD.n7186 VDD.n7185 155.102
R14430 VDD.n7179 VDD.n7178 155.102
R14431 VDD.n7207 VDD.n7206 155.102
R14432 VDD.n7200 VDD.n7199 155.102
R14433 VDD.n7228 VDD.n7227 155.102
R14434 VDD.n7221 VDD.n7220 155.102
R14435 VDD.n7249 VDD.n7248 155.102
R14436 VDD.n7242 VDD.n7241 155.102
R14437 VDD.n7270 VDD.n7269 155.102
R14438 VDD.n7263 VDD.n7262 155.102
R14439 VDD.n413 VDD.t100 154.846
R14440 VDD.n414 VDD.t209 154.846
R14441 VDD.n198 VDD.n193 153.601
R14442 VDD.n196 VDD.n192 153.601
R14443 VDD.n241 VDD.n192 153.601
R14444 VDD.n242 VDD.n193 153.601
R14445 VDD.n220 VDD.n173 153.601
R14446 VDD.n219 VDD.n171 153.601
R14447 VDD.n372 VDD.n171 153.601
R14448 VDD.n373 VDD.n173 153.601
R14449 VDD.n290 VDD.n284 153.601
R14450 VDD.n281 VDD.n279 153.601
R14451 VDD.n286 VDD.n279 153.601
R14452 VDD.n290 VDD.n289 153.601
R14453 VDD.n368 VDD.n272 153.601
R14454 VDD.n276 VDD.n275 153.601
R14455 VDD.n276 VDD.n271 153.601
R14456 VDD.n369 VDD.n368 153.601
R14457 VDD.n363 VDD.n357 153.601
R14458 VDD.n354 VDD.n352 153.601
R14459 VDD.n359 VDD.n352 153.601
R14460 VDD.n363 VDD.n362 153.601
R14461 VDD.n347 VDD.n341 153.601
R14462 VDD.n338 VDD.n336 153.601
R14463 VDD.n343 VDD.n336 153.601
R14464 VDD.n347 VDD.n346 153.601
R14465 VDD.n324 VDD.n318 153.601
R14466 VDD.n315 VDD.n313 153.601
R14467 VDD.n320 VDD.n313 153.601
R14468 VDD.n324 VDD.n323 153.601
R14469 VDD.n308 VDD.n302 153.601
R14470 VDD.n299 VDD.n297 153.601
R14471 VDD.n304 VDD.n297 153.601
R14472 VDD.n308 VDD.n307 153.601
R14473 VDD.n258 VDD.n251 153.601
R14474 VDD.n255 VDD.n254 153.601
R14475 VDD.n255 VDD.n250 153.601
R14476 VDD.n259 VDD.n258 153.601
R14477 VDD.n382 VDD.n235 153.601
R14478 VDD.n232 VDD.n230 153.601
R14479 VDD.n237 VDD.n230 153.601
R14480 VDD.n382 VDD.n381 153.601
R14481 VDD.n264 VDD.n227 153.601
R14482 VDD.n389 VDD.n228 153.601
R14483 VDD.n392 VDD.n227 153.601
R14484 VDD.n390 VDD.n389 153.601
R14485 VDD.n446 VDD.n441 153.601
R14486 VDD.n444 VDD.n440 153.601
R14487 VDD.n489 VDD.n440 153.601
R14488 VDD.n490 VDD.n441 153.601
R14489 VDD.n468 VDD.n421 153.601
R14490 VDD.n467 VDD.n419 153.601
R14491 VDD.n620 VDD.n419 153.601
R14492 VDD.n621 VDD.n421 153.601
R14493 VDD.n538 VDD.n532 153.601
R14494 VDD.n529 VDD.n527 153.601
R14495 VDD.n534 VDD.n527 153.601
R14496 VDD.n538 VDD.n537 153.601
R14497 VDD.n616 VDD.n520 153.601
R14498 VDD.n524 VDD.n523 153.601
R14499 VDD.n524 VDD.n519 153.601
R14500 VDD.n617 VDD.n616 153.601
R14501 VDD.n611 VDD.n605 153.601
R14502 VDD.n602 VDD.n600 153.601
R14503 VDD.n607 VDD.n600 153.601
R14504 VDD.n611 VDD.n610 153.601
R14505 VDD.n595 VDD.n589 153.601
R14506 VDD.n586 VDD.n584 153.601
R14507 VDD.n591 VDD.n584 153.601
R14508 VDD.n595 VDD.n594 153.601
R14509 VDD.n572 VDD.n566 153.601
R14510 VDD.n563 VDD.n561 153.601
R14511 VDD.n568 VDD.n561 153.601
R14512 VDD.n572 VDD.n571 153.601
R14513 VDD.n556 VDD.n550 153.601
R14514 VDD.n547 VDD.n545 153.601
R14515 VDD.n552 VDD.n545 153.601
R14516 VDD.n556 VDD.n555 153.601
R14517 VDD.n506 VDD.n499 153.601
R14518 VDD.n503 VDD.n502 153.601
R14519 VDD.n503 VDD.n498 153.601
R14520 VDD.n507 VDD.n506 153.601
R14521 VDD.n630 VDD.n483 153.601
R14522 VDD.n480 VDD.n478 153.601
R14523 VDD.n485 VDD.n478 153.601
R14524 VDD.n630 VDD.n629 153.601
R14525 VDD.n512 VDD.n475 153.601
R14526 VDD.n637 VDD.n476 153.601
R14527 VDD.n640 VDD.n475 153.601
R14528 VDD.n638 VDD.n637 153.601
R14529 VDD.n705 VDD.n700 153.601
R14530 VDD.n703 VDD.n699 153.601
R14531 VDD.n748 VDD.n699 153.601
R14532 VDD.n749 VDD.n700 153.601
R14533 VDD.n727 VDD.n680 153.601
R14534 VDD.n726 VDD.n678 153.601
R14535 VDD.n879 VDD.n678 153.601
R14536 VDD.n880 VDD.n680 153.601
R14537 VDD.n797 VDD.n791 153.601
R14538 VDD.n788 VDD.n786 153.601
R14539 VDD.n793 VDD.n786 153.601
R14540 VDD.n797 VDD.n796 153.601
R14541 VDD.n875 VDD.n779 153.601
R14542 VDD.n783 VDD.n782 153.601
R14543 VDD.n783 VDD.n778 153.601
R14544 VDD.n876 VDD.n875 153.601
R14545 VDD.n870 VDD.n864 153.601
R14546 VDD.n861 VDD.n859 153.601
R14547 VDD.n866 VDD.n859 153.601
R14548 VDD.n870 VDD.n869 153.601
R14549 VDD.n854 VDD.n848 153.601
R14550 VDD.n845 VDD.n843 153.601
R14551 VDD.n850 VDD.n843 153.601
R14552 VDD.n854 VDD.n853 153.601
R14553 VDD.n831 VDD.n825 153.601
R14554 VDD.n822 VDD.n820 153.601
R14555 VDD.n827 VDD.n820 153.601
R14556 VDD.n831 VDD.n830 153.601
R14557 VDD.n815 VDD.n809 153.601
R14558 VDD.n806 VDD.n804 153.601
R14559 VDD.n811 VDD.n804 153.601
R14560 VDD.n815 VDD.n814 153.601
R14561 VDD.n765 VDD.n758 153.601
R14562 VDD.n762 VDD.n761 153.601
R14563 VDD.n762 VDD.n757 153.601
R14564 VDD.n766 VDD.n765 153.601
R14565 VDD.n889 VDD.n742 153.601
R14566 VDD.n739 VDD.n737 153.601
R14567 VDD.n744 VDD.n737 153.601
R14568 VDD.n889 VDD.n888 153.601
R14569 VDD.n771 VDD.n734 153.601
R14570 VDD.n896 VDD.n735 153.601
R14571 VDD.n899 VDD.n734 153.601
R14572 VDD.n897 VDD.n896 153.601
R14573 VDD.n964 VDD.n959 153.601
R14574 VDD.n962 VDD.n958 153.601
R14575 VDD.n1007 VDD.n958 153.601
R14576 VDD.n1008 VDD.n959 153.601
R14577 VDD.n986 VDD.n939 153.601
R14578 VDD.n985 VDD.n937 153.601
R14579 VDD.n1138 VDD.n937 153.601
R14580 VDD.n1139 VDD.n939 153.601
R14581 VDD.n1056 VDD.n1050 153.601
R14582 VDD.n1047 VDD.n1045 153.601
R14583 VDD.n1052 VDD.n1045 153.601
R14584 VDD.n1056 VDD.n1055 153.601
R14585 VDD.n1134 VDD.n1038 153.601
R14586 VDD.n1042 VDD.n1041 153.601
R14587 VDD.n1042 VDD.n1037 153.601
R14588 VDD.n1135 VDD.n1134 153.601
R14589 VDD.n1129 VDD.n1123 153.601
R14590 VDD.n1120 VDD.n1118 153.601
R14591 VDD.n1125 VDD.n1118 153.601
R14592 VDD.n1129 VDD.n1128 153.601
R14593 VDD.n1113 VDD.n1107 153.601
R14594 VDD.n1104 VDD.n1102 153.601
R14595 VDD.n1109 VDD.n1102 153.601
R14596 VDD.n1113 VDD.n1112 153.601
R14597 VDD.n1090 VDD.n1084 153.601
R14598 VDD.n1081 VDD.n1079 153.601
R14599 VDD.n1086 VDD.n1079 153.601
R14600 VDD.n1090 VDD.n1089 153.601
R14601 VDD.n1074 VDD.n1068 153.601
R14602 VDD.n1065 VDD.n1063 153.601
R14603 VDD.n1070 VDD.n1063 153.601
R14604 VDD.n1074 VDD.n1073 153.601
R14605 VDD.n1024 VDD.n1017 153.601
R14606 VDD.n1021 VDD.n1020 153.601
R14607 VDD.n1021 VDD.n1016 153.601
R14608 VDD.n1025 VDD.n1024 153.601
R14609 VDD.n1148 VDD.n1001 153.601
R14610 VDD.n998 VDD.n996 153.601
R14611 VDD.n1003 VDD.n996 153.601
R14612 VDD.n1148 VDD.n1147 153.601
R14613 VDD.n1030 VDD.n993 153.601
R14614 VDD.n1155 VDD.n994 153.601
R14615 VDD.n1158 VDD.n993 153.601
R14616 VDD.n1156 VDD.n1155 153.601
R14617 VDD.n1223 VDD.n1218 153.601
R14618 VDD.n1221 VDD.n1217 153.601
R14619 VDD.n1266 VDD.n1217 153.601
R14620 VDD.n1267 VDD.n1218 153.601
R14621 VDD.n1245 VDD.n1198 153.601
R14622 VDD.n1244 VDD.n1196 153.601
R14623 VDD.n1397 VDD.n1196 153.601
R14624 VDD.n1398 VDD.n1198 153.601
R14625 VDD.n1315 VDD.n1309 153.601
R14626 VDD.n1306 VDD.n1304 153.601
R14627 VDD.n1311 VDD.n1304 153.601
R14628 VDD.n1315 VDD.n1314 153.601
R14629 VDD.n1393 VDD.n1297 153.601
R14630 VDD.n1301 VDD.n1300 153.601
R14631 VDD.n1301 VDD.n1296 153.601
R14632 VDD.n1394 VDD.n1393 153.601
R14633 VDD.n1388 VDD.n1382 153.601
R14634 VDD.n1379 VDD.n1377 153.601
R14635 VDD.n1384 VDD.n1377 153.601
R14636 VDD.n1388 VDD.n1387 153.601
R14637 VDD.n1372 VDD.n1366 153.601
R14638 VDD.n1363 VDD.n1361 153.601
R14639 VDD.n1368 VDD.n1361 153.601
R14640 VDD.n1372 VDD.n1371 153.601
R14641 VDD.n1349 VDD.n1343 153.601
R14642 VDD.n1340 VDD.n1338 153.601
R14643 VDD.n1345 VDD.n1338 153.601
R14644 VDD.n1349 VDD.n1348 153.601
R14645 VDD.n1333 VDD.n1327 153.601
R14646 VDD.n1324 VDD.n1322 153.601
R14647 VDD.n1329 VDD.n1322 153.601
R14648 VDD.n1333 VDD.n1332 153.601
R14649 VDD.n1283 VDD.n1276 153.601
R14650 VDD.n1280 VDD.n1279 153.601
R14651 VDD.n1280 VDD.n1275 153.601
R14652 VDD.n1284 VDD.n1283 153.601
R14653 VDD.n1407 VDD.n1260 153.601
R14654 VDD.n1257 VDD.n1255 153.601
R14655 VDD.n1262 VDD.n1255 153.601
R14656 VDD.n1407 VDD.n1406 153.601
R14657 VDD.n1289 VDD.n1252 153.601
R14658 VDD.n1414 VDD.n1253 153.601
R14659 VDD.n1417 VDD.n1252 153.601
R14660 VDD.n1415 VDD.n1414 153.601
R14661 VDD.n1482 VDD.n1477 153.601
R14662 VDD.n1480 VDD.n1476 153.601
R14663 VDD.n1525 VDD.n1476 153.601
R14664 VDD.n1526 VDD.n1477 153.601
R14665 VDD.n1504 VDD.n1457 153.601
R14666 VDD.n1503 VDD.n1455 153.601
R14667 VDD.n1656 VDD.n1455 153.601
R14668 VDD.n1657 VDD.n1457 153.601
R14669 VDD.n1574 VDD.n1568 153.601
R14670 VDD.n1565 VDD.n1563 153.601
R14671 VDD.n1570 VDD.n1563 153.601
R14672 VDD.n1574 VDD.n1573 153.601
R14673 VDD.n1652 VDD.n1556 153.601
R14674 VDD.n1560 VDD.n1559 153.601
R14675 VDD.n1560 VDD.n1555 153.601
R14676 VDD.n1653 VDD.n1652 153.601
R14677 VDD.n1647 VDD.n1641 153.601
R14678 VDD.n1638 VDD.n1636 153.601
R14679 VDD.n1643 VDD.n1636 153.601
R14680 VDD.n1647 VDD.n1646 153.601
R14681 VDD.n1631 VDD.n1625 153.601
R14682 VDD.n1622 VDD.n1620 153.601
R14683 VDD.n1627 VDD.n1620 153.601
R14684 VDD.n1631 VDD.n1630 153.601
R14685 VDD.n1608 VDD.n1602 153.601
R14686 VDD.n1599 VDD.n1597 153.601
R14687 VDD.n1604 VDD.n1597 153.601
R14688 VDD.n1608 VDD.n1607 153.601
R14689 VDD.n1592 VDD.n1586 153.601
R14690 VDD.n1583 VDD.n1581 153.601
R14691 VDD.n1588 VDD.n1581 153.601
R14692 VDD.n1592 VDD.n1591 153.601
R14693 VDD.n1542 VDD.n1535 153.601
R14694 VDD.n1539 VDD.n1538 153.601
R14695 VDD.n1539 VDD.n1534 153.601
R14696 VDD.n1543 VDD.n1542 153.601
R14697 VDD.n1666 VDD.n1519 153.601
R14698 VDD.n1516 VDD.n1514 153.601
R14699 VDD.n1521 VDD.n1514 153.601
R14700 VDD.n1666 VDD.n1665 153.601
R14701 VDD.n1548 VDD.n1511 153.601
R14702 VDD.n1673 VDD.n1512 153.601
R14703 VDD.n1676 VDD.n1511 153.601
R14704 VDD.n1674 VDD.n1673 153.601
R14705 VDD.n1741 VDD.n1736 153.601
R14706 VDD.n1739 VDD.n1735 153.601
R14707 VDD.n1784 VDD.n1735 153.601
R14708 VDD.n1785 VDD.n1736 153.601
R14709 VDD.n1763 VDD.n1716 153.601
R14710 VDD.n1762 VDD.n1714 153.601
R14711 VDD.n1915 VDD.n1714 153.601
R14712 VDD.n1916 VDD.n1716 153.601
R14713 VDD.n1833 VDD.n1827 153.601
R14714 VDD.n1824 VDD.n1822 153.601
R14715 VDD.n1829 VDD.n1822 153.601
R14716 VDD.n1833 VDD.n1832 153.601
R14717 VDD.n1911 VDD.n1815 153.601
R14718 VDD.n1819 VDD.n1818 153.601
R14719 VDD.n1819 VDD.n1814 153.601
R14720 VDD.n1912 VDD.n1911 153.601
R14721 VDD.n1906 VDD.n1900 153.601
R14722 VDD.n1897 VDD.n1895 153.601
R14723 VDD.n1902 VDD.n1895 153.601
R14724 VDD.n1906 VDD.n1905 153.601
R14725 VDD.n1890 VDD.n1884 153.601
R14726 VDD.n1881 VDD.n1879 153.601
R14727 VDD.n1886 VDD.n1879 153.601
R14728 VDD.n1890 VDD.n1889 153.601
R14729 VDD.n1867 VDD.n1861 153.601
R14730 VDD.n1858 VDD.n1856 153.601
R14731 VDD.n1863 VDD.n1856 153.601
R14732 VDD.n1867 VDD.n1866 153.601
R14733 VDD.n1851 VDD.n1845 153.601
R14734 VDD.n1842 VDD.n1840 153.601
R14735 VDD.n1847 VDD.n1840 153.601
R14736 VDD.n1851 VDD.n1850 153.601
R14737 VDD.n1801 VDD.n1794 153.601
R14738 VDD.n1798 VDD.n1797 153.601
R14739 VDD.n1798 VDD.n1793 153.601
R14740 VDD.n1802 VDD.n1801 153.601
R14741 VDD.n1925 VDD.n1778 153.601
R14742 VDD.n1775 VDD.n1773 153.601
R14743 VDD.n1780 VDD.n1773 153.601
R14744 VDD.n1925 VDD.n1924 153.601
R14745 VDD.n1807 VDD.n1770 153.601
R14746 VDD.n1932 VDD.n1771 153.601
R14747 VDD.n1935 VDD.n1770 153.601
R14748 VDD.n1933 VDD.n1932 153.601
R14749 VDD.n2000 VDD.n1995 153.601
R14750 VDD.n1998 VDD.n1994 153.601
R14751 VDD.n2043 VDD.n1994 153.601
R14752 VDD.n2044 VDD.n1995 153.601
R14753 VDD.n2022 VDD.n1975 153.601
R14754 VDD.n2021 VDD.n1973 153.601
R14755 VDD.n2174 VDD.n1973 153.601
R14756 VDD.n2175 VDD.n1975 153.601
R14757 VDD.n2092 VDD.n2086 153.601
R14758 VDD.n2083 VDD.n2081 153.601
R14759 VDD.n2088 VDD.n2081 153.601
R14760 VDD.n2092 VDD.n2091 153.601
R14761 VDD.n2170 VDD.n2074 153.601
R14762 VDD.n2078 VDD.n2077 153.601
R14763 VDD.n2078 VDD.n2073 153.601
R14764 VDD.n2171 VDD.n2170 153.601
R14765 VDD.n2165 VDD.n2159 153.601
R14766 VDD.n2156 VDD.n2154 153.601
R14767 VDD.n2161 VDD.n2154 153.601
R14768 VDD.n2165 VDD.n2164 153.601
R14769 VDD.n2149 VDD.n2143 153.601
R14770 VDD.n2140 VDD.n2138 153.601
R14771 VDD.n2145 VDD.n2138 153.601
R14772 VDD.n2149 VDD.n2148 153.601
R14773 VDD.n2126 VDD.n2120 153.601
R14774 VDD.n2117 VDD.n2115 153.601
R14775 VDD.n2122 VDD.n2115 153.601
R14776 VDD.n2126 VDD.n2125 153.601
R14777 VDD.n2110 VDD.n2104 153.601
R14778 VDD.n2101 VDD.n2099 153.601
R14779 VDD.n2106 VDD.n2099 153.601
R14780 VDD.n2110 VDD.n2109 153.601
R14781 VDD.n2060 VDD.n2053 153.601
R14782 VDD.n2057 VDD.n2056 153.601
R14783 VDD.n2057 VDD.n2052 153.601
R14784 VDD.n2061 VDD.n2060 153.601
R14785 VDD.n2184 VDD.n2037 153.601
R14786 VDD.n2034 VDD.n2032 153.601
R14787 VDD.n2039 VDD.n2032 153.601
R14788 VDD.n2184 VDD.n2183 153.601
R14789 VDD.n2066 VDD.n2029 153.601
R14790 VDD.n2191 VDD.n2030 153.601
R14791 VDD.n2194 VDD.n2029 153.601
R14792 VDD.n2192 VDD.n2191 153.601
R14793 VDD.n2259 VDD.n2254 153.601
R14794 VDD.n2257 VDD.n2253 153.601
R14795 VDD.n2302 VDD.n2253 153.601
R14796 VDD.n2303 VDD.n2254 153.601
R14797 VDD.n2281 VDD.n2234 153.601
R14798 VDD.n2280 VDD.n2232 153.601
R14799 VDD.n2433 VDD.n2232 153.601
R14800 VDD.n2434 VDD.n2234 153.601
R14801 VDD.n2351 VDD.n2345 153.601
R14802 VDD.n2342 VDD.n2340 153.601
R14803 VDD.n2347 VDD.n2340 153.601
R14804 VDD.n2351 VDD.n2350 153.601
R14805 VDD.n2429 VDD.n2333 153.601
R14806 VDD.n2337 VDD.n2336 153.601
R14807 VDD.n2337 VDD.n2332 153.601
R14808 VDD.n2430 VDD.n2429 153.601
R14809 VDD.n2424 VDD.n2418 153.601
R14810 VDD.n2415 VDD.n2413 153.601
R14811 VDD.n2420 VDD.n2413 153.601
R14812 VDD.n2424 VDD.n2423 153.601
R14813 VDD.n2408 VDD.n2402 153.601
R14814 VDD.n2399 VDD.n2397 153.601
R14815 VDD.n2404 VDD.n2397 153.601
R14816 VDD.n2408 VDD.n2407 153.601
R14817 VDD.n2385 VDD.n2379 153.601
R14818 VDD.n2376 VDD.n2374 153.601
R14819 VDD.n2381 VDD.n2374 153.601
R14820 VDD.n2385 VDD.n2384 153.601
R14821 VDD.n2369 VDD.n2363 153.601
R14822 VDD.n2360 VDD.n2358 153.601
R14823 VDD.n2365 VDD.n2358 153.601
R14824 VDD.n2369 VDD.n2368 153.601
R14825 VDD.n2319 VDD.n2312 153.601
R14826 VDD.n2316 VDD.n2315 153.601
R14827 VDD.n2316 VDD.n2311 153.601
R14828 VDD.n2320 VDD.n2319 153.601
R14829 VDD.n2443 VDD.n2296 153.601
R14830 VDD.n2293 VDD.n2291 153.601
R14831 VDD.n2298 VDD.n2291 153.601
R14832 VDD.n2443 VDD.n2442 153.601
R14833 VDD.n2325 VDD.n2288 153.601
R14834 VDD.n2450 VDD.n2289 153.601
R14835 VDD.n2453 VDD.n2288 153.601
R14836 VDD.n2451 VDD.n2450 153.601
R14837 VDD.n2518 VDD.n2513 153.601
R14838 VDD.n2516 VDD.n2512 153.601
R14839 VDD.n2561 VDD.n2512 153.601
R14840 VDD.n2562 VDD.n2513 153.601
R14841 VDD.n2540 VDD.n2493 153.601
R14842 VDD.n2539 VDD.n2491 153.601
R14843 VDD.n2692 VDD.n2491 153.601
R14844 VDD.n2693 VDD.n2493 153.601
R14845 VDD.n2610 VDD.n2604 153.601
R14846 VDD.n2601 VDD.n2599 153.601
R14847 VDD.n2606 VDD.n2599 153.601
R14848 VDD.n2610 VDD.n2609 153.601
R14849 VDD.n2688 VDD.n2592 153.601
R14850 VDD.n2596 VDD.n2595 153.601
R14851 VDD.n2596 VDD.n2591 153.601
R14852 VDD.n2689 VDD.n2688 153.601
R14853 VDD.n2683 VDD.n2677 153.601
R14854 VDD.n2674 VDD.n2672 153.601
R14855 VDD.n2679 VDD.n2672 153.601
R14856 VDD.n2683 VDD.n2682 153.601
R14857 VDD.n2667 VDD.n2661 153.601
R14858 VDD.n2658 VDD.n2656 153.601
R14859 VDD.n2663 VDD.n2656 153.601
R14860 VDD.n2667 VDD.n2666 153.601
R14861 VDD.n2644 VDD.n2638 153.601
R14862 VDD.n2635 VDD.n2633 153.601
R14863 VDD.n2640 VDD.n2633 153.601
R14864 VDD.n2644 VDD.n2643 153.601
R14865 VDD.n2628 VDD.n2622 153.601
R14866 VDD.n2619 VDD.n2617 153.601
R14867 VDD.n2624 VDD.n2617 153.601
R14868 VDD.n2628 VDD.n2627 153.601
R14869 VDD.n2578 VDD.n2571 153.601
R14870 VDD.n2575 VDD.n2574 153.601
R14871 VDD.n2575 VDD.n2570 153.601
R14872 VDD.n2579 VDD.n2578 153.601
R14873 VDD.n2702 VDD.n2555 153.601
R14874 VDD.n2552 VDD.n2550 153.601
R14875 VDD.n2557 VDD.n2550 153.601
R14876 VDD.n2702 VDD.n2701 153.601
R14877 VDD.n2584 VDD.n2547 153.601
R14878 VDD.n2709 VDD.n2548 153.601
R14879 VDD.n2712 VDD.n2547 153.601
R14880 VDD.n2710 VDD.n2709 153.601
R14881 VDD.n2777 VDD.n2772 153.601
R14882 VDD.n2775 VDD.n2771 153.601
R14883 VDD.n2820 VDD.n2771 153.601
R14884 VDD.n2821 VDD.n2772 153.601
R14885 VDD.n2799 VDD.n2752 153.601
R14886 VDD.n2798 VDD.n2750 153.601
R14887 VDD.n2951 VDD.n2750 153.601
R14888 VDD.n2952 VDD.n2752 153.601
R14889 VDD.n2869 VDD.n2863 153.601
R14890 VDD.n2860 VDD.n2858 153.601
R14891 VDD.n2865 VDD.n2858 153.601
R14892 VDD.n2869 VDD.n2868 153.601
R14893 VDD.n2947 VDD.n2851 153.601
R14894 VDD.n2855 VDD.n2854 153.601
R14895 VDD.n2855 VDD.n2850 153.601
R14896 VDD.n2948 VDD.n2947 153.601
R14897 VDD.n2942 VDD.n2936 153.601
R14898 VDD.n2933 VDD.n2931 153.601
R14899 VDD.n2938 VDD.n2931 153.601
R14900 VDD.n2942 VDD.n2941 153.601
R14901 VDD.n2926 VDD.n2920 153.601
R14902 VDD.n2917 VDD.n2915 153.601
R14903 VDD.n2922 VDD.n2915 153.601
R14904 VDD.n2926 VDD.n2925 153.601
R14905 VDD.n2903 VDD.n2897 153.601
R14906 VDD.n2894 VDD.n2892 153.601
R14907 VDD.n2899 VDD.n2892 153.601
R14908 VDD.n2903 VDD.n2902 153.601
R14909 VDD.n2887 VDD.n2881 153.601
R14910 VDD.n2878 VDD.n2876 153.601
R14911 VDD.n2883 VDD.n2876 153.601
R14912 VDD.n2887 VDD.n2886 153.601
R14913 VDD.n2837 VDD.n2830 153.601
R14914 VDD.n2834 VDD.n2833 153.601
R14915 VDD.n2834 VDD.n2829 153.601
R14916 VDD.n2838 VDD.n2837 153.601
R14917 VDD.n2961 VDD.n2814 153.601
R14918 VDD.n2811 VDD.n2809 153.601
R14919 VDD.n2816 VDD.n2809 153.601
R14920 VDD.n2961 VDD.n2960 153.601
R14921 VDD.n2843 VDD.n2806 153.601
R14922 VDD.n2968 VDD.n2807 153.601
R14923 VDD.n2971 VDD.n2806 153.601
R14924 VDD.n2969 VDD.n2968 153.601
R14925 VDD.n3036 VDD.n3031 153.601
R14926 VDD.n3034 VDD.n3030 153.601
R14927 VDD.n3079 VDD.n3030 153.601
R14928 VDD.n3080 VDD.n3031 153.601
R14929 VDD.n3058 VDD.n3011 153.601
R14930 VDD.n3057 VDD.n3009 153.601
R14931 VDD.n3210 VDD.n3009 153.601
R14932 VDD.n3211 VDD.n3011 153.601
R14933 VDD.n3128 VDD.n3122 153.601
R14934 VDD.n3119 VDD.n3117 153.601
R14935 VDD.n3124 VDD.n3117 153.601
R14936 VDD.n3128 VDD.n3127 153.601
R14937 VDD.n3206 VDD.n3110 153.601
R14938 VDD.n3114 VDD.n3113 153.601
R14939 VDD.n3114 VDD.n3109 153.601
R14940 VDD.n3207 VDD.n3206 153.601
R14941 VDD.n3201 VDD.n3195 153.601
R14942 VDD.n3192 VDD.n3190 153.601
R14943 VDD.n3197 VDD.n3190 153.601
R14944 VDD.n3201 VDD.n3200 153.601
R14945 VDD.n3185 VDD.n3179 153.601
R14946 VDD.n3176 VDD.n3174 153.601
R14947 VDD.n3181 VDD.n3174 153.601
R14948 VDD.n3185 VDD.n3184 153.601
R14949 VDD.n3162 VDD.n3156 153.601
R14950 VDD.n3153 VDD.n3151 153.601
R14951 VDD.n3158 VDD.n3151 153.601
R14952 VDD.n3162 VDD.n3161 153.601
R14953 VDD.n3146 VDD.n3140 153.601
R14954 VDD.n3137 VDD.n3135 153.601
R14955 VDD.n3142 VDD.n3135 153.601
R14956 VDD.n3146 VDD.n3145 153.601
R14957 VDD.n3096 VDD.n3089 153.601
R14958 VDD.n3093 VDD.n3092 153.601
R14959 VDD.n3093 VDD.n3088 153.601
R14960 VDD.n3097 VDD.n3096 153.601
R14961 VDD.n3220 VDD.n3073 153.601
R14962 VDD.n3070 VDD.n3068 153.601
R14963 VDD.n3075 VDD.n3068 153.601
R14964 VDD.n3220 VDD.n3219 153.601
R14965 VDD.n3102 VDD.n3065 153.601
R14966 VDD.n3227 VDD.n3066 153.601
R14967 VDD.n3230 VDD.n3065 153.601
R14968 VDD.n3228 VDD.n3227 153.601
R14969 VDD.n3295 VDD.n3290 153.601
R14970 VDD.n3293 VDD.n3289 153.601
R14971 VDD.n3338 VDD.n3289 153.601
R14972 VDD.n3339 VDD.n3290 153.601
R14973 VDD.n3317 VDD.n3270 153.601
R14974 VDD.n3316 VDD.n3268 153.601
R14975 VDD.n3469 VDD.n3268 153.601
R14976 VDD.n3470 VDD.n3270 153.601
R14977 VDD.n3387 VDD.n3381 153.601
R14978 VDD.n3378 VDD.n3376 153.601
R14979 VDD.n3383 VDD.n3376 153.601
R14980 VDD.n3387 VDD.n3386 153.601
R14981 VDD.n3465 VDD.n3369 153.601
R14982 VDD.n3373 VDD.n3372 153.601
R14983 VDD.n3373 VDD.n3368 153.601
R14984 VDD.n3466 VDD.n3465 153.601
R14985 VDD.n3460 VDD.n3454 153.601
R14986 VDD.n3451 VDD.n3449 153.601
R14987 VDD.n3456 VDD.n3449 153.601
R14988 VDD.n3460 VDD.n3459 153.601
R14989 VDD.n3444 VDD.n3438 153.601
R14990 VDD.n3435 VDD.n3433 153.601
R14991 VDD.n3440 VDD.n3433 153.601
R14992 VDD.n3444 VDD.n3443 153.601
R14993 VDD.n3421 VDD.n3415 153.601
R14994 VDD.n3412 VDD.n3410 153.601
R14995 VDD.n3417 VDD.n3410 153.601
R14996 VDD.n3421 VDD.n3420 153.601
R14997 VDD.n3405 VDD.n3399 153.601
R14998 VDD.n3396 VDD.n3394 153.601
R14999 VDD.n3401 VDD.n3394 153.601
R15000 VDD.n3405 VDD.n3404 153.601
R15001 VDD.n3355 VDD.n3348 153.601
R15002 VDD.n3352 VDD.n3351 153.601
R15003 VDD.n3352 VDD.n3347 153.601
R15004 VDD.n3356 VDD.n3355 153.601
R15005 VDD.n3479 VDD.n3332 153.601
R15006 VDD.n3329 VDD.n3327 153.601
R15007 VDD.n3334 VDD.n3327 153.601
R15008 VDD.n3479 VDD.n3478 153.601
R15009 VDD.n3361 VDD.n3324 153.601
R15010 VDD.n3486 VDD.n3325 153.601
R15011 VDD.n3489 VDD.n3324 153.601
R15012 VDD.n3487 VDD.n3486 153.601
R15013 VDD.n3554 VDD.n3549 153.601
R15014 VDD.n3552 VDD.n3548 153.601
R15015 VDD.n3597 VDD.n3548 153.601
R15016 VDD.n3598 VDD.n3549 153.601
R15017 VDD.n3576 VDD.n3529 153.601
R15018 VDD.n3575 VDD.n3527 153.601
R15019 VDD.n3728 VDD.n3527 153.601
R15020 VDD.n3729 VDD.n3529 153.601
R15021 VDD.n3646 VDD.n3640 153.601
R15022 VDD.n3637 VDD.n3635 153.601
R15023 VDD.n3642 VDD.n3635 153.601
R15024 VDD.n3646 VDD.n3645 153.601
R15025 VDD.n3724 VDD.n3628 153.601
R15026 VDD.n3632 VDD.n3631 153.601
R15027 VDD.n3632 VDD.n3627 153.601
R15028 VDD.n3725 VDD.n3724 153.601
R15029 VDD.n3719 VDD.n3713 153.601
R15030 VDD.n3710 VDD.n3708 153.601
R15031 VDD.n3715 VDD.n3708 153.601
R15032 VDD.n3719 VDD.n3718 153.601
R15033 VDD.n3703 VDD.n3697 153.601
R15034 VDD.n3694 VDD.n3692 153.601
R15035 VDD.n3699 VDD.n3692 153.601
R15036 VDD.n3703 VDD.n3702 153.601
R15037 VDD.n3680 VDD.n3674 153.601
R15038 VDD.n3671 VDD.n3669 153.601
R15039 VDD.n3676 VDD.n3669 153.601
R15040 VDD.n3680 VDD.n3679 153.601
R15041 VDD.n3664 VDD.n3658 153.601
R15042 VDD.n3655 VDD.n3653 153.601
R15043 VDD.n3660 VDD.n3653 153.601
R15044 VDD.n3664 VDD.n3663 153.601
R15045 VDD.n3614 VDD.n3607 153.601
R15046 VDD.n3611 VDD.n3610 153.601
R15047 VDD.n3611 VDD.n3606 153.601
R15048 VDD.n3615 VDD.n3614 153.601
R15049 VDD.n3738 VDD.n3591 153.601
R15050 VDD.n3588 VDD.n3586 153.601
R15051 VDD.n3593 VDD.n3586 153.601
R15052 VDD.n3738 VDD.n3737 153.601
R15053 VDD.n3620 VDD.n3583 153.601
R15054 VDD.n3745 VDD.n3584 153.601
R15055 VDD.n3748 VDD.n3583 153.601
R15056 VDD.n3746 VDD.n3745 153.601
R15057 VDD.n3813 VDD.n3808 153.601
R15058 VDD.n3811 VDD.n3807 153.601
R15059 VDD.n3856 VDD.n3807 153.601
R15060 VDD.n3857 VDD.n3808 153.601
R15061 VDD.n3835 VDD.n3788 153.601
R15062 VDD.n3834 VDD.n3786 153.601
R15063 VDD.n3987 VDD.n3786 153.601
R15064 VDD.n3988 VDD.n3788 153.601
R15065 VDD.n3905 VDD.n3899 153.601
R15066 VDD.n3896 VDD.n3894 153.601
R15067 VDD.n3901 VDD.n3894 153.601
R15068 VDD.n3905 VDD.n3904 153.601
R15069 VDD.n3983 VDD.n3887 153.601
R15070 VDD.n3891 VDD.n3890 153.601
R15071 VDD.n3891 VDD.n3886 153.601
R15072 VDD.n3984 VDD.n3983 153.601
R15073 VDD.n3978 VDD.n3972 153.601
R15074 VDD.n3969 VDD.n3967 153.601
R15075 VDD.n3974 VDD.n3967 153.601
R15076 VDD.n3978 VDD.n3977 153.601
R15077 VDD.n3962 VDD.n3956 153.601
R15078 VDD.n3953 VDD.n3951 153.601
R15079 VDD.n3958 VDD.n3951 153.601
R15080 VDD.n3962 VDD.n3961 153.601
R15081 VDD.n3939 VDD.n3933 153.601
R15082 VDD.n3930 VDD.n3928 153.601
R15083 VDD.n3935 VDD.n3928 153.601
R15084 VDD.n3939 VDD.n3938 153.601
R15085 VDD.n3923 VDD.n3917 153.601
R15086 VDD.n3914 VDD.n3912 153.601
R15087 VDD.n3919 VDD.n3912 153.601
R15088 VDD.n3923 VDD.n3922 153.601
R15089 VDD.n3873 VDD.n3866 153.601
R15090 VDD.n3870 VDD.n3869 153.601
R15091 VDD.n3870 VDD.n3865 153.601
R15092 VDD.n3874 VDD.n3873 153.601
R15093 VDD.n3997 VDD.n3850 153.601
R15094 VDD.n3847 VDD.n3845 153.601
R15095 VDD.n3852 VDD.n3845 153.601
R15096 VDD.n3997 VDD.n3996 153.601
R15097 VDD.n3879 VDD.n3842 153.601
R15098 VDD.n4004 VDD.n3843 153.601
R15099 VDD.n4007 VDD.n3842 153.601
R15100 VDD.n4005 VDD.n4004 153.601
R15101 VDD.n4072 VDD.n4067 153.601
R15102 VDD.n4070 VDD.n4066 153.601
R15103 VDD.n4115 VDD.n4066 153.601
R15104 VDD.n4116 VDD.n4067 153.601
R15105 VDD.n4094 VDD.n4047 153.601
R15106 VDD.n4093 VDD.n4045 153.601
R15107 VDD.n4246 VDD.n4045 153.601
R15108 VDD.n4247 VDD.n4047 153.601
R15109 VDD.n4164 VDD.n4158 153.601
R15110 VDD.n4155 VDD.n4153 153.601
R15111 VDD.n4160 VDD.n4153 153.601
R15112 VDD.n4164 VDD.n4163 153.601
R15113 VDD.n4242 VDD.n4146 153.601
R15114 VDD.n4150 VDD.n4149 153.601
R15115 VDD.n4150 VDD.n4145 153.601
R15116 VDD.n4243 VDD.n4242 153.601
R15117 VDD.n4237 VDD.n4231 153.601
R15118 VDD.n4228 VDD.n4226 153.601
R15119 VDD.n4233 VDD.n4226 153.601
R15120 VDD.n4237 VDD.n4236 153.601
R15121 VDD.n4221 VDD.n4215 153.601
R15122 VDD.n4212 VDD.n4210 153.601
R15123 VDD.n4217 VDD.n4210 153.601
R15124 VDD.n4221 VDD.n4220 153.601
R15125 VDD.n4198 VDD.n4192 153.601
R15126 VDD.n4189 VDD.n4187 153.601
R15127 VDD.n4194 VDD.n4187 153.601
R15128 VDD.n4198 VDD.n4197 153.601
R15129 VDD.n4182 VDD.n4176 153.601
R15130 VDD.n4173 VDD.n4171 153.601
R15131 VDD.n4178 VDD.n4171 153.601
R15132 VDD.n4182 VDD.n4181 153.601
R15133 VDD.n4132 VDD.n4125 153.601
R15134 VDD.n4129 VDD.n4128 153.601
R15135 VDD.n4129 VDD.n4124 153.601
R15136 VDD.n4133 VDD.n4132 153.601
R15137 VDD.n4256 VDD.n4109 153.601
R15138 VDD.n4106 VDD.n4104 153.601
R15139 VDD.n4111 VDD.n4104 153.601
R15140 VDD.n4256 VDD.n4255 153.601
R15141 VDD.n4138 VDD.n4101 153.601
R15142 VDD.n4263 VDD.n4102 153.601
R15143 VDD.n4266 VDD.n4101 153.601
R15144 VDD.n4264 VDD.n4263 153.601
R15145 VDD.n4331 VDD.n4326 153.601
R15146 VDD.n4329 VDD.n4325 153.601
R15147 VDD.n4374 VDD.n4325 153.601
R15148 VDD.n4375 VDD.n4326 153.601
R15149 VDD.n4353 VDD.n4306 153.601
R15150 VDD.n4352 VDD.n4304 153.601
R15151 VDD.n4505 VDD.n4304 153.601
R15152 VDD.n4506 VDD.n4306 153.601
R15153 VDD.n4423 VDD.n4417 153.601
R15154 VDD.n4414 VDD.n4412 153.601
R15155 VDD.n4419 VDD.n4412 153.601
R15156 VDD.n4423 VDD.n4422 153.601
R15157 VDD.n4501 VDD.n4405 153.601
R15158 VDD.n4409 VDD.n4408 153.601
R15159 VDD.n4409 VDD.n4404 153.601
R15160 VDD.n4502 VDD.n4501 153.601
R15161 VDD.n4496 VDD.n4490 153.601
R15162 VDD.n4487 VDD.n4485 153.601
R15163 VDD.n4492 VDD.n4485 153.601
R15164 VDD.n4496 VDD.n4495 153.601
R15165 VDD.n4480 VDD.n4474 153.601
R15166 VDD.n4471 VDD.n4469 153.601
R15167 VDD.n4476 VDD.n4469 153.601
R15168 VDD.n4480 VDD.n4479 153.601
R15169 VDD.n4457 VDD.n4451 153.601
R15170 VDD.n4448 VDD.n4446 153.601
R15171 VDD.n4453 VDD.n4446 153.601
R15172 VDD.n4457 VDD.n4456 153.601
R15173 VDD.n4441 VDD.n4435 153.601
R15174 VDD.n4432 VDD.n4430 153.601
R15175 VDD.n4437 VDD.n4430 153.601
R15176 VDD.n4441 VDD.n4440 153.601
R15177 VDD.n4391 VDD.n4384 153.601
R15178 VDD.n4388 VDD.n4387 153.601
R15179 VDD.n4388 VDD.n4383 153.601
R15180 VDD.n4392 VDD.n4391 153.601
R15181 VDD.n4515 VDD.n4368 153.601
R15182 VDD.n4365 VDD.n4363 153.601
R15183 VDD.n4370 VDD.n4363 153.601
R15184 VDD.n4515 VDD.n4514 153.601
R15185 VDD.n4397 VDD.n4360 153.601
R15186 VDD.n4522 VDD.n4361 153.601
R15187 VDD.n4525 VDD.n4360 153.601
R15188 VDD.n4523 VDD.n4522 153.601
R15189 VDD.n7094 VDD.n5043 153.601
R15190 VDD.n5049 VDD.n5044 153.601
R15191 VDD.n7095 VDD.n7094 153.601
R15192 VDD.n7088 VDD.n5044 153.601
R15193 VDD.n7084 VDD.n5054 153.601
R15194 VDD.n5059 VDD.n5055 153.601
R15195 VDD.n7085 VDD.n7084 153.601
R15196 VDD.n7078 VDD.n5055 153.601
R15197 VDD.n7074 VDD.n5064 153.601
R15198 VDD.n5072 VDD.n5065 153.601
R15199 VDD.n7075 VDD.n7074 153.601
R15200 VDD.n7068 VDD.n5065 153.601
R15201 VDD.n7064 VDD.n5077 153.601
R15202 VDD.n5083 VDD.n5078 153.601
R15203 VDD.n7065 VDD.n7064 153.601
R15204 VDD.n7058 VDD.n5078 153.601
R15205 VDD.n7054 VDD.n5088 153.601
R15206 VDD.n5093 VDD.n5089 153.601
R15207 VDD.n7055 VDD.n7054 153.601
R15208 VDD.n7048 VDD.n5089 153.601
R15209 VDD.n7044 VDD.n5098 153.601
R15210 VDD.n5106 VDD.n5099 153.601
R15211 VDD.n7045 VDD.n7044 153.601
R15212 VDD.n7038 VDD.n5099 153.601
R15213 VDD.n7027 VDD.n5114 153.601
R15214 VDD.n5121 VDD.n5115 153.601
R15215 VDD.n7028 VDD.n7027 153.601
R15216 VDD.n7021 VDD.n5115 153.601
R15217 VDD.n7017 VDD.n5126 153.601
R15218 VDD.n5134 VDD.n5127 153.601
R15219 VDD.n7018 VDD.n7017 153.601
R15220 VDD.n7011 VDD.n5127 153.601
R15221 VDD.n7007 VDD.n5139 153.601
R15222 VDD.n5145 VDD.n5140 153.601
R15223 VDD.n7008 VDD.n7007 153.601
R15224 VDD.n7001 VDD.n5140 153.601
R15225 VDD.n6997 VDD.n5150 153.601
R15226 VDD.n5155 VDD.n5151 153.601
R15227 VDD.n6998 VDD.n6997 153.601
R15228 VDD.n6991 VDD.n5151 153.601
R15229 VDD.n6987 VDD.n5160 153.601
R15230 VDD.n5168 VDD.n5161 153.601
R15231 VDD.n6988 VDD.n6987 153.601
R15232 VDD.n6981 VDD.n5161 153.601
R15233 VDD.n6959 VDD.n5176 153.601
R15234 VDD.n6958 VDD.n5174 153.601
R15235 VDD.n6968 VDD.n5176 153.601
R15236 VDD.n6967 VDD.n5174 153.601
R15237 VDD.n6953 VDD.n5183 153.601
R15238 VDD.n5187 VDD.n5184 153.601
R15239 VDD.n6954 VDD.n6953 153.601
R15240 VDD.n6947 VDD.n5184 153.601
R15241 VDD.n6943 VDD.n5192 153.601
R15242 VDD.n5200 VDD.n5193 153.601
R15243 VDD.n6944 VDD.n6943 153.601
R15244 VDD.n6937 VDD.n5193 153.601
R15245 VDD.n6933 VDD.n5205 153.601
R15246 VDD.n5211 VDD.n5206 153.601
R15247 VDD.n6934 VDD.n6933 153.601
R15248 VDD.n6927 VDD.n5206 153.601
R15249 VDD.n6923 VDD.n5216 153.601
R15250 VDD.n5221 VDD.n5217 153.601
R15251 VDD.n6924 VDD.n6923 153.601
R15252 VDD.n6917 VDD.n5217 153.601
R15253 VDD.n6913 VDD.n5226 153.601
R15254 VDD.n5234 VDD.n5227 153.601
R15255 VDD.n6914 VDD.n6913 153.601
R15256 VDD.n6907 VDD.n5227 153.601
R15257 VDD.n6896 VDD.n5242 153.601
R15258 VDD.n5249 VDD.n5243 153.601
R15259 VDD.n6897 VDD.n6896 153.601
R15260 VDD.n6890 VDD.n5243 153.601
R15261 VDD.n6886 VDD.n5254 153.601
R15262 VDD.n5262 VDD.n5255 153.601
R15263 VDD.n6887 VDD.n6886 153.601
R15264 VDD.n6880 VDD.n5255 153.601
R15265 VDD.n6876 VDD.n5267 153.601
R15266 VDD.n5273 VDD.n5268 153.601
R15267 VDD.n6877 VDD.n6876 153.601
R15268 VDD.n6870 VDD.n5268 153.601
R15269 VDD.n6866 VDD.n5278 153.601
R15270 VDD.n5283 VDD.n5279 153.601
R15271 VDD.n6867 VDD.n6866 153.601
R15272 VDD.n6860 VDD.n5279 153.601
R15273 VDD.n6856 VDD.n5288 153.601
R15274 VDD.n5296 VDD.n5289 153.601
R15275 VDD.n6857 VDD.n6856 153.601
R15276 VDD.n6850 VDD.n5289 153.601
R15277 VDD.n6828 VDD.n5304 153.601
R15278 VDD.n6827 VDD.n5302 153.601
R15279 VDD.n6837 VDD.n5304 153.601
R15280 VDD.n6836 VDD.n5302 153.601
R15281 VDD.n6822 VDD.n5311 153.601
R15282 VDD.n5315 VDD.n5312 153.601
R15283 VDD.n6823 VDD.n6822 153.601
R15284 VDD.n6816 VDD.n5312 153.601
R15285 VDD.n6812 VDD.n5320 153.601
R15286 VDD.n5328 VDD.n5321 153.601
R15287 VDD.n6813 VDD.n6812 153.601
R15288 VDD.n6806 VDD.n5321 153.601
R15289 VDD.n6802 VDD.n5333 153.601
R15290 VDD.n5339 VDD.n5334 153.601
R15291 VDD.n6803 VDD.n6802 153.601
R15292 VDD.n6796 VDD.n5334 153.601
R15293 VDD.n6792 VDD.n5344 153.601
R15294 VDD.n5349 VDD.n5345 153.601
R15295 VDD.n6793 VDD.n6792 153.601
R15296 VDD.n6786 VDD.n5345 153.601
R15297 VDD.n6782 VDD.n5354 153.601
R15298 VDD.n5362 VDD.n5355 153.601
R15299 VDD.n6783 VDD.n6782 153.601
R15300 VDD.n6776 VDD.n5355 153.601
R15301 VDD.n6765 VDD.n5370 153.601
R15302 VDD.n5377 VDD.n5371 153.601
R15303 VDD.n6766 VDD.n6765 153.601
R15304 VDD.n6759 VDD.n5371 153.601
R15305 VDD.n6755 VDD.n5382 153.601
R15306 VDD.n5390 VDD.n5383 153.601
R15307 VDD.n6756 VDD.n6755 153.601
R15308 VDD.n6749 VDD.n5383 153.601
R15309 VDD.n6745 VDD.n5395 153.601
R15310 VDD.n5401 VDD.n5396 153.601
R15311 VDD.n6746 VDD.n6745 153.601
R15312 VDD.n6739 VDD.n5396 153.601
R15313 VDD.n6735 VDD.n5406 153.601
R15314 VDD.n5411 VDD.n5407 153.601
R15315 VDD.n6736 VDD.n6735 153.601
R15316 VDD.n6729 VDD.n5407 153.601
R15317 VDD.n6725 VDD.n5416 153.601
R15318 VDD.n5424 VDD.n5417 153.601
R15319 VDD.n6726 VDD.n6725 153.601
R15320 VDD.n6719 VDD.n5417 153.601
R15321 VDD.n6697 VDD.n5432 153.601
R15322 VDD.n6696 VDD.n5430 153.601
R15323 VDD.n6706 VDD.n5432 153.601
R15324 VDD.n6705 VDD.n5430 153.601
R15325 VDD.n6691 VDD.n5439 153.601
R15326 VDD.n5443 VDD.n5440 153.601
R15327 VDD.n6692 VDD.n6691 153.601
R15328 VDD.n6685 VDD.n5440 153.601
R15329 VDD.n6681 VDD.n5448 153.601
R15330 VDD.n5456 VDD.n5449 153.601
R15331 VDD.n6682 VDD.n6681 153.601
R15332 VDD.n6675 VDD.n5449 153.601
R15333 VDD.n6671 VDD.n5461 153.601
R15334 VDD.n5467 VDD.n5462 153.601
R15335 VDD.n6672 VDD.n6671 153.601
R15336 VDD.n6665 VDD.n5462 153.601
R15337 VDD.n6661 VDD.n5472 153.601
R15338 VDD.n5477 VDD.n5473 153.601
R15339 VDD.n6662 VDD.n6661 153.601
R15340 VDD.n6655 VDD.n5473 153.601
R15341 VDD.n6651 VDD.n5482 153.601
R15342 VDD.n5490 VDD.n5483 153.601
R15343 VDD.n6652 VDD.n6651 153.601
R15344 VDD.n6645 VDD.n5483 153.601
R15345 VDD.n6634 VDD.n5498 153.601
R15346 VDD.n5505 VDD.n5499 153.601
R15347 VDD.n6635 VDD.n6634 153.601
R15348 VDD.n6628 VDD.n5499 153.601
R15349 VDD.n6624 VDD.n5510 153.601
R15350 VDD.n5518 VDD.n5511 153.601
R15351 VDD.n6625 VDD.n6624 153.601
R15352 VDD.n6618 VDD.n5511 153.601
R15353 VDD.n6614 VDD.n5523 153.601
R15354 VDD.n5529 VDD.n5524 153.601
R15355 VDD.n6615 VDD.n6614 153.601
R15356 VDD.n6608 VDD.n5524 153.601
R15357 VDD.n6604 VDD.n5534 153.601
R15358 VDD.n5539 VDD.n5535 153.601
R15359 VDD.n6605 VDD.n6604 153.601
R15360 VDD.n6598 VDD.n5535 153.601
R15361 VDD.n6594 VDD.n5544 153.601
R15362 VDD.n5552 VDD.n5545 153.601
R15363 VDD.n6595 VDD.n6594 153.601
R15364 VDD.n6588 VDD.n5545 153.601
R15365 VDD.n6566 VDD.n5560 153.601
R15366 VDD.n6565 VDD.n5558 153.601
R15367 VDD.n6575 VDD.n5560 153.601
R15368 VDD.n6574 VDD.n5558 153.601
R15369 VDD.n6560 VDD.n5567 153.601
R15370 VDD.n5571 VDD.n5568 153.601
R15371 VDD.n6561 VDD.n6560 153.601
R15372 VDD.n6554 VDD.n5568 153.601
R15373 VDD.n6550 VDD.n5576 153.601
R15374 VDD.n5584 VDD.n5577 153.601
R15375 VDD.n6551 VDD.n6550 153.601
R15376 VDD.n6544 VDD.n5577 153.601
R15377 VDD.n6540 VDD.n5589 153.601
R15378 VDD.n5595 VDD.n5590 153.601
R15379 VDD.n6541 VDD.n6540 153.601
R15380 VDD.n6534 VDD.n5590 153.601
R15381 VDD.n6530 VDD.n5600 153.601
R15382 VDD.n5605 VDD.n5601 153.601
R15383 VDD.n6531 VDD.n6530 153.601
R15384 VDD.n6524 VDD.n5601 153.601
R15385 VDD.n6520 VDD.n5610 153.601
R15386 VDD.n5618 VDD.n5611 153.601
R15387 VDD.n6521 VDD.n6520 153.601
R15388 VDD.n6514 VDD.n5611 153.601
R15389 VDD.n6503 VDD.n5626 153.601
R15390 VDD.n5633 VDD.n5627 153.601
R15391 VDD.n6504 VDD.n6503 153.601
R15392 VDD.n6497 VDD.n5627 153.601
R15393 VDD.n6493 VDD.n5638 153.601
R15394 VDD.n5646 VDD.n5639 153.601
R15395 VDD.n6494 VDD.n6493 153.601
R15396 VDD.n6487 VDD.n5639 153.601
R15397 VDD.n6483 VDD.n5651 153.601
R15398 VDD.n5657 VDD.n5652 153.601
R15399 VDD.n6484 VDD.n6483 153.601
R15400 VDD.n6477 VDD.n5652 153.601
R15401 VDD.n6473 VDD.n5662 153.601
R15402 VDD.n5667 VDD.n5663 153.601
R15403 VDD.n6474 VDD.n6473 153.601
R15404 VDD.n6467 VDD.n5663 153.601
R15405 VDD.n6463 VDD.n5672 153.601
R15406 VDD.n5680 VDD.n5673 153.601
R15407 VDD.n6464 VDD.n6463 153.601
R15408 VDD.n6457 VDD.n5673 153.601
R15409 VDD.n6435 VDD.n5688 153.601
R15410 VDD.n6434 VDD.n5686 153.601
R15411 VDD.n6444 VDD.n5688 153.601
R15412 VDD.n6443 VDD.n5686 153.601
R15413 VDD.n6429 VDD.n5695 153.601
R15414 VDD.n5699 VDD.n5696 153.601
R15415 VDD.n6430 VDD.n6429 153.601
R15416 VDD.n6423 VDD.n5696 153.601
R15417 VDD.n6419 VDD.n5704 153.601
R15418 VDD.n5712 VDD.n5705 153.601
R15419 VDD.n6420 VDD.n6419 153.601
R15420 VDD.n6413 VDD.n5705 153.601
R15421 VDD.n6409 VDD.n5717 153.601
R15422 VDD.n5723 VDD.n5718 153.601
R15423 VDD.n6410 VDD.n6409 153.601
R15424 VDD.n6403 VDD.n5718 153.601
R15425 VDD.n6399 VDD.n5728 153.601
R15426 VDD.n5733 VDD.n5729 153.601
R15427 VDD.n6400 VDD.n6399 153.601
R15428 VDD.n6393 VDD.n5729 153.601
R15429 VDD.n6389 VDD.n5738 153.601
R15430 VDD.n5746 VDD.n5739 153.601
R15431 VDD.n6390 VDD.n6389 153.601
R15432 VDD.n6383 VDD.n5739 153.601
R15433 VDD.n6372 VDD.n5754 153.601
R15434 VDD.n5761 VDD.n5755 153.601
R15435 VDD.n6373 VDD.n6372 153.601
R15436 VDD.n6366 VDD.n5755 153.601
R15437 VDD.n6362 VDD.n5766 153.601
R15438 VDD.n5774 VDD.n5767 153.601
R15439 VDD.n6363 VDD.n6362 153.601
R15440 VDD.n6356 VDD.n5767 153.601
R15441 VDD.n6352 VDD.n5779 153.601
R15442 VDD.n5785 VDD.n5780 153.601
R15443 VDD.n6353 VDD.n6352 153.601
R15444 VDD.n6346 VDD.n5780 153.601
R15445 VDD.n6342 VDD.n5790 153.601
R15446 VDD.n5795 VDD.n5791 153.601
R15447 VDD.n6343 VDD.n6342 153.601
R15448 VDD.n6336 VDD.n5791 153.601
R15449 VDD.n6332 VDD.n5800 153.601
R15450 VDD.n5808 VDD.n5801 153.601
R15451 VDD.n6333 VDD.n6332 153.601
R15452 VDD.n6326 VDD.n5801 153.601
R15453 VDD.n6304 VDD.n5816 153.601
R15454 VDD.n6303 VDD.n5814 153.601
R15455 VDD.n6313 VDD.n5816 153.601
R15456 VDD.n6312 VDD.n5814 153.601
R15457 VDD.n6298 VDD.n5823 153.601
R15458 VDD.n5827 VDD.n5824 153.601
R15459 VDD.n6299 VDD.n6298 153.601
R15460 VDD.n6292 VDD.n5824 153.601
R15461 VDD.n6288 VDD.n5832 153.601
R15462 VDD.n5840 VDD.n5833 153.601
R15463 VDD.n6289 VDD.n6288 153.601
R15464 VDD.n6282 VDD.n5833 153.601
R15465 VDD.n6278 VDD.n5845 153.601
R15466 VDD.n5851 VDD.n5846 153.601
R15467 VDD.n6279 VDD.n6278 153.601
R15468 VDD.n6272 VDD.n5846 153.601
R15469 VDD.n6268 VDD.n5856 153.601
R15470 VDD.n5861 VDD.n5857 153.601
R15471 VDD.n6269 VDD.n6268 153.601
R15472 VDD.n6262 VDD.n5857 153.601
R15473 VDD.n6258 VDD.n5866 153.601
R15474 VDD.n5874 VDD.n5867 153.601
R15475 VDD.n6259 VDD.n6258 153.601
R15476 VDD.n6252 VDD.n5867 153.601
R15477 VDD.n6241 VDD.n5882 153.601
R15478 VDD.n5889 VDD.n5883 153.601
R15479 VDD.n6242 VDD.n6241 153.601
R15480 VDD.n6235 VDD.n5883 153.601
R15481 VDD.n6231 VDD.n5894 153.601
R15482 VDD.n5902 VDD.n5895 153.601
R15483 VDD.n6232 VDD.n6231 153.601
R15484 VDD.n6225 VDD.n5895 153.601
R15485 VDD.n6221 VDD.n5907 153.601
R15486 VDD.n5913 VDD.n5908 153.601
R15487 VDD.n6222 VDD.n6221 153.601
R15488 VDD.n6215 VDD.n5908 153.601
R15489 VDD.n6211 VDD.n5918 153.601
R15490 VDD.n5923 VDD.n5919 153.601
R15491 VDD.n6212 VDD.n6211 153.601
R15492 VDD.n6205 VDD.n5919 153.601
R15493 VDD.n6201 VDD.n5928 153.601
R15494 VDD.n5936 VDD.n5929 153.601
R15495 VDD.n6202 VDD.n6201 153.601
R15496 VDD.n6195 VDD.n5929 153.601
R15497 VDD.n6173 VDD.n5944 153.601
R15498 VDD.n6172 VDD.n5942 153.601
R15499 VDD.n6182 VDD.n5944 153.601
R15500 VDD.n6181 VDD.n5942 153.601
R15501 VDD.n6167 VDD.n5951 153.601
R15502 VDD.n5955 VDD.n5952 153.601
R15503 VDD.n6168 VDD.n6167 153.601
R15504 VDD.n6161 VDD.n5952 153.601
R15505 VDD.n6157 VDD.n5960 153.601
R15506 VDD.n5968 VDD.n5961 153.601
R15507 VDD.n6158 VDD.n6157 153.601
R15508 VDD.n6151 VDD.n5961 153.601
R15509 VDD.n6147 VDD.n5973 153.601
R15510 VDD.n5979 VDD.n5974 153.601
R15511 VDD.n6148 VDD.n6147 153.601
R15512 VDD.n6141 VDD.n5974 153.601
R15513 VDD.n6137 VDD.n5984 153.601
R15514 VDD.n5989 VDD.n5985 153.601
R15515 VDD.n6138 VDD.n6137 153.601
R15516 VDD.n6131 VDD.n5985 153.601
R15517 VDD.n6127 VDD.n5994 153.601
R15518 VDD.n6002 VDD.n5995 153.601
R15519 VDD.n6128 VDD.n6127 153.601
R15520 VDD.n6121 VDD.n5995 153.601
R15521 VDD.n6110 VDD.n6010 153.601
R15522 VDD.n6017 VDD.n6011 153.601
R15523 VDD.n6111 VDD.n6110 153.601
R15524 VDD.n6104 VDD.n6011 153.601
R15525 VDD.n6100 VDD.n6022 153.601
R15526 VDD.n6030 VDD.n6023 153.601
R15527 VDD.n6101 VDD.n6100 153.601
R15528 VDD.n6094 VDD.n6023 153.601
R15529 VDD.n6090 VDD.n6035 153.601
R15530 VDD.n6041 VDD.n6036 153.601
R15531 VDD.n6091 VDD.n6090 153.601
R15532 VDD.n6084 VDD.n6036 153.601
R15533 VDD.n6080 VDD.n6046 153.601
R15534 VDD.n6051 VDD.n6047 153.601
R15535 VDD.n6081 VDD.n6080 153.601
R15536 VDD.n6074 VDD.n6047 153.601
R15537 VDD.n6070 VDD.n6056 153.601
R15538 VDD.n6060 VDD.n6057 153.601
R15539 VDD.n6071 VDD.n6070 153.601
R15540 VDD.n6061 VDD.n6057 153.601
R15541 VDD.t100 VDD.n412 151.594
R15542 VDD.n664 VDD.t144 150.56
R15543 VDD.n660 VDD.t105 150.56
R15544 VDD.n923 VDD.t125 150.56
R15545 VDD.n919 VDD.t207 150.56
R15546 VDD.n1182 VDD.t185 150.56
R15547 VDD.n1178 VDD.t177 150.56
R15548 VDD.n1441 VDD.t132 150.56
R15549 VDD.n1437 VDD.t98 150.56
R15550 VDD.n1700 VDD.t149 150.56
R15551 VDD.n1696 VDD.t108 150.56
R15552 VDD.n1959 VDD.t166 150.56
R15553 VDD.n1955 VDD.t139 150.56
R15554 VDD.n2218 VDD.t158 150.56
R15555 VDD.n2214 VDD.t118 150.56
R15556 VDD.n2477 VDD.t164 150.56
R15557 VDD.n2473 VDD.t130 150.56
R15558 VDD.n2736 VDD.t162 150.56
R15559 VDD.n2732 VDD.t128 150.56
R15560 VDD.n2995 VDD.t172 150.56
R15561 VDD.n2991 VDD.t142 150.56
R15562 VDD.n3254 VDD.t179 150.56
R15563 VDD.n3250 VDD.t168 150.56
R15564 VDD.n3513 VDD.t137 150.56
R15565 VDD.n3509 VDD.t103 150.56
R15566 VDD.n3772 VDD.t153 150.56
R15567 VDD.n3768 VDD.t113 150.56
R15568 VDD.n4031 VDD.t115 150.56
R15569 VDD.n4027 VDD.t203 150.56
R15570 VDD.n4290 VDD.t194 150.56
R15571 VDD.n4286 VDD.t181 150.56
R15572 VDD.n4549 VDD.t183 150.56
R15573 VDD.n4545 VDD.t174 150.56
R15574 VDD.n162 VDD.t196 150.273
R15575 VDD.n158 VDD.t189 150.273
R15576 VDD.t209 VDD.n153 150.273
R15577 VDD.t122 VDD.n672 150.273
R15578 VDD.t201 VDD.n931 150.273
R15579 VDD.t110 VDD.n1190 150.273
R15580 VDD.t146 VDD.n1449 150.273
R15581 VDD.t120 VDD.n1708 150.273
R15582 VDD.t155 VDD.n1967 150.273
R15583 VDD.t212 VDD.n2226 150.273
R15584 VDD.t160 VDD.n2485 150.273
R15585 VDD.t170 VDD.n2744 150.273
R15586 VDD.t205 VDD.n3003 150.273
R15587 VDD.t134 VDD.n3262 150.273
R15588 VDD.t151 VDD.n3521 150.273
R15589 VDD.t198 VDD.n3780 150.273
R15590 VDD.t187 VDD.n4039 150.273
R15591 VDD.t192 VDD.n4298 150.273
R15592 VDD.n6096 VDD.n6093 143.812
R15593 VDD.n6114 VDD.n6113 143.812
R15594 VDD.n6123 VDD.n6120 143.812
R15595 VDD.n6153 VDD.n6150 143.812
R15596 VDD.n6178 VDD.n6177 143.812
R15597 VDD.n6197 VDD.n6194 143.812
R15598 VDD.n6227 VDD.n6224 143.812
R15599 VDD.n6245 VDD.n6244 143.812
R15600 VDD.n6254 VDD.n6251 143.812
R15601 VDD.n6284 VDD.n6281 143.812
R15602 VDD.n6309 VDD.n6308 143.812
R15603 VDD.n6328 VDD.n6325 143.812
R15604 VDD.n6358 VDD.n6355 143.812
R15605 VDD.n6376 VDD.n6375 143.812
R15606 VDD.n6385 VDD.n6382 143.812
R15607 VDD.n6415 VDD.n6412 143.812
R15608 VDD.n6440 VDD.n6439 143.812
R15609 VDD.n6459 VDD.n6456 143.812
R15610 VDD.n6489 VDD.n6486 143.812
R15611 VDD.n6507 VDD.n6506 143.812
R15612 VDD.n6516 VDD.n6513 143.812
R15613 VDD.n6546 VDD.n6543 143.812
R15614 VDD.n6571 VDD.n6570 143.812
R15615 VDD.n6590 VDD.n6587 143.812
R15616 VDD.n6620 VDD.n6617 143.812
R15617 VDD.n6638 VDD.n6637 143.812
R15618 VDD.n6647 VDD.n6644 143.812
R15619 VDD.n6677 VDD.n6674 143.812
R15620 VDD.n6702 VDD.n6701 143.812
R15621 VDD.n6721 VDD.n6718 143.812
R15622 VDD.n6751 VDD.n6748 143.812
R15623 VDD.n6769 VDD.n6768 143.812
R15624 VDD.n6778 VDD.n6775 143.812
R15625 VDD.n6808 VDD.n6805 143.812
R15626 VDD.n6833 VDD.n6832 143.812
R15627 VDD.n6852 VDD.n6849 143.812
R15628 VDD.n6882 VDD.n6879 143.812
R15629 VDD.n6900 VDD.n6899 143.812
R15630 VDD.n6909 VDD.n6906 143.812
R15631 VDD.n6939 VDD.n6936 143.812
R15632 VDD.n6964 VDD.n6963 143.812
R15633 VDD.n6983 VDD.n6980 143.812
R15634 VDD.n7013 VDD.n7010 143.812
R15635 VDD.n7031 VDD.n7030 143.812
R15636 VDD.n7040 VDD.n7037 143.812
R15637 VDD.n7070 VDD.n7067 143.812
R15638 VDD.n7099 VDD.n7097 143.812
R15639 VDD.n7101 VDD.n7100 125.284
R15640 VDD.n6063 VDD.t523 123.344
R15641 VDD.n6073 VDD.t523 123.344
R15642 VDD.n6076 VDD.t371 123.344
R15643 VDD.n6083 VDD.t371 123.344
R15644 VDD.n6086 VDD.t356 123.344
R15645 VDD.n6093 VDD.t356 123.344
R15646 VDD.n6096 VDD.t316 123.344
R15647 VDD.n6103 VDD.t316 123.344
R15648 VDD.n6106 VDD.t326 123.344
R15649 VDD.n6113 VDD.t326 123.344
R15650 VDD.n6114 VDD.t460 123.344
R15651 VDD.n6120 VDD.t460 123.344
R15652 VDD.n6123 VDD.t4 123.344
R15653 VDD.n6130 VDD.t4 123.344
R15654 VDD.n6133 VDD.t618 123.344
R15655 VDD.n6140 VDD.t618 123.344
R15656 VDD.n6143 VDD.t388 123.344
R15657 VDD.n6150 VDD.t388 123.344
R15658 VDD.n6153 VDD.t458 123.344
R15659 VDD.n6160 VDD.t458 123.344
R15660 VDD.n6163 VDD.t20 123.344
R15661 VDD.n6170 VDD.t20 123.344
R15662 VDD.t474 VDD.n6171 123.344
R15663 VDD.t474 VDD.n6178 123.344
R15664 VDD.n6177 VDD.t716 123.344
R15665 VDD.n6194 VDD.t716 123.344
R15666 VDD.n6197 VDD.t27 123.344
R15667 VDD.n6204 VDD.t27 123.344
R15668 VDD.n6207 VDD.t81 123.344
R15669 VDD.n6214 VDD.t81 123.344
R15670 VDD.n6217 VDD.t540 123.344
R15671 VDD.n6224 VDD.t540 123.344
R15672 VDD.n6227 VDD.t395 123.344
R15673 VDD.n6234 VDD.t395 123.344
R15674 VDD.n6237 VDD.t282 123.344
R15675 VDD.n6244 VDD.t282 123.344
R15676 VDD.n6245 VDD.t839 123.344
R15677 VDD.n6251 VDD.t839 123.344
R15678 VDD.n6254 VDD.t280 123.344
R15679 VDD.n6261 VDD.t280 123.344
R15680 VDD.n6264 VDD.t547 123.344
R15681 VDD.n6271 VDD.t547 123.344
R15682 VDD.n6274 VDD.t538 123.344
R15683 VDD.n6281 VDD.t538 123.344
R15684 VDD.n6284 VDD.t836 123.344
R15685 VDD.n6291 VDD.t836 123.344
R15686 VDD.n6294 VDD.t542 123.344
R15687 VDD.n6301 VDD.t542 123.344
R15688 VDD.t536 VDD.n6302 123.344
R15689 VDD.t536 VDD.n6309 123.344
R15690 VDD.n6308 VDD.t720 123.344
R15691 VDD.n6325 VDD.t720 123.344
R15692 VDD.n6328 VDD.t385 123.344
R15693 VDD.n6335 VDD.t385 123.344
R15694 VDD.n6338 VDD.t804 123.344
R15695 VDD.n6345 VDD.t804 123.344
R15696 VDD.n6348 VDD.t390 123.344
R15697 VDD.n6355 VDD.t390 123.344
R15698 VDD.n6358 VDD.t64 123.344
R15699 VDD.n6365 VDD.t64 123.344
R15700 VDD.n6368 VDD.t0 123.344
R15701 VDD.n6375 VDD.t0 123.344
R15702 VDD.n6376 VDD.t735 123.344
R15703 VDD.n6382 VDD.t735 123.344
R15704 VDD.n6385 VDD.t2 123.344
R15705 VDD.n6392 VDD.t2 123.344
R15706 VDD.n6395 VDD.t349 123.344
R15707 VDD.n6402 VDD.t349 123.344
R15708 VDD.n6405 VDD.t561 123.344
R15709 VDD.n6412 VDD.t561 123.344
R15710 VDD.n6415 VDD.t862 123.344
R15711 VDD.n6422 VDD.t862 123.344
R15712 VDD.n6425 VDD.t277 123.344
R15713 VDD.n6432 VDD.t277 123.344
R15714 VDD.t285 VDD.n6433 123.344
R15715 VDD.t285 VDD.n6440 123.344
R15716 VDD.n6439 VDD.t450 123.344
R15717 VDD.n6456 VDD.t450 123.344
R15718 VDD.n6459 VDD.t495 123.344
R15719 VDD.n6466 VDD.t495 123.344
R15720 VDD.n6469 VDD.t347 123.344
R15721 VDD.n6476 VDD.t347 123.344
R15722 VDD.n6479 VDD.t639 123.344
R15723 VDD.n6486 VDD.t639 123.344
R15724 VDD.n6489 VDD.t503 123.344
R15725 VDD.n6496 VDD.t503 123.344
R15726 VDD.n6499 VDD.t430 123.344
R15727 VDD.n6506 VDD.t430 123.344
R15728 VDD.n6507 VDD.t899 123.344
R15729 VDD.n6513 VDD.t899 123.344
R15730 VDD.n6516 VDD.t428 123.344
R15731 VDD.n6523 VDD.t428 123.344
R15732 VDD.n6526 VDD.t78 123.344
R15733 VDD.n6533 VDD.t78 123.344
R15734 VDD.n6536 VDD.t637 123.344
R15735 VDD.n6543 VDD.t637 123.344
R15736 VDD.n6546 VDD.t257 123.344
R15737 VDD.n6553 VDD.t257 123.344
R15738 VDD.n6556 VDD.t18 123.344
R15739 VDD.n6563 VDD.t18 123.344
R15740 VDD.t563 VDD.n6564 123.344
R15741 VDD.t563 VDD.n6571 123.344
R15742 VDD.n6570 VDD.t16 123.344
R15743 VDD.n6587 VDD.t16 123.344
R15744 VDD.n6590 VDD.t70 123.344
R15745 VDD.n6597 VDD.t70 123.344
R15746 VDD.n6600 VDD.t400 123.344
R15747 VDD.n6607 VDD.t400 123.344
R15748 VDD.n6610 VDD.t635 123.344
R15749 VDD.n6617 VDD.t635 123.344
R15750 VDD.n6620 VDD.t625 123.344
R15751 VDD.n6627 VDD.t625 123.344
R15752 VDD.n6630 VDD.t306 123.344
R15753 VDD.n6637 VDD.t306 123.344
R15754 VDD.n6638 VDD.t40 123.344
R15755 VDD.n6644 VDD.t40 123.344
R15756 VDD.n6647 VDD.t420 123.344
R15757 VDD.n6654 VDD.t420 123.344
R15758 VDD.n6657 VDD.t465 123.344
R15759 VDD.n6664 VDD.t465 123.344
R15760 VDD.n6667 VDD.t352 123.344
R15761 VDD.n6674 VDD.t352 123.344
R15762 VDD.n6677 VDD.t37 123.344
R15763 VDD.n6684 VDD.t37 123.344
R15764 VDD.n6687 VDD.t68 123.344
R15765 VDD.n6694 VDD.t68 123.344
R15766 VDD.t364 VDD.n6695 123.344
R15767 VDD.t364 VDD.n6702 123.344
R15768 VDD.n6701 VDD.t718 123.344
R15769 VDD.n6718 VDD.t718 123.344
R15770 VDD.n6721 VDD.t411 123.344
R15771 VDD.n6728 VDD.t411 123.344
R15772 VDD.n6731 VDD.t287 123.344
R15773 VDD.n6738 VDD.t287 123.344
R15774 VDD.n6741 VDD.t568 123.344
R15775 VDD.n6748 VDD.t568 123.344
R15776 VDD.n6751 VDD.t439 123.344
R15777 VDD.n6758 VDD.t439 123.344
R15778 VDD.n6761 VDD.t215 123.344
R15779 VDD.n6768 VDD.t215 123.344
R15780 VDD.n6769 VDD.t485 123.344
R15781 VDD.n6775 VDD.t485 123.344
R15782 VDD.n6778 VDD.t74 123.344
R15783 VDD.n6785 VDD.t74 123.344
R15784 VDD.n6788 VDD.t604 123.344
R15785 VDD.n6795 VDD.t604 123.344
R15786 VDD.n6798 VDD.t358 123.344
R15787 VDD.n6805 VDD.t358 123.344
R15788 VDD.n6808 VDD.t482 123.344
R15789 VDD.n6815 VDD.t482 123.344
R15790 VDD.n6818 VDD.t94 123.344
R15791 VDD.n6825 VDD.t94 123.344
R15792 VDD.t493 VDD.n6826 123.344
R15793 VDD.t493 VDD.n6833 123.344
R15794 VDD.n6832 VDD.t275 123.344
R15795 VDD.n6849 VDD.t275 123.344
R15796 VDD.n6852 VDD.t308 123.344
R15797 VDD.n6859 VDD.t308 123.344
R15798 VDD.n6862 VDD.t418 123.344
R15799 VDD.n6869 VDD.t418 123.344
R15800 VDD.n6872 VDD.t90 123.344
R15801 VDD.n6879 VDD.t90 123.344
R15802 VDD.n6882 VDD.t442 123.344
R15803 VDD.n6889 VDD.t442 123.344
R15804 VDD.n6892 VDD.t501 123.344
R15805 VDD.n6899 VDD.t501 123.344
R15806 VDD.n6900 VDD.t376 123.344
R15807 VDD.n6906 VDD.t376 123.344
R15808 VDD.n6909 VDD.t261 123.344
R15809 VDD.n6916 VDD.t261 123.344
R15810 VDD.n6919 VDD.t335 123.344
R15811 VDD.n6926 VDD.t335 123.344
R15812 VDD.n6929 VDD.t566 123.344
R15813 VDD.n6936 VDD.t566 123.344
R15814 VDD.n6939 VDD.t343 123.344
R15815 VDD.n6946 VDD.t343 123.344
R15816 VDD.n6949 VDD.t487 123.344
R15817 VDD.n6956 VDD.t487 123.344
R15818 VDD.t478 VDD.n6957 123.344
R15819 VDD.t478 VDD.n6964 123.344
R15820 VDD.n6963 VDD.t452 123.344
R15821 VDD.n6980 VDD.t452 123.344
R15822 VDD.n6983 VDD.t425 123.344
R15823 VDD.n6990 VDD.t425 123.344
R15824 VDD.n6993 VDD.t506 123.344
R15825 VDD.n7000 VDD.t506 123.344
R15826 VDD.n7003 VDD.t763 123.344
R15827 VDD.n7010 VDD.t763 123.344
R15828 VDD.n7013 VDD.t529 123.344
R15829 VDD.n7020 VDD.t529 123.344
R15830 VDD.n7023 VDD.t222 123.344
R15831 VDD.n7030 VDD.t222 123.344
R15832 VDD.n7031 VDD.t614 123.344
R15833 VDD.n7037 VDD.t614 123.344
R15834 VDD.n7040 VDD.t303 123.344
R15835 VDD.n7047 VDD.t303 123.344
R15836 VDD.n7050 VDD.t62 123.344
R15837 VDD.n7057 VDD.t62 123.344
R15838 VDD.n7060 VDD.t408 123.344
R15839 VDD.n7067 VDD.t408 123.344
R15840 VDD.n7070 VDD.t611 123.344
R15841 VDD.n7077 VDD.t611 123.344
R15842 VDD.n7080 VDD.t628 123.344
R15843 VDD.n7087 VDD.t628 123.344
R15844 VDD.n7090 VDD.t643 123.344
R15845 VDD.n7097 VDD.t643 123.344
R15846 VDD.t755 VDD.n7099 123.344
R15847 VDD.n7304 VDD.n7303 99.0123
R15848 VDD.n7305 VDD.n7304 99.0123
R15849 VDD.n6076 VDD.n6073 75.5806
R15850 VDD.n6086 VDD.n6083 75.5806
R15851 VDD.n6106 VDD.n6103 75.5806
R15852 VDD.n6133 VDD.n6130 75.5806
R15853 VDD.n6143 VDD.n6140 75.5806
R15854 VDD.n6163 VDD.n6160 75.5806
R15855 VDD.n6171 VDD.n6170 75.5806
R15856 VDD.n6207 VDD.n6204 75.5806
R15857 VDD.n6217 VDD.n6214 75.5806
R15858 VDD.n6237 VDD.n6234 75.5806
R15859 VDD.n6264 VDD.n6261 75.5806
R15860 VDD.n6274 VDD.n6271 75.5806
R15861 VDD.n6294 VDD.n6291 75.5806
R15862 VDD.n6302 VDD.n6301 75.5806
R15863 VDD.n6338 VDD.n6335 75.5806
R15864 VDD.n6348 VDD.n6345 75.5806
R15865 VDD.n6368 VDD.n6365 75.5806
R15866 VDD.n6395 VDD.n6392 75.5806
R15867 VDD.n6405 VDD.n6402 75.5806
R15868 VDD.n6425 VDD.n6422 75.5806
R15869 VDD.n6433 VDD.n6432 75.5806
R15870 VDD.n6469 VDD.n6466 75.5806
R15871 VDD.n6479 VDD.n6476 75.5806
R15872 VDD.n6499 VDD.n6496 75.5806
R15873 VDD.n6526 VDD.n6523 75.5806
R15874 VDD.n6536 VDD.n6533 75.5806
R15875 VDD.n6556 VDD.n6553 75.5806
R15876 VDD.n6564 VDD.n6563 75.5806
R15877 VDD.n6600 VDD.n6597 75.5806
R15878 VDD.n6610 VDD.n6607 75.5806
R15879 VDD.n6630 VDD.n6627 75.5806
R15880 VDD.n6657 VDD.n6654 75.5806
R15881 VDD.n6667 VDD.n6664 75.5806
R15882 VDD.n6687 VDD.n6684 75.5806
R15883 VDD.n6695 VDD.n6694 75.5806
R15884 VDD.n6731 VDD.n6728 75.5806
R15885 VDD.n6741 VDD.n6738 75.5806
R15886 VDD.n6761 VDD.n6758 75.5806
R15887 VDD.n6788 VDD.n6785 75.5806
R15888 VDD.n6798 VDD.n6795 75.5806
R15889 VDD.n6818 VDD.n6815 75.5806
R15890 VDD.n6826 VDD.n6825 75.5806
R15891 VDD.n6862 VDD.n6859 75.5806
R15892 VDD.n6872 VDD.n6869 75.5806
R15893 VDD.n6892 VDD.n6889 75.5806
R15894 VDD.n6919 VDD.n6916 75.5806
R15895 VDD.n6929 VDD.n6926 75.5806
R15896 VDD.n6949 VDD.n6946 75.5806
R15897 VDD.n6957 VDD.n6956 75.5806
R15898 VDD.n6993 VDD.n6990 75.5806
R15899 VDD.n7003 VDD.n7000 75.5806
R15900 VDD.n7023 VDD.n7020 75.5806
R15901 VDD.n7050 VDD.n7047 75.5806
R15902 VDD.n7060 VDD.n7057 75.5806
R15903 VDD.n7080 VDD.n7077 75.5806
R15904 VDD.n7090 VDD.n7087 75.5806
R15905 VDD.n153 VDD.t967 74.951
R15906 VDD.n672 VDD.t929 74.951
R15907 VDD.n931 VDD.t943 74.951
R15908 VDD.n1190 VDD.t924 74.951
R15909 VDD.n1449 VDD.t966 74.951
R15910 VDD.n1708 VDD.t935 74.951
R15911 VDD.n1967 VDD.t963 74.951
R15912 VDD.n2226 VDD.t961 74.951
R15913 VDD.n2485 VDD.t939 74.951
R15914 VDD.n2744 VDD.t959 74.951
R15915 VDD.n3003 VDD.t974 74.951
R15916 VDD.n3262 VDD.t969 74.951
R15917 VDD.n3521 VDD.t965 74.951
R15918 VDD.n3780 VDD.t946 74.951
R15919 VDD.n4039 VDD.t958 74.951
R15920 VDD.n4298 VDD.t962 74.951
R15921 VDD.n161 VDD.t947 74.4891
R15922 VDD.n157 VDD.t954 74.4891
R15923 VDD.n412 VDD.t964 73.6304
R15924 VDD.n665 VDD.t948 73.6304
R15925 VDD.n661 VDD.t955 73.6304
R15926 VDD.n924 VDD.t933 73.6304
R15927 VDD.n920 VDD.t949 73.6304
R15928 VDD.n1183 VDD.t970 73.6304
R15929 VDD.n1179 VDD.t930 73.6304
R15930 VDD.n1442 VDD.t931 73.6304
R15931 VDD.n1438 VDD.t944 73.6304
R15932 VDD.n1701 VDD.t925 73.6304
R15933 VDD.n1697 VDD.t940 73.6304
R15934 VDD.n1960 VDD.t926 73.6304
R15935 VDD.n1956 VDD.t941 73.6304
R15936 VDD.n2219 VDD.t973 73.6304
R15937 VDD.n2215 VDD.t936 73.6304
R15938 VDD.n2478 VDD.t938 73.6304
R15939 VDD.n2474 VDD.t952 73.6304
R15940 VDD.n2737 VDD.t971 73.6304
R15941 VDD.n2733 VDD.t932 73.6304
R15942 VDD.n2996 VDD.t968 73.6304
R15943 VDD.n2992 VDD.t927 73.6304
R15944 VDD.n3255 VDD.t972 73.6304
R15945 VDD.n3251 VDD.t934 73.6304
R15946 VDD.n3514 VDD.t928 73.6304
R15947 VDD.n3510 VDD.t942 73.6304
R15948 VDD.n3773 VDD.t937 73.6304
R15949 VDD.n3769 VDD.t950 73.6304
R15950 VDD.n4032 VDD.t957 73.6304
R15951 VDD.n4028 VDD.t960 73.6304
R15952 VDD.n4291 VDD.t951 73.6304
R15953 VDD.n4287 VDD.t956 73.6304
R15954 VDD.n4550 VDD.t945 73.6304
R15955 VDD.n4546 VDD.t953 73.6304
R15956 VDD VDD.t775 69.9004
R15957 VDD VDD.t448 69.9004
R15958 VDD VDD.t853 69.9004
R15959 VDD VDD.t789 69.9004
R15960 VDD VDD.t361 69.9004
R15961 VDD VDD.t382 69.9004
R15962 VDD VDD.t893 69.9004
R15963 VDD VDD.t508 69.9004
R15964 VDD VDD.n7106 65.5111
R15965 VDD.n7295 VDD.n7294 54.1632
R15966 VDD.n671 VDD 39.9701
R15967 VDD.n670 VDD 38.0684
R15968 VDD.n378 VDD.t190 37.5148
R15969 VDD.n403 VDD.t190 37.5148
R15970 VDD.t101 VDD.n182 37.5148
R15971 VDD.t101 VDD.n223 37.5148
R15972 VDD.n626 VDD.t210 37.5148
R15973 VDD.n651 VDD.t210 37.5148
R15974 VDD.t106 VDD.n430 37.5148
R15975 VDD.t106 VDD.n471 37.5148
R15976 VDD.n885 VDD.t123 37.5148
R15977 VDD.n910 VDD.t123 37.5148
R15978 VDD.t126 VDD.n689 37.5148
R15979 VDD.t126 VDD.n730 37.5148
R15980 VDD.n1144 VDD.t12 37.5148
R15981 VDD.n1169 VDD.t12 37.5148
R15982 VDD.t51 VDD.n948 37.5148
R15983 VDD.t51 VDD.n989 37.5148
R15984 VDD.n1403 VDD.t111 37.5148
R15985 VDD.n1428 VDD.t111 37.5148
R15986 VDD.t53 VDD.n1207 37.5148
R15987 VDD.t53 VDD.n1248 37.5148
R15988 VDD.n1662 VDD.t147 37.5148
R15989 VDD.n1687 VDD.t147 37.5148
R15990 VDD.t46 VDD.n1466 37.5148
R15991 VDD.t46 VDD.n1507 37.5148
R15992 VDD.n1921 VDD.t22 37.5148
R15993 VDD.n1946 VDD.t22 37.5148
R15994 VDD.t140 VDD.n1725 37.5148
R15995 VDD.t140 VDD.n1766 37.5148
R15996 VDD.n2180 VDD.t156 37.5148
R15997 VDD.n2205 VDD.t156 37.5148
R15998 VDD.t35 VDD.n1984 37.5148
R15999 VDD.t35 VDD.n2025 37.5148
R16000 VDD.n2439 VDD.t213 37.5148
R16001 VDD.n2464 VDD.t213 37.5148
R16002 VDD.t29 VDD.n2243 37.5148
R16003 VDD.t29 VDD.n2284 37.5148
R16004 VDD.n2698 VDD.t72 37.5148
R16005 VDD.n2723 VDD.t72 37.5148
R16006 VDD.t83 VDD.n2502 37.5148
R16007 VDD.t83 VDD.n2543 37.5148
R16008 VDD.n2957 VDD.t57 37.5148
R16009 VDD.n2982 VDD.t57 37.5148
R16010 VDD.t10 VDD.n2761 37.5148
R16011 VDD.t10 VDD.n2802 37.5148
R16012 VDD.n3216 VDD.t48 37.5148
R16013 VDD.n3241 VDD.t48 37.5148
R16014 VDD.t55 VDD.n3020 37.5148
R16015 VDD.t55 VDD.n3061 37.5148
R16016 VDD.n3475 VDD.t135 37.5148
R16017 VDD.n3500 VDD.t135 37.5148
R16018 VDD.t92 VDD.n3279 37.5148
R16019 VDD.t92 VDD.n3320 37.5148
R16020 VDD.n3734 VDD.t24 37.5148
R16021 VDD.n3759 VDD.t24 37.5148
R16022 VDD.t14 VDD.n3538 37.5148
R16023 VDD.t14 VDD.n3579 37.5148
R16024 VDD.n3993 VDD.t199 37.5148
R16025 VDD.n4018 VDD.t199 37.5148
R16026 VDD.t116 VDD.n3797 37.5148
R16027 VDD.t116 VDD.n3838 37.5148
R16028 VDD.n4252 VDD.t8 37.5148
R16029 VDD.n4277 VDD.t8 37.5148
R16030 VDD.t6 VDD.n4056 37.5148
R16031 VDD.t6 VDD.n4097 37.5148
R16032 VDD.n4511 VDD.t76 37.5148
R16033 VDD.n4536 VDD.t76 37.5148
R16034 VDD.t175 VDD.n4315 37.5148
R16035 VDD.t175 VDD.n4356 37.5148
R16036 VDD.n930 VDD 37.1783
R16037 VDD.n266 VDD.n265 37.0005
R16038 VDD.n378 VDD.n266 37.0005
R16039 VDD.n379 VDD.n236 37.0005
R16040 VDD.n379 VDD.n378 37.0005
R16041 VDD.n383 VDD.n183 37.0005
R16042 VDD.n403 VDD.n183 37.0005
R16043 VDD.n383 VDD.n231 37.0005
R16044 VDD.n231 VDD.n182 37.0005
R16045 VDD.n234 VDD.n233 37.0005
R16046 VDD.n233 VDD.n223 37.0005
R16047 VDD.n261 VDD.n260 37.0005
R16048 VDD.n378 VDD.n261 37.0005
R16049 VDD.n257 VDD.n180 37.0005
R16050 VDD.n403 VDD.n180 37.0005
R16051 VDD.n257 VDD.n256 37.0005
R16052 VDD.n256 VDD.n182 37.0005
R16053 VDD.n253 VDD.n252 37.0005
R16054 VDD.n252 VDD.n223 37.0005
R16055 VDD.n305 VDD.n267 37.0005
R16056 VDD.n378 VDD.n267 37.0005
R16057 VDD.n309 VDD.n184 37.0005
R16058 VDD.n403 VDD.n184 37.0005
R16059 VDD.n309 VDD.n298 37.0005
R16060 VDD.n298 VDD.n182 37.0005
R16061 VDD.n301 VDD.n300 37.0005
R16062 VDD.n300 VDD.n223 37.0005
R16063 VDD.n321 VDD.n247 37.0005
R16064 VDD.n378 VDD.n247 37.0005
R16065 VDD.n325 VDD.n179 37.0005
R16066 VDD.n403 VDD.n179 37.0005
R16067 VDD.n325 VDD.n314 37.0005
R16068 VDD.n314 VDD.n182 37.0005
R16069 VDD.n317 VDD.n316 37.0005
R16070 VDD.n316 VDD.n223 37.0005
R16071 VDD.n332 VDD.n328 37.0005
R16072 VDD.n328 VDD.n182 37.0005
R16073 VDD.n330 VDD.n329 37.0005
R16074 VDD.n329 VDD.n223 37.0005
R16075 VDD.n344 VDD.n268 37.0005
R16076 VDD.n378 VDD.n268 37.0005
R16077 VDD.n348 VDD.n185 37.0005
R16078 VDD.n403 VDD.n185 37.0005
R16079 VDD.n348 VDD.n337 37.0005
R16080 VDD.n337 VDD.n182 37.0005
R16081 VDD.n340 VDD.n339 37.0005
R16082 VDD.n339 VDD.n223 37.0005
R16083 VDD.n360 VDD.n246 37.0005
R16084 VDD.n378 VDD.n246 37.0005
R16085 VDD.n364 VDD.n178 37.0005
R16086 VDD.n403 VDD.n178 37.0005
R16087 VDD.n364 VDD.n353 37.0005
R16088 VDD.n353 VDD.n182 37.0005
R16089 VDD.n356 VDD.n355 37.0005
R16090 VDD.n355 VDD.n223 37.0005
R16091 VDD.n371 VDD.n370 37.0005
R16092 VDD.n378 VDD.n371 37.0005
R16093 VDD.n367 VDD.n186 37.0005
R16094 VDD.n403 VDD.n186 37.0005
R16095 VDD.n367 VDD.n277 37.0005
R16096 VDD.n277 VDD.n182 37.0005
R16097 VDD.n274 VDD.n273 37.0005
R16098 VDD.n273 VDD.n223 37.0005
R16099 VDD.n287 VDD.n245 37.0005
R16100 VDD.n378 VDD.n245 37.0005
R16101 VDD.n291 VDD.n177 37.0005
R16102 VDD.n403 VDD.n177 37.0005
R16103 VDD.n291 VDD.n280 37.0005
R16104 VDD.n280 VDD.n182 37.0005
R16105 VDD.n283 VDD.n282 37.0005
R16106 VDD.n282 VDD.n223 37.0005
R16107 VDD.n375 VDD.n374 37.0005
R16108 VDD.n378 VDD.n375 37.0005
R16109 VDD.n405 VDD.n404 37.0005
R16110 VDD.n404 VDD.n403 37.0005
R16111 VDD.n405 VDD.n172 37.0005
R16112 VDD.n182 VDD.n172 37.0005
R16113 VDD.n222 VDD.n221 37.0005
R16114 VDD.n223 VDD.n222 37.0005
R16115 VDD.n244 VDD.n243 37.0005
R16116 VDD.n378 VDD.n244 37.0005
R16117 VDD.n396 VDD.n176 37.0005
R16118 VDD.n403 VDD.n176 37.0005
R16119 VDD.n396 VDD.n395 37.0005
R16120 VDD.n395 VDD.n182 37.0005
R16121 VDD.n197 VDD.n195 37.0005
R16122 VDD.n223 VDD.n195 37.0005
R16123 VDD.n377 VDD.n376 37.0005
R16124 VDD.n378 VDD.n377 37.0005
R16125 VDD.n402 VDD.n401 37.0005
R16126 VDD.n403 VDD.n402 37.0005
R16127 VDD.n391 VDD.n226 37.0005
R16128 VDD.n226 VDD.n223 37.0005
R16129 VDD.n388 VDD.n181 37.0005
R16130 VDD.n403 VDD.n181 37.0005
R16131 VDD.n388 VDD.n225 37.0005
R16132 VDD.n225 VDD.n182 37.0005
R16133 VDD.n514 VDD.n513 37.0005
R16134 VDD.n626 VDD.n514 37.0005
R16135 VDD.n627 VDD.n484 37.0005
R16136 VDD.n627 VDD.n626 37.0005
R16137 VDD.n631 VDD.n431 37.0005
R16138 VDD.n651 VDD.n431 37.0005
R16139 VDD.n631 VDD.n479 37.0005
R16140 VDD.n479 VDD.n430 37.0005
R16141 VDD.n482 VDD.n481 37.0005
R16142 VDD.n481 VDD.n471 37.0005
R16143 VDD.n509 VDD.n508 37.0005
R16144 VDD.n626 VDD.n509 37.0005
R16145 VDD.n505 VDD.n428 37.0005
R16146 VDD.n651 VDD.n428 37.0005
R16147 VDD.n505 VDD.n504 37.0005
R16148 VDD.n504 VDD.n430 37.0005
R16149 VDD.n501 VDD.n500 37.0005
R16150 VDD.n500 VDD.n471 37.0005
R16151 VDD.n553 VDD.n515 37.0005
R16152 VDD.n626 VDD.n515 37.0005
R16153 VDD.n557 VDD.n432 37.0005
R16154 VDD.n651 VDD.n432 37.0005
R16155 VDD.n557 VDD.n546 37.0005
R16156 VDD.n546 VDD.n430 37.0005
R16157 VDD.n549 VDD.n548 37.0005
R16158 VDD.n548 VDD.n471 37.0005
R16159 VDD.n569 VDD.n495 37.0005
R16160 VDD.n626 VDD.n495 37.0005
R16161 VDD.n573 VDD.n427 37.0005
R16162 VDD.n651 VDD.n427 37.0005
R16163 VDD.n573 VDD.n562 37.0005
R16164 VDD.n562 VDD.n430 37.0005
R16165 VDD.n565 VDD.n564 37.0005
R16166 VDD.n564 VDD.n471 37.0005
R16167 VDD.n580 VDD.n576 37.0005
R16168 VDD.n576 VDD.n430 37.0005
R16169 VDD.n578 VDD.n577 37.0005
R16170 VDD.n577 VDD.n471 37.0005
R16171 VDD.n592 VDD.n516 37.0005
R16172 VDD.n626 VDD.n516 37.0005
R16173 VDD.n596 VDD.n433 37.0005
R16174 VDD.n651 VDD.n433 37.0005
R16175 VDD.n596 VDD.n585 37.0005
R16176 VDD.n585 VDD.n430 37.0005
R16177 VDD.n588 VDD.n587 37.0005
R16178 VDD.n587 VDD.n471 37.0005
R16179 VDD.n608 VDD.n494 37.0005
R16180 VDD.n626 VDD.n494 37.0005
R16181 VDD.n612 VDD.n426 37.0005
R16182 VDD.n651 VDD.n426 37.0005
R16183 VDD.n612 VDD.n601 37.0005
R16184 VDD.n601 VDD.n430 37.0005
R16185 VDD.n604 VDD.n603 37.0005
R16186 VDD.n603 VDD.n471 37.0005
R16187 VDD.n619 VDD.n618 37.0005
R16188 VDD.n626 VDD.n619 37.0005
R16189 VDD.n615 VDD.n434 37.0005
R16190 VDD.n651 VDD.n434 37.0005
R16191 VDD.n615 VDD.n525 37.0005
R16192 VDD.n525 VDD.n430 37.0005
R16193 VDD.n522 VDD.n521 37.0005
R16194 VDD.n521 VDD.n471 37.0005
R16195 VDD.n535 VDD.n493 37.0005
R16196 VDD.n626 VDD.n493 37.0005
R16197 VDD.n539 VDD.n425 37.0005
R16198 VDD.n651 VDD.n425 37.0005
R16199 VDD.n539 VDD.n528 37.0005
R16200 VDD.n528 VDD.n430 37.0005
R16201 VDD.n531 VDD.n530 37.0005
R16202 VDD.n530 VDD.n471 37.0005
R16203 VDD.n623 VDD.n622 37.0005
R16204 VDD.n626 VDD.n623 37.0005
R16205 VDD.n653 VDD.n652 37.0005
R16206 VDD.n652 VDD.n651 37.0005
R16207 VDD.n653 VDD.n420 37.0005
R16208 VDD.n430 VDD.n420 37.0005
R16209 VDD.n470 VDD.n469 37.0005
R16210 VDD.n471 VDD.n470 37.0005
R16211 VDD.n492 VDD.n491 37.0005
R16212 VDD.n626 VDD.n492 37.0005
R16213 VDD.n644 VDD.n424 37.0005
R16214 VDD.n651 VDD.n424 37.0005
R16215 VDD.n644 VDD.n643 37.0005
R16216 VDD.n643 VDD.n430 37.0005
R16217 VDD.n445 VDD.n443 37.0005
R16218 VDD.n471 VDD.n443 37.0005
R16219 VDD.n625 VDD.n624 37.0005
R16220 VDD.n626 VDD.n625 37.0005
R16221 VDD.n650 VDD.n649 37.0005
R16222 VDD.n651 VDD.n650 37.0005
R16223 VDD.n639 VDD.n474 37.0005
R16224 VDD.n474 VDD.n471 37.0005
R16225 VDD.n636 VDD.n429 37.0005
R16226 VDD.n651 VDD.n429 37.0005
R16227 VDD.n636 VDD.n473 37.0005
R16228 VDD.n473 VDD.n430 37.0005
R16229 VDD.n773 VDD.n772 37.0005
R16230 VDD.n885 VDD.n773 37.0005
R16231 VDD.n886 VDD.n743 37.0005
R16232 VDD.n886 VDD.n885 37.0005
R16233 VDD.n890 VDD.n690 37.0005
R16234 VDD.n910 VDD.n690 37.0005
R16235 VDD.n890 VDD.n738 37.0005
R16236 VDD.n738 VDD.n689 37.0005
R16237 VDD.n741 VDD.n740 37.0005
R16238 VDD.n740 VDD.n730 37.0005
R16239 VDD.n768 VDD.n767 37.0005
R16240 VDD.n885 VDD.n768 37.0005
R16241 VDD.n764 VDD.n687 37.0005
R16242 VDD.n910 VDD.n687 37.0005
R16243 VDD.n764 VDD.n763 37.0005
R16244 VDD.n763 VDD.n689 37.0005
R16245 VDD.n760 VDD.n759 37.0005
R16246 VDD.n759 VDD.n730 37.0005
R16247 VDD.n812 VDD.n774 37.0005
R16248 VDD.n885 VDD.n774 37.0005
R16249 VDD.n816 VDD.n691 37.0005
R16250 VDD.n910 VDD.n691 37.0005
R16251 VDD.n816 VDD.n805 37.0005
R16252 VDD.n805 VDD.n689 37.0005
R16253 VDD.n808 VDD.n807 37.0005
R16254 VDD.n807 VDD.n730 37.0005
R16255 VDD.n828 VDD.n754 37.0005
R16256 VDD.n885 VDD.n754 37.0005
R16257 VDD.n832 VDD.n686 37.0005
R16258 VDD.n910 VDD.n686 37.0005
R16259 VDD.n832 VDD.n821 37.0005
R16260 VDD.n821 VDD.n689 37.0005
R16261 VDD.n824 VDD.n823 37.0005
R16262 VDD.n823 VDD.n730 37.0005
R16263 VDD.n839 VDD.n835 37.0005
R16264 VDD.n835 VDD.n689 37.0005
R16265 VDD.n837 VDD.n836 37.0005
R16266 VDD.n836 VDD.n730 37.0005
R16267 VDD.n851 VDD.n775 37.0005
R16268 VDD.n885 VDD.n775 37.0005
R16269 VDD.n855 VDD.n692 37.0005
R16270 VDD.n910 VDD.n692 37.0005
R16271 VDD.n855 VDD.n844 37.0005
R16272 VDD.n844 VDD.n689 37.0005
R16273 VDD.n847 VDD.n846 37.0005
R16274 VDD.n846 VDD.n730 37.0005
R16275 VDD.n867 VDD.n753 37.0005
R16276 VDD.n885 VDD.n753 37.0005
R16277 VDD.n871 VDD.n685 37.0005
R16278 VDD.n910 VDD.n685 37.0005
R16279 VDD.n871 VDD.n860 37.0005
R16280 VDD.n860 VDD.n689 37.0005
R16281 VDD.n863 VDD.n862 37.0005
R16282 VDD.n862 VDD.n730 37.0005
R16283 VDD.n878 VDD.n877 37.0005
R16284 VDD.n885 VDD.n878 37.0005
R16285 VDD.n874 VDD.n693 37.0005
R16286 VDD.n910 VDD.n693 37.0005
R16287 VDD.n874 VDD.n784 37.0005
R16288 VDD.n784 VDD.n689 37.0005
R16289 VDD.n781 VDD.n780 37.0005
R16290 VDD.n780 VDD.n730 37.0005
R16291 VDD.n794 VDD.n752 37.0005
R16292 VDD.n885 VDD.n752 37.0005
R16293 VDD.n798 VDD.n684 37.0005
R16294 VDD.n910 VDD.n684 37.0005
R16295 VDD.n798 VDD.n787 37.0005
R16296 VDD.n787 VDD.n689 37.0005
R16297 VDD.n790 VDD.n789 37.0005
R16298 VDD.n789 VDD.n730 37.0005
R16299 VDD.n882 VDD.n881 37.0005
R16300 VDD.n885 VDD.n882 37.0005
R16301 VDD.n912 VDD.n911 37.0005
R16302 VDD.n911 VDD.n910 37.0005
R16303 VDD.n912 VDD.n679 37.0005
R16304 VDD.n689 VDD.n679 37.0005
R16305 VDD.n729 VDD.n728 37.0005
R16306 VDD.n730 VDD.n729 37.0005
R16307 VDD.n751 VDD.n750 37.0005
R16308 VDD.n885 VDD.n751 37.0005
R16309 VDD.n903 VDD.n683 37.0005
R16310 VDD.n910 VDD.n683 37.0005
R16311 VDD.n903 VDD.n902 37.0005
R16312 VDD.n902 VDD.n689 37.0005
R16313 VDD.n704 VDD.n702 37.0005
R16314 VDD.n730 VDD.n702 37.0005
R16315 VDD.n884 VDD.n883 37.0005
R16316 VDD.n885 VDD.n884 37.0005
R16317 VDD.n909 VDD.n908 37.0005
R16318 VDD.n910 VDD.n909 37.0005
R16319 VDD.n898 VDD.n733 37.0005
R16320 VDD.n733 VDD.n730 37.0005
R16321 VDD.n895 VDD.n688 37.0005
R16322 VDD.n910 VDD.n688 37.0005
R16323 VDD.n895 VDD.n732 37.0005
R16324 VDD.n732 VDD.n689 37.0005
R16325 VDD.n1032 VDD.n1031 37.0005
R16326 VDD.n1144 VDD.n1032 37.0005
R16327 VDD.n1145 VDD.n1002 37.0005
R16328 VDD.n1145 VDD.n1144 37.0005
R16329 VDD.n1149 VDD.n949 37.0005
R16330 VDD.n1169 VDD.n949 37.0005
R16331 VDD.n1149 VDD.n997 37.0005
R16332 VDD.n997 VDD.n948 37.0005
R16333 VDD.n1000 VDD.n999 37.0005
R16334 VDD.n999 VDD.n989 37.0005
R16335 VDD.n1027 VDD.n1026 37.0005
R16336 VDD.n1144 VDD.n1027 37.0005
R16337 VDD.n1023 VDD.n946 37.0005
R16338 VDD.n1169 VDD.n946 37.0005
R16339 VDD.n1023 VDD.n1022 37.0005
R16340 VDD.n1022 VDD.n948 37.0005
R16341 VDD.n1019 VDD.n1018 37.0005
R16342 VDD.n1018 VDD.n989 37.0005
R16343 VDD.n1071 VDD.n1033 37.0005
R16344 VDD.n1144 VDD.n1033 37.0005
R16345 VDD.n1075 VDD.n950 37.0005
R16346 VDD.n1169 VDD.n950 37.0005
R16347 VDD.n1075 VDD.n1064 37.0005
R16348 VDD.n1064 VDD.n948 37.0005
R16349 VDD.n1067 VDD.n1066 37.0005
R16350 VDD.n1066 VDD.n989 37.0005
R16351 VDD.n1087 VDD.n1013 37.0005
R16352 VDD.n1144 VDD.n1013 37.0005
R16353 VDD.n1091 VDD.n945 37.0005
R16354 VDD.n1169 VDD.n945 37.0005
R16355 VDD.n1091 VDD.n1080 37.0005
R16356 VDD.n1080 VDD.n948 37.0005
R16357 VDD.n1083 VDD.n1082 37.0005
R16358 VDD.n1082 VDD.n989 37.0005
R16359 VDD.n1098 VDD.n1094 37.0005
R16360 VDD.n1094 VDD.n948 37.0005
R16361 VDD.n1096 VDD.n1095 37.0005
R16362 VDD.n1095 VDD.n989 37.0005
R16363 VDD.n1110 VDD.n1034 37.0005
R16364 VDD.n1144 VDD.n1034 37.0005
R16365 VDD.n1114 VDD.n951 37.0005
R16366 VDD.n1169 VDD.n951 37.0005
R16367 VDD.n1114 VDD.n1103 37.0005
R16368 VDD.n1103 VDD.n948 37.0005
R16369 VDD.n1106 VDD.n1105 37.0005
R16370 VDD.n1105 VDD.n989 37.0005
R16371 VDD.n1126 VDD.n1012 37.0005
R16372 VDD.n1144 VDD.n1012 37.0005
R16373 VDD.n1130 VDD.n944 37.0005
R16374 VDD.n1169 VDD.n944 37.0005
R16375 VDD.n1130 VDD.n1119 37.0005
R16376 VDD.n1119 VDD.n948 37.0005
R16377 VDD.n1122 VDD.n1121 37.0005
R16378 VDD.n1121 VDD.n989 37.0005
R16379 VDD.n1137 VDD.n1136 37.0005
R16380 VDD.n1144 VDD.n1137 37.0005
R16381 VDD.n1133 VDD.n952 37.0005
R16382 VDD.n1169 VDD.n952 37.0005
R16383 VDD.n1133 VDD.n1043 37.0005
R16384 VDD.n1043 VDD.n948 37.0005
R16385 VDD.n1040 VDD.n1039 37.0005
R16386 VDD.n1039 VDD.n989 37.0005
R16387 VDD.n1053 VDD.n1011 37.0005
R16388 VDD.n1144 VDD.n1011 37.0005
R16389 VDD.n1057 VDD.n943 37.0005
R16390 VDD.n1169 VDD.n943 37.0005
R16391 VDD.n1057 VDD.n1046 37.0005
R16392 VDD.n1046 VDD.n948 37.0005
R16393 VDD.n1049 VDD.n1048 37.0005
R16394 VDD.n1048 VDD.n989 37.0005
R16395 VDD.n1141 VDD.n1140 37.0005
R16396 VDD.n1144 VDD.n1141 37.0005
R16397 VDD.n1171 VDD.n1170 37.0005
R16398 VDD.n1170 VDD.n1169 37.0005
R16399 VDD.n1171 VDD.n938 37.0005
R16400 VDD.n948 VDD.n938 37.0005
R16401 VDD.n988 VDD.n987 37.0005
R16402 VDD.n989 VDD.n988 37.0005
R16403 VDD.n1010 VDD.n1009 37.0005
R16404 VDD.n1144 VDD.n1010 37.0005
R16405 VDD.n1162 VDD.n942 37.0005
R16406 VDD.n1169 VDD.n942 37.0005
R16407 VDD.n1162 VDD.n1161 37.0005
R16408 VDD.n1161 VDD.n948 37.0005
R16409 VDD.n963 VDD.n961 37.0005
R16410 VDD.n989 VDD.n961 37.0005
R16411 VDD.n1143 VDD.n1142 37.0005
R16412 VDD.n1144 VDD.n1143 37.0005
R16413 VDD.n1168 VDD.n1167 37.0005
R16414 VDD.n1169 VDD.n1168 37.0005
R16415 VDD.n1157 VDD.n992 37.0005
R16416 VDD.n992 VDD.n989 37.0005
R16417 VDD.n1154 VDD.n947 37.0005
R16418 VDD.n1169 VDD.n947 37.0005
R16419 VDD.n1154 VDD.n991 37.0005
R16420 VDD.n991 VDD.n948 37.0005
R16421 VDD.n1291 VDD.n1290 37.0005
R16422 VDD.n1403 VDD.n1291 37.0005
R16423 VDD.n1404 VDD.n1261 37.0005
R16424 VDD.n1404 VDD.n1403 37.0005
R16425 VDD.n1408 VDD.n1208 37.0005
R16426 VDD.n1428 VDD.n1208 37.0005
R16427 VDD.n1408 VDD.n1256 37.0005
R16428 VDD.n1256 VDD.n1207 37.0005
R16429 VDD.n1259 VDD.n1258 37.0005
R16430 VDD.n1258 VDD.n1248 37.0005
R16431 VDD.n1286 VDD.n1285 37.0005
R16432 VDD.n1403 VDD.n1286 37.0005
R16433 VDD.n1282 VDD.n1205 37.0005
R16434 VDD.n1428 VDD.n1205 37.0005
R16435 VDD.n1282 VDD.n1281 37.0005
R16436 VDD.n1281 VDD.n1207 37.0005
R16437 VDD.n1278 VDD.n1277 37.0005
R16438 VDD.n1277 VDD.n1248 37.0005
R16439 VDD.n1330 VDD.n1292 37.0005
R16440 VDD.n1403 VDD.n1292 37.0005
R16441 VDD.n1334 VDD.n1209 37.0005
R16442 VDD.n1428 VDD.n1209 37.0005
R16443 VDD.n1334 VDD.n1323 37.0005
R16444 VDD.n1323 VDD.n1207 37.0005
R16445 VDD.n1326 VDD.n1325 37.0005
R16446 VDD.n1325 VDD.n1248 37.0005
R16447 VDD.n1346 VDD.n1272 37.0005
R16448 VDD.n1403 VDD.n1272 37.0005
R16449 VDD.n1350 VDD.n1204 37.0005
R16450 VDD.n1428 VDD.n1204 37.0005
R16451 VDD.n1350 VDD.n1339 37.0005
R16452 VDD.n1339 VDD.n1207 37.0005
R16453 VDD.n1342 VDD.n1341 37.0005
R16454 VDD.n1341 VDD.n1248 37.0005
R16455 VDD.n1357 VDD.n1353 37.0005
R16456 VDD.n1353 VDD.n1207 37.0005
R16457 VDD.n1355 VDD.n1354 37.0005
R16458 VDD.n1354 VDD.n1248 37.0005
R16459 VDD.n1369 VDD.n1293 37.0005
R16460 VDD.n1403 VDD.n1293 37.0005
R16461 VDD.n1373 VDD.n1210 37.0005
R16462 VDD.n1428 VDD.n1210 37.0005
R16463 VDD.n1373 VDD.n1362 37.0005
R16464 VDD.n1362 VDD.n1207 37.0005
R16465 VDD.n1365 VDD.n1364 37.0005
R16466 VDD.n1364 VDD.n1248 37.0005
R16467 VDD.n1385 VDD.n1271 37.0005
R16468 VDD.n1403 VDD.n1271 37.0005
R16469 VDD.n1389 VDD.n1203 37.0005
R16470 VDD.n1428 VDD.n1203 37.0005
R16471 VDD.n1389 VDD.n1378 37.0005
R16472 VDD.n1378 VDD.n1207 37.0005
R16473 VDD.n1381 VDD.n1380 37.0005
R16474 VDD.n1380 VDD.n1248 37.0005
R16475 VDD.n1396 VDD.n1395 37.0005
R16476 VDD.n1403 VDD.n1396 37.0005
R16477 VDD.n1392 VDD.n1211 37.0005
R16478 VDD.n1428 VDD.n1211 37.0005
R16479 VDD.n1392 VDD.n1302 37.0005
R16480 VDD.n1302 VDD.n1207 37.0005
R16481 VDD.n1299 VDD.n1298 37.0005
R16482 VDD.n1298 VDD.n1248 37.0005
R16483 VDD.n1312 VDD.n1270 37.0005
R16484 VDD.n1403 VDD.n1270 37.0005
R16485 VDD.n1316 VDD.n1202 37.0005
R16486 VDD.n1428 VDD.n1202 37.0005
R16487 VDD.n1316 VDD.n1305 37.0005
R16488 VDD.n1305 VDD.n1207 37.0005
R16489 VDD.n1308 VDD.n1307 37.0005
R16490 VDD.n1307 VDD.n1248 37.0005
R16491 VDD.n1400 VDD.n1399 37.0005
R16492 VDD.n1403 VDD.n1400 37.0005
R16493 VDD.n1430 VDD.n1429 37.0005
R16494 VDD.n1429 VDD.n1428 37.0005
R16495 VDD.n1430 VDD.n1197 37.0005
R16496 VDD.n1207 VDD.n1197 37.0005
R16497 VDD.n1247 VDD.n1246 37.0005
R16498 VDD.n1248 VDD.n1247 37.0005
R16499 VDD.n1269 VDD.n1268 37.0005
R16500 VDD.n1403 VDD.n1269 37.0005
R16501 VDD.n1421 VDD.n1201 37.0005
R16502 VDD.n1428 VDD.n1201 37.0005
R16503 VDD.n1421 VDD.n1420 37.0005
R16504 VDD.n1420 VDD.n1207 37.0005
R16505 VDD.n1222 VDD.n1220 37.0005
R16506 VDD.n1248 VDD.n1220 37.0005
R16507 VDD.n1402 VDD.n1401 37.0005
R16508 VDD.n1403 VDD.n1402 37.0005
R16509 VDD.n1427 VDD.n1426 37.0005
R16510 VDD.n1428 VDD.n1427 37.0005
R16511 VDD.n1416 VDD.n1251 37.0005
R16512 VDD.n1251 VDD.n1248 37.0005
R16513 VDD.n1413 VDD.n1206 37.0005
R16514 VDD.n1428 VDD.n1206 37.0005
R16515 VDD.n1413 VDD.n1250 37.0005
R16516 VDD.n1250 VDD.n1207 37.0005
R16517 VDD.n1550 VDD.n1549 37.0005
R16518 VDD.n1662 VDD.n1550 37.0005
R16519 VDD.n1663 VDD.n1520 37.0005
R16520 VDD.n1663 VDD.n1662 37.0005
R16521 VDD.n1667 VDD.n1467 37.0005
R16522 VDD.n1687 VDD.n1467 37.0005
R16523 VDD.n1667 VDD.n1515 37.0005
R16524 VDD.n1515 VDD.n1466 37.0005
R16525 VDD.n1518 VDD.n1517 37.0005
R16526 VDD.n1517 VDD.n1507 37.0005
R16527 VDD.n1545 VDD.n1544 37.0005
R16528 VDD.n1662 VDD.n1545 37.0005
R16529 VDD.n1541 VDD.n1464 37.0005
R16530 VDD.n1687 VDD.n1464 37.0005
R16531 VDD.n1541 VDD.n1540 37.0005
R16532 VDD.n1540 VDD.n1466 37.0005
R16533 VDD.n1537 VDD.n1536 37.0005
R16534 VDD.n1536 VDD.n1507 37.0005
R16535 VDD.n1589 VDD.n1551 37.0005
R16536 VDD.n1662 VDD.n1551 37.0005
R16537 VDD.n1593 VDD.n1468 37.0005
R16538 VDD.n1687 VDD.n1468 37.0005
R16539 VDD.n1593 VDD.n1582 37.0005
R16540 VDD.n1582 VDD.n1466 37.0005
R16541 VDD.n1585 VDD.n1584 37.0005
R16542 VDD.n1584 VDD.n1507 37.0005
R16543 VDD.n1605 VDD.n1531 37.0005
R16544 VDD.n1662 VDD.n1531 37.0005
R16545 VDD.n1609 VDD.n1463 37.0005
R16546 VDD.n1687 VDD.n1463 37.0005
R16547 VDD.n1609 VDD.n1598 37.0005
R16548 VDD.n1598 VDD.n1466 37.0005
R16549 VDD.n1601 VDD.n1600 37.0005
R16550 VDD.n1600 VDD.n1507 37.0005
R16551 VDD.n1616 VDD.n1612 37.0005
R16552 VDD.n1612 VDD.n1466 37.0005
R16553 VDD.n1614 VDD.n1613 37.0005
R16554 VDD.n1613 VDD.n1507 37.0005
R16555 VDD.n1628 VDD.n1552 37.0005
R16556 VDD.n1662 VDD.n1552 37.0005
R16557 VDD.n1632 VDD.n1469 37.0005
R16558 VDD.n1687 VDD.n1469 37.0005
R16559 VDD.n1632 VDD.n1621 37.0005
R16560 VDD.n1621 VDD.n1466 37.0005
R16561 VDD.n1624 VDD.n1623 37.0005
R16562 VDD.n1623 VDD.n1507 37.0005
R16563 VDD.n1644 VDD.n1530 37.0005
R16564 VDD.n1662 VDD.n1530 37.0005
R16565 VDD.n1648 VDD.n1462 37.0005
R16566 VDD.n1687 VDD.n1462 37.0005
R16567 VDD.n1648 VDD.n1637 37.0005
R16568 VDD.n1637 VDD.n1466 37.0005
R16569 VDD.n1640 VDD.n1639 37.0005
R16570 VDD.n1639 VDD.n1507 37.0005
R16571 VDD.n1655 VDD.n1654 37.0005
R16572 VDD.n1662 VDD.n1655 37.0005
R16573 VDD.n1651 VDD.n1470 37.0005
R16574 VDD.n1687 VDD.n1470 37.0005
R16575 VDD.n1651 VDD.n1561 37.0005
R16576 VDD.n1561 VDD.n1466 37.0005
R16577 VDD.n1558 VDD.n1557 37.0005
R16578 VDD.n1557 VDD.n1507 37.0005
R16579 VDD.n1571 VDD.n1529 37.0005
R16580 VDD.n1662 VDD.n1529 37.0005
R16581 VDD.n1575 VDD.n1461 37.0005
R16582 VDD.n1687 VDD.n1461 37.0005
R16583 VDD.n1575 VDD.n1564 37.0005
R16584 VDD.n1564 VDD.n1466 37.0005
R16585 VDD.n1567 VDD.n1566 37.0005
R16586 VDD.n1566 VDD.n1507 37.0005
R16587 VDD.n1659 VDD.n1658 37.0005
R16588 VDD.n1662 VDD.n1659 37.0005
R16589 VDD.n1689 VDD.n1688 37.0005
R16590 VDD.n1688 VDD.n1687 37.0005
R16591 VDD.n1689 VDD.n1456 37.0005
R16592 VDD.n1466 VDD.n1456 37.0005
R16593 VDD.n1506 VDD.n1505 37.0005
R16594 VDD.n1507 VDD.n1506 37.0005
R16595 VDD.n1528 VDD.n1527 37.0005
R16596 VDD.n1662 VDD.n1528 37.0005
R16597 VDD.n1680 VDD.n1460 37.0005
R16598 VDD.n1687 VDD.n1460 37.0005
R16599 VDD.n1680 VDD.n1679 37.0005
R16600 VDD.n1679 VDD.n1466 37.0005
R16601 VDD.n1481 VDD.n1479 37.0005
R16602 VDD.n1507 VDD.n1479 37.0005
R16603 VDD.n1661 VDD.n1660 37.0005
R16604 VDD.n1662 VDD.n1661 37.0005
R16605 VDD.n1686 VDD.n1685 37.0005
R16606 VDD.n1687 VDD.n1686 37.0005
R16607 VDD.n1675 VDD.n1510 37.0005
R16608 VDD.n1510 VDD.n1507 37.0005
R16609 VDD.n1672 VDD.n1465 37.0005
R16610 VDD.n1687 VDD.n1465 37.0005
R16611 VDD.n1672 VDD.n1509 37.0005
R16612 VDD.n1509 VDD.n1466 37.0005
R16613 VDD.n1809 VDD.n1808 37.0005
R16614 VDD.n1921 VDD.n1809 37.0005
R16615 VDD.n1922 VDD.n1779 37.0005
R16616 VDD.n1922 VDD.n1921 37.0005
R16617 VDD.n1926 VDD.n1726 37.0005
R16618 VDD.n1946 VDD.n1726 37.0005
R16619 VDD.n1926 VDD.n1774 37.0005
R16620 VDD.n1774 VDD.n1725 37.0005
R16621 VDD.n1777 VDD.n1776 37.0005
R16622 VDD.n1776 VDD.n1766 37.0005
R16623 VDD.n1804 VDD.n1803 37.0005
R16624 VDD.n1921 VDD.n1804 37.0005
R16625 VDD.n1800 VDD.n1723 37.0005
R16626 VDD.n1946 VDD.n1723 37.0005
R16627 VDD.n1800 VDD.n1799 37.0005
R16628 VDD.n1799 VDD.n1725 37.0005
R16629 VDD.n1796 VDD.n1795 37.0005
R16630 VDD.n1795 VDD.n1766 37.0005
R16631 VDD.n1848 VDD.n1810 37.0005
R16632 VDD.n1921 VDD.n1810 37.0005
R16633 VDD.n1852 VDD.n1727 37.0005
R16634 VDD.n1946 VDD.n1727 37.0005
R16635 VDD.n1852 VDD.n1841 37.0005
R16636 VDD.n1841 VDD.n1725 37.0005
R16637 VDD.n1844 VDD.n1843 37.0005
R16638 VDD.n1843 VDD.n1766 37.0005
R16639 VDD.n1864 VDD.n1790 37.0005
R16640 VDD.n1921 VDD.n1790 37.0005
R16641 VDD.n1868 VDD.n1722 37.0005
R16642 VDD.n1946 VDD.n1722 37.0005
R16643 VDD.n1868 VDD.n1857 37.0005
R16644 VDD.n1857 VDD.n1725 37.0005
R16645 VDD.n1860 VDD.n1859 37.0005
R16646 VDD.n1859 VDD.n1766 37.0005
R16647 VDD.n1875 VDD.n1871 37.0005
R16648 VDD.n1871 VDD.n1725 37.0005
R16649 VDD.n1873 VDD.n1872 37.0005
R16650 VDD.n1872 VDD.n1766 37.0005
R16651 VDD.n1887 VDD.n1811 37.0005
R16652 VDD.n1921 VDD.n1811 37.0005
R16653 VDD.n1891 VDD.n1728 37.0005
R16654 VDD.n1946 VDD.n1728 37.0005
R16655 VDD.n1891 VDD.n1880 37.0005
R16656 VDD.n1880 VDD.n1725 37.0005
R16657 VDD.n1883 VDD.n1882 37.0005
R16658 VDD.n1882 VDD.n1766 37.0005
R16659 VDD.n1903 VDD.n1789 37.0005
R16660 VDD.n1921 VDD.n1789 37.0005
R16661 VDD.n1907 VDD.n1721 37.0005
R16662 VDD.n1946 VDD.n1721 37.0005
R16663 VDD.n1907 VDD.n1896 37.0005
R16664 VDD.n1896 VDD.n1725 37.0005
R16665 VDD.n1899 VDD.n1898 37.0005
R16666 VDD.n1898 VDD.n1766 37.0005
R16667 VDD.n1914 VDD.n1913 37.0005
R16668 VDD.n1921 VDD.n1914 37.0005
R16669 VDD.n1910 VDD.n1729 37.0005
R16670 VDD.n1946 VDD.n1729 37.0005
R16671 VDD.n1910 VDD.n1820 37.0005
R16672 VDD.n1820 VDD.n1725 37.0005
R16673 VDD.n1817 VDD.n1816 37.0005
R16674 VDD.n1816 VDD.n1766 37.0005
R16675 VDD.n1830 VDD.n1788 37.0005
R16676 VDD.n1921 VDD.n1788 37.0005
R16677 VDD.n1834 VDD.n1720 37.0005
R16678 VDD.n1946 VDD.n1720 37.0005
R16679 VDD.n1834 VDD.n1823 37.0005
R16680 VDD.n1823 VDD.n1725 37.0005
R16681 VDD.n1826 VDD.n1825 37.0005
R16682 VDD.n1825 VDD.n1766 37.0005
R16683 VDD.n1918 VDD.n1917 37.0005
R16684 VDD.n1921 VDD.n1918 37.0005
R16685 VDD.n1948 VDD.n1947 37.0005
R16686 VDD.n1947 VDD.n1946 37.0005
R16687 VDD.n1948 VDD.n1715 37.0005
R16688 VDD.n1725 VDD.n1715 37.0005
R16689 VDD.n1765 VDD.n1764 37.0005
R16690 VDD.n1766 VDD.n1765 37.0005
R16691 VDD.n1787 VDD.n1786 37.0005
R16692 VDD.n1921 VDD.n1787 37.0005
R16693 VDD.n1939 VDD.n1719 37.0005
R16694 VDD.n1946 VDD.n1719 37.0005
R16695 VDD.n1939 VDD.n1938 37.0005
R16696 VDD.n1938 VDD.n1725 37.0005
R16697 VDD.n1740 VDD.n1738 37.0005
R16698 VDD.n1766 VDD.n1738 37.0005
R16699 VDD.n1920 VDD.n1919 37.0005
R16700 VDD.n1921 VDD.n1920 37.0005
R16701 VDD.n1945 VDD.n1944 37.0005
R16702 VDD.n1946 VDD.n1945 37.0005
R16703 VDD.n1934 VDD.n1769 37.0005
R16704 VDD.n1769 VDD.n1766 37.0005
R16705 VDD.n1931 VDD.n1724 37.0005
R16706 VDD.n1946 VDD.n1724 37.0005
R16707 VDD.n1931 VDD.n1768 37.0005
R16708 VDD.n1768 VDD.n1725 37.0005
R16709 VDD.n2068 VDD.n2067 37.0005
R16710 VDD.n2180 VDD.n2068 37.0005
R16711 VDD.n2181 VDD.n2038 37.0005
R16712 VDD.n2181 VDD.n2180 37.0005
R16713 VDD.n2185 VDD.n1985 37.0005
R16714 VDD.n2205 VDD.n1985 37.0005
R16715 VDD.n2185 VDD.n2033 37.0005
R16716 VDD.n2033 VDD.n1984 37.0005
R16717 VDD.n2036 VDD.n2035 37.0005
R16718 VDD.n2035 VDD.n2025 37.0005
R16719 VDD.n2063 VDD.n2062 37.0005
R16720 VDD.n2180 VDD.n2063 37.0005
R16721 VDD.n2059 VDD.n1982 37.0005
R16722 VDD.n2205 VDD.n1982 37.0005
R16723 VDD.n2059 VDD.n2058 37.0005
R16724 VDD.n2058 VDD.n1984 37.0005
R16725 VDD.n2055 VDD.n2054 37.0005
R16726 VDD.n2054 VDD.n2025 37.0005
R16727 VDD.n2107 VDD.n2069 37.0005
R16728 VDD.n2180 VDD.n2069 37.0005
R16729 VDD.n2111 VDD.n1986 37.0005
R16730 VDD.n2205 VDD.n1986 37.0005
R16731 VDD.n2111 VDD.n2100 37.0005
R16732 VDD.n2100 VDD.n1984 37.0005
R16733 VDD.n2103 VDD.n2102 37.0005
R16734 VDD.n2102 VDD.n2025 37.0005
R16735 VDD.n2123 VDD.n2049 37.0005
R16736 VDD.n2180 VDD.n2049 37.0005
R16737 VDD.n2127 VDD.n1981 37.0005
R16738 VDD.n2205 VDD.n1981 37.0005
R16739 VDD.n2127 VDD.n2116 37.0005
R16740 VDD.n2116 VDD.n1984 37.0005
R16741 VDD.n2119 VDD.n2118 37.0005
R16742 VDD.n2118 VDD.n2025 37.0005
R16743 VDD.n2134 VDD.n2130 37.0005
R16744 VDD.n2130 VDD.n1984 37.0005
R16745 VDD.n2132 VDD.n2131 37.0005
R16746 VDD.n2131 VDD.n2025 37.0005
R16747 VDD.n2146 VDD.n2070 37.0005
R16748 VDD.n2180 VDD.n2070 37.0005
R16749 VDD.n2150 VDD.n1987 37.0005
R16750 VDD.n2205 VDD.n1987 37.0005
R16751 VDD.n2150 VDD.n2139 37.0005
R16752 VDD.n2139 VDD.n1984 37.0005
R16753 VDD.n2142 VDD.n2141 37.0005
R16754 VDD.n2141 VDD.n2025 37.0005
R16755 VDD.n2162 VDD.n2048 37.0005
R16756 VDD.n2180 VDD.n2048 37.0005
R16757 VDD.n2166 VDD.n1980 37.0005
R16758 VDD.n2205 VDD.n1980 37.0005
R16759 VDD.n2166 VDD.n2155 37.0005
R16760 VDD.n2155 VDD.n1984 37.0005
R16761 VDD.n2158 VDD.n2157 37.0005
R16762 VDD.n2157 VDD.n2025 37.0005
R16763 VDD.n2173 VDD.n2172 37.0005
R16764 VDD.n2180 VDD.n2173 37.0005
R16765 VDD.n2169 VDD.n1988 37.0005
R16766 VDD.n2205 VDD.n1988 37.0005
R16767 VDD.n2169 VDD.n2079 37.0005
R16768 VDD.n2079 VDD.n1984 37.0005
R16769 VDD.n2076 VDD.n2075 37.0005
R16770 VDD.n2075 VDD.n2025 37.0005
R16771 VDD.n2089 VDD.n2047 37.0005
R16772 VDD.n2180 VDD.n2047 37.0005
R16773 VDD.n2093 VDD.n1979 37.0005
R16774 VDD.n2205 VDD.n1979 37.0005
R16775 VDD.n2093 VDD.n2082 37.0005
R16776 VDD.n2082 VDD.n1984 37.0005
R16777 VDD.n2085 VDD.n2084 37.0005
R16778 VDD.n2084 VDD.n2025 37.0005
R16779 VDD.n2177 VDD.n2176 37.0005
R16780 VDD.n2180 VDD.n2177 37.0005
R16781 VDD.n2207 VDD.n2206 37.0005
R16782 VDD.n2206 VDD.n2205 37.0005
R16783 VDD.n2207 VDD.n1974 37.0005
R16784 VDD.n1984 VDD.n1974 37.0005
R16785 VDD.n2024 VDD.n2023 37.0005
R16786 VDD.n2025 VDD.n2024 37.0005
R16787 VDD.n2046 VDD.n2045 37.0005
R16788 VDD.n2180 VDD.n2046 37.0005
R16789 VDD.n2198 VDD.n1978 37.0005
R16790 VDD.n2205 VDD.n1978 37.0005
R16791 VDD.n2198 VDD.n2197 37.0005
R16792 VDD.n2197 VDD.n1984 37.0005
R16793 VDD.n1999 VDD.n1997 37.0005
R16794 VDD.n2025 VDD.n1997 37.0005
R16795 VDD.n2179 VDD.n2178 37.0005
R16796 VDD.n2180 VDD.n2179 37.0005
R16797 VDD.n2204 VDD.n2203 37.0005
R16798 VDD.n2205 VDD.n2204 37.0005
R16799 VDD.n2193 VDD.n2028 37.0005
R16800 VDD.n2028 VDD.n2025 37.0005
R16801 VDD.n2190 VDD.n1983 37.0005
R16802 VDD.n2205 VDD.n1983 37.0005
R16803 VDD.n2190 VDD.n2027 37.0005
R16804 VDD.n2027 VDD.n1984 37.0005
R16805 VDD.n2327 VDD.n2326 37.0005
R16806 VDD.n2439 VDD.n2327 37.0005
R16807 VDD.n2440 VDD.n2297 37.0005
R16808 VDD.n2440 VDD.n2439 37.0005
R16809 VDD.n2444 VDD.n2244 37.0005
R16810 VDD.n2464 VDD.n2244 37.0005
R16811 VDD.n2444 VDD.n2292 37.0005
R16812 VDD.n2292 VDD.n2243 37.0005
R16813 VDD.n2295 VDD.n2294 37.0005
R16814 VDD.n2294 VDD.n2284 37.0005
R16815 VDD.n2322 VDD.n2321 37.0005
R16816 VDD.n2439 VDD.n2322 37.0005
R16817 VDD.n2318 VDD.n2241 37.0005
R16818 VDD.n2464 VDD.n2241 37.0005
R16819 VDD.n2318 VDD.n2317 37.0005
R16820 VDD.n2317 VDD.n2243 37.0005
R16821 VDD.n2314 VDD.n2313 37.0005
R16822 VDD.n2313 VDD.n2284 37.0005
R16823 VDD.n2366 VDD.n2328 37.0005
R16824 VDD.n2439 VDD.n2328 37.0005
R16825 VDD.n2370 VDD.n2245 37.0005
R16826 VDD.n2464 VDD.n2245 37.0005
R16827 VDD.n2370 VDD.n2359 37.0005
R16828 VDD.n2359 VDD.n2243 37.0005
R16829 VDD.n2362 VDD.n2361 37.0005
R16830 VDD.n2361 VDD.n2284 37.0005
R16831 VDD.n2382 VDD.n2308 37.0005
R16832 VDD.n2439 VDD.n2308 37.0005
R16833 VDD.n2386 VDD.n2240 37.0005
R16834 VDD.n2464 VDD.n2240 37.0005
R16835 VDD.n2386 VDD.n2375 37.0005
R16836 VDD.n2375 VDD.n2243 37.0005
R16837 VDD.n2378 VDD.n2377 37.0005
R16838 VDD.n2377 VDD.n2284 37.0005
R16839 VDD.n2393 VDD.n2389 37.0005
R16840 VDD.n2389 VDD.n2243 37.0005
R16841 VDD.n2391 VDD.n2390 37.0005
R16842 VDD.n2390 VDD.n2284 37.0005
R16843 VDD.n2405 VDD.n2329 37.0005
R16844 VDD.n2439 VDD.n2329 37.0005
R16845 VDD.n2409 VDD.n2246 37.0005
R16846 VDD.n2464 VDD.n2246 37.0005
R16847 VDD.n2409 VDD.n2398 37.0005
R16848 VDD.n2398 VDD.n2243 37.0005
R16849 VDD.n2401 VDD.n2400 37.0005
R16850 VDD.n2400 VDD.n2284 37.0005
R16851 VDD.n2421 VDD.n2307 37.0005
R16852 VDD.n2439 VDD.n2307 37.0005
R16853 VDD.n2425 VDD.n2239 37.0005
R16854 VDD.n2464 VDD.n2239 37.0005
R16855 VDD.n2425 VDD.n2414 37.0005
R16856 VDD.n2414 VDD.n2243 37.0005
R16857 VDD.n2417 VDD.n2416 37.0005
R16858 VDD.n2416 VDD.n2284 37.0005
R16859 VDD.n2432 VDD.n2431 37.0005
R16860 VDD.n2439 VDD.n2432 37.0005
R16861 VDD.n2428 VDD.n2247 37.0005
R16862 VDD.n2464 VDD.n2247 37.0005
R16863 VDD.n2428 VDD.n2338 37.0005
R16864 VDD.n2338 VDD.n2243 37.0005
R16865 VDD.n2335 VDD.n2334 37.0005
R16866 VDD.n2334 VDD.n2284 37.0005
R16867 VDD.n2348 VDD.n2306 37.0005
R16868 VDD.n2439 VDD.n2306 37.0005
R16869 VDD.n2352 VDD.n2238 37.0005
R16870 VDD.n2464 VDD.n2238 37.0005
R16871 VDD.n2352 VDD.n2341 37.0005
R16872 VDD.n2341 VDD.n2243 37.0005
R16873 VDD.n2344 VDD.n2343 37.0005
R16874 VDD.n2343 VDD.n2284 37.0005
R16875 VDD.n2436 VDD.n2435 37.0005
R16876 VDD.n2439 VDD.n2436 37.0005
R16877 VDD.n2466 VDD.n2465 37.0005
R16878 VDD.n2465 VDD.n2464 37.0005
R16879 VDD.n2466 VDD.n2233 37.0005
R16880 VDD.n2243 VDD.n2233 37.0005
R16881 VDD.n2283 VDD.n2282 37.0005
R16882 VDD.n2284 VDD.n2283 37.0005
R16883 VDD.n2305 VDD.n2304 37.0005
R16884 VDD.n2439 VDD.n2305 37.0005
R16885 VDD.n2457 VDD.n2237 37.0005
R16886 VDD.n2464 VDD.n2237 37.0005
R16887 VDD.n2457 VDD.n2456 37.0005
R16888 VDD.n2456 VDD.n2243 37.0005
R16889 VDD.n2258 VDD.n2256 37.0005
R16890 VDD.n2284 VDD.n2256 37.0005
R16891 VDD.n2438 VDD.n2437 37.0005
R16892 VDD.n2439 VDD.n2438 37.0005
R16893 VDD.n2463 VDD.n2462 37.0005
R16894 VDD.n2464 VDD.n2463 37.0005
R16895 VDD.n2452 VDD.n2287 37.0005
R16896 VDD.n2287 VDD.n2284 37.0005
R16897 VDD.n2449 VDD.n2242 37.0005
R16898 VDD.n2464 VDD.n2242 37.0005
R16899 VDD.n2449 VDD.n2286 37.0005
R16900 VDD.n2286 VDD.n2243 37.0005
R16901 VDD.n2586 VDD.n2585 37.0005
R16902 VDD.n2698 VDD.n2586 37.0005
R16903 VDD.n2699 VDD.n2556 37.0005
R16904 VDD.n2699 VDD.n2698 37.0005
R16905 VDD.n2703 VDD.n2503 37.0005
R16906 VDD.n2723 VDD.n2503 37.0005
R16907 VDD.n2703 VDD.n2551 37.0005
R16908 VDD.n2551 VDD.n2502 37.0005
R16909 VDD.n2554 VDD.n2553 37.0005
R16910 VDD.n2553 VDD.n2543 37.0005
R16911 VDD.n2581 VDD.n2580 37.0005
R16912 VDD.n2698 VDD.n2581 37.0005
R16913 VDD.n2577 VDD.n2500 37.0005
R16914 VDD.n2723 VDD.n2500 37.0005
R16915 VDD.n2577 VDD.n2576 37.0005
R16916 VDD.n2576 VDD.n2502 37.0005
R16917 VDD.n2573 VDD.n2572 37.0005
R16918 VDD.n2572 VDD.n2543 37.0005
R16919 VDD.n2625 VDD.n2587 37.0005
R16920 VDD.n2698 VDD.n2587 37.0005
R16921 VDD.n2629 VDD.n2504 37.0005
R16922 VDD.n2723 VDD.n2504 37.0005
R16923 VDD.n2629 VDD.n2618 37.0005
R16924 VDD.n2618 VDD.n2502 37.0005
R16925 VDD.n2621 VDD.n2620 37.0005
R16926 VDD.n2620 VDD.n2543 37.0005
R16927 VDD.n2641 VDD.n2567 37.0005
R16928 VDD.n2698 VDD.n2567 37.0005
R16929 VDD.n2645 VDD.n2499 37.0005
R16930 VDD.n2723 VDD.n2499 37.0005
R16931 VDD.n2645 VDD.n2634 37.0005
R16932 VDD.n2634 VDD.n2502 37.0005
R16933 VDD.n2637 VDD.n2636 37.0005
R16934 VDD.n2636 VDD.n2543 37.0005
R16935 VDD.n2652 VDD.n2648 37.0005
R16936 VDD.n2648 VDD.n2502 37.0005
R16937 VDD.n2650 VDD.n2649 37.0005
R16938 VDD.n2649 VDD.n2543 37.0005
R16939 VDD.n2664 VDD.n2588 37.0005
R16940 VDD.n2698 VDD.n2588 37.0005
R16941 VDD.n2668 VDD.n2505 37.0005
R16942 VDD.n2723 VDD.n2505 37.0005
R16943 VDD.n2668 VDD.n2657 37.0005
R16944 VDD.n2657 VDD.n2502 37.0005
R16945 VDD.n2660 VDD.n2659 37.0005
R16946 VDD.n2659 VDD.n2543 37.0005
R16947 VDD.n2680 VDD.n2566 37.0005
R16948 VDD.n2698 VDD.n2566 37.0005
R16949 VDD.n2684 VDD.n2498 37.0005
R16950 VDD.n2723 VDD.n2498 37.0005
R16951 VDD.n2684 VDD.n2673 37.0005
R16952 VDD.n2673 VDD.n2502 37.0005
R16953 VDD.n2676 VDD.n2675 37.0005
R16954 VDD.n2675 VDD.n2543 37.0005
R16955 VDD.n2691 VDD.n2690 37.0005
R16956 VDD.n2698 VDD.n2691 37.0005
R16957 VDD.n2687 VDD.n2506 37.0005
R16958 VDD.n2723 VDD.n2506 37.0005
R16959 VDD.n2687 VDD.n2597 37.0005
R16960 VDD.n2597 VDD.n2502 37.0005
R16961 VDD.n2594 VDD.n2593 37.0005
R16962 VDD.n2593 VDD.n2543 37.0005
R16963 VDD.n2607 VDD.n2565 37.0005
R16964 VDD.n2698 VDD.n2565 37.0005
R16965 VDD.n2611 VDD.n2497 37.0005
R16966 VDD.n2723 VDD.n2497 37.0005
R16967 VDD.n2611 VDD.n2600 37.0005
R16968 VDD.n2600 VDD.n2502 37.0005
R16969 VDD.n2603 VDD.n2602 37.0005
R16970 VDD.n2602 VDD.n2543 37.0005
R16971 VDD.n2695 VDD.n2694 37.0005
R16972 VDD.n2698 VDD.n2695 37.0005
R16973 VDD.n2725 VDD.n2724 37.0005
R16974 VDD.n2724 VDD.n2723 37.0005
R16975 VDD.n2725 VDD.n2492 37.0005
R16976 VDD.n2502 VDD.n2492 37.0005
R16977 VDD.n2542 VDD.n2541 37.0005
R16978 VDD.n2543 VDD.n2542 37.0005
R16979 VDD.n2564 VDD.n2563 37.0005
R16980 VDD.n2698 VDD.n2564 37.0005
R16981 VDD.n2716 VDD.n2496 37.0005
R16982 VDD.n2723 VDD.n2496 37.0005
R16983 VDD.n2716 VDD.n2715 37.0005
R16984 VDD.n2715 VDD.n2502 37.0005
R16985 VDD.n2517 VDD.n2515 37.0005
R16986 VDD.n2543 VDD.n2515 37.0005
R16987 VDD.n2697 VDD.n2696 37.0005
R16988 VDD.n2698 VDD.n2697 37.0005
R16989 VDD.n2722 VDD.n2721 37.0005
R16990 VDD.n2723 VDD.n2722 37.0005
R16991 VDD.n2711 VDD.n2546 37.0005
R16992 VDD.n2546 VDD.n2543 37.0005
R16993 VDD.n2708 VDD.n2501 37.0005
R16994 VDD.n2723 VDD.n2501 37.0005
R16995 VDD.n2708 VDD.n2545 37.0005
R16996 VDD.n2545 VDD.n2502 37.0005
R16997 VDD.n2845 VDD.n2844 37.0005
R16998 VDD.n2957 VDD.n2845 37.0005
R16999 VDD.n2958 VDD.n2815 37.0005
R17000 VDD.n2958 VDD.n2957 37.0005
R17001 VDD.n2962 VDD.n2762 37.0005
R17002 VDD.n2982 VDD.n2762 37.0005
R17003 VDD.n2962 VDD.n2810 37.0005
R17004 VDD.n2810 VDD.n2761 37.0005
R17005 VDD.n2813 VDD.n2812 37.0005
R17006 VDD.n2812 VDD.n2802 37.0005
R17007 VDD.n2840 VDD.n2839 37.0005
R17008 VDD.n2957 VDD.n2840 37.0005
R17009 VDD.n2836 VDD.n2759 37.0005
R17010 VDD.n2982 VDD.n2759 37.0005
R17011 VDD.n2836 VDD.n2835 37.0005
R17012 VDD.n2835 VDD.n2761 37.0005
R17013 VDD.n2832 VDD.n2831 37.0005
R17014 VDD.n2831 VDD.n2802 37.0005
R17015 VDD.n2884 VDD.n2846 37.0005
R17016 VDD.n2957 VDD.n2846 37.0005
R17017 VDD.n2888 VDD.n2763 37.0005
R17018 VDD.n2982 VDD.n2763 37.0005
R17019 VDD.n2888 VDD.n2877 37.0005
R17020 VDD.n2877 VDD.n2761 37.0005
R17021 VDD.n2880 VDD.n2879 37.0005
R17022 VDD.n2879 VDD.n2802 37.0005
R17023 VDD.n2900 VDD.n2826 37.0005
R17024 VDD.n2957 VDD.n2826 37.0005
R17025 VDD.n2904 VDD.n2758 37.0005
R17026 VDD.n2982 VDD.n2758 37.0005
R17027 VDD.n2904 VDD.n2893 37.0005
R17028 VDD.n2893 VDD.n2761 37.0005
R17029 VDD.n2896 VDD.n2895 37.0005
R17030 VDD.n2895 VDD.n2802 37.0005
R17031 VDD.n2911 VDD.n2907 37.0005
R17032 VDD.n2907 VDD.n2761 37.0005
R17033 VDD.n2909 VDD.n2908 37.0005
R17034 VDD.n2908 VDD.n2802 37.0005
R17035 VDD.n2923 VDD.n2847 37.0005
R17036 VDD.n2957 VDD.n2847 37.0005
R17037 VDD.n2927 VDD.n2764 37.0005
R17038 VDD.n2982 VDD.n2764 37.0005
R17039 VDD.n2927 VDD.n2916 37.0005
R17040 VDD.n2916 VDD.n2761 37.0005
R17041 VDD.n2919 VDD.n2918 37.0005
R17042 VDD.n2918 VDD.n2802 37.0005
R17043 VDD.n2939 VDD.n2825 37.0005
R17044 VDD.n2957 VDD.n2825 37.0005
R17045 VDD.n2943 VDD.n2757 37.0005
R17046 VDD.n2982 VDD.n2757 37.0005
R17047 VDD.n2943 VDD.n2932 37.0005
R17048 VDD.n2932 VDD.n2761 37.0005
R17049 VDD.n2935 VDD.n2934 37.0005
R17050 VDD.n2934 VDD.n2802 37.0005
R17051 VDD.n2950 VDD.n2949 37.0005
R17052 VDD.n2957 VDD.n2950 37.0005
R17053 VDD.n2946 VDD.n2765 37.0005
R17054 VDD.n2982 VDD.n2765 37.0005
R17055 VDD.n2946 VDD.n2856 37.0005
R17056 VDD.n2856 VDD.n2761 37.0005
R17057 VDD.n2853 VDD.n2852 37.0005
R17058 VDD.n2852 VDD.n2802 37.0005
R17059 VDD.n2866 VDD.n2824 37.0005
R17060 VDD.n2957 VDD.n2824 37.0005
R17061 VDD.n2870 VDD.n2756 37.0005
R17062 VDD.n2982 VDD.n2756 37.0005
R17063 VDD.n2870 VDD.n2859 37.0005
R17064 VDD.n2859 VDD.n2761 37.0005
R17065 VDD.n2862 VDD.n2861 37.0005
R17066 VDD.n2861 VDD.n2802 37.0005
R17067 VDD.n2954 VDD.n2953 37.0005
R17068 VDD.n2957 VDD.n2954 37.0005
R17069 VDD.n2984 VDD.n2983 37.0005
R17070 VDD.n2983 VDD.n2982 37.0005
R17071 VDD.n2984 VDD.n2751 37.0005
R17072 VDD.n2761 VDD.n2751 37.0005
R17073 VDD.n2801 VDD.n2800 37.0005
R17074 VDD.n2802 VDD.n2801 37.0005
R17075 VDD.n2823 VDD.n2822 37.0005
R17076 VDD.n2957 VDD.n2823 37.0005
R17077 VDD.n2975 VDD.n2755 37.0005
R17078 VDD.n2982 VDD.n2755 37.0005
R17079 VDD.n2975 VDD.n2974 37.0005
R17080 VDD.n2974 VDD.n2761 37.0005
R17081 VDD.n2776 VDD.n2774 37.0005
R17082 VDD.n2802 VDD.n2774 37.0005
R17083 VDD.n2956 VDD.n2955 37.0005
R17084 VDD.n2957 VDD.n2956 37.0005
R17085 VDD.n2981 VDD.n2980 37.0005
R17086 VDD.n2982 VDD.n2981 37.0005
R17087 VDD.n2970 VDD.n2805 37.0005
R17088 VDD.n2805 VDD.n2802 37.0005
R17089 VDD.n2967 VDD.n2760 37.0005
R17090 VDD.n2982 VDD.n2760 37.0005
R17091 VDD.n2967 VDD.n2804 37.0005
R17092 VDD.n2804 VDD.n2761 37.0005
R17093 VDD.n3104 VDD.n3103 37.0005
R17094 VDD.n3216 VDD.n3104 37.0005
R17095 VDD.n3217 VDD.n3074 37.0005
R17096 VDD.n3217 VDD.n3216 37.0005
R17097 VDD.n3221 VDD.n3021 37.0005
R17098 VDD.n3241 VDD.n3021 37.0005
R17099 VDD.n3221 VDD.n3069 37.0005
R17100 VDD.n3069 VDD.n3020 37.0005
R17101 VDD.n3072 VDD.n3071 37.0005
R17102 VDD.n3071 VDD.n3061 37.0005
R17103 VDD.n3099 VDD.n3098 37.0005
R17104 VDD.n3216 VDD.n3099 37.0005
R17105 VDD.n3095 VDD.n3018 37.0005
R17106 VDD.n3241 VDD.n3018 37.0005
R17107 VDD.n3095 VDD.n3094 37.0005
R17108 VDD.n3094 VDD.n3020 37.0005
R17109 VDD.n3091 VDD.n3090 37.0005
R17110 VDD.n3090 VDD.n3061 37.0005
R17111 VDD.n3143 VDD.n3105 37.0005
R17112 VDD.n3216 VDD.n3105 37.0005
R17113 VDD.n3147 VDD.n3022 37.0005
R17114 VDD.n3241 VDD.n3022 37.0005
R17115 VDD.n3147 VDD.n3136 37.0005
R17116 VDD.n3136 VDD.n3020 37.0005
R17117 VDD.n3139 VDD.n3138 37.0005
R17118 VDD.n3138 VDD.n3061 37.0005
R17119 VDD.n3159 VDD.n3085 37.0005
R17120 VDD.n3216 VDD.n3085 37.0005
R17121 VDD.n3163 VDD.n3017 37.0005
R17122 VDD.n3241 VDD.n3017 37.0005
R17123 VDD.n3163 VDD.n3152 37.0005
R17124 VDD.n3152 VDD.n3020 37.0005
R17125 VDD.n3155 VDD.n3154 37.0005
R17126 VDD.n3154 VDD.n3061 37.0005
R17127 VDD.n3170 VDD.n3166 37.0005
R17128 VDD.n3166 VDD.n3020 37.0005
R17129 VDD.n3168 VDD.n3167 37.0005
R17130 VDD.n3167 VDD.n3061 37.0005
R17131 VDD.n3182 VDD.n3106 37.0005
R17132 VDD.n3216 VDD.n3106 37.0005
R17133 VDD.n3186 VDD.n3023 37.0005
R17134 VDD.n3241 VDD.n3023 37.0005
R17135 VDD.n3186 VDD.n3175 37.0005
R17136 VDD.n3175 VDD.n3020 37.0005
R17137 VDD.n3178 VDD.n3177 37.0005
R17138 VDD.n3177 VDD.n3061 37.0005
R17139 VDD.n3198 VDD.n3084 37.0005
R17140 VDD.n3216 VDD.n3084 37.0005
R17141 VDD.n3202 VDD.n3016 37.0005
R17142 VDD.n3241 VDD.n3016 37.0005
R17143 VDD.n3202 VDD.n3191 37.0005
R17144 VDD.n3191 VDD.n3020 37.0005
R17145 VDD.n3194 VDD.n3193 37.0005
R17146 VDD.n3193 VDD.n3061 37.0005
R17147 VDD.n3209 VDD.n3208 37.0005
R17148 VDD.n3216 VDD.n3209 37.0005
R17149 VDD.n3205 VDD.n3024 37.0005
R17150 VDD.n3241 VDD.n3024 37.0005
R17151 VDD.n3205 VDD.n3115 37.0005
R17152 VDD.n3115 VDD.n3020 37.0005
R17153 VDD.n3112 VDD.n3111 37.0005
R17154 VDD.n3111 VDD.n3061 37.0005
R17155 VDD.n3125 VDD.n3083 37.0005
R17156 VDD.n3216 VDD.n3083 37.0005
R17157 VDD.n3129 VDD.n3015 37.0005
R17158 VDD.n3241 VDD.n3015 37.0005
R17159 VDD.n3129 VDD.n3118 37.0005
R17160 VDD.n3118 VDD.n3020 37.0005
R17161 VDD.n3121 VDD.n3120 37.0005
R17162 VDD.n3120 VDD.n3061 37.0005
R17163 VDD.n3213 VDD.n3212 37.0005
R17164 VDD.n3216 VDD.n3213 37.0005
R17165 VDD.n3243 VDD.n3242 37.0005
R17166 VDD.n3242 VDD.n3241 37.0005
R17167 VDD.n3243 VDD.n3010 37.0005
R17168 VDD.n3020 VDD.n3010 37.0005
R17169 VDD.n3060 VDD.n3059 37.0005
R17170 VDD.n3061 VDD.n3060 37.0005
R17171 VDD.n3082 VDD.n3081 37.0005
R17172 VDD.n3216 VDD.n3082 37.0005
R17173 VDD.n3234 VDD.n3014 37.0005
R17174 VDD.n3241 VDD.n3014 37.0005
R17175 VDD.n3234 VDD.n3233 37.0005
R17176 VDD.n3233 VDD.n3020 37.0005
R17177 VDD.n3035 VDD.n3033 37.0005
R17178 VDD.n3061 VDD.n3033 37.0005
R17179 VDD.n3215 VDD.n3214 37.0005
R17180 VDD.n3216 VDD.n3215 37.0005
R17181 VDD.n3240 VDD.n3239 37.0005
R17182 VDD.n3241 VDD.n3240 37.0005
R17183 VDD.n3229 VDD.n3064 37.0005
R17184 VDD.n3064 VDD.n3061 37.0005
R17185 VDD.n3226 VDD.n3019 37.0005
R17186 VDD.n3241 VDD.n3019 37.0005
R17187 VDD.n3226 VDD.n3063 37.0005
R17188 VDD.n3063 VDD.n3020 37.0005
R17189 VDD.n3363 VDD.n3362 37.0005
R17190 VDD.n3475 VDD.n3363 37.0005
R17191 VDD.n3476 VDD.n3333 37.0005
R17192 VDD.n3476 VDD.n3475 37.0005
R17193 VDD.n3480 VDD.n3280 37.0005
R17194 VDD.n3500 VDD.n3280 37.0005
R17195 VDD.n3480 VDD.n3328 37.0005
R17196 VDD.n3328 VDD.n3279 37.0005
R17197 VDD.n3331 VDD.n3330 37.0005
R17198 VDD.n3330 VDD.n3320 37.0005
R17199 VDD.n3358 VDD.n3357 37.0005
R17200 VDD.n3475 VDD.n3358 37.0005
R17201 VDD.n3354 VDD.n3277 37.0005
R17202 VDD.n3500 VDD.n3277 37.0005
R17203 VDD.n3354 VDD.n3353 37.0005
R17204 VDD.n3353 VDD.n3279 37.0005
R17205 VDD.n3350 VDD.n3349 37.0005
R17206 VDD.n3349 VDD.n3320 37.0005
R17207 VDD.n3402 VDD.n3364 37.0005
R17208 VDD.n3475 VDD.n3364 37.0005
R17209 VDD.n3406 VDD.n3281 37.0005
R17210 VDD.n3500 VDD.n3281 37.0005
R17211 VDD.n3406 VDD.n3395 37.0005
R17212 VDD.n3395 VDD.n3279 37.0005
R17213 VDD.n3398 VDD.n3397 37.0005
R17214 VDD.n3397 VDD.n3320 37.0005
R17215 VDD.n3418 VDD.n3344 37.0005
R17216 VDD.n3475 VDD.n3344 37.0005
R17217 VDD.n3422 VDD.n3276 37.0005
R17218 VDD.n3500 VDD.n3276 37.0005
R17219 VDD.n3422 VDD.n3411 37.0005
R17220 VDD.n3411 VDD.n3279 37.0005
R17221 VDD.n3414 VDD.n3413 37.0005
R17222 VDD.n3413 VDD.n3320 37.0005
R17223 VDD.n3429 VDD.n3425 37.0005
R17224 VDD.n3425 VDD.n3279 37.0005
R17225 VDD.n3427 VDD.n3426 37.0005
R17226 VDD.n3426 VDD.n3320 37.0005
R17227 VDD.n3441 VDD.n3365 37.0005
R17228 VDD.n3475 VDD.n3365 37.0005
R17229 VDD.n3445 VDD.n3282 37.0005
R17230 VDD.n3500 VDD.n3282 37.0005
R17231 VDD.n3445 VDD.n3434 37.0005
R17232 VDD.n3434 VDD.n3279 37.0005
R17233 VDD.n3437 VDD.n3436 37.0005
R17234 VDD.n3436 VDD.n3320 37.0005
R17235 VDD.n3457 VDD.n3343 37.0005
R17236 VDD.n3475 VDD.n3343 37.0005
R17237 VDD.n3461 VDD.n3275 37.0005
R17238 VDD.n3500 VDD.n3275 37.0005
R17239 VDD.n3461 VDD.n3450 37.0005
R17240 VDD.n3450 VDD.n3279 37.0005
R17241 VDD.n3453 VDD.n3452 37.0005
R17242 VDD.n3452 VDD.n3320 37.0005
R17243 VDD.n3468 VDD.n3467 37.0005
R17244 VDD.n3475 VDD.n3468 37.0005
R17245 VDD.n3464 VDD.n3283 37.0005
R17246 VDD.n3500 VDD.n3283 37.0005
R17247 VDD.n3464 VDD.n3374 37.0005
R17248 VDD.n3374 VDD.n3279 37.0005
R17249 VDD.n3371 VDD.n3370 37.0005
R17250 VDD.n3370 VDD.n3320 37.0005
R17251 VDD.n3384 VDD.n3342 37.0005
R17252 VDD.n3475 VDD.n3342 37.0005
R17253 VDD.n3388 VDD.n3274 37.0005
R17254 VDD.n3500 VDD.n3274 37.0005
R17255 VDD.n3388 VDD.n3377 37.0005
R17256 VDD.n3377 VDD.n3279 37.0005
R17257 VDD.n3380 VDD.n3379 37.0005
R17258 VDD.n3379 VDD.n3320 37.0005
R17259 VDD.n3472 VDD.n3471 37.0005
R17260 VDD.n3475 VDD.n3472 37.0005
R17261 VDD.n3502 VDD.n3501 37.0005
R17262 VDD.n3501 VDD.n3500 37.0005
R17263 VDD.n3502 VDD.n3269 37.0005
R17264 VDD.n3279 VDD.n3269 37.0005
R17265 VDD.n3319 VDD.n3318 37.0005
R17266 VDD.n3320 VDD.n3319 37.0005
R17267 VDD.n3341 VDD.n3340 37.0005
R17268 VDD.n3475 VDD.n3341 37.0005
R17269 VDD.n3493 VDD.n3273 37.0005
R17270 VDD.n3500 VDD.n3273 37.0005
R17271 VDD.n3493 VDD.n3492 37.0005
R17272 VDD.n3492 VDD.n3279 37.0005
R17273 VDD.n3294 VDD.n3292 37.0005
R17274 VDD.n3320 VDD.n3292 37.0005
R17275 VDD.n3474 VDD.n3473 37.0005
R17276 VDD.n3475 VDD.n3474 37.0005
R17277 VDD.n3499 VDD.n3498 37.0005
R17278 VDD.n3500 VDD.n3499 37.0005
R17279 VDD.n3488 VDD.n3323 37.0005
R17280 VDD.n3323 VDD.n3320 37.0005
R17281 VDD.n3485 VDD.n3278 37.0005
R17282 VDD.n3500 VDD.n3278 37.0005
R17283 VDD.n3485 VDD.n3322 37.0005
R17284 VDD.n3322 VDD.n3279 37.0005
R17285 VDD.n3622 VDD.n3621 37.0005
R17286 VDD.n3734 VDD.n3622 37.0005
R17287 VDD.n3735 VDD.n3592 37.0005
R17288 VDD.n3735 VDD.n3734 37.0005
R17289 VDD.n3739 VDD.n3539 37.0005
R17290 VDD.n3759 VDD.n3539 37.0005
R17291 VDD.n3739 VDD.n3587 37.0005
R17292 VDD.n3587 VDD.n3538 37.0005
R17293 VDD.n3590 VDD.n3589 37.0005
R17294 VDD.n3589 VDD.n3579 37.0005
R17295 VDD.n3617 VDD.n3616 37.0005
R17296 VDD.n3734 VDD.n3617 37.0005
R17297 VDD.n3613 VDD.n3536 37.0005
R17298 VDD.n3759 VDD.n3536 37.0005
R17299 VDD.n3613 VDD.n3612 37.0005
R17300 VDD.n3612 VDD.n3538 37.0005
R17301 VDD.n3609 VDD.n3608 37.0005
R17302 VDD.n3608 VDD.n3579 37.0005
R17303 VDD.n3661 VDD.n3623 37.0005
R17304 VDD.n3734 VDD.n3623 37.0005
R17305 VDD.n3665 VDD.n3540 37.0005
R17306 VDD.n3759 VDD.n3540 37.0005
R17307 VDD.n3665 VDD.n3654 37.0005
R17308 VDD.n3654 VDD.n3538 37.0005
R17309 VDD.n3657 VDD.n3656 37.0005
R17310 VDD.n3656 VDD.n3579 37.0005
R17311 VDD.n3677 VDD.n3603 37.0005
R17312 VDD.n3734 VDD.n3603 37.0005
R17313 VDD.n3681 VDD.n3535 37.0005
R17314 VDD.n3759 VDD.n3535 37.0005
R17315 VDD.n3681 VDD.n3670 37.0005
R17316 VDD.n3670 VDD.n3538 37.0005
R17317 VDD.n3673 VDD.n3672 37.0005
R17318 VDD.n3672 VDD.n3579 37.0005
R17319 VDD.n3688 VDD.n3684 37.0005
R17320 VDD.n3684 VDD.n3538 37.0005
R17321 VDD.n3686 VDD.n3685 37.0005
R17322 VDD.n3685 VDD.n3579 37.0005
R17323 VDD.n3700 VDD.n3624 37.0005
R17324 VDD.n3734 VDD.n3624 37.0005
R17325 VDD.n3704 VDD.n3541 37.0005
R17326 VDD.n3759 VDD.n3541 37.0005
R17327 VDD.n3704 VDD.n3693 37.0005
R17328 VDD.n3693 VDD.n3538 37.0005
R17329 VDD.n3696 VDD.n3695 37.0005
R17330 VDD.n3695 VDD.n3579 37.0005
R17331 VDD.n3716 VDD.n3602 37.0005
R17332 VDD.n3734 VDD.n3602 37.0005
R17333 VDD.n3720 VDD.n3534 37.0005
R17334 VDD.n3759 VDD.n3534 37.0005
R17335 VDD.n3720 VDD.n3709 37.0005
R17336 VDD.n3709 VDD.n3538 37.0005
R17337 VDD.n3712 VDD.n3711 37.0005
R17338 VDD.n3711 VDD.n3579 37.0005
R17339 VDD.n3727 VDD.n3726 37.0005
R17340 VDD.n3734 VDD.n3727 37.0005
R17341 VDD.n3723 VDD.n3542 37.0005
R17342 VDD.n3759 VDD.n3542 37.0005
R17343 VDD.n3723 VDD.n3633 37.0005
R17344 VDD.n3633 VDD.n3538 37.0005
R17345 VDD.n3630 VDD.n3629 37.0005
R17346 VDD.n3629 VDD.n3579 37.0005
R17347 VDD.n3643 VDD.n3601 37.0005
R17348 VDD.n3734 VDD.n3601 37.0005
R17349 VDD.n3647 VDD.n3533 37.0005
R17350 VDD.n3759 VDD.n3533 37.0005
R17351 VDD.n3647 VDD.n3636 37.0005
R17352 VDD.n3636 VDD.n3538 37.0005
R17353 VDD.n3639 VDD.n3638 37.0005
R17354 VDD.n3638 VDD.n3579 37.0005
R17355 VDD.n3731 VDD.n3730 37.0005
R17356 VDD.n3734 VDD.n3731 37.0005
R17357 VDD.n3761 VDD.n3760 37.0005
R17358 VDD.n3760 VDD.n3759 37.0005
R17359 VDD.n3761 VDD.n3528 37.0005
R17360 VDD.n3538 VDD.n3528 37.0005
R17361 VDD.n3578 VDD.n3577 37.0005
R17362 VDD.n3579 VDD.n3578 37.0005
R17363 VDD.n3600 VDD.n3599 37.0005
R17364 VDD.n3734 VDD.n3600 37.0005
R17365 VDD.n3752 VDD.n3532 37.0005
R17366 VDD.n3759 VDD.n3532 37.0005
R17367 VDD.n3752 VDD.n3751 37.0005
R17368 VDD.n3751 VDD.n3538 37.0005
R17369 VDD.n3553 VDD.n3551 37.0005
R17370 VDD.n3579 VDD.n3551 37.0005
R17371 VDD.n3733 VDD.n3732 37.0005
R17372 VDD.n3734 VDD.n3733 37.0005
R17373 VDD.n3758 VDD.n3757 37.0005
R17374 VDD.n3759 VDD.n3758 37.0005
R17375 VDD.n3747 VDD.n3582 37.0005
R17376 VDD.n3582 VDD.n3579 37.0005
R17377 VDD.n3744 VDD.n3537 37.0005
R17378 VDD.n3759 VDD.n3537 37.0005
R17379 VDD.n3744 VDD.n3581 37.0005
R17380 VDD.n3581 VDD.n3538 37.0005
R17381 VDD.n3881 VDD.n3880 37.0005
R17382 VDD.n3993 VDD.n3881 37.0005
R17383 VDD.n3994 VDD.n3851 37.0005
R17384 VDD.n3994 VDD.n3993 37.0005
R17385 VDD.n3998 VDD.n3798 37.0005
R17386 VDD.n4018 VDD.n3798 37.0005
R17387 VDD.n3998 VDD.n3846 37.0005
R17388 VDD.n3846 VDD.n3797 37.0005
R17389 VDD.n3849 VDD.n3848 37.0005
R17390 VDD.n3848 VDD.n3838 37.0005
R17391 VDD.n3876 VDD.n3875 37.0005
R17392 VDD.n3993 VDD.n3876 37.0005
R17393 VDD.n3872 VDD.n3795 37.0005
R17394 VDD.n4018 VDD.n3795 37.0005
R17395 VDD.n3872 VDD.n3871 37.0005
R17396 VDD.n3871 VDD.n3797 37.0005
R17397 VDD.n3868 VDD.n3867 37.0005
R17398 VDD.n3867 VDD.n3838 37.0005
R17399 VDD.n3920 VDD.n3882 37.0005
R17400 VDD.n3993 VDD.n3882 37.0005
R17401 VDD.n3924 VDD.n3799 37.0005
R17402 VDD.n4018 VDD.n3799 37.0005
R17403 VDD.n3924 VDD.n3913 37.0005
R17404 VDD.n3913 VDD.n3797 37.0005
R17405 VDD.n3916 VDD.n3915 37.0005
R17406 VDD.n3915 VDD.n3838 37.0005
R17407 VDD.n3936 VDD.n3862 37.0005
R17408 VDD.n3993 VDD.n3862 37.0005
R17409 VDD.n3940 VDD.n3794 37.0005
R17410 VDD.n4018 VDD.n3794 37.0005
R17411 VDD.n3940 VDD.n3929 37.0005
R17412 VDD.n3929 VDD.n3797 37.0005
R17413 VDD.n3932 VDD.n3931 37.0005
R17414 VDD.n3931 VDD.n3838 37.0005
R17415 VDD.n3947 VDD.n3943 37.0005
R17416 VDD.n3943 VDD.n3797 37.0005
R17417 VDD.n3945 VDD.n3944 37.0005
R17418 VDD.n3944 VDD.n3838 37.0005
R17419 VDD.n3959 VDD.n3883 37.0005
R17420 VDD.n3993 VDD.n3883 37.0005
R17421 VDD.n3963 VDD.n3800 37.0005
R17422 VDD.n4018 VDD.n3800 37.0005
R17423 VDD.n3963 VDD.n3952 37.0005
R17424 VDD.n3952 VDD.n3797 37.0005
R17425 VDD.n3955 VDD.n3954 37.0005
R17426 VDD.n3954 VDD.n3838 37.0005
R17427 VDD.n3975 VDD.n3861 37.0005
R17428 VDD.n3993 VDD.n3861 37.0005
R17429 VDD.n3979 VDD.n3793 37.0005
R17430 VDD.n4018 VDD.n3793 37.0005
R17431 VDD.n3979 VDD.n3968 37.0005
R17432 VDD.n3968 VDD.n3797 37.0005
R17433 VDD.n3971 VDD.n3970 37.0005
R17434 VDD.n3970 VDD.n3838 37.0005
R17435 VDD.n3986 VDD.n3985 37.0005
R17436 VDD.n3993 VDD.n3986 37.0005
R17437 VDD.n3982 VDD.n3801 37.0005
R17438 VDD.n4018 VDD.n3801 37.0005
R17439 VDD.n3982 VDD.n3892 37.0005
R17440 VDD.n3892 VDD.n3797 37.0005
R17441 VDD.n3889 VDD.n3888 37.0005
R17442 VDD.n3888 VDD.n3838 37.0005
R17443 VDD.n3902 VDD.n3860 37.0005
R17444 VDD.n3993 VDD.n3860 37.0005
R17445 VDD.n3906 VDD.n3792 37.0005
R17446 VDD.n4018 VDD.n3792 37.0005
R17447 VDD.n3906 VDD.n3895 37.0005
R17448 VDD.n3895 VDD.n3797 37.0005
R17449 VDD.n3898 VDD.n3897 37.0005
R17450 VDD.n3897 VDD.n3838 37.0005
R17451 VDD.n3990 VDD.n3989 37.0005
R17452 VDD.n3993 VDD.n3990 37.0005
R17453 VDD.n4020 VDD.n4019 37.0005
R17454 VDD.n4019 VDD.n4018 37.0005
R17455 VDD.n4020 VDD.n3787 37.0005
R17456 VDD.n3797 VDD.n3787 37.0005
R17457 VDD.n3837 VDD.n3836 37.0005
R17458 VDD.n3838 VDD.n3837 37.0005
R17459 VDD.n3859 VDD.n3858 37.0005
R17460 VDD.n3993 VDD.n3859 37.0005
R17461 VDD.n4011 VDD.n3791 37.0005
R17462 VDD.n4018 VDD.n3791 37.0005
R17463 VDD.n4011 VDD.n4010 37.0005
R17464 VDD.n4010 VDD.n3797 37.0005
R17465 VDD.n3812 VDD.n3810 37.0005
R17466 VDD.n3838 VDD.n3810 37.0005
R17467 VDD.n3992 VDD.n3991 37.0005
R17468 VDD.n3993 VDD.n3992 37.0005
R17469 VDD.n4017 VDD.n4016 37.0005
R17470 VDD.n4018 VDD.n4017 37.0005
R17471 VDD.n4006 VDD.n3841 37.0005
R17472 VDD.n3841 VDD.n3838 37.0005
R17473 VDD.n4003 VDD.n3796 37.0005
R17474 VDD.n4018 VDD.n3796 37.0005
R17475 VDD.n4003 VDD.n3840 37.0005
R17476 VDD.n3840 VDD.n3797 37.0005
R17477 VDD.n4140 VDD.n4139 37.0005
R17478 VDD.n4252 VDD.n4140 37.0005
R17479 VDD.n4253 VDD.n4110 37.0005
R17480 VDD.n4253 VDD.n4252 37.0005
R17481 VDD.n4257 VDD.n4057 37.0005
R17482 VDD.n4277 VDD.n4057 37.0005
R17483 VDD.n4257 VDD.n4105 37.0005
R17484 VDD.n4105 VDD.n4056 37.0005
R17485 VDD.n4108 VDD.n4107 37.0005
R17486 VDD.n4107 VDD.n4097 37.0005
R17487 VDD.n4135 VDD.n4134 37.0005
R17488 VDD.n4252 VDD.n4135 37.0005
R17489 VDD.n4131 VDD.n4054 37.0005
R17490 VDD.n4277 VDD.n4054 37.0005
R17491 VDD.n4131 VDD.n4130 37.0005
R17492 VDD.n4130 VDD.n4056 37.0005
R17493 VDD.n4127 VDD.n4126 37.0005
R17494 VDD.n4126 VDD.n4097 37.0005
R17495 VDD.n4179 VDD.n4141 37.0005
R17496 VDD.n4252 VDD.n4141 37.0005
R17497 VDD.n4183 VDD.n4058 37.0005
R17498 VDD.n4277 VDD.n4058 37.0005
R17499 VDD.n4183 VDD.n4172 37.0005
R17500 VDD.n4172 VDD.n4056 37.0005
R17501 VDD.n4175 VDD.n4174 37.0005
R17502 VDD.n4174 VDD.n4097 37.0005
R17503 VDD.n4195 VDD.n4121 37.0005
R17504 VDD.n4252 VDD.n4121 37.0005
R17505 VDD.n4199 VDD.n4053 37.0005
R17506 VDD.n4277 VDD.n4053 37.0005
R17507 VDD.n4199 VDD.n4188 37.0005
R17508 VDD.n4188 VDD.n4056 37.0005
R17509 VDD.n4191 VDD.n4190 37.0005
R17510 VDD.n4190 VDD.n4097 37.0005
R17511 VDD.n4206 VDD.n4202 37.0005
R17512 VDD.n4202 VDD.n4056 37.0005
R17513 VDD.n4204 VDD.n4203 37.0005
R17514 VDD.n4203 VDD.n4097 37.0005
R17515 VDD.n4218 VDD.n4142 37.0005
R17516 VDD.n4252 VDD.n4142 37.0005
R17517 VDD.n4222 VDD.n4059 37.0005
R17518 VDD.n4277 VDD.n4059 37.0005
R17519 VDD.n4222 VDD.n4211 37.0005
R17520 VDD.n4211 VDD.n4056 37.0005
R17521 VDD.n4214 VDD.n4213 37.0005
R17522 VDD.n4213 VDD.n4097 37.0005
R17523 VDD.n4234 VDD.n4120 37.0005
R17524 VDD.n4252 VDD.n4120 37.0005
R17525 VDD.n4238 VDD.n4052 37.0005
R17526 VDD.n4277 VDD.n4052 37.0005
R17527 VDD.n4238 VDD.n4227 37.0005
R17528 VDD.n4227 VDD.n4056 37.0005
R17529 VDD.n4230 VDD.n4229 37.0005
R17530 VDD.n4229 VDD.n4097 37.0005
R17531 VDD.n4245 VDD.n4244 37.0005
R17532 VDD.n4252 VDD.n4245 37.0005
R17533 VDD.n4241 VDD.n4060 37.0005
R17534 VDD.n4277 VDD.n4060 37.0005
R17535 VDD.n4241 VDD.n4151 37.0005
R17536 VDD.n4151 VDD.n4056 37.0005
R17537 VDD.n4148 VDD.n4147 37.0005
R17538 VDD.n4147 VDD.n4097 37.0005
R17539 VDD.n4161 VDD.n4119 37.0005
R17540 VDD.n4252 VDD.n4119 37.0005
R17541 VDD.n4165 VDD.n4051 37.0005
R17542 VDD.n4277 VDD.n4051 37.0005
R17543 VDD.n4165 VDD.n4154 37.0005
R17544 VDD.n4154 VDD.n4056 37.0005
R17545 VDD.n4157 VDD.n4156 37.0005
R17546 VDD.n4156 VDD.n4097 37.0005
R17547 VDD.n4249 VDD.n4248 37.0005
R17548 VDD.n4252 VDD.n4249 37.0005
R17549 VDD.n4279 VDD.n4278 37.0005
R17550 VDD.n4278 VDD.n4277 37.0005
R17551 VDD.n4279 VDD.n4046 37.0005
R17552 VDD.n4056 VDD.n4046 37.0005
R17553 VDD.n4096 VDD.n4095 37.0005
R17554 VDD.n4097 VDD.n4096 37.0005
R17555 VDD.n4118 VDD.n4117 37.0005
R17556 VDD.n4252 VDD.n4118 37.0005
R17557 VDD.n4270 VDD.n4050 37.0005
R17558 VDD.n4277 VDD.n4050 37.0005
R17559 VDD.n4270 VDD.n4269 37.0005
R17560 VDD.n4269 VDD.n4056 37.0005
R17561 VDD.n4071 VDD.n4069 37.0005
R17562 VDD.n4097 VDD.n4069 37.0005
R17563 VDD.n4251 VDD.n4250 37.0005
R17564 VDD.n4252 VDD.n4251 37.0005
R17565 VDD.n4276 VDD.n4275 37.0005
R17566 VDD.n4277 VDD.n4276 37.0005
R17567 VDD.n4265 VDD.n4100 37.0005
R17568 VDD.n4100 VDD.n4097 37.0005
R17569 VDD.n4262 VDD.n4055 37.0005
R17570 VDD.n4277 VDD.n4055 37.0005
R17571 VDD.n4262 VDD.n4099 37.0005
R17572 VDD.n4099 VDD.n4056 37.0005
R17573 VDD.n4399 VDD.n4398 37.0005
R17574 VDD.n4511 VDD.n4399 37.0005
R17575 VDD.n4512 VDD.n4369 37.0005
R17576 VDD.n4512 VDD.n4511 37.0005
R17577 VDD.n4516 VDD.n4316 37.0005
R17578 VDD.n4536 VDD.n4316 37.0005
R17579 VDD.n4516 VDD.n4364 37.0005
R17580 VDD.n4364 VDD.n4315 37.0005
R17581 VDD.n4367 VDD.n4366 37.0005
R17582 VDD.n4366 VDD.n4356 37.0005
R17583 VDD.n4394 VDD.n4393 37.0005
R17584 VDD.n4511 VDD.n4394 37.0005
R17585 VDD.n4390 VDD.n4313 37.0005
R17586 VDD.n4536 VDD.n4313 37.0005
R17587 VDD.n4390 VDD.n4389 37.0005
R17588 VDD.n4389 VDD.n4315 37.0005
R17589 VDD.n4386 VDD.n4385 37.0005
R17590 VDD.n4385 VDD.n4356 37.0005
R17591 VDD.n4438 VDD.n4400 37.0005
R17592 VDD.n4511 VDD.n4400 37.0005
R17593 VDD.n4442 VDD.n4317 37.0005
R17594 VDD.n4536 VDD.n4317 37.0005
R17595 VDD.n4442 VDD.n4431 37.0005
R17596 VDD.n4431 VDD.n4315 37.0005
R17597 VDD.n4434 VDD.n4433 37.0005
R17598 VDD.n4433 VDD.n4356 37.0005
R17599 VDD.n4454 VDD.n4380 37.0005
R17600 VDD.n4511 VDD.n4380 37.0005
R17601 VDD.n4458 VDD.n4312 37.0005
R17602 VDD.n4536 VDD.n4312 37.0005
R17603 VDD.n4458 VDD.n4447 37.0005
R17604 VDD.n4447 VDD.n4315 37.0005
R17605 VDD.n4450 VDD.n4449 37.0005
R17606 VDD.n4449 VDD.n4356 37.0005
R17607 VDD.n4465 VDD.n4461 37.0005
R17608 VDD.n4461 VDD.n4315 37.0005
R17609 VDD.n4463 VDD.n4462 37.0005
R17610 VDD.n4462 VDD.n4356 37.0005
R17611 VDD.n4477 VDD.n4401 37.0005
R17612 VDD.n4511 VDD.n4401 37.0005
R17613 VDD.n4481 VDD.n4318 37.0005
R17614 VDD.n4536 VDD.n4318 37.0005
R17615 VDD.n4481 VDD.n4470 37.0005
R17616 VDD.n4470 VDD.n4315 37.0005
R17617 VDD.n4473 VDD.n4472 37.0005
R17618 VDD.n4472 VDD.n4356 37.0005
R17619 VDD.n4493 VDD.n4379 37.0005
R17620 VDD.n4511 VDD.n4379 37.0005
R17621 VDD.n4497 VDD.n4311 37.0005
R17622 VDD.n4536 VDD.n4311 37.0005
R17623 VDD.n4497 VDD.n4486 37.0005
R17624 VDD.n4486 VDD.n4315 37.0005
R17625 VDD.n4489 VDD.n4488 37.0005
R17626 VDD.n4488 VDD.n4356 37.0005
R17627 VDD.n4504 VDD.n4503 37.0005
R17628 VDD.n4511 VDD.n4504 37.0005
R17629 VDD.n4500 VDD.n4319 37.0005
R17630 VDD.n4536 VDD.n4319 37.0005
R17631 VDD.n4500 VDD.n4410 37.0005
R17632 VDD.n4410 VDD.n4315 37.0005
R17633 VDD.n4407 VDD.n4406 37.0005
R17634 VDD.n4406 VDD.n4356 37.0005
R17635 VDD.n4420 VDD.n4378 37.0005
R17636 VDD.n4511 VDD.n4378 37.0005
R17637 VDD.n4424 VDD.n4310 37.0005
R17638 VDD.n4536 VDD.n4310 37.0005
R17639 VDD.n4424 VDD.n4413 37.0005
R17640 VDD.n4413 VDD.n4315 37.0005
R17641 VDD.n4416 VDD.n4415 37.0005
R17642 VDD.n4415 VDD.n4356 37.0005
R17643 VDD.n4508 VDD.n4507 37.0005
R17644 VDD.n4511 VDD.n4508 37.0005
R17645 VDD.n4538 VDD.n4537 37.0005
R17646 VDD.n4537 VDD.n4536 37.0005
R17647 VDD.n4538 VDD.n4305 37.0005
R17648 VDD.n4315 VDD.n4305 37.0005
R17649 VDD.n4355 VDD.n4354 37.0005
R17650 VDD.n4356 VDD.n4355 37.0005
R17651 VDD.n4377 VDD.n4376 37.0005
R17652 VDD.n4511 VDD.n4377 37.0005
R17653 VDD.n4529 VDD.n4309 37.0005
R17654 VDD.n4536 VDD.n4309 37.0005
R17655 VDD.n4529 VDD.n4528 37.0005
R17656 VDD.n4528 VDD.n4315 37.0005
R17657 VDD.n4330 VDD.n4328 37.0005
R17658 VDD.n4356 VDD.n4328 37.0005
R17659 VDD.n4510 VDD.n4509 37.0005
R17660 VDD.n4511 VDD.n4510 37.0005
R17661 VDD.n4535 VDD.n4534 37.0005
R17662 VDD.n4536 VDD.n4535 37.0005
R17663 VDD.n4524 VDD.n4359 37.0005
R17664 VDD.n4359 VDD.n4356 37.0005
R17665 VDD.n4521 VDD.n4314 37.0005
R17666 VDD.n4536 VDD.n4314 37.0005
R17667 VDD.n4521 VDD.n4358 37.0005
R17668 VDD.n4358 VDD.n4315 37.0005
R17669 VDD.n4563 VDD.n4561 37.0005
R17670 VDD.n4561 VDD.t819 37.0005
R17671 VDD.n5023 VDD.n4562 37.0005
R17672 VDD.n4562 VDD.t819 37.0005
R17673 VDD.n5032 VDD.n5031 37.0005
R17674 VDD.n5031 VDD.t796 37.0005
R17675 VDD.n5029 VDD.n5028 37.0005
R17676 VDD.n5016 VDD.n4565 37.0005
R17677 VDD.n4565 VDD.t332 37.0005
R17678 VDD.n5012 VDD.n4564 37.0005
R17679 VDD.n5007 VDD.n5006 37.0005
R17680 VDD.n5006 VDD.t269 37.0005
R17681 VDD.n5004 VDD.n5003 37.0005
R17682 VDD.n4998 VDD.n4573 37.0005
R17683 VDD.n4573 VDD.t468 37.0005
R17684 VDD.n4994 VDD.n4572 37.0005
R17685 VDD.n4582 VDD.n4580 37.0005
R17686 VDD.n4580 VDD.t252 37.0005
R17687 VDD.n4982 VDD.n4581 37.0005
R17688 VDD.n4581 VDD.t252 37.0005
R17689 VDD.n4991 VDD.n4990 37.0005
R17690 VDD.n4990 VDD.t583 37.0005
R17691 VDD.n4988 VDD.n4987 37.0005
R17692 VDD.n4975 VDD.n4584 37.0005
R17693 VDD.n4584 VDD.t585 37.0005
R17694 VDD.n4971 VDD.n4583 37.0005
R17695 VDD.n4966 VDD.n4965 37.0005
R17696 VDD.n4965 VDD.t703 37.0005
R17697 VDD.n4963 VDD.n4962 37.0005
R17698 VDD.n4957 VDD.n4592 37.0005
R17699 VDD.n4592 VDD.t888 37.0005
R17700 VDD.n4953 VDD.n4591 37.0005
R17701 VDD.n4601 VDD.n4599 37.0005
R17702 VDD.n4599 VDD.t292 37.0005
R17703 VDD.n4941 VDD.n4600 37.0005
R17704 VDD.n4600 VDD.t292 37.0005
R17705 VDD.n4950 VDD.n4949 37.0005
R17706 VDD.n4949 VDD.t598 37.0005
R17707 VDD.n4947 VDD.n4946 37.0005
R17708 VDD.n4934 VDD.n4603 37.0005
R17709 VDD.n4603 VDD.t549 37.0005
R17710 VDD.n4930 VDD.n4602 37.0005
R17711 VDD.n4925 VDD.n4924 37.0005
R17712 VDD.n4924 VDD.t732 37.0005
R17713 VDD.n4922 VDD.n4921 37.0005
R17714 VDD.n4916 VDD.n4611 37.0005
R17715 VDD.n4611 VDD.t31 37.0005
R17716 VDD.n4912 VDD.n4610 37.0005
R17717 VDD.n4620 VDD.n4618 37.0005
R17718 VDD.n4618 VDD.t828 37.0005
R17719 VDD.n4900 VDD.n4619 37.0005
R17720 VDD.n4619 VDD.t828 37.0005
R17721 VDD.n4909 VDD.n4908 37.0005
R17722 VDD.n4908 VDD.t891 37.0005
R17723 VDD.n4906 VDD.n4905 37.0005
R17724 VDD.n4893 VDD.n4622 37.0005
R17725 VDD.n4622 VDD.t526 37.0005
R17726 VDD.n4889 VDD.n4621 37.0005
R17727 VDD.n4884 VDD.n4883 37.0005
R17728 VDD.n4883 VDD.t454 37.0005
R17729 VDD.n4881 VDD.n4880 37.0005
R17730 VDD.n4875 VDD.n4630 37.0005
R17731 VDD.n4630 VDD.t59 37.0005
R17732 VDD.n4871 VDD.n4629 37.0005
R17733 VDD.n4639 VDD.n4637 37.0005
R17734 VDD.n4637 VDD.t744 37.0005
R17735 VDD.n4859 VDD.n4638 37.0005
R17736 VDD.n4638 VDD.t744 37.0005
R17737 VDD.n4868 VDD.n4867 37.0005
R17738 VDD.n4867 VDD.t594 37.0005
R17739 VDD.n4865 VDD.n4864 37.0005
R17740 VDD.n4852 VDD.n4641 37.0005
R17741 VDD.n4641 VDD.t596 37.0005
R17742 VDD.n4848 VDD.n4640 37.0005
R17743 VDD.n4843 VDD.n4842 37.0005
R17744 VDD.n4842 VDD.t368 37.0005
R17745 VDD.n4840 VDD.n4839 37.0005
R17746 VDD.n4834 VDD.n4649 37.0005
R17747 VDD.n4649 VDD.t553 37.0005
R17748 VDD.n4830 VDD.n4648 37.0005
R17749 VDD.n4658 VDD.n4656 37.0005
R17750 VDD.n4656 VDD.t822 37.0005
R17751 VDD.n4818 VDD.n4657 37.0005
R17752 VDD.n4657 VDD.t822 37.0005
R17753 VDD.n4827 VDD.n4826 37.0005
R17754 VDD.n4826 VDD.t296 37.0005
R17755 VDD.n4824 VDD.n4823 37.0005
R17756 VDD.n4811 VDD.n4660 37.0005
R17757 VDD.n4660 VDD.t645 37.0005
R17758 VDD.n4807 VDD.n4659 37.0005
R17759 VDD.n4802 VDD.n4801 37.0005
R17760 VDD.n4801 VDD.t794 37.0005
R17761 VDD.n4799 VDD.n4798 37.0005
R17762 VDD.n4793 VDD.n4668 37.0005
R17763 VDD.n4668 VDD.t87 37.0005
R17764 VDD.n4789 VDD.n4667 37.0005
R17765 VDD.n4677 VDD.n4675 37.0005
R17766 VDD.n4675 VDD.t224 37.0005
R17767 VDD.n4777 VDD.n4676 37.0005
R17768 VDD.n4676 VDD.t224 37.0005
R17769 VDD.n4786 VDD.n4785 37.0005
R17770 VDD.n4785 VDD.t422 37.0005
R17771 VDD.n4783 VDD.n4782 37.0005
R17772 VDD.n4770 VDD.n4679 37.0005
R17773 VDD.n4679 VDD.t725 37.0005
R17774 VDD.n4766 VDD.n4678 37.0005
R17775 VDD.n4761 VDD.n4760 37.0005
R17776 VDD.n4760 VDD.t878 37.0005
R17777 VDD.n4758 VDD.n4757 37.0005
R17778 VDD.n4752 VDD.n4687 37.0005
R17779 VDD.n4687 VDD.t747 37.0005
R17780 VDD.n4748 VDD.n4686 37.0005
R17781 VDD.n4696 VDD.n4694 37.0005
R17782 VDD.n4694 VDD.t812 37.0005
R17783 VDD.n4736 VDD.n4695 37.0005
R17784 VDD.n4695 VDD.t812 37.0005
R17785 VDD.n4745 VDD.n4744 37.0005
R17786 VDD.n4744 VDD.t842 37.0005
R17787 VDD.n4742 VDD.n4741 37.0005
R17788 VDD.n4729 VDD.n4698 37.0005
R17789 VDD.n4698 VDD.t869 37.0005
R17790 VDD.n4725 VDD.n4697 37.0005
R17791 VDD.n4720 VDD.n4719 37.0005
R17792 VDD.n4719 VDD.t571 37.0005
R17793 VDD.n4717 VDD.n4716 37.0005
R17794 VDD.n4711 VDD.n4706 37.0005
R17795 VDD.n4706 VDD.t340 37.0005
R17796 VDD.n4707 VDD.n4705 37.0005
R17797 VDD.n6059 VDD.n6058 37.0005
R17798 VDD.n6058 VDD.t523 37.0005
R17799 VDD.n6079 VDD.n6078 37.0005
R17800 VDD.n6078 VDD.t371 37.0005
R17801 VDD.n6050 VDD.n6049 37.0005
R17802 VDD.n6049 VDD.t371 37.0005
R17803 VDD.n6089 VDD.n6088 37.0005
R17804 VDD.n6088 VDD.t356 37.0005
R17805 VDD.n6040 VDD.n6039 37.0005
R17806 VDD.n6039 VDD.t356 37.0005
R17807 VDD.n6099 VDD.n6098 37.0005
R17808 VDD.n6098 VDD.t316 37.0005
R17809 VDD.n6029 VDD.n6028 37.0005
R17810 VDD.n6028 VDD.t316 37.0005
R17811 VDD.n6109 VDD.n6108 37.0005
R17812 VDD.n6108 VDD.t326 37.0005
R17813 VDD.n6016 VDD.n6015 37.0005
R17814 VDD.n6015 VDD.t326 37.0005
R17815 VDD.n6005 VDD.n6003 37.0005
R17816 VDD.n6003 VDD.t460 37.0005
R17817 VDD.n6117 VDD.n6004 37.0005
R17818 VDD.n6004 VDD.t460 37.0005
R17819 VDD.n6126 VDD.n6125 37.0005
R17820 VDD.n6125 VDD.t4 37.0005
R17821 VDD.n6001 VDD.n6000 37.0005
R17822 VDD.n6000 VDD.t4 37.0005
R17823 VDD.n6136 VDD.n6135 37.0005
R17824 VDD.n6135 VDD.t618 37.0005
R17825 VDD.n5988 VDD.n5987 37.0005
R17826 VDD.n5987 VDD.t618 37.0005
R17827 VDD.n6146 VDD.n6145 37.0005
R17828 VDD.n6145 VDD.t388 37.0005
R17829 VDD.n5978 VDD.n5977 37.0005
R17830 VDD.n5977 VDD.t388 37.0005
R17831 VDD.n6156 VDD.n6155 37.0005
R17832 VDD.n6155 VDD.t458 37.0005
R17833 VDD.n5967 VDD.n5966 37.0005
R17834 VDD.n5966 VDD.t458 37.0005
R17835 VDD.n6166 VDD.n6165 37.0005
R17836 VDD.n6165 VDD.t20 37.0005
R17837 VDD.n5954 VDD.n5953 37.0005
R17838 VDD.n5953 VDD.t20 37.0005
R17839 VDD.n6186 VDD.n6185 37.0005
R17840 VDD.n6185 VDD.t474 37.0005
R17841 VDD.n6175 VDD.n6174 37.0005
R17842 VDD.t474 VDD.n6175 37.0005
R17843 VDD.n6200 VDD.n6199 37.0005
R17844 VDD.n6199 VDD.t27 37.0005
R17845 VDD.n5935 VDD.n5934 37.0005
R17846 VDD.n5934 VDD.t27 37.0005
R17847 VDD.n6210 VDD.n6209 37.0005
R17848 VDD.n6209 VDD.t81 37.0005
R17849 VDD.n5922 VDD.n5921 37.0005
R17850 VDD.n5921 VDD.t81 37.0005
R17851 VDD.n6220 VDD.n6219 37.0005
R17852 VDD.n6219 VDD.t540 37.0005
R17853 VDD.n5912 VDD.n5911 37.0005
R17854 VDD.n5911 VDD.t540 37.0005
R17855 VDD.n6230 VDD.n6229 37.0005
R17856 VDD.n6229 VDD.t395 37.0005
R17857 VDD.n5901 VDD.n5900 37.0005
R17858 VDD.n5900 VDD.t395 37.0005
R17859 VDD.n6240 VDD.n6239 37.0005
R17860 VDD.n6239 VDD.t282 37.0005
R17861 VDD.n5888 VDD.n5887 37.0005
R17862 VDD.n5887 VDD.t282 37.0005
R17863 VDD.n5877 VDD.n5875 37.0005
R17864 VDD.n5875 VDD.t839 37.0005
R17865 VDD.n6248 VDD.n5876 37.0005
R17866 VDD.n5876 VDD.t839 37.0005
R17867 VDD.n6257 VDD.n6256 37.0005
R17868 VDD.n6256 VDD.t280 37.0005
R17869 VDD.n5873 VDD.n5872 37.0005
R17870 VDD.n5872 VDD.t280 37.0005
R17871 VDD.n6267 VDD.n6266 37.0005
R17872 VDD.n6266 VDD.t547 37.0005
R17873 VDD.n5860 VDD.n5859 37.0005
R17874 VDD.n5859 VDD.t547 37.0005
R17875 VDD.n6277 VDD.n6276 37.0005
R17876 VDD.n6276 VDD.t538 37.0005
R17877 VDD.n5850 VDD.n5849 37.0005
R17878 VDD.n5849 VDD.t538 37.0005
R17879 VDD.n6287 VDD.n6286 37.0005
R17880 VDD.n6286 VDD.t836 37.0005
R17881 VDD.n5839 VDD.n5838 37.0005
R17882 VDD.n5838 VDD.t836 37.0005
R17883 VDD.n6297 VDD.n6296 37.0005
R17884 VDD.n6296 VDD.t542 37.0005
R17885 VDD.n5826 VDD.n5825 37.0005
R17886 VDD.n5825 VDD.t542 37.0005
R17887 VDD.n6317 VDD.n6316 37.0005
R17888 VDD.n6316 VDD.t536 37.0005
R17889 VDD.n6306 VDD.n6305 37.0005
R17890 VDD.t536 VDD.n6306 37.0005
R17891 VDD.n6331 VDD.n6330 37.0005
R17892 VDD.n6330 VDD.t385 37.0005
R17893 VDD.n5807 VDD.n5806 37.0005
R17894 VDD.n5806 VDD.t385 37.0005
R17895 VDD.n6341 VDD.n6340 37.0005
R17896 VDD.n6340 VDD.t804 37.0005
R17897 VDD.n5794 VDD.n5793 37.0005
R17898 VDD.n5793 VDD.t804 37.0005
R17899 VDD.n6351 VDD.n6350 37.0005
R17900 VDD.n6350 VDD.t390 37.0005
R17901 VDD.n5784 VDD.n5783 37.0005
R17902 VDD.n5783 VDD.t390 37.0005
R17903 VDD.n6361 VDD.n6360 37.0005
R17904 VDD.n6360 VDD.t64 37.0005
R17905 VDD.n5773 VDD.n5772 37.0005
R17906 VDD.n5772 VDD.t64 37.0005
R17907 VDD.n6371 VDD.n6370 37.0005
R17908 VDD.n6370 VDD.t0 37.0005
R17909 VDD.n5760 VDD.n5759 37.0005
R17910 VDD.n5759 VDD.t0 37.0005
R17911 VDD.n5749 VDD.n5747 37.0005
R17912 VDD.n5747 VDD.t735 37.0005
R17913 VDD.n6379 VDD.n5748 37.0005
R17914 VDD.n5748 VDD.t735 37.0005
R17915 VDD.n6388 VDD.n6387 37.0005
R17916 VDD.n6387 VDD.t2 37.0005
R17917 VDD.n5745 VDD.n5744 37.0005
R17918 VDD.n5744 VDD.t2 37.0005
R17919 VDD.n6398 VDD.n6397 37.0005
R17920 VDD.n6397 VDD.t349 37.0005
R17921 VDD.n5732 VDD.n5731 37.0005
R17922 VDD.n5731 VDD.t349 37.0005
R17923 VDD.n6408 VDD.n6407 37.0005
R17924 VDD.n6407 VDD.t561 37.0005
R17925 VDD.n5722 VDD.n5721 37.0005
R17926 VDD.n5721 VDD.t561 37.0005
R17927 VDD.n6418 VDD.n6417 37.0005
R17928 VDD.n6417 VDD.t862 37.0005
R17929 VDD.n5711 VDD.n5710 37.0005
R17930 VDD.n5710 VDD.t862 37.0005
R17931 VDD.n6428 VDD.n6427 37.0005
R17932 VDD.n6427 VDD.t277 37.0005
R17933 VDD.n5698 VDD.n5697 37.0005
R17934 VDD.n5697 VDD.t277 37.0005
R17935 VDD.n6448 VDD.n6447 37.0005
R17936 VDD.n6447 VDD.t285 37.0005
R17937 VDD.n6437 VDD.n6436 37.0005
R17938 VDD.t285 VDD.n6437 37.0005
R17939 VDD.n6462 VDD.n6461 37.0005
R17940 VDD.n6461 VDD.t495 37.0005
R17941 VDD.n5679 VDD.n5678 37.0005
R17942 VDD.n5678 VDD.t495 37.0005
R17943 VDD.n6472 VDD.n6471 37.0005
R17944 VDD.n6471 VDD.t347 37.0005
R17945 VDD.n5666 VDD.n5665 37.0005
R17946 VDD.n5665 VDD.t347 37.0005
R17947 VDD.n6482 VDD.n6481 37.0005
R17948 VDD.n6481 VDD.t639 37.0005
R17949 VDD.n5656 VDD.n5655 37.0005
R17950 VDD.n5655 VDD.t639 37.0005
R17951 VDD.n6492 VDD.n6491 37.0005
R17952 VDD.n6491 VDD.t503 37.0005
R17953 VDD.n5645 VDD.n5644 37.0005
R17954 VDD.n5644 VDD.t503 37.0005
R17955 VDD.n6502 VDD.n6501 37.0005
R17956 VDD.n6501 VDD.t430 37.0005
R17957 VDD.n5632 VDD.n5631 37.0005
R17958 VDD.n5631 VDD.t430 37.0005
R17959 VDD.n5621 VDD.n5619 37.0005
R17960 VDD.n5619 VDD.t899 37.0005
R17961 VDD.n6510 VDD.n5620 37.0005
R17962 VDD.n5620 VDD.t899 37.0005
R17963 VDD.n6519 VDD.n6518 37.0005
R17964 VDD.n6518 VDD.t428 37.0005
R17965 VDD.n5617 VDD.n5616 37.0005
R17966 VDD.n5616 VDD.t428 37.0005
R17967 VDD.n6529 VDD.n6528 37.0005
R17968 VDD.n6528 VDD.t78 37.0005
R17969 VDD.n5604 VDD.n5603 37.0005
R17970 VDD.n5603 VDD.t78 37.0005
R17971 VDD.n6539 VDD.n6538 37.0005
R17972 VDD.n6538 VDD.t637 37.0005
R17973 VDD.n5594 VDD.n5593 37.0005
R17974 VDD.n5593 VDD.t637 37.0005
R17975 VDD.n6549 VDD.n6548 37.0005
R17976 VDD.n6548 VDD.t257 37.0005
R17977 VDD.n5583 VDD.n5582 37.0005
R17978 VDD.n5582 VDD.t257 37.0005
R17979 VDD.n6559 VDD.n6558 37.0005
R17980 VDD.n6558 VDD.t18 37.0005
R17981 VDD.n5570 VDD.n5569 37.0005
R17982 VDD.n5569 VDD.t18 37.0005
R17983 VDD.n6579 VDD.n6578 37.0005
R17984 VDD.n6578 VDD.t563 37.0005
R17985 VDD.n6568 VDD.n6567 37.0005
R17986 VDD.t563 VDD.n6568 37.0005
R17987 VDD.n6593 VDD.n6592 37.0005
R17988 VDD.n6592 VDD.t70 37.0005
R17989 VDD.n5551 VDD.n5550 37.0005
R17990 VDD.n5550 VDD.t70 37.0005
R17991 VDD.n6603 VDD.n6602 37.0005
R17992 VDD.n6602 VDD.t400 37.0005
R17993 VDD.n5538 VDD.n5537 37.0005
R17994 VDD.n5537 VDD.t400 37.0005
R17995 VDD.n6613 VDD.n6612 37.0005
R17996 VDD.n6612 VDD.t635 37.0005
R17997 VDD.n5528 VDD.n5527 37.0005
R17998 VDD.n5527 VDD.t635 37.0005
R17999 VDD.n6623 VDD.n6622 37.0005
R18000 VDD.n6622 VDD.t625 37.0005
R18001 VDD.n5517 VDD.n5516 37.0005
R18002 VDD.n5516 VDD.t625 37.0005
R18003 VDD.n6633 VDD.n6632 37.0005
R18004 VDD.n6632 VDD.t306 37.0005
R18005 VDD.n5504 VDD.n5503 37.0005
R18006 VDD.n5503 VDD.t306 37.0005
R18007 VDD.n5493 VDD.n5491 37.0005
R18008 VDD.n5491 VDD.t40 37.0005
R18009 VDD.n6641 VDD.n5492 37.0005
R18010 VDD.n5492 VDD.t40 37.0005
R18011 VDD.n6650 VDD.n6649 37.0005
R18012 VDD.n6649 VDD.t420 37.0005
R18013 VDD.n5489 VDD.n5488 37.0005
R18014 VDD.n5488 VDD.t420 37.0005
R18015 VDD.n6660 VDD.n6659 37.0005
R18016 VDD.n6659 VDD.t465 37.0005
R18017 VDD.n5476 VDD.n5475 37.0005
R18018 VDD.n5475 VDD.t465 37.0005
R18019 VDD.n6670 VDD.n6669 37.0005
R18020 VDD.n6669 VDD.t352 37.0005
R18021 VDD.n5466 VDD.n5465 37.0005
R18022 VDD.n5465 VDD.t352 37.0005
R18023 VDD.n6680 VDD.n6679 37.0005
R18024 VDD.n6679 VDD.t37 37.0005
R18025 VDD.n5455 VDD.n5454 37.0005
R18026 VDD.n5454 VDD.t37 37.0005
R18027 VDD.n6690 VDD.n6689 37.0005
R18028 VDD.n6689 VDD.t68 37.0005
R18029 VDD.n5442 VDD.n5441 37.0005
R18030 VDD.n5441 VDD.t68 37.0005
R18031 VDD.n6710 VDD.n6709 37.0005
R18032 VDD.n6709 VDD.t364 37.0005
R18033 VDD.n6699 VDD.n6698 37.0005
R18034 VDD.t364 VDD.n6699 37.0005
R18035 VDD.n6724 VDD.n6723 37.0005
R18036 VDD.n6723 VDD.t411 37.0005
R18037 VDD.n5423 VDD.n5422 37.0005
R18038 VDD.n5422 VDD.t411 37.0005
R18039 VDD.n6734 VDD.n6733 37.0005
R18040 VDD.n6733 VDD.t287 37.0005
R18041 VDD.n5410 VDD.n5409 37.0005
R18042 VDD.n5409 VDD.t287 37.0005
R18043 VDD.n6744 VDD.n6743 37.0005
R18044 VDD.n6743 VDD.t568 37.0005
R18045 VDD.n5400 VDD.n5399 37.0005
R18046 VDD.n5399 VDD.t568 37.0005
R18047 VDD.n6754 VDD.n6753 37.0005
R18048 VDD.n6753 VDD.t439 37.0005
R18049 VDD.n5389 VDD.n5388 37.0005
R18050 VDD.n5388 VDD.t439 37.0005
R18051 VDD.n6764 VDD.n6763 37.0005
R18052 VDD.n6763 VDD.t215 37.0005
R18053 VDD.n5376 VDD.n5375 37.0005
R18054 VDD.n5375 VDD.t215 37.0005
R18055 VDD.n5365 VDD.n5363 37.0005
R18056 VDD.n5363 VDD.t485 37.0005
R18057 VDD.n6772 VDD.n5364 37.0005
R18058 VDD.n5364 VDD.t485 37.0005
R18059 VDD.n6781 VDD.n6780 37.0005
R18060 VDD.n6780 VDD.t74 37.0005
R18061 VDD.n5361 VDD.n5360 37.0005
R18062 VDD.n5360 VDD.t74 37.0005
R18063 VDD.n6791 VDD.n6790 37.0005
R18064 VDD.n6790 VDD.t604 37.0005
R18065 VDD.n5348 VDD.n5347 37.0005
R18066 VDD.n5347 VDD.t604 37.0005
R18067 VDD.n6801 VDD.n6800 37.0005
R18068 VDD.n6800 VDD.t358 37.0005
R18069 VDD.n5338 VDD.n5337 37.0005
R18070 VDD.n5337 VDD.t358 37.0005
R18071 VDD.n6811 VDD.n6810 37.0005
R18072 VDD.n6810 VDD.t482 37.0005
R18073 VDD.n5327 VDD.n5326 37.0005
R18074 VDD.n5326 VDD.t482 37.0005
R18075 VDD.n6821 VDD.n6820 37.0005
R18076 VDD.n6820 VDD.t94 37.0005
R18077 VDD.n5314 VDD.n5313 37.0005
R18078 VDD.n5313 VDD.t94 37.0005
R18079 VDD.n6841 VDD.n6840 37.0005
R18080 VDD.n6840 VDD.t493 37.0005
R18081 VDD.n6830 VDD.n6829 37.0005
R18082 VDD.t493 VDD.n6830 37.0005
R18083 VDD.n6855 VDD.n6854 37.0005
R18084 VDD.n6854 VDD.t308 37.0005
R18085 VDD.n5295 VDD.n5294 37.0005
R18086 VDD.n5294 VDD.t308 37.0005
R18087 VDD.n6865 VDD.n6864 37.0005
R18088 VDD.n6864 VDD.t418 37.0005
R18089 VDD.n5282 VDD.n5281 37.0005
R18090 VDD.n5281 VDD.t418 37.0005
R18091 VDD.n6875 VDD.n6874 37.0005
R18092 VDD.n6874 VDD.t90 37.0005
R18093 VDD.n5272 VDD.n5271 37.0005
R18094 VDD.n5271 VDD.t90 37.0005
R18095 VDD.n6885 VDD.n6884 37.0005
R18096 VDD.n6884 VDD.t442 37.0005
R18097 VDD.n5261 VDD.n5260 37.0005
R18098 VDD.n5260 VDD.t442 37.0005
R18099 VDD.n6895 VDD.n6894 37.0005
R18100 VDD.n6894 VDD.t501 37.0005
R18101 VDD.n5248 VDD.n5247 37.0005
R18102 VDD.n5247 VDD.t501 37.0005
R18103 VDD.n5237 VDD.n5235 37.0005
R18104 VDD.n5235 VDD.t376 37.0005
R18105 VDD.n6903 VDD.n5236 37.0005
R18106 VDD.n5236 VDD.t376 37.0005
R18107 VDD.n6912 VDD.n6911 37.0005
R18108 VDD.n6911 VDD.t261 37.0005
R18109 VDD.n5233 VDD.n5232 37.0005
R18110 VDD.n5232 VDD.t261 37.0005
R18111 VDD.n6922 VDD.n6921 37.0005
R18112 VDD.n6921 VDD.t335 37.0005
R18113 VDD.n5220 VDD.n5219 37.0005
R18114 VDD.n5219 VDD.t335 37.0005
R18115 VDD.n6932 VDD.n6931 37.0005
R18116 VDD.n6931 VDD.t566 37.0005
R18117 VDD.n5210 VDD.n5209 37.0005
R18118 VDD.n5209 VDD.t566 37.0005
R18119 VDD.n6942 VDD.n6941 37.0005
R18120 VDD.n6941 VDD.t343 37.0005
R18121 VDD.n5199 VDD.n5198 37.0005
R18122 VDD.n5198 VDD.t343 37.0005
R18123 VDD.n6952 VDD.n6951 37.0005
R18124 VDD.n6951 VDD.t487 37.0005
R18125 VDD.n5186 VDD.n5185 37.0005
R18126 VDD.n5185 VDD.t487 37.0005
R18127 VDD.n6972 VDD.n6971 37.0005
R18128 VDD.n6971 VDD.t478 37.0005
R18129 VDD.n6961 VDD.n6960 37.0005
R18130 VDD.t478 VDD.n6961 37.0005
R18131 VDD.n6986 VDD.n6985 37.0005
R18132 VDD.n6985 VDD.t425 37.0005
R18133 VDD.n5167 VDD.n5166 37.0005
R18134 VDD.n5166 VDD.t425 37.0005
R18135 VDD.n6996 VDD.n6995 37.0005
R18136 VDD.n6995 VDD.t506 37.0005
R18137 VDD.n5154 VDD.n5153 37.0005
R18138 VDD.n5153 VDD.t506 37.0005
R18139 VDD.n7006 VDD.n7005 37.0005
R18140 VDD.n7005 VDD.t763 37.0005
R18141 VDD.n5144 VDD.n5143 37.0005
R18142 VDD.n5143 VDD.t763 37.0005
R18143 VDD.n7016 VDD.n7015 37.0005
R18144 VDD.n7015 VDD.t529 37.0005
R18145 VDD.n5133 VDD.n5132 37.0005
R18146 VDD.n5132 VDD.t529 37.0005
R18147 VDD.n7026 VDD.n7025 37.0005
R18148 VDD.n7025 VDD.t222 37.0005
R18149 VDD.n5120 VDD.n5119 37.0005
R18150 VDD.n5119 VDD.t222 37.0005
R18151 VDD.n5109 VDD.n5107 37.0005
R18152 VDD.n5107 VDD.t614 37.0005
R18153 VDD.n7034 VDD.n5108 37.0005
R18154 VDD.n5108 VDD.t614 37.0005
R18155 VDD.n7043 VDD.n7042 37.0005
R18156 VDD.n7042 VDD.t303 37.0005
R18157 VDD.n5105 VDD.n5104 37.0005
R18158 VDD.n5104 VDD.t303 37.0005
R18159 VDD.n7053 VDD.n7052 37.0005
R18160 VDD.n7052 VDD.t62 37.0005
R18161 VDD.n5092 VDD.n5091 37.0005
R18162 VDD.n5091 VDD.t62 37.0005
R18163 VDD.n7063 VDD.n7062 37.0005
R18164 VDD.n7062 VDD.t408 37.0005
R18165 VDD.n5082 VDD.n5081 37.0005
R18166 VDD.n5081 VDD.t408 37.0005
R18167 VDD.n7073 VDD.n7072 37.0005
R18168 VDD.n7072 VDD.t611 37.0005
R18169 VDD.n5071 VDD.n5070 37.0005
R18170 VDD.n5070 VDD.t611 37.0005
R18171 VDD.n7083 VDD.n7082 37.0005
R18172 VDD.n7082 VDD.t628 37.0005
R18173 VDD.n5058 VDD.n5057 37.0005
R18174 VDD.n5057 VDD.t628 37.0005
R18175 VDD.n7093 VDD.n7092 37.0005
R18176 VDD.n7092 VDD.t643 37.0005
R18177 VDD.n5048 VDD.n5047 37.0005
R18178 VDD.n5047 VDD.t643 37.0005
R18179 VDD.n6045 VDD.n6043 37.0005
R18180 VDD.n6043 VDD.t371 37.0005
R18181 VDD.n6079 VDD.n6044 37.0005
R18182 VDD.n6044 VDD.t371 37.0005
R18183 VDD.n6034 VDD.n6032 37.0005
R18184 VDD.n6032 VDD.t356 37.0005
R18185 VDD.n6089 VDD.n6033 37.0005
R18186 VDD.n6033 VDD.t356 37.0005
R18187 VDD.n6021 VDD.n6019 37.0005
R18188 VDD.n6019 VDD.t316 37.0005
R18189 VDD.n6099 VDD.n6020 37.0005
R18190 VDD.n6020 VDD.t316 37.0005
R18191 VDD.n6009 VDD.n6007 37.0005
R18192 VDD.n6007 VDD.t326 37.0005
R18193 VDD.n6109 VDD.n6008 37.0005
R18194 VDD.n6008 VDD.t326 37.0005
R18195 VDD.n5993 VDD.n5991 37.0005
R18196 VDD.n5991 VDD.t4 37.0005
R18197 VDD.n6126 VDD.n5992 37.0005
R18198 VDD.n5992 VDD.t4 37.0005
R18199 VDD.n5983 VDD.n5981 37.0005
R18200 VDD.n5981 VDD.t618 37.0005
R18201 VDD.n6136 VDD.n5982 37.0005
R18202 VDD.n5982 VDD.t618 37.0005
R18203 VDD.n5972 VDD.n5970 37.0005
R18204 VDD.n5970 VDD.t388 37.0005
R18205 VDD.n6146 VDD.n5971 37.0005
R18206 VDD.n5971 VDD.t388 37.0005
R18207 VDD.n5959 VDD.n5957 37.0005
R18208 VDD.n5957 VDD.t458 37.0005
R18209 VDD.n6156 VDD.n5958 37.0005
R18210 VDD.n5958 VDD.t458 37.0005
R18211 VDD.n5950 VDD.n5948 37.0005
R18212 VDD.n5948 VDD.t20 37.0005
R18213 VDD.n6166 VDD.n5949 37.0005
R18214 VDD.n5949 VDD.t20 37.0005
R18215 VDD.n6184 VDD.n6183 37.0005
R18216 VDD.t474 VDD.n6184 37.0005
R18217 VDD.n6186 VDD.n5943 37.0005
R18218 VDD.t474 VDD.n5943 37.0005
R18219 VDD.n5939 VDD.n5937 37.0005
R18220 VDD.n5937 VDD.t716 37.0005
R18221 VDD.n6191 VDD.n5938 37.0005
R18222 VDD.n5938 VDD.t716 37.0005
R18223 VDD.n5927 VDD.n5925 37.0005
R18224 VDD.n5925 VDD.t27 37.0005
R18225 VDD.n6200 VDD.n5926 37.0005
R18226 VDD.n5926 VDD.t27 37.0005
R18227 VDD.n5917 VDD.n5915 37.0005
R18228 VDD.n5915 VDD.t81 37.0005
R18229 VDD.n6210 VDD.n5916 37.0005
R18230 VDD.n5916 VDD.t81 37.0005
R18231 VDD.n5906 VDD.n5904 37.0005
R18232 VDD.n5904 VDD.t540 37.0005
R18233 VDD.n6220 VDD.n5905 37.0005
R18234 VDD.n5905 VDD.t540 37.0005
R18235 VDD.n5893 VDD.n5891 37.0005
R18236 VDD.n5891 VDD.t395 37.0005
R18237 VDD.n6230 VDD.n5892 37.0005
R18238 VDD.n5892 VDD.t395 37.0005
R18239 VDD.n5881 VDD.n5879 37.0005
R18240 VDD.n5879 VDD.t282 37.0005
R18241 VDD.n6240 VDD.n5880 37.0005
R18242 VDD.n5880 VDD.t282 37.0005
R18243 VDD.n5865 VDD.n5863 37.0005
R18244 VDD.n5863 VDD.t280 37.0005
R18245 VDD.n6257 VDD.n5864 37.0005
R18246 VDD.n5864 VDD.t280 37.0005
R18247 VDD.n5855 VDD.n5853 37.0005
R18248 VDD.n5853 VDD.t547 37.0005
R18249 VDD.n6267 VDD.n5854 37.0005
R18250 VDD.n5854 VDD.t547 37.0005
R18251 VDD.n5844 VDD.n5842 37.0005
R18252 VDD.n5842 VDD.t538 37.0005
R18253 VDD.n6277 VDD.n5843 37.0005
R18254 VDD.n5843 VDD.t538 37.0005
R18255 VDD.n5831 VDD.n5829 37.0005
R18256 VDD.n5829 VDD.t836 37.0005
R18257 VDD.n6287 VDD.n5830 37.0005
R18258 VDD.n5830 VDD.t836 37.0005
R18259 VDD.n5822 VDD.n5820 37.0005
R18260 VDD.n5820 VDD.t542 37.0005
R18261 VDD.n6297 VDD.n5821 37.0005
R18262 VDD.n5821 VDD.t542 37.0005
R18263 VDD.n6315 VDD.n6314 37.0005
R18264 VDD.t536 VDD.n6315 37.0005
R18265 VDD.n6317 VDD.n5815 37.0005
R18266 VDD.t536 VDD.n5815 37.0005
R18267 VDD.n5811 VDD.n5809 37.0005
R18268 VDD.n5809 VDD.t720 37.0005
R18269 VDD.n6322 VDD.n5810 37.0005
R18270 VDD.n5810 VDD.t720 37.0005
R18271 VDD.n5799 VDD.n5797 37.0005
R18272 VDD.n5797 VDD.t385 37.0005
R18273 VDD.n6331 VDD.n5798 37.0005
R18274 VDD.n5798 VDD.t385 37.0005
R18275 VDD.n5789 VDD.n5787 37.0005
R18276 VDD.n5787 VDD.t804 37.0005
R18277 VDD.n6341 VDD.n5788 37.0005
R18278 VDD.n5788 VDD.t804 37.0005
R18279 VDD.n5778 VDD.n5776 37.0005
R18280 VDD.n5776 VDD.t390 37.0005
R18281 VDD.n6351 VDD.n5777 37.0005
R18282 VDD.n5777 VDD.t390 37.0005
R18283 VDD.n5765 VDD.n5763 37.0005
R18284 VDD.n5763 VDD.t64 37.0005
R18285 VDD.n6361 VDD.n5764 37.0005
R18286 VDD.n5764 VDD.t64 37.0005
R18287 VDD.n5753 VDD.n5751 37.0005
R18288 VDD.n5751 VDD.t0 37.0005
R18289 VDD.n6371 VDD.n5752 37.0005
R18290 VDD.n5752 VDD.t0 37.0005
R18291 VDD.n5737 VDD.n5735 37.0005
R18292 VDD.n5735 VDD.t2 37.0005
R18293 VDD.n6388 VDD.n5736 37.0005
R18294 VDD.n5736 VDD.t2 37.0005
R18295 VDD.n5727 VDD.n5725 37.0005
R18296 VDD.n5725 VDD.t349 37.0005
R18297 VDD.n6398 VDD.n5726 37.0005
R18298 VDD.n5726 VDD.t349 37.0005
R18299 VDD.n5716 VDD.n5714 37.0005
R18300 VDD.n5714 VDD.t561 37.0005
R18301 VDD.n6408 VDD.n5715 37.0005
R18302 VDD.n5715 VDD.t561 37.0005
R18303 VDD.n5703 VDD.n5701 37.0005
R18304 VDD.n5701 VDD.t862 37.0005
R18305 VDD.n6418 VDD.n5702 37.0005
R18306 VDD.n5702 VDD.t862 37.0005
R18307 VDD.n5694 VDD.n5692 37.0005
R18308 VDD.n5692 VDD.t277 37.0005
R18309 VDD.n6428 VDD.n5693 37.0005
R18310 VDD.n5693 VDD.t277 37.0005
R18311 VDD.n6446 VDD.n6445 37.0005
R18312 VDD.t285 VDD.n6446 37.0005
R18313 VDD.n6448 VDD.n5687 37.0005
R18314 VDD.t285 VDD.n5687 37.0005
R18315 VDD.n5683 VDD.n5681 37.0005
R18316 VDD.n5681 VDD.t450 37.0005
R18317 VDD.n6453 VDD.n5682 37.0005
R18318 VDD.n5682 VDD.t450 37.0005
R18319 VDD.n5671 VDD.n5669 37.0005
R18320 VDD.n5669 VDD.t495 37.0005
R18321 VDD.n6462 VDD.n5670 37.0005
R18322 VDD.n5670 VDD.t495 37.0005
R18323 VDD.n5661 VDD.n5659 37.0005
R18324 VDD.n5659 VDD.t347 37.0005
R18325 VDD.n6472 VDD.n5660 37.0005
R18326 VDD.n5660 VDD.t347 37.0005
R18327 VDD.n5650 VDD.n5648 37.0005
R18328 VDD.n5648 VDD.t639 37.0005
R18329 VDD.n6482 VDD.n5649 37.0005
R18330 VDD.n5649 VDD.t639 37.0005
R18331 VDD.n5637 VDD.n5635 37.0005
R18332 VDD.n5635 VDD.t503 37.0005
R18333 VDD.n6492 VDD.n5636 37.0005
R18334 VDD.n5636 VDD.t503 37.0005
R18335 VDD.n5625 VDD.n5623 37.0005
R18336 VDD.n5623 VDD.t430 37.0005
R18337 VDD.n6502 VDD.n5624 37.0005
R18338 VDD.n5624 VDD.t430 37.0005
R18339 VDD.n5609 VDD.n5607 37.0005
R18340 VDD.n5607 VDD.t428 37.0005
R18341 VDD.n6519 VDD.n5608 37.0005
R18342 VDD.n5608 VDD.t428 37.0005
R18343 VDD.n5599 VDD.n5597 37.0005
R18344 VDD.n5597 VDD.t78 37.0005
R18345 VDD.n6529 VDD.n5598 37.0005
R18346 VDD.n5598 VDD.t78 37.0005
R18347 VDD.n5588 VDD.n5586 37.0005
R18348 VDD.n5586 VDD.t637 37.0005
R18349 VDD.n6539 VDD.n5587 37.0005
R18350 VDD.n5587 VDD.t637 37.0005
R18351 VDD.n5575 VDD.n5573 37.0005
R18352 VDD.n5573 VDD.t257 37.0005
R18353 VDD.n6549 VDD.n5574 37.0005
R18354 VDD.n5574 VDD.t257 37.0005
R18355 VDD.n5566 VDD.n5564 37.0005
R18356 VDD.n5564 VDD.t18 37.0005
R18357 VDD.n6559 VDD.n5565 37.0005
R18358 VDD.n5565 VDD.t18 37.0005
R18359 VDD.n6577 VDD.n6576 37.0005
R18360 VDD.t563 VDD.n6577 37.0005
R18361 VDD.n6579 VDD.n5559 37.0005
R18362 VDD.t563 VDD.n5559 37.0005
R18363 VDD.n5555 VDD.n5553 37.0005
R18364 VDD.n5553 VDD.t16 37.0005
R18365 VDD.n6584 VDD.n5554 37.0005
R18366 VDD.n5554 VDD.t16 37.0005
R18367 VDD.n5543 VDD.n5541 37.0005
R18368 VDD.n5541 VDD.t70 37.0005
R18369 VDD.n6593 VDD.n5542 37.0005
R18370 VDD.n5542 VDD.t70 37.0005
R18371 VDD.n5533 VDD.n5531 37.0005
R18372 VDD.n5531 VDD.t400 37.0005
R18373 VDD.n6603 VDD.n5532 37.0005
R18374 VDD.n5532 VDD.t400 37.0005
R18375 VDD.n5522 VDD.n5520 37.0005
R18376 VDD.n5520 VDD.t635 37.0005
R18377 VDD.n6613 VDD.n5521 37.0005
R18378 VDD.n5521 VDD.t635 37.0005
R18379 VDD.n5509 VDD.n5507 37.0005
R18380 VDD.n5507 VDD.t625 37.0005
R18381 VDD.n6623 VDD.n5508 37.0005
R18382 VDD.n5508 VDD.t625 37.0005
R18383 VDD.n5497 VDD.n5495 37.0005
R18384 VDD.n5495 VDD.t306 37.0005
R18385 VDD.n6633 VDD.n5496 37.0005
R18386 VDD.n5496 VDD.t306 37.0005
R18387 VDD.n5481 VDD.n5479 37.0005
R18388 VDD.n5479 VDD.t420 37.0005
R18389 VDD.n6650 VDD.n5480 37.0005
R18390 VDD.n5480 VDD.t420 37.0005
R18391 VDD.n5471 VDD.n5469 37.0005
R18392 VDD.n5469 VDD.t465 37.0005
R18393 VDD.n6660 VDD.n5470 37.0005
R18394 VDD.n5470 VDD.t465 37.0005
R18395 VDD.n5460 VDD.n5458 37.0005
R18396 VDD.n5458 VDD.t352 37.0005
R18397 VDD.n6670 VDD.n5459 37.0005
R18398 VDD.n5459 VDD.t352 37.0005
R18399 VDD.n5447 VDD.n5445 37.0005
R18400 VDD.n5445 VDD.t37 37.0005
R18401 VDD.n6680 VDD.n5446 37.0005
R18402 VDD.n5446 VDD.t37 37.0005
R18403 VDD.n5438 VDD.n5436 37.0005
R18404 VDD.n5436 VDD.t68 37.0005
R18405 VDD.n6690 VDD.n5437 37.0005
R18406 VDD.n5437 VDD.t68 37.0005
R18407 VDD.n6708 VDD.n6707 37.0005
R18408 VDD.t364 VDD.n6708 37.0005
R18409 VDD.n6710 VDD.n5431 37.0005
R18410 VDD.t364 VDD.n5431 37.0005
R18411 VDD.n5427 VDD.n5425 37.0005
R18412 VDD.n5425 VDD.t718 37.0005
R18413 VDD.n6715 VDD.n5426 37.0005
R18414 VDD.n5426 VDD.t718 37.0005
R18415 VDD.n5415 VDD.n5413 37.0005
R18416 VDD.n5413 VDD.t411 37.0005
R18417 VDD.n6724 VDD.n5414 37.0005
R18418 VDD.n5414 VDD.t411 37.0005
R18419 VDD.n5405 VDD.n5403 37.0005
R18420 VDD.n5403 VDD.t287 37.0005
R18421 VDD.n6734 VDD.n5404 37.0005
R18422 VDD.n5404 VDD.t287 37.0005
R18423 VDD.n5394 VDD.n5392 37.0005
R18424 VDD.n5392 VDD.t568 37.0005
R18425 VDD.n6744 VDD.n5393 37.0005
R18426 VDD.n5393 VDD.t568 37.0005
R18427 VDD.n5381 VDD.n5379 37.0005
R18428 VDD.n5379 VDD.t439 37.0005
R18429 VDD.n6754 VDD.n5380 37.0005
R18430 VDD.n5380 VDD.t439 37.0005
R18431 VDD.n5369 VDD.n5367 37.0005
R18432 VDD.n5367 VDD.t215 37.0005
R18433 VDD.n6764 VDD.n5368 37.0005
R18434 VDD.n5368 VDD.t215 37.0005
R18435 VDD.n5353 VDD.n5351 37.0005
R18436 VDD.n5351 VDD.t74 37.0005
R18437 VDD.n6781 VDD.n5352 37.0005
R18438 VDD.n5352 VDD.t74 37.0005
R18439 VDD.n5343 VDD.n5341 37.0005
R18440 VDD.n5341 VDD.t604 37.0005
R18441 VDD.n6791 VDD.n5342 37.0005
R18442 VDD.n5342 VDD.t604 37.0005
R18443 VDD.n5332 VDD.n5330 37.0005
R18444 VDD.n5330 VDD.t358 37.0005
R18445 VDD.n6801 VDD.n5331 37.0005
R18446 VDD.n5331 VDD.t358 37.0005
R18447 VDD.n5319 VDD.n5317 37.0005
R18448 VDD.n5317 VDD.t482 37.0005
R18449 VDD.n6811 VDD.n5318 37.0005
R18450 VDD.n5318 VDD.t482 37.0005
R18451 VDD.n5310 VDD.n5308 37.0005
R18452 VDD.n5308 VDD.t94 37.0005
R18453 VDD.n6821 VDD.n5309 37.0005
R18454 VDD.n5309 VDD.t94 37.0005
R18455 VDD.n6839 VDD.n6838 37.0005
R18456 VDD.t493 VDD.n6839 37.0005
R18457 VDD.n6841 VDD.n5303 37.0005
R18458 VDD.t493 VDD.n5303 37.0005
R18459 VDD.n5299 VDD.n5297 37.0005
R18460 VDD.n5297 VDD.t275 37.0005
R18461 VDD.n6846 VDD.n5298 37.0005
R18462 VDD.n5298 VDD.t275 37.0005
R18463 VDD.n5287 VDD.n5285 37.0005
R18464 VDD.n5285 VDD.t308 37.0005
R18465 VDD.n6855 VDD.n5286 37.0005
R18466 VDD.n5286 VDD.t308 37.0005
R18467 VDD.n5277 VDD.n5275 37.0005
R18468 VDD.n5275 VDD.t418 37.0005
R18469 VDD.n6865 VDD.n5276 37.0005
R18470 VDD.n5276 VDD.t418 37.0005
R18471 VDD.n5266 VDD.n5264 37.0005
R18472 VDD.n5264 VDD.t90 37.0005
R18473 VDD.n6875 VDD.n5265 37.0005
R18474 VDD.n5265 VDD.t90 37.0005
R18475 VDD.n5253 VDD.n5251 37.0005
R18476 VDD.n5251 VDD.t442 37.0005
R18477 VDD.n6885 VDD.n5252 37.0005
R18478 VDD.n5252 VDD.t442 37.0005
R18479 VDD.n5241 VDD.n5239 37.0005
R18480 VDD.n5239 VDD.t501 37.0005
R18481 VDD.n6895 VDD.n5240 37.0005
R18482 VDD.n5240 VDD.t501 37.0005
R18483 VDD.n5225 VDD.n5223 37.0005
R18484 VDD.n5223 VDD.t261 37.0005
R18485 VDD.n6912 VDD.n5224 37.0005
R18486 VDD.n5224 VDD.t261 37.0005
R18487 VDD.n5215 VDD.n5213 37.0005
R18488 VDD.n5213 VDD.t335 37.0005
R18489 VDD.n6922 VDD.n5214 37.0005
R18490 VDD.n5214 VDD.t335 37.0005
R18491 VDD.n5204 VDD.n5202 37.0005
R18492 VDD.n5202 VDD.t566 37.0005
R18493 VDD.n6932 VDD.n5203 37.0005
R18494 VDD.n5203 VDD.t566 37.0005
R18495 VDD.n5191 VDD.n5189 37.0005
R18496 VDD.n5189 VDD.t343 37.0005
R18497 VDD.n6942 VDD.n5190 37.0005
R18498 VDD.n5190 VDD.t343 37.0005
R18499 VDD.n5182 VDD.n5180 37.0005
R18500 VDD.n5180 VDD.t487 37.0005
R18501 VDD.n6952 VDD.n5181 37.0005
R18502 VDD.n5181 VDD.t487 37.0005
R18503 VDD.n6970 VDD.n6969 37.0005
R18504 VDD.t478 VDD.n6970 37.0005
R18505 VDD.n6972 VDD.n5175 37.0005
R18506 VDD.t478 VDD.n5175 37.0005
R18507 VDD.n5171 VDD.n5169 37.0005
R18508 VDD.n5169 VDD.t452 37.0005
R18509 VDD.n6977 VDD.n5170 37.0005
R18510 VDD.n5170 VDD.t452 37.0005
R18511 VDD.n5159 VDD.n5157 37.0005
R18512 VDD.n5157 VDD.t425 37.0005
R18513 VDD.n6986 VDD.n5158 37.0005
R18514 VDD.n5158 VDD.t425 37.0005
R18515 VDD.n5149 VDD.n5147 37.0005
R18516 VDD.n5147 VDD.t506 37.0005
R18517 VDD.n6996 VDD.n5148 37.0005
R18518 VDD.n5148 VDD.t506 37.0005
R18519 VDD.n5138 VDD.n5136 37.0005
R18520 VDD.n5136 VDD.t763 37.0005
R18521 VDD.n7006 VDD.n5137 37.0005
R18522 VDD.n5137 VDD.t763 37.0005
R18523 VDD.n5125 VDD.n5123 37.0005
R18524 VDD.n5123 VDD.t529 37.0005
R18525 VDD.n7016 VDD.n5124 37.0005
R18526 VDD.n5124 VDD.t529 37.0005
R18527 VDD.n5113 VDD.n5111 37.0005
R18528 VDD.n5111 VDD.t222 37.0005
R18529 VDD.n7026 VDD.n5112 37.0005
R18530 VDD.n5112 VDD.t222 37.0005
R18531 VDD.n5097 VDD.n5095 37.0005
R18532 VDD.n5095 VDD.t303 37.0005
R18533 VDD.n7043 VDD.n5096 37.0005
R18534 VDD.n5096 VDD.t303 37.0005
R18535 VDD.n5087 VDD.n5085 37.0005
R18536 VDD.n5085 VDD.t62 37.0005
R18537 VDD.n7053 VDD.n5086 37.0005
R18538 VDD.n5086 VDD.t62 37.0005
R18539 VDD.n5076 VDD.n5074 37.0005
R18540 VDD.n5074 VDD.t408 37.0005
R18541 VDD.n7063 VDD.n5075 37.0005
R18542 VDD.n5075 VDD.t408 37.0005
R18543 VDD.n5063 VDD.n5061 37.0005
R18544 VDD.n5061 VDD.t611 37.0005
R18545 VDD.n7073 VDD.n5062 37.0005
R18546 VDD.n5062 VDD.t611 37.0005
R18547 VDD.n5053 VDD.n5051 37.0005
R18548 VDD.n5051 VDD.t628 37.0005
R18549 VDD.n7083 VDD.n5052 37.0005
R18550 VDD.n5052 VDD.t628 37.0005
R18551 VDD.n5042 VDD.n5040 37.0005
R18552 VDD.n5040 VDD.t643 37.0005
R18553 VDD.n7093 VDD.n5041 37.0005
R18554 VDD.n5041 VDD.t643 37.0005
R18555 VDD.n5038 VDD.n5037 37.0005
R18556 VDD.t755 VDD.n5038 37.0005
R18557 VDD.n7103 VDD.n5036 37.0005
R18558 VDD.n6055 VDD.n6053 37.0005
R18559 VDD.n6053 VDD.t523 37.0005
R18560 VDD.n6069 VDD.n6065 37.0005
R18561 VDD.n6065 VDD.t523 37.0005
R18562 VDD.n6069 VDD.n6054 37.0005
R18563 VDD.n6054 VDD.t523 37.0005
R18564 VDD.n143 VDD.n141 37.0005
R18565 VDD.n141 VDD.t776 37.0005
R18566 VDD.n7119 VDD.n142 37.0005
R18567 VDD.n142 VDD.t776 37.0005
R18568 VDD.n7108 VDD.n144 37.0005
R18569 VDD.n144 VDD.t915 37.0005
R18570 VDD.n7112 VDD.n145 37.0005
R18571 VDD.n138 VDD.n137 37.0005
R18572 VDD.t773 VDD.n138 37.0005
R18573 VDD.n7126 VDD.n136 37.0005
R18574 VDD.n124 VDD.n122 37.0005
R18575 VDD.n122 VDD.t905 37.0005
R18576 VDD.n7140 VDD.n123 37.0005
R18577 VDD.n123 VDD.t905 37.0005
R18578 VDD.n7129 VDD.n125 37.0005
R18579 VDD.n125 VDD.t880 37.0005
R18580 VDD.n7133 VDD.n126 37.0005
R18581 VDD.n119 VDD.n118 37.0005
R18582 VDD.t903 VDD.n119 37.0005
R18583 VDD.n7147 VDD.n117 37.0005
R18584 VDD.n105 VDD.n103 37.0005
R18585 VDD.n103 VDD.t866 37.0005
R18586 VDD.n7161 VDD.n104 37.0005
R18587 VDD.n104 VDD.t866 37.0005
R18588 VDD.n7150 VDD.n106 37.0005
R18589 VDD.n106 VDD.t544 37.0005
R18590 VDD.n7154 VDD.n107 37.0005
R18591 VDD.n100 VDD.n99 37.0005
R18592 VDD.t855 VDD.n100 37.0005
R18593 VDD.n7168 VDD.n98 37.0005
R18594 VDD.n86 VDD.n84 37.0005
R18595 VDD.n84 VDD.t790 37.0005
R18596 VDD.n7182 VDD.n85 37.0005
R18597 VDD.n85 VDD.t790 37.0005
R18598 VDD.n7171 VDD.n87 37.0005
R18599 VDD.n87 VDD.t96 37.0005
R18600 VDD.n7175 VDD.n88 37.0005
R18601 VDD.n81 VDD.n80 37.0005
R18602 VDD.t298 VDD.n81 37.0005
R18603 VDD.n7189 VDD.n79 37.0005
R18604 VDD.n67 VDD.n65 37.0005
R18605 VDD.n65 VDD.t713 37.0005
R18606 VDD.n7203 VDD.n66 37.0005
R18607 VDD.n66 VDD.t713 37.0005
R18608 VDD.n7192 VDD.n68 37.0005
R18609 VDD.n68 VDD.t402 37.0005
R18610 VDD.n7196 VDD.n69 37.0005
R18611 VDD.n62 VDD.n61 37.0005
R18612 VDD.t714 VDD.n62 37.0005
R18613 VDD.n7210 VDD.n60 37.0005
R18614 VDD.n48 VDD.n46 37.0005
R18615 VDD.n46 VDD.t427 37.0005
R18616 VDD.n7224 VDD.n47 37.0005
R18617 VDD.n47 VDD.t427 37.0005
R18618 VDD.n7213 VDD.n49 37.0005
R18619 VDD.n49 VDD.t630 37.0005
R18620 VDD.n7217 VDD.n50 37.0005
R18621 VDD.n43 VDD.n42 37.0005
R18622 VDD.t383 VDD.n43 37.0005
R18623 VDD.n7231 VDD.n41 37.0005
R18624 VDD.n29 VDD.n27 37.0005
R18625 VDD.n27 VDD.t894 37.0005
R18626 VDD.n7245 VDD.n28 37.0005
R18627 VDD.n28 VDD.t894 37.0005
R18628 VDD.n7234 VDD.n30 37.0005
R18629 VDD.n30 VDD.t301 37.0005
R18630 VDD.n7238 VDD.n31 37.0005
R18631 VDD.n24 VDD.n23 37.0005
R18632 VDD.t895 VDD.n24 37.0005
R18633 VDD.n7252 VDD.n22 37.0005
R18634 VDD.n10 VDD.n8 37.0005
R18635 VDD.n8 VDD.t911 37.0005
R18636 VDD.n7266 VDD.n9 37.0005
R18637 VDD.n9 VDD.t911 37.0005
R18638 VDD.n7255 VDD.n11 37.0005
R18639 VDD.n11 VDD.t314 37.0005
R18640 VDD.n7259 VDD.n12 37.0005
R18641 VDD.n5 VDD.n4 37.0005
R18642 VDD.t509 VDD.n5 37.0005
R18643 VDD.n7273 VDD.n3 37.0005
R18644 VDD.n7291 VDD.n7285 37.0005
R18645 VDD.n7287 VDD.n7284 37.0005
R18646 VDD.n7284 VDD.t883 37.0005
R18647 VDD.n7306 VDD.n7305 37.0005
R18648 VDD.t44 VDD.n7306 37.0005
R18649 VDD.n7303 VDD.n7302 37.0005
R18650 VDD.n7302 VDD.t42 37.0005
R18651 VDD.n7308 VDD.n7307 37.0005
R18652 VDD.n7307 VDD.t44 37.0005
R18653 VDD.n7300 VDD.n7279 37.0005
R18654 VDD.n7301 VDD.n7300 36.7882
R18655 VDD.n7275 VDD.n7274 36.5657
R18656 VDD.n929 VDD 35.5304
R18657 VDD.n1189 VDD 34.3865
R18658 VDD.n7332 VDD.n7331 34.3156
R18659 VDD.n1188 VDD 32.9924
R18660 VDD.n7100 VDD.n5036 31.6493
R18661 VDD.n1448 VDD 31.5947
R18662 VDD.n7330 VDD.n7311 31.0857
R18663 VDD.n1447 VDD 30.4544
R18664 VDD.n166 VDD.n156 28.8139
R18665 VDD.n1707 VDD 28.8029
R18666 VDD.n5030 VDD.n5029 28.7118
R18667 VDD.n5013 VDD.n4564 28.7118
R18668 VDD.n5005 VDD.n5004 28.7118
R18669 VDD.n4995 VDD.n4572 28.7118
R18670 VDD.n4989 VDD.n4988 28.7118
R18671 VDD.n4972 VDD.n4583 28.7118
R18672 VDD.n4964 VDD.n4963 28.7118
R18673 VDD.n4954 VDD.n4591 28.7118
R18674 VDD.n4948 VDD.n4947 28.7118
R18675 VDD.n4931 VDD.n4602 28.7118
R18676 VDD.n4923 VDD.n4922 28.7118
R18677 VDD.n4913 VDD.n4610 28.7118
R18678 VDD.n4907 VDD.n4906 28.7118
R18679 VDD.n4890 VDD.n4621 28.7118
R18680 VDD.n4882 VDD.n4881 28.7118
R18681 VDD.n4872 VDD.n4629 28.7118
R18682 VDD.n4866 VDD.n4865 28.7118
R18683 VDD.n4849 VDD.n4640 28.7118
R18684 VDD.n4841 VDD.n4840 28.7118
R18685 VDD.n4831 VDD.n4648 28.7118
R18686 VDD.n4825 VDD.n4824 28.7118
R18687 VDD.n4808 VDD.n4659 28.7118
R18688 VDD.n4800 VDD.n4799 28.7118
R18689 VDD.n4790 VDD.n4667 28.7118
R18690 VDD.n4784 VDD.n4783 28.7118
R18691 VDD.n4767 VDD.n4678 28.7118
R18692 VDD.n4759 VDD.n4758 28.7118
R18693 VDD.n4749 VDD.n4686 28.7118
R18694 VDD.n4743 VDD.n4742 28.7118
R18695 VDD.n4726 VDD.n4697 28.7118
R18696 VDD.n4718 VDD.n4717 28.7118
R18697 VDD.n4708 VDD.n4705 28.7118
R18698 VDD.n7109 VDD.n145 28.7118
R18699 VDD.n140 VDD.n136 28.7118
R18700 VDD.n7130 VDD.n126 28.7118
R18701 VDD.n121 VDD.n117 28.7118
R18702 VDD.n7151 VDD.n107 28.7118
R18703 VDD.n102 VDD.n98 28.7118
R18704 VDD.n7172 VDD.n88 28.7118
R18705 VDD.n83 VDD.n79 28.7118
R18706 VDD.n7193 VDD.n69 28.7118
R18707 VDD.n64 VDD.n60 28.7118
R18708 VDD.n7214 VDD.n50 28.7118
R18709 VDD.n45 VDD.n41 28.7118
R18710 VDD.n7235 VDD.n31 28.7118
R18711 VDD.n26 VDD.n22 28.7118
R18712 VDD.n7256 VDD.n12 28.7118
R18713 VDD.n7 VDD.n3 28.7118
R18714 VDD.n5034 VDD 28.2279
R18715 VDD.n1706 VDD 27.9164
R18716 VDD.n1966 VDD 26.0111
R18717 VDD.n403 VDD.n182 25.5883
R18718 VDD.n651 VDD.n430 25.5883
R18719 VDD.n910 VDD.n689 25.5883
R18720 VDD.n1169 VDD.n948 25.5883
R18721 VDD.n1428 VDD.n1207 25.5883
R18722 VDD.n1687 VDD.n1466 25.5883
R18723 VDD.n1946 VDD.n1725 25.5883
R18724 VDD.n2205 VDD.n1984 25.5883
R18725 VDD.n2464 VDD.n2243 25.5883
R18726 VDD.n2723 VDD.n2502 25.5883
R18727 VDD.n2982 VDD.n2761 25.5883
R18728 VDD.n3241 VDD.n3020 25.5883
R18729 VDD.n3500 VDD.n3279 25.5883
R18730 VDD.n3759 VDD.n3538 25.5883
R18731 VDD.n4018 VDD.n3797 25.5883
R18732 VDD.n4277 VDD.n4056 25.5883
R18733 VDD.n4536 VDD.n4315 25.5883
R18734 VDD.n1965 VDD 25.3784
R18735 VDD.n7301 VDD.n7299 24.6676
R18736 VDD.t42 VDD.n7283 23.5846
R18737 VDD.t44 VDD.n7283 23.5846
R18738 VDD.t44 VDD.n7295 23.5846
R18739 VDD.n7294 VDD.t883 23.5846
R18740 VDD.n2225 VDD 23.2193
R18741 VDD.n264 VDD.n262 23.1255
R18742 VDD.n262 VDD.t190 23.1255
R18743 VDD.n263 VDD.n228 23.1255
R18744 VDD.n263 VDD.t190 23.1255
R18745 VDD.n238 VDD.n237 23.1255
R18746 VDD.n238 VDD.t190 23.1255
R18747 VDD.n381 VDD.n380 23.1255
R18748 VDD.n380 VDD.t190 23.1255
R18749 VDD.n232 VDD.n217 23.1255
R18750 VDD.t101 VDD.n217 23.1255
R18751 VDD.n235 VDD.n218 23.1255
R18752 VDD.t101 VDD.n218 23.1255
R18753 VDD.n250 VDD.n248 23.1255
R18754 VDD.n248 VDD.t190 23.1255
R18755 VDD.n259 VDD.n249 23.1255
R18756 VDD.n249 VDD.t190 23.1255
R18757 VDD.n254 VDD.n215 23.1255
R18758 VDD.t101 VDD.n215 23.1255
R18759 VDD.n251 VDD.n216 23.1255
R18760 VDD.t101 VDD.n216 23.1255
R18761 VDD.n304 VDD.n303 23.1255
R18762 VDD.n303 VDD.t190 23.1255
R18763 VDD.n307 VDD.n306 23.1255
R18764 VDD.n306 VDD.t190 23.1255
R18765 VDD.n299 VDD.n213 23.1255
R18766 VDD.t101 VDD.n213 23.1255
R18767 VDD.n302 VDD.n214 23.1255
R18768 VDD.t101 VDD.n214 23.1255
R18769 VDD.n320 VDD.n319 23.1255
R18770 VDD.n319 VDD.t190 23.1255
R18771 VDD.n323 VDD.n322 23.1255
R18772 VDD.n322 VDD.t190 23.1255
R18773 VDD.n315 VDD.n211 23.1255
R18774 VDD.t101 VDD.n211 23.1255
R18775 VDD.n318 VDD.n212 23.1255
R18776 VDD.t101 VDD.n212 23.1255
R18777 VDD.n327 VDD.n209 23.1255
R18778 VDD.t101 VDD.n209 23.1255
R18779 VDD.n331 VDD.n210 23.1255
R18780 VDD.t101 VDD.n210 23.1255
R18781 VDD.n343 VDD.n342 23.1255
R18782 VDD.n342 VDD.t190 23.1255
R18783 VDD.n346 VDD.n345 23.1255
R18784 VDD.n345 VDD.t190 23.1255
R18785 VDD.n338 VDD.n207 23.1255
R18786 VDD.t101 VDD.n207 23.1255
R18787 VDD.n341 VDD.n208 23.1255
R18788 VDD.t101 VDD.n208 23.1255
R18789 VDD.n359 VDD.n358 23.1255
R18790 VDD.n358 VDD.t190 23.1255
R18791 VDD.n362 VDD.n361 23.1255
R18792 VDD.n361 VDD.t190 23.1255
R18793 VDD.n354 VDD.n205 23.1255
R18794 VDD.t101 VDD.n205 23.1255
R18795 VDD.n357 VDD.n206 23.1255
R18796 VDD.t101 VDD.n206 23.1255
R18797 VDD.n271 VDD.n269 23.1255
R18798 VDD.n269 VDD.t190 23.1255
R18799 VDD.n369 VDD.n270 23.1255
R18800 VDD.n270 VDD.t190 23.1255
R18801 VDD.n275 VDD.n203 23.1255
R18802 VDD.t101 VDD.n203 23.1255
R18803 VDD.n272 VDD.n204 23.1255
R18804 VDD.t101 VDD.n204 23.1255
R18805 VDD.n286 VDD.n285 23.1255
R18806 VDD.n285 VDD.t190 23.1255
R18807 VDD.n289 VDD.n288 23.1255
R18808 VDD.n288 VDD.t190 23.1255
R18809 VDD.n281 VDD.n201 23.1255
R18810 VDD.t101 VDD.n201 23.1255
R18811 VDD.n284 VDD.n202 23.1255
R18812 VDD.t101 VDD.n202 23.1255
R18813 VDD.n372 VDD.n174 23.1255
R18814 VDD.t190 VDD.n174 23.1255
R18815 VDD.n373 VDD.n175 23.1255
R18816 VDD.t190 VDD.n175 23.1255
R18817 VDD.n219 VDD.n199 23.1255
R18818 VDD.t101 VDD.n199 23.1255
R18819 VDD.n220 VDD.n200 23.1255
R18820 VDD.t101 VDD.n200 23.1255
R18821 VDD.n241 VDD.n239 23.1255
R18822 VDD.n239 VDD.t190 23.1255
R18823 VDD.n242 VDD.n240 23.1255
R18824 VDD.n240 VDD.t190 23.1255
R18825 VDD.n196 VDD.n194 23.1255
R18826 VDD.t101 VDD.n194 23.1255
R18827 VDD.n394 VDD.n198 23.1255
R18828 VDD.n394 VDD.t101 23.1255
R18829 VDD.n189 VDD.n187 23.1255
R18830 VDD.n187 VDD.t190 23.1255
R18831 VDD.n190 VDD.n188 23.1255
R18832 VDD.n188 VDD.t190 23.1255
R18833 VDD.n393 VDD.n392 23.1255
R18834 VDD.t101 VDD.n393 23.1255
R18835 VDD.n390 VDD.n224 23.1255
R18836 VDD.t101 VDD.n224 23.1255
R18837 VDD.n512 VDD.n510 23.1255
R18838 VDD.n510 VDD.t210 23.1255
R18839 VDD.n511 VDD.n476 23.1255
R18840 VDD.n511 VDD.t210 23.1255
R18841 VDD.n486 VDD.n485 23.1255
R18842 VDD.n486 VDD.t210 23.1255
R18843 VDD.n629 VDD.n628 23.1255
R18844 VDD.n628 VDD.t210 23.1255
R18845 VDD.n480 VDD.n465 23.1255
R18846 VDD.t106 VDD.n465 23.1255
R18847 VDD.n483 VDD.n466 23.1255
R18848 VDD.t106 VDD.n466 23.1255
R18849 VDD.n498 VDD.n496 23.1255
R18850 VDD.n496 VDD.t210 23.1255
R18851 VDD.n507 VDD.n497 23.1255
R18852 VDD.n497 VDD.t210 23.1255
R18853 VDD.n502 VDD.n463 23.1255
R18854 VDD.t106 VDD.n463 23.1255
R18855 VDD.n499 VDD.n464 23.1255
R18856 VDD.t106 VDD.n464 23.1255
R18857 VDD.n552 VDD.n551 23.1255
R18858 VDD.n551 VDD.t210 23.1255
R18859 VDD.n555 VDD.n554 23.1255
R18860 VDD.n554 VDD.t210 23.1255
R18861 VDD.n547 VDD.n461 23.1255
R18862 VDD.t106 VDD.n461 23.1255
R18863 VDD.n550 VDD.n462 23.1255
R18864 VDD.t106 VDD.n462 23.1255
R18865 VDD.n568 VDD.n567 23.1255
R18866 VDD.n567 VDD.t210 23.1255
R18867 VDD.n571 VDD.n570 23.1255
R18868 VDD.n570 VDD.t210 23.1255
R18869 VDD.n563 VDD.n459 23.1255
R18870 VDD.t106 VDD.n459 23.1255
R18871 VDD.n566 VDD.n460 23.1255
R18872 VDD.t106 VDD.n460 23.1255
R18873 VDD.n575 VDD.n457 23.1255
R18874 VDD.t106 VDD.n457 23.1255
R18875 VDD.n579 VDD.n458 23.1255
R18876 VDD.t106 VDD.n458 23.1255
R18877 VDD.n591 VDD.n590 23.1255
R18878 VDD.n590 VDD.t210 23.1255
R18879 VDD.n594 VDD.n593 23.1255
R18880 VDD.n593 VDD.t210 23.1255
R18881 VDD.n586 VDD.n455 23.1255
R18882 VDD.t106 VDD.n455 23.1255
R18883 VDD.n589 VDD.n456 23.1255
R18884 VDD.t106 VDD.n456 23.1255
R18885 VDD.n607 VDD.n606 23.1255
R18886 VDD.n606 VDD.t210 23.1255
R18887 VDD.n610 VDD.n609 23.1255
R18888 VDD.n609 VDD.t210 23.1255
R18889 VDD.n602 VDD.n453 23.1255
R18890 VDD.t106 VDD.n453 23.1255
R18891 VDD.n605 VDD.n454 23.1255
R18892 VDD.t106 VDD.n454 23.1255
R18893 VDD.n519 VDD.n517 23.1255
R18894 VDD.n517 VDD.t210 23.1255
R18895 VDD.n617 VDD.n518 23.1255
R18896 VDD.n518 VDD.t210 23.1255
R18897 VDD.n523 VDD.n451 23.1255
R18898 VDD.t106 VDD.n451 23.1255
R18899 VDD.n520 VDD.n452 23.1255
R18900 VDD.t106 VDD.n452 23.1255
R18901 VDD.n534 VDD.n533 23.1255
R18902 VDD.n533 VDD.t210 23.1255
R18903 VDD.n537 VDD.n536 23.1255
R18904 VDD.n536 VDD.t210 23.1255
R18905 VDD.n529 VDD.n449 23.1255
R18906 VDD.t106 VDD.n449 23.1255
R18907 VDD.n532 VDD.n450 23.1255
R18908 VDD.t106 VDD.n450 23.1255
R18909 VDD.n620 VDD.n422 23.1255
R18910 VDD.t210 VDD.n422 23.1255
R18911 VDD.n621 VDD.n423 23.1255
R18912 VDD.t210 VDD.n423 23.1255
R18913 VDD.n467 VDD.n447 23.1255
R18914 VDD.t106 VDD.n447 23.1255
R18915 VDD.n468 VDD.n448 23.1255
R18916 VDD.t106 VDD.n448 23.1255
R18917 VDD.n489 VDD.n487 23.1255
R18918 VDD.n487 VDD.t210 23.1255
R18919 VDD.n490 VDD.n488 23.1255
R18920 VDD.n488 VDD.t210 23.1255
R18921 VDD.n444 VDD.n442 23.1255
R18922 VDD.t106 VDD.n442 23.1255
R18923 VDD.n642 VDD.n446 23.1255
R18924 VDD.n642 VDD.t106 23.1255
R18925 VDD.n437 VDD.n435 23.1255
R18926 VDD.n435 VDD.t210 23.1255
R18927 VDD.n438 VDD.n436 23.1255
R18928 VDD.n436 VDD.t210 23.1255
R18929 VDD.n641 VDD.n640 23.1255
R18930 VDD.t106 VDD.n641 23.1255
R18931 VDD.n638 VDD.n472 23.1255
R18932 VDD.t106 VDD.n472 23.1255
R18933 VDD.n771 VDD.n769 23.1255
R18934 VDD.n769 VDD.t123 23.1255
R18935 VDD.n770 VDD.n735 23.1255
R18936 VDD.n770 VDD.t123 23.1255
R18937 VDD.n745 VDD.n744 23.1255
R18938 VDD.n745 VDD.t123 23.1255
R18939 VDD.n888 VDD.n887 23.1255
R18940 VDD.n887 VDD.t123 23.1255
R18941 VDD.n739 VDD.n724 23.1255
R18942 VDD.t126 VDD.n724 23.1255
R18943 VDD.n742 VDD.n725 23.1255
R18944 VDD.t126 VDD.n725 23.1255
R18945 VDD.n757 VDD.n755 23.1255
R18946 VDD.n755 VDD.t123 23.1255
R18947 VDD.n766 VDD.n756 23.1255
R18948 VDD.n756 VDD.t123 23.1255
R18949 VDD.n761 VDD.n722 23.1255
R18950 VDD.t126 VDD.n722 23.1255
R18951 VDD.n758 VDD.n723 23.1255
R18952 VDD.t126 VDD.n723 23.1255
R18953 VDD.n811 VDD.n810 23.1255
R18954 VDD.n810 VDD.t123 23.1255
R18955 VDD.n814 VDD.n813 23.1255
R18956 VDD.n813 VDD.t123 23.1255
R18957 VDD.n806 VDD.n720 23.1255
R18958 VDD.t126 VDD.n720 23.1255
R18959 VDD.n809 VDD.n721 23.1255
R18960 VDD.t126 VDD.n721 23.1255
R18961 VDD.n827 VDD.n826 23.1255
R18962 VDD.n826 VDD.t123 23.1255
R18963 VDD.n830 VDD.n829 23.1255
R18964 VDD.n829 VDD.t123 23.1255
R18965 VDD.n822 VDD.n718 23.1255
R18966 VDD.t126 VDD.n718 23.1255
R18967 VDD.n825 VDD.n719 23.1255
R18968 VDD.t126 VDD.n719 23.1255
R18969 VDD.n834 VDD.n716 23.1255
R18970 VDD.t126 VDD.n716 23.1255
R18971 VDD.n838 VDD.n717 23.1255
R18972 VDD.t126 VDD.n717 23.1255
R18973 VDD.n850 VDD.n849 23.1255
R18974 VDD.n849 VDD.t123 23.1255
R18975 VDD.n853 VDD.n852 23.1255
R18976 VDD.n852 VDD.t123 23.1255
R18977 VDD.n845 VDD.n714 23.1255
R18978 VDD.t126 VDD.n714 23.1255
R18979 VDD.n848 VDD.n715 23.1255
R18980 VDD.t126 VDD.n715 23.1255
R18981 VDD.n866 VDD.n865 23.1255
R18982 VDD.n865 VDD.t123 23.1255
R18983 VDD.n869 VDD.n868 23.1255
R18984 VDD.n868 VDD.t123 23.1255
R18985 VDD.n861 VDD.n712 23.1255
R18986 VDD.t126 VDD.n712 23.1255
R18987 VDD.n864 VDD.n713 23.1255
R18988 VDD.t126 VDD.n713 23.1255
R18989 VDD.n778 VDD.n776 23.1255
R18990 VDD.n776 VDD.t123 23.1255
R18991 VDD.n876 VDD.n777 23.1255
R18992 VDD.n777 VDD.t123 23.1255
R18993 VDD.n782 VDD.n710 23.1255
R18994 VDD.t126 VDD.n710 23.1255
R18995 VDD.n779 VDD.n711 23.1255
R18996 VDD.t126 VDD.n711 23.1255
R18997 VDD.n793 VDD.n792 23.1255
R18998 VDD.n792 VDD.t123 23.1255
R18999 VDD.n796 VDD.n795 23.1255
R19000 VDD.n795 VDD.t123 23.1255
R19001 VDD.n788 VDD.n708 23.1255
R19002 VDD.t126 VDD.n708 23.1255
R19003 VDD.n791 VDD.n709 23.1255
R19004 VDD.t126 VDD.n709 23.1255
R19005 VDD.n879 VDD.n681 23.1255
R19006 VDD.t123 VDD.n681 23.1255
R19007 VDD.n880 VDD.n682 23.1255
R19008 VDD.t123 VDD.n682 23.1255
R19009 VDD.n726 VDD.n706 23.1255
R19010 VDD.t126 VDD.n706 23.1255
R19011 VDD.n727 VDD.n707 23.1255
R19012 VDD.t126 VDD.n707 23.1255
R19013 VDD.n748 VDD.n746 23.1255
R19014 VDD.n746 VDD.t123 23.1255
R19015 VDD.n749 VDD.n747 23.1255
R19016 VDD.n747 VDD.t123 23.1255
R19017 VDD.n703 VDD.n701 23.1255
R19018 VDD.t126 VDD.n701 23.1255
R19019 VDD.n901 VDD.n705 23.1255
R19020 VDD.n901 VDD.t126 23.1255
R19021 VDD.n696 VDD.n694 23.1255
R19022 VDD.n694 VDD.t123 23.1255
R19023 VDD.n697 VDD.n695 23.1255
R19024 VDD.n695 VDD.t123 23.1255
R19025 VDD.n900 VDD.n899 23.1255
R19026 VDD.t126 VDD.n900 23.1255
R19027 VDD.n897 VDD.n731 23.1255
R19028 VDD.t126 VDD.n731 23.1255
R19029 VDD.n1030 VDD.n1028 23.1255
R19030 VDD.n1028 VDD.t12 23.1255
R19031 VDD.n1029 VDD.n994 23.1255
R19032 VDD.n1029 VDD.t12 23.1255
R19033 VDD.n1004 VDD.n1003 23.1255
R19034 VDD.n1004 VDD.t12 23.1255
R19035 VDD.n1147 VDD.n1146 23.1255
R19036 VDD.n1146 VDD.t12 23.1255
R19037 VDD.n998 VDD.n983 23.1255
R19038 VDD.t51 VDD.n983 23.1255
R19039 VDD.n1001 VDD.n984 23.1255
R19040 VDD.t51 VDD.n984 23.1255
R19041 VDD.n1016 VDD.n1014 23.1255
R19042 VDD.n1014 VDD.t12 23.1255
R19043 VDD.n1025 VDD.n1015 23.1255
R19044 VDD.n1015 VDD.t12 23.1255
R19045 VDD.n1020 VDD.n981 23.1255
R19046 VDD.t51 VDD.n981 23.1255
R19047 VDD.n1017 VDD.n982 23.1255
R19048 VDD.t51 VDD.n982 23.1255
R19049 VDD.n1070 VDD.n1069 23.1255
R19050 VDD.n1069 VDD.t12 23.1255
R19051 VDD.n1073 VDD.n1072 23.1255
R19052 VDD.n1072 VDD.t12 23.1255
R19053 VDD.n1065 VDD.n979 23.1255
R19054 VDD.t51 VDD.n979 23.1255
R19055 VDD.n1068 VDD.n980 23.1255
R19056 VDD.t51 VDD.n980 23.1255
R19057 VDD.n1086 VDD.n1085 23.1255
R19058 VDD.n1085 VDD.t12 23.1255
R19059 VDD.n1089 VDD.n1088 23.1255
R19060 VDD.n1088 VDD.t12 23.1255
R19061 VDD.n1081 VDD.n977 23.1255
R19062 VDD.t51 VDD.n977 23.1255
R19063 VDD.n1084 VDD.n978 23.1255
R19064 VDD.t51 VDD.n978 23.1255
R19065 VDD.n1093 VDD.n975 23.1255
R19066 VDD.t51 VDD.n975 23.1255
R19067 VDD.n1097 VDD.n976 23.1255
R19068 VDD.t51 VDD.n976 23.1255
R19069 VDD.n1109 VDD.n1108 23.1255
R19070 VDD.n1108 VDD.t12 23.1255
R19071 VDD.n1112 VDD.n1111 23.1255
R19072 VDD.n1111 VDD.t12 23.1255
R19073 VDD.n1104 VDD.n973 23.1255
R19074 VDD.t51 VDD.n973 23.1255
R19075 VDD.n1107 VDD.n974 23.1255
R19076 VDD.t51 VDD.n974 23.1255
R19077 VDD.n1125 VDD.n1124 23.1255
R19078 VDD.n1124 VDD.t12 23.1255
R19079 VDD.n1128 VDD.n1127 23.1255
R19080 VDD.n1127 VDD.t12 23.1255
R19081 VDD.n1120 VDD.n971 23.1255
R19082 VDD.t51 VDD.n971 23.1255
R19083 VDD.n1123 VDD.n972 23.1255
R19084 VDD.t51 VDD.n972 23.1255
R19085 VDD.n1037 VDD.n1035 23.1255
R19086 VDD.n1035 VDD.t12 23.1255
R19087 VDD.n1135 VDD.n1036 23.1255
R19088 VDD.n1036 VDD.t12 23.1255
R19089 VDD.n1041 VDD.n969 23.1255
R19090 VDD.t51 VDD.n969 23.1255
R19091 VDD.n1038 VDD.n970 23.1255
R19092 VDD.t51 VDD.n970 23.1255
R19093 VDD.n1052 VDD.n1051 23.1255
R19094 VDD.n1051 VDD.t12 23.1255
R19095 VDD.n1055 VDD.n1054 23.1255
R19096 VDD.n1054 VDD.t12 23.1255
R19097 VDD.n1047 VDD.n967 23.1255
R19098 VDD.t51 VDD.n967 23.1255
R19099 VDD.n1050 VDD.n968 23.1255
R19100 VDD.t51 VDD.n968 23.1255
R19101 VDD.n1138 VDD.n940 23.1255
R19102 VDD.t12 VDD.n940 23.1255
R19103 VDD.n1139 VDD.n941 23.1255
R19104 VDD.t12 VDD.n941 23.1255
R19105 VDD.n985 VDD.n965 23.1255
R19106 VDD.t51 VDD.n965 23.1255
R19107 VDD.n986 VDD.n966 23.1255
R19108 VDD.t51 VDD.n966 23.1255
R19109 VDD.n1007 VDD.n1005 23.1255
R19110 VDD.n1005 VDD.t12 23.1255
R19111 VDD.n1008 VDD.n1006 23.1255
R19112 VDD.n1006 VDD.t12 23.1255
R19113 VDD.n962 VDD.n960 23.1255
R19114 VDD.t51 VDD.n960 23.1255
R19115 VDD.n1160 VDD.n964 23.1255
R19116 VDD.n1160 VDD.t51 23.1255
R19117 VDD.n955 VDD.n953 23.1255
R19118 VDD.n953 VDD.t12 23.1255
R19119 VDD.n956 VDD.n954 23.1255
R19120 VDD.n954 VDD.t12 23.1255
R19121 VDD.n1159 VDD.n1158 23.1255
R19122 VDD.t51 VDD.n1159 23.1255
R19123 VDD.n1156 VDD.n990 23.1255
R19124 VDD.t51 VDD.n990 23.1255
R19125 VDD.n1289 VDD.n1287 23.1255
R19126 VDD.n1287 VDD.t111 23.1255
R19127 VDD.n1288 VDD.n1253 23.1255
R19128 VDD.n1288 VDD.t111 23.1255
R19129 VDD.n1263 VDD.n1262 23.1255
R19130 VDD.n1263 VDD.t111 23.1255
R19131 VDD.n1406 VDD.n1405 23.1255
R19132 VDD.n1405 VDD.t111 23.1255
R19133 VDD.n1257 VDD.n1242 23.1255
R19134 VDD.t53 VDD.n1242 23.1255
R19135 VDD.n1260 VDD.n1243 23.1255
R19136 VDD.t53 VDD.n1243 23.1255
R19137 VDD.n1275 VDD.n1273 23.1255
R19138 VDD.n1273 VDD.t111 23.1255
R19139 VDD.n1284 VDD.n1274 23.1255
R19140 VDD.n1274 VDD.t111 23.1255
R19141 VDD.n1279 VDD.n1240 23.1255
R19142 VDD.t53 VDD.n1240 23.1255
R19143 VDD.n1276 VDD.n1241 23.1255
R19144 VDD.t53 VDD.n1241 23.1255
R19145 VDD.n1329 VDD.n1328 23.1255
R19146 VDD.n1328 VDD.t111 23.1255
R19147 VDD.n1332 VDD.n1331 23.1255
R19148 VDD.n1331 VDD.t111 23.1255
R19149 VDD.n1324 VDD.n1238 23.1255
R19150 VDD.t53 VDD.n1238 23.1255
R19151 VDD.n1327 VDD.n1239 23.1255
R19152 VDD.t53 VDD.n1239 23.1255
R19153 VDD.n1345 VDD.n1344 23.1255
R19154 VDD.n1344 VDD.t111 23.1255
R19155 VDD.n1348 VDD.n1347 23.1255
R19156 VDD.n1347 VDD.t111 23.1255
R19157 VDD.n1340 VDD.n1236 23.1255
R19158 VDD.t53 VDD.n1236 23.1255
R19159 VDD.n1343 VDD.n1237 23.1255
R19160 VDD.t53 VDD.n1237 23.1255
R19161 VDD.n1352 VDD.n1234 23.1255
R19162 VDD.t53 VDD.n1234 23.1255
R19163 VDD.n1356 VDD.n1235 23.1255
R19164 VDD.t53 VDD.n1235 23.1255
R19165 VDD.n1368 VDD.n1367 23.1255
R19166 VDD.n1367 VDD.t111 23.1255
R19167 VDD.n1371 VDD.n1370 23.1255
R19168 VDD.n1370 VDD.t111 23.1255
R19169 VDD.n1363 VDD.n1232 23.1255
R19170 VDD.t53 VDD.n1232 23.1255
R19171 VDD.n1366 VDD.n1233 23.1255
R19172 VDD.t53 VDD.n1233 23.1255
R19173 VDD.n1384 VDD.n1383 23.1255
R19174 VDD.n1383 VDD.t111 23.1255
R19175 VDD.n1387 VDD.n1386 23.1255
R19176 VDD.n1386 VDD.t111 23.1255
R19177 VDD.n1379 VDD.n1230 23.1255
R19178 VDD.t53 VDD.n1230 23.1255
R19179 VDD.n1382 VDD.n1231 23.1255
R19180 VDD.t53 VDD.n1231 23.1255
R19181 VDD.n1296 VDD.n1294 23.1255
R19182 VDD.n1294 VDD.t111 23.1255
R19183 VDD.n1394 VDD.n1295 23.1255
R19184 VDD.n1295 VDD.t111 23.1255
R19185 VDD.n1300 VDD.n1228 23.1255
R19186 VDD.t53 VDD.n1228 23.1255
R19187 VDD.n1297 VDD.n1229 23.1255
R19188 VDD.t53 VDD.n1229 23.1255
R19189 VDD.n1311 VDD.n1310 23.1255
R19190 VDD.n1310 VDD.t111 23.1255
R19191 VDD.n1314 VDD.n1313 23.1255
R19192 VDD.n1313 VDD.t111 23.1255
R19193 VDD.n1306 VDD.n1226 23.1255
R19194 VDD.t53 VDD.n1226 23.1255
R19195 VDD.n1309 VDD.n1227 23.1255
R19196 VDD.t53 VDD.n1227 23.1255
R19197 VDD.n1397 VDD.n1199 23.1255
R19198 VDD.t111 VDD.n1199 23.1255
R19199 VDD.n1398 VDD.n1200 23.1255
R19200 VDD.t111 VDD.n1200 23.1255
R19201 VDD.n1244 VDD.n1224 23.1255
R19202 VDD.t53 VDD.n1224 23.1255
R19203 VDD.n1245 VDD.n1225 23.1255
R19204 VDD.t53 VDD.n1225 23.1255
R19205 VDD.n1266 VDD.n1264 23.1255
R19206 VDD.n1264 VDD.t111 23.1255
R19207 VDD.n1267 VDD.n1265 23.1255
R19208 VDD.n1265 VDD.t111 23.1255
R19209 VDD.n1221 VDD.n1219 23.1255
R19210 VDD.t53 VDD.n1219 23.1255
R19211 VDD.n1419 VDD.n1223 23.1255
R19212 VDD.n1419 VDD.t53 23.1255
R19213 VDD.n1214 VDD.n1212 23.1255
R19214 VDD.n1212 VDD.t111 23.1255
R19215 VDD.n1215 VDD.n1213 23.1255
R19216 VDD.n1213 VDD.t111 23.1255
R19217 VDD.n1418 VDD.n1417 23.1255
R19218 VDD.t53 VDD.n1418 23.1255
R19219 VDD.n1415 VDD.n1249 23.1255
R19220 VDD.t53 VDD.n1249 23.1255
R19221 VDD.n1548 VDD.n1546 23.1255
R19222 VDD.n1546 VDD.t147 23.1255
R19223 VDD.n1547 VDD.n1512 23.1255
R19224 VDD.n1547 VDD.t147 23.1255
R19225 VDD.n1522 VDD.n1521 23.1255
R19226 VDD.n1522 VDD.t147 23.1255
R19227 VDD.n1665 VDD.n1664 23.1255
R19228 VDD.n1664 VDD.t147 23.1255
R19229 VDD.n1516 VDD.n1501 23.1255
R19230 VDD.t46 VDD.n1501 23.1255
R19231 VDD.n1519 VDD.n1502 23.1255
R19232 VDD.t46 VDD.n1502 23.1255
R19233 VDD.n1534 VDD.n1532 23.1255
R19234 VDD.n1532 VDD.t147 23.1255
R19235 VDD.n1543 VDD.n1533 23.1255
R19236 VDD.n1533 VDD.t147 23.1255
R19237 VDD.n1538 VDD.n1499 23.1255
R19238 VDD.t46 VDD.n1499 23.1255
R19239 VDD.n1535 VDD.n1500 23.1255
R19240 VDD.t46 VDD.n1500 23.1255
R19241 VDD.n1588 VDD.n1587 23.1255
R19242 VDD.n1587 VDD.t147 23.1255
R19243 VDD.n1591 VDD.n1590 23.1255
R19244 VDD.n1590 VDD.t147 23.1255
R19245 VDD.n1583 VDD.n1497 23.1255
R19246 VDD.t46 VDD.n1497 23.1255
R19247 VDD.n1586 VDD.n1498 23.1255
R19248 VDD.t46 VDD.n1498 23.1255
R19249 VDD.n1604 VDD.n1603 23.1255
R19250 VDD.n1603 VDD.t147 23.1255
R19251 VDD.n1607 VDD.n1606 23.1255
R19252 VDD.n1606 VDD.t147 23.1255
R19253 VDD.n1599 VDD.n1495 23.1255
R19254 VDD.t46 VDD.n1495 23.1255
R19255 VDD.n1602 VDD.n1496 23.1255
R19256 VDD.t46 VDD.n1496 23.1255
R19257 VDD.n1611 VDD.n1493 23.1255
R19258 VDD.t46 VDD.n1493 23.1255
R19259 VDD.n1615 VDD.n1494 23.1255
R19260 VDD.t46 VDD.n1494 23.1255
R19261 VDD.n1627 VDD.n1626 23.1255
R19262 VDD.n1626 VDD.t147 23.1255
R19263 VDD.n1630 VDD.n1629 23.1255
R19264 VDD.n1629 VDD.t147 23.1255
R19265 VDD.n1622 VDD.n1491 23.1255
R19266 VDD.t46 VDD.n1491 23.1255
R19267 VDD.n1625 VDD.n1492 23.1255
R19268 VDD.t46 VDD.n1492 23.1255
R19269 VDD.n1643 VDD.n1642 23.1255
R19270 VDD.n1642 VDD.t147 23.1255
R19271 VDD.n1646 VDD.n1645 23.1255
R19272 VDD.n1645 VDD.t147 23.1255
R19273 VDD.n1638 VDD.n1489 23.1255
R19274 VDD.t46 VDD.n1489 23.1255
R19275 VDD.n1641 VDD.n1490 23.1255
R19276 VDD.t46 VDD.n1490 23.1255
R19277 VDD.n1555 VDD.n1553 23.1255
R19278 VDD.n1553 VDD.t147 23.1255
R19279 VDD.n1653 VDD.n1554 23.1255
R19280 VDD.n1554 VDD.t147 23.1255
R19281 VDD.n1559 VDD.n1487 23.1255
R19282 VDD.t46 VDD.n1487 23.1255
R19283 VDD.n1556 VDD.n1488 23.1255
R19284 VDD.t46 VDD.n1488 23.1255
R19285 VDD.n1570 VDD.n1569 23.1255
R19286 VDD.n1569 VDD.t147 23.1255
R19287 VDD.n1573 VDD.n1572 23.1255
R19288 VDD.n1572 VDD.t147 23.1255
R19289 VDD.n1565 VDD.n1485 23.1255
R19290 VDD.t46 VDD.n1485 23.1255
R19291 VDD.n1568 VDD.n1486 23.1255
R19292 VDD.t46 VDD.n1486 23.1255
R19293 VDD.n1656 VDD.n1458 23.1255
R19294 VDD.t147 VDD.n1458 23.1255
R19295 VDD.n1657 VDD.n1459 23.1255
R19296 VDD.t147 VDD.n1459 23.1255
R19297 VDD.n1503 VDD.n1483 23.1255
R19298 VDD.t46 VDD.n1483 23.1255
R19299 VDD.n1504 VDD.n1484 23.1255
R19300 VDD.t46 VDD.n1484 23.1255
R19301 VDD.n1525 VDD.n1523 23.1255
R19302 VDD.n1523 VDD.t147 23.1255
R19303 VDD.n1526 VDD.n1524 23.1255
R19304 VDD.n1524 VDD.t147 23.1255
R19305 VDD.n1480 VDD.n1478 23.1255
R19306 VDD.t46 VDD.n1478 23.1255
R19307 VDD.n1678 VDD.n1482 23.1255
R19308 VDD.n1678 VDD.t46 23.1255
R19309 VDD.n1473 VDD.n1471 23.1255
R19310 VDD.n1471 VDD.t147 23.1255
R19311 VDD.n1474 VDD.n1472 23.1255
R19312 VDD.n1472 VDD.t147 23.1255
R19313 VDD.n1677 VDD.n1676 23.1255
R19314 VDD.t46 VDD.n1677 23.1255
R19315 VDD.n1674 VDD.n1508 23.1255
R19316 VDD.t46 VDD.n1508 23.1255
R19317 VDD.n1807 VDD.n1805 23.1255
R19318 VDD.n1805 VDD.t22 23.1255
R19319 VDD.n1806 VDD.n1771 23.1255
R19320 VDD.n1806 VDD.t22 23.1255
R19321 VDD.n1781 VDD.n1780 23.1255
R19322 VDD.n1781 VDD.t22 23.1255
R19323 VDD.n1924 VDD.n1923 23.1255
R19324 VDD.n1923 VDD.t22 23.1255
R19325 VDD.n1775 VDD.n1760 23.1255
R19326 VDD.t140 VDD.n1760 23.1255
R19327 VDD.n1778 VDD.n1761 23.1255
R19328 VDD.t140 VDD.n1761 23.1255
R19329 VDD.n1793 VDD.n1791 23.1255
R19330 VDD.n1791 VDD.t22 23.1255
R19331 VDD.n1802 VDD.n1792 23.1255
R19332 VDD.n1792 VDD.t22 23.1255
R19333 VDD.n1797 VDD.n1758 23.1255
R19334 VDD.t140 VDD.n1758 23.1255
R19335 VDD.n1794 VDD.n1759 23.1255
R19336 VDD.t140 VDD.n1759 23.1255
R19337 VDD.n1847 VDD.n1846 23.1255
R19338 VDD.n1846 VDD.t22 23.1255
R19339 VDD.n1850 VDD.n1849 23.1255
R19340 VDD.n1849 VDD.t22 23.1255
R19341 VDD.n1842 VDD.n1756 23.1255
R19342 VDD.t140 VDD.n1756 23.1255
R19343 VDD.n1845 VDD.n1757 23.1255
R19344 VDD.t140 VDD.n1757 23.1255
R19345 VDD.n1863 VDD.n1862 23.1255
R19346 VDD.n1862 VDD.t22 23.1255
R19347 VDD.n1866 VDD.n1865 23.1255
R19348 VDD.n1865 VDD.t22 23.1255
R19349 VDD.n1858 VDD.n1754 23.1255
R19350 VDD.t140 VDD.n1754 23.1255
R19351 VDD.n1861 VDD.n1755 23.1255
R19352 VDD.t140 VDD.n1755 23.1255
R19353 VDD.n1870 VDD.n1752 23.1255
R19354 VDD.t140 VDD.n1752 23.1255
R19355 VDD.n1874 VDD.n1753 23.1255
R19356 VDD.t140 VDD.n1753 23.1255
R19357 VDD.n1886 VDD.n1885 23.1255
R19358 VDD.n1885 VDD.t22 23.1255
R19359 VDD.n1889 VDD.n1888 23.1255
R19360 VDD.n1888 VDD.t22 23.1255
R19361 VDD.n1881 VDD.n1750 23.1255
R19362 VDD.t140 VDD.n1750 23.1255
R19363 VDD.n1884 VDD.n1751 23.1255
R19364 VDD.t140 VDD.n1751 23.1255
R19365 VDD.n1902 VDD.n1901 23.1255
R19366 VDD.n1901 VDD.t22 23.1255
R19367 VDD.n1905 VDD.n1904 23.1255
R19368 VDD.n1904 VDD.t22 23.1255
R19369 VDD.n1897 VDD.n1748 23.1255
R19370 VDD.t140 VDD.n1748 23.1255
R19371 VDD.n1900 VDD.n1749 23.1255
R19372 VDD.t140 VDD.n1749 23.1255
R19373 VDD.n1814 VDD.n1812 23.1255
R19374 VDD.n1812 VDD.t22 23.1255
R19375 VDD.n1912 VDD.n1813 23.1255
R19376 VDD.n1813 VDD.t22 23.1255
R19377 VDD.n1818 VDD.n1746 23.1255
R19378 VDD.t140 VDD.n1746 23.1255
R19379 VDD.n1815 VDD.n1747 23.1255
R19380 VDD.t140 VDD.n1747 23.1255
R19381 VDD.n1829 VDD.n1828 23.1255
R19382 VDD.n1828 VDD.t22 23.1255
R19383 VDD.n1832 VDD.n1831 23.1255
R19384 VDD.n1831 VDD.t22 23.1255
R19385 VDD.n1824 VDD.n1744 23.1255
R19386 VDD.t140 VDD.n1744 23.1255
R19387 VDD.n1827 VDD.n1745 23.1255
R19388 VDD.t140 VDD.n1745 23.1255
R19389 VDD.n1915 VDD.n1717 23.1255
R19390 VDD.t22 VDD.n1717 23.1255
R19391 VDD.n1916 VDD.n1718 23.1255
R19392 VDD.t22 VDD.n1718 23.1255
R19393 VDD.n1762 VDD.n1742 23.1255
R19394 VDD.t140 VDD.n1742 23.1255
R19395 VDD.n1763 VDD.n1743 23.1255
R19396 VDD.t140 VDD.n1743 23.1255
R19397 VDD.n1784 VDD.n1782 23.1255
R19398 VDD.n1782 VDD.t22 23.1255
R19399 VDD.n1785 VDD.n1783 23.1255
R19400 VDD.n1783 VDD.t22 23.1255
R19401 VDD.n1739 VDD.n1737 23.1255
R19402 VDD.t140 VDD.n1737 23.1255
R19403 VDD.n1937 VDD.n1741 23.1255
R19404 VDD.n1937 VDD.t140 23.1255
R19405 VDD.n1732 VDD.n1730 23.1255
R19406 VDD.n1730 VDD.t22 23.1255
R19407 VDD.n1733 VDD.n1731 23.1255
R19408 VDD.n1731 VDD.t22 23.1255
R19409 VDD.n1936 VDD.n1935 23.1255
R19410 VDD.t140 VDD.n1936 23.1255
R19411 VDD.n1933 VDD.n1767 23.1255
R19412 VDD.t140 VDD.n1767 23.1255
R19413 VDD.n2066 VDD.n2064 23.1255
R19414 VDD.n2064 VDD.t156 23.1255
R19415 VDD.n2065 VDD.n2030 23.1255
R19416 VDD.n2065 VDD.t156 23.1255
R19417 VDD.n2040 VDD.n2039 23.1255
R19418 VDD.n2040 VDD.t156 23.1255
R19419 VDD.n2183 VDD.n2182 23.1255
R19420 VDD.n2182 VDD.t156 23.1255
R19421 VDD.n2034 VDD.n2019 23.1255
R19422 VDD.t35 VDD.n2019 23.1255
R19423 VDD.n2037 VDD.n2020 23.1255
R19424 VDD.t35 VDD.n2020 23.1255
R19425 VDD.n2052 VDD.n2050 23.1255
R19426 VDD.n2050 VDD.t156 23.1255
R19427 VDD.n2061 VDD.n2051 23.1255
R19428 VDD.n2051 VDD.t156 23.1255
R19429 VDD.n2056 VDD.n2017 23.1255
R19430 VDD.t35 VDD.n2017 23.1255
R19431 VDD.n2053 VDD.n2018 23.1255
R19432 VDD.t35 VDD.n2018 23.1255
R19433 VDD.n2106 VDD.n2105 23.1255
R19434 VDD.n2105 VDD.t156 23.1255
R19435 VDD.n2109 VDD.n2108 23.1255
R19436 VDD.n2108 VDD.t156 23.1255
R19437 VDD.n2101 VDD.n2015 23.1255
R19438 VDD.t35 VDD.n2015 23.1255
R19439 VDD.n2104 VDD.n2016 23.1255
R19440 VDD.t35 VDD.n2016 23.1255
R19441 VDD.n2122 VDD.n2121 23.1255
R19442 VDD.n2121 VDD.t156 23.1255
R19443 VDD.n2125 VDD.n2124 23.1255
R19444 VDD.n2124 VDD.t156 23.1255
R19445 VDD.n2117 VDD.n2013 23.1255
R19446 VDD.t35 VDD.n2013 23.1255
R19447 VDD.n2120 VDD.n2014 23.1255
R19448 VDD.t35 VDD.n2014 23.1255
R19449 VDD.n2129 VDD.n2011 23.1255
R19450 VDD.t35 VDD.n2011 23.1255
R19451 VDD.n2133 VDD.n2012 23.1255
R19452 VDD.t35 VDD.n2012 23.1255
R19453 VDD.n2145 VDD.n2144 23.1255
R19454 VDD.n2144 VDD.t156 23.1255
R19455 VDD.n2148 VDD.n2147 23.1255
R19456 VDD.n2147 VDD.t156 23.1255
R19457 VDD.n2140 VDD.n2009 23.1255
R19458 VDD.t35 VDD.n2009 23.1255
R19459 VDD.n2143 VDD.n2010 23.1255
R19460 VDD.t35 VDD.n2010 23.1255
R19461 VDD.n2161 VDD.n2160 23.1255
R19462 VDD.n2160 VDD.t156 23.1255
R19463 VDD.n2164 VDD.n2163 23.1255
R19464 VDD.n2163 VDD.t156 23.1255
R19465 VDD.n2156 VDD.n2007 23.1255
R19466 VDD.t35 VDD.n2007 23.1255
R19467 VDD.n2159 VDD.n2008 23.1255
R19468 VDD.t35 VDD.n2008 23.1255
R19469 VDD.n2073 VDD.n2071 23.1255
R19470 VDD.n2071 VDD.t156 23.1255
R19471 VDD.n2171 VDD.n2072 23.1255
R19472 VDD.n2072 VDD.t156 23.1255
R19473 VDD.n2077 VDD.n2005 23.1255
R19474 VDD.t35 VDD.n2005 23.1255
R19475 VDD.n2074 VDD.n2006 23.1255
R19476 VDD.t35 VDD.n2006 23.1255
R19477 VDD.n2088 VDD.n2087 23.1255
R19478 VDD.n2087 VDD.t156 23.1255
R19479 VDD.n2091 VDD.n2090 23.1255
R19480 VDD.n2090 VDD.t156 23.1255
R19481 VDD.n2083 VDD.n2003 23.1255
R19482 VDD.t35 VDD.n2003 23.1255
R19483 VDD.n2086 VDD.n2004 23.1255
R19484 VDD.t35 VDD.n2004 23.1255
R19485 VDD.n2174 VDD.n1976 23.1255
R19486 VDD.t156 VDD.n1976 23.1255
R19487 VDD.n2175 VDD.n1977 23.1255
R19488 VDD.t156 VDD.n1977 23.1255
R19489 VDD.n2021 VDD.n2001 23.1255
R19490 VDD.t35 VDD.n2001 23.1255
R19491 VDD.n2022 VDD.n2002 23.1255
R19492 VDD.t35 VDD.n2002 23.1255
R19493 VDD.n2043 VDD.n2041 23.1255
R19494 VDD.n2041 VDD.t156 23.1255
R19495 VDD.n2044 VDD.n2042 23.1255
R19496 VDD.n2042 VDD.t156 23.1255
R19497 VDD.n1998 VDD.n1996 23.1255
R19498 VDD.t35 VDD.n1996 23.1255
R19499 VDD.n2196 VDD.n2000 23.1255
R19500 VDD.n2196 VDD.t35 23.1255
R19501 VDD.n1991 VDD.n1989 23.1255
R19502 VDD.n1989 VDD.t156 23.1255
R19503 VDD.n1992 VDD.n1990 23.1255
R19504 VDD.n1990 VDD.t156 23.1255
R19505 VDD.n2195 VDD.n2194 23.1255
R19506 VDD.t35 VDD.n2195 23.1255
R19507 VDD.n2192 VDD.n2026 23.1255
R19508 VDD.t35 VDD.n2026 23.1255
R19509 VDD.n2325 VDD.n2323 23.1255
R19510 VDD.n2323 VDD.t213 23.1255
R19511 VDD.n2324 VDD.n2289 23.1255
R19512 VDD.n2324 VDD.t213 23.1255
R19513 VDD.n2299 VDD.n2298 23.1255
R19514 VDD.n2299 VDD.t213 23.1255
R19515 VDD.n2442 VDD.n2441 23.1255
R19516 VDD.n2441 VDD.t213 23.1255
R19517 VDD.n2293 VDD.n2278 23.1255
R19518 VDD.t29 VDD.n2278 23.1255
R19519 VDD.n2296 VDD.n2279 23.1255
R19520 VDD.t29 VDD.n2279 23.1255
R19521 VDD.n2311 VDD.n2309 23.1255
R19522 VDD.n2309 VDD.t213 23.1255
R19523 VDD.n2320 VDD.n2310 23.1255
R19524 VDD.n2310 VDD.t213 23.1255
R19525 VDD.n2315 VDD.n2276 23.1255
R19526 VDD.t29 VDD.n2276 23.1255
R19527 VDD.n2312 VDD.n2277 23.1255
R19528 VDD.t29 VDD.n2277 23.1255
R19529 VDD.n2365 VDD.n2364 23.1255
R19530 VDD.n2364 VDD.t213 23.1255
R19531 VDD.n2368 VDD.n2367 23.1255
R19532 VDD.n2367 VDD.t213 23.1255
R19533 VDD.n2360 VDD.n2274 23.1255
R19534 VDD.t29 VDD.n2274 23.1255
R19535 VDD.n2363 VDD.n2275 23.1255
R19536 VDD.t29 VDD.n2275 23.1255
R19537 VDD.n2381 VDD.n2380 23.1255
R19538 VDD.n2380 VDD.t213 23.1255
R19539 VDD.n2384 VDD.n2383 23.1255
R19540 VDD.n2383 VDD.t213 23.1255
R19541 VDD.n2376 VDD.n2272 23.1255
R19542 VDD.t29 VDD.n2272 23.1255
R19543 VDD.n2379 VDD.n2273 23.1255
R19544 VDD.t29 VDD.n2273 23.1255
R19545 VDD.n2388 VDD.n2270 23.1255
R19546 VDD.t29 VDD.n2270 23.1255
R19547 VDD.n2392 VDD.n2271 23.1255
R19548 VDD.t29 VDD.n2271 23.1255
R19549 VDD.n2404 VDD.n2403 23.1255
R19550 VDD.n2403 VDD.t213 23.1255
R19551 VDD.n2407 VDD.n2406 23.1255
R19552 VDD.n2406 VDD.t213 23.1255
R19553 VDD.n2399 VDD.n2268 23.1255
R19554 VDD.t29 VDD.n2268 23.1255
R19555 VDD.n2402 VDD.n2269 23.1255
R19556 VDD.t29 VDD.n2269 23.1255
R19557 VDD.n2420 VDD.n2419 23.1255
R19558 VDD.n2419 VDD.t213 23.1255
R19559 VDD.n2423 VDD.n2422 23.1255
R19560 VDD.n2422 VDD.t213 23.1255
R19561 VDD.n2415 VDD.n2266 23.1255
R19562 VDD.t29 VDD.n2266 23.1255
R19563 VDD.n2418 VDD.n2267 23.1255
R19564 VDD.t29 VDD.n2267 23.1255
R19565 VDD.n2332 VDD.n2330 23.1255
R19566 VDD.n2330 VDD.t213 23.1255
R19567 VDD.n2430 VDD.n2331 23.1255
R19568 VDD.n2331 VDD.t213 23.1255
R19569 VDD.n2336 VDD.n2264 23.1255
R19570 VDD.t29 VDD.n2264 23.1255
R19571 VDD.n2333 VDD.n2265 23.1255
R19572 VDD.t29 VDD.n2265 23.1255
R19573 VDD.n2347 VDD.n2346 23.1255
R19574 VDD.n2346 VDD.t213 23.1255
R19575 VDD.n2350 VDD.n2349 23.1255
R19576 VDD.n2349 VDD.t213 23.1255
R19577 VDD.n2342 VDD.n2262 23.1255
R19578 VDD.t29 VDD.n2262 23.1255
R19579 VDD.n2345 VDD.n2263 23.1255
R19580 VDD.t29 VDD.n2263 23.1255
R19581 VDD.n2433 VDD.n2235 23.1255
R19582 VDD.t213 VDD.n2235 23.1255
R19583 VDD.n2434 VDD.n2236 23.1255
R19584 VDD.t213 VDD.n2236 23.1255
R19585 VDD.n2280 VDD.n2260 23.1255
R19586 VDD.t29 VDD.n2260 23.1255
R19587 VDD.n2281 VDD.n2261 23.1255
R19588 VDD.t29 VDD.n2261 23.1255
R19589 VDD.n2302 VDD.n2300 23.1255
R19590 VDD.n2300 VDD.t213 23.1255
R19591 VDD.n2303 VDD.n2301 23.1255
R19592 VDD.n2301 VDD.t213 23.1255
R19593 VDD.n2257 VDD.n2255 23.1255
R19594 VDD.t29 VDD.n2255 23.1255
R19595 VDD.n2455 VDD.n2259 23.1255
R19596 VDD.n2455 VDD.t29 23.1255
R19597 VDD.n2250 VDD.n2248 23.1255
R19598 VDD.n2248 VDD.t213 23.1255
R19599 VDD.n2251 VDD.n2249 23.1255
R19600 VDD.n2249 VDD.t213 23.1255
R19601 VDD.n2454 VDD.n2453 23.1255
R19602 VDD.t29 VDD.n2454 23.1255
R19603 VDD.n2451 VDD.n2285 23.1255
R19604 VDD.t29 VDD.n2285 23.1255
R19605 VDD.n2584 VDD.n2582 23.1255
R19606 VDD.n2582 VDD.t72 23.1255
R19607 VDD.n2583 VDD.n2548 23.1255
R19608 VDD.n2583 VDD.t72 23.1255
R19609 VDD.n2558 VDD.n2557 23.1255
R19610 VDD.n2558 VDD.t72 23.1255
R19611 VDD.n2701 VDD.n2700 23.1255
R19612 VDD.n2700 VDD.t72 23.1255
R19613 VDD.n2552 VDD.n2537 23.1255
R19614 VDD.t83 VDD.n2537 23.1255
R19615 VDD.n2555 VDD.n2538 23.1255
R19616 VDD.t83 VDD.n2538 23.1255
R19617 VDD.n2570 VDD.n2568 23.1255
R19618 VDD.n2568 VDD.t72 23.1255
R19619 VDD.n2579 VDD.n2569 23.1255
R19620 VDD.n2569 VDD.t72 23.1255
R19621 VDD.n2574 VDD.n2535 23.1255
R19622 VDD.t83 VDD.n2535 23.1255
R19623 VDD.n2571 VDD.n2536 23.1255
R19624 VDD.t83 VDD.n2536 23.1255
R19625 VDD.n2624 VDD.n2623 23.1255
R19626 VDD.n2623 VDD.t72 23.1255
R19627 VDD.n2627 VDD.n2626 23.1255
R19628 VDD.n2626 VDD.t72 23.1255
R19629 VDD.n2619 VDD.n2533 23.1255
R19630 VDD.t83 VDD.n2533 23.1255
R19631 VDD.n2622 VDD.n2534 23.1255
R19632 VDD.t83 VDD.n2534 23.1255
R19633 VDD.n2640 VDD.n2639 23.1255
R19634 VDD.n2639 VDD.t72 23.1255
R19635 VDD.n2643 VDD.n2642 23.1255
R19636 VDD.n2642 VDD.t72 23.1255
R19637 VDD.n2635 VDD.n2531 23.1255
R19638 VDD.t83 VDD.n2531 23.1255
R19639 VDD.n2638 VDD.n2532 23.1255
R19640 VDD.t83 VDD.n2532 23.1255
R19641 VDD.n2647 VDD.n2529 23.1255
R19642 VDD.t83 VDD.n2529 23.1255
R19643 VDD.n2651 VDD.n2530 23.1255
R19644 VDD.t83 VDD.n2530 23.1255
R19645 VDD.n2663 VDD.n2662 23.1255
R19646 VDD.n2662 VDD.t72 23.1255
R19647 VDD.n2666 VDD.n2665 23.1255
R19648 VDD.n2665 VDD.t72 23.1255
R19649 VDD.n2658 VDD.n2527 23.1255
R19650 VDD.t83 VDD.n2527 23.1255
R19651 VDD.n2661 VDD.n2528 23.1255
R19652 VDD.t83 VDD.n2528 23.1255
R19653 VDD.n2679 VDD.n2678 23.1255
R19654 VDD.n2678 VDD.t72 23.1255
R19655 VDD.n2682 VDD.n2681 23.1255
R19656 VDD.n2681 VDD.t72 23.1255
R19657 VDD.n2674 VDD.n2525 23.1255
R19658 VDD.t83 VDD.n2525 23.1255
R19659 VDD.n2677 VDD.n2526 23.1255
R19660 VDD.t83 VDD.n2526 23.1255
R19661 VDD.n2591 VDD.n2589 23.1255
R19662 VDD.n2589 VDD.t72 23.1255
R19663 VDD.n2689 VDD.n2590 23.1255
R19664 VDD.n2590 VDD.t72 23.1255
R19665 VDD.n2595 VDD.n2523 23.1255
R19666 VDD.t83 VDD.n2523 23.1255
R19667 VDD.n2592 VDD.n2524 23.1255
R19668 VDD.t83 VDD.n2524 23.1255
R19669 VDD.n2606 VDD.n2605 23.1255
R19670 VDD.n2605 VDD.t72 23.1255
R19671 VDD.n2609 VDD.n2608 23.1255
R19672 VDD.n2608 VDD.t72 23.1255
R19673 VDD.n2601 VDD.n2521 23.1255
R19674 VDD.t83 VDD.n2521 23.1255
R19675 VDD.n2604 VDD.n2522 23.1255
R19676 VDD.t83 VDD.n2522 23.1255
R19677 VDD.n2692 VDD.n2494 23.1255
R19678 VDD.t72 VDD.n2494 23.1255
R19679 VDD.n2693 VDD.n2495 23.1255
R19680 VDD.t72 VDD.n2495 23.1255
R19681 VDD.n2539 VDD.n2519 23.1255
R19682 VDD.t83 VDD.n2519 23.1255
R19683 VDD.n2540 VDD.n2520 23.1255
R19684 VDD.t83 VDD.n2520 23.1255
R19685 VDD.n2561 VDD.n2559 23.1255
R19686 VDD.n2559 VDD.t72 23.1255
R19687 VDD.n2562 VDD.n2560 23.1255
R19688 VDD.n2560 VDD.t72 23.1255
R19689 VDD.n2516 VDD.n2514 23.1255
R19690 VDD.t83 VDD.n2514 23.1255
R19691 VDD.n2714 VDD.n2518 23.1255
R19692 VDD.n2714 VDD.t83 23.1255
R19693 VDD.n2509 VDD.n2507 23.1255
R19694 VDD.n2507 VDD.t72 23.1255
R19695 VDD.n2510 VDD.n2508 23.1255
R19696 VDD.n2508 VDD.t72 23.1255
R19697 VDD.n2713 VDD.n2712 23.1255
R19698 VDD.t83 VDD.n2713 23.1255
R19699 VDD.n2710 VDD.n2544 23.1255
R19700 VDD.t83 VDD.n2544 23.1255
R19701 VDD.n2843 VDD.n2841 23.1255
R19702 VDD.n2841 VDD.t57 23.1255
R19703 VDD.n2842 VDD.n2807 23.1255
R19704 VDD.n2842 VDD.t57 23.1255
R19705 VDD.n2817 VDD.n2816 23.1255
R19706 VDD.n2817 VDD.t57 23.1255
R19707 VDD.n2960 VDD.n2959 23.1255
R19708 VDD.n2959 VDD.t57 23.1255
R19709 VDD.n2811 VDD.n2796 23.1255
R19710 VDD.t10 VDD.n2796 23.1255
R19711 VDD.n2814 VDD.n2797 23.1255
R19712 VDD.t10 VDD.n2797 23.1255
R19713 VDD.n2829 VDD.n2827 23.1255
R19714 VDD.n2827 VDD.t57 23.1255
R19715 VDD.n2838 VDD.n2828 23.1255
R19716 VDD.n2828 VDD.t57 23.1255
R19717 VDD.n2833 VDD.n2794 23.1255
R19718 VDD.t10 VDD.n2794 23.1255
R19719 VDD.n2830 VDD.n2795 23.1255
R19720 VDD.t10 VDD.n2795 23.1255
R19721 VDD.n2883 VDD.n2882 23.1255
R19722 VDD.n2882 VDD.t57 23.1255
R19723 VDD.n2886 VDD.n2885 23.1255
R19724 VDD.n2885 VDD.t57 23.1255
R19725 VDD.n2878 VDD.n2792 23.1255
R19726 VDD.t10 VDD.n2792 23.1255
R19727 VDD.n2881 VDD.n2793 23.1255
R19728 VDD.t10 VDD.n2793 23.1255
R19729 VDD.n2899 VDD.n2898 23.1255
R19730 VDD.n2898 VDD.t57 23.1255
R19731 VDD.n2902 VDD.n2901 23.1255
R19732 VDD.n2901 VDD.t57 23.1255
R19733 VDD.n2894 VDD.n2790 23.1255
R19734 VDD.t10 VDD.n2790 23.1255
R19735 VDD.n2897 VDD.n2791 23.1255
R19736 VDD.t10 VDD.n2791 23.1255
R19737 VDD.n2906 VDD.n2788 23.1255
R19738 VDD.t10 VDD.n2788 23.1255
R19739 VDD.n2910 VDD.n2789 23.1255
R19740 VDD.t10 VDD.n2789 23.1255
R19741 VDD.n2922 VDD.n2921 23.1255
R19742 VDD.n2921 VDD.t57 23.1255
R19743 VDD.n2925 VDD.n2924 23.1255
R19744 VDD.n2924 VDD.t57 23.1255
R19745 VDD.n2917 VDD.n2786 23.1255
R19746 VDD.t10 VDD.n2786 23.1255
R19747 VDD.n2920 VDD.n2787 23.1255
R19748 VDD.t10 VDD.n2787 23.1255
R19749 VDD.n2938 VDD.n2937 23.1255
R19750 VDD.n2937 VDD.t57 23.1255
R19751 VDD.n2941 VDD.n2940 23.1255
R19752 VDD.n2940 VDD.t57 23.1255
R19753 VDD.n2933 VDD.n2784 23.1255
R19754 VDD.t10 VDD.n2784 23.1255
R19755 VDD.n2936 VDD.n2785 23.1255
R19756 VDD.t10 VDD.n2785 23.1255
R19757 VDD.n2850 VDD.n2848 23.1255
R19758 VDD.n2848 VDD.t57 23.1255
R19759 VDD.n2948 VDD.n2849 23.1255
R19760 VDD.n2849 VDD.t57 23.1255
R19761 VDD.n2854 VDD.n2782 23.1255
R19762 VDD.t10 VDD.n2782 23.1255
R19763 VDD.n2851 VDD.n2783 23.1255
R19764 VDD.t10 VDD.n2783 23.1255
R19765 VDD.n2865 VDD.n2864 23.1255
R19766 VDD.n2864 VDD.t57 23.1255
R19767 VDD.n2868 VDD.n2867 23.1255
R19768 VDD.n2867 VDD.t57 23.1255
R19769 VDD.n2860 VDD.n2780 23.1255
R19770 VDD.t10 VDD.n2780 23.1255
R19771 VDD.n2863 VDD.n2781 23.1255
R19772 VDD.t10 VDD.n2781 23.1255
R19773 VDD.n2951 VDD.n2753 23.1255
R19774 VDD.t57 VDD.n2753 23.1255
R19775 VDD.n2952 VDD.n2754 23.1255
R19776 VDD.t57 VDD.n2754 23.1255
R19777 VDD.n2798 VDD.n2778 23.1255
R19778 VDD.t10 VDD.n2778 23.1255
R19779 VDD.n2799 VDD.n2779 23.1255
R19780 VDD.t10 VDD.n2779 23.1255
R19781 VDD.n2820 VDD.n2818 23.1255
R19782 VDD.n2818 VDD.t57 23.1255
R19783 VDD.n2821 VDD.n2819 23.1255
R19784 VDD.n2819 VDD.t57 23.1255
R19785 VDD.n2775 VDD.n2773 23.1255
R19786 VDD.t10 VDD.n2773 23.1255
R19787 VDD.n2973 VDD.n2777 23.1255
R19788 VDD.n2973 VDD.t10 23.1255
R19789 VDD.n2768 VDD.n2766 23.1255
R19790 VDD.n2766 VDD.t57 23.1255
R19791 VDD.n2769 VDD.n2767 23.1255
R19792 VDD.n2767 VDD.t57 23.1255
R19793 VDD.n2972 VDD.n2971 23.1255
R19794 VDD.t10 VDD.n2972 23.1255
R19795 VDD.n2969 VDD.n2803 23.1255
R19796 VDD.t10 VDD.n2803 23.1255
R19797 VDD.n3102 VDD.n3100 23.1255
R19798 VDD.n3100 VDD.t48 23.1255
R19799 VDD.n3101 VDD.n3066 23.1255
R19800 VDD.n3101 VDD.t48 23.1255
R19801 VDD.n3076 VDD.n3075 23.1255
R19802 VDD.n3076 VDD.t48 23.1255
R19803 VDD.n3219 VDD.n3218 23.1255
R19804 VDD.n3218 VDD.t48 23.1255
R19805 VDD.n3070 VDD.n3055 23.1255
R19806 VDD.t55 VDD.n3055 23.1255
R19807 VDD.n3073 VDD.n3056 23.1255
R19808 VDD.t55 VDD.n3056 23.1255
R19809 VDD.n3088 VDD.n3086 23.1255
R19810 VDD.n3086 VDD.t48 23.1255
R19811 VDD.n3097 VDD.n3087 23.1255
R19812 VDD.n3087 VDD.t48 23.1255
R19813 VDD.n3092 VDD.n3053 23.1255
R19814 VDD.t55 VDD.n3053 23.1255
R19815 VDD.n3089 VDD.n3054 23.1255
R19816 VDD.t55 VDD.n3054 23.1255
R19817 VDD.n3142 VDD.n3141 23.1255
R19818 VDD.n3141 VDD.t48 23.1255
R19819 VDD.n3145 VDD.n3144 23.1255
R19820 VDD.n3144 VDD.t48 23.1255
R19821 VDD.n3137 VDD.n3051 23.1255
R19822 VDD.t55 VDD.n3051 23.1255
R19823 VDD.n3140 VDD.n3052 23.1255
R19824 VDD.t55 VDD.n3052 23.1255
R19825 VDD.n3158 VDD.n3157 23.1255
R19826 VDD.n3157 VDD.t48 23.1255
R19827 VDD.n3161 VDD.n3160 23.1255
R19828 VDD.n3160 VDD.t48 23.1255
R19829 VDD.n3153 VDD.n3049 23.1255
R19830 VDD.t55 VDD.n3049 23.1255
R19831 VDD.n3156 VDD.n3050 23.1255
R19832 VDD.t55 VDD.n3050 23.1255
R19833 VDD.n3165 VDD.n3047 23.1255
R19834 VDD.t55 VDD.n3047 23.1255
R19835 VDD.n3169 VDD.n3048 23.1255
R19836 VDD.t55 VDD.n3048 23.1255
R19837 VDD.n3181 VDD.n3180 23.1255
R19838 VDD.n3180 VDD.t48 23.1255
R19839 VDD.n3184 VDD.n3183 23.1255
R19840 VDD.n3183 VDD.t48 23.1255
R19841 VDD.n3176 VDD.n3045 23.1255
R19842 VDD.t55 VDD.n3045 23.1255
R19843 VDD.n3179 VDD.n3046 23.1255
R19844 VDD.t55 VDD.n3046 23.1255
R19845 VDD.n3197 VDD.n3196 23.1255
R19846 VDD.n3196 VDD.t48 23.1255
R19847 VDD.n3200 VDD.n3199 23.1255
R19848 VDD.n3199 VDD.t48 23.1255
R19849 VDD.n3192 VDD.n3043 23.1255
R19850 VDD.t55 VDD.n3043 23.1255
R19851 VDD.n3195 VDD.n3044 23.1255
R19852 VDD.t55 VDD.n3044 23.1255
R19853 VDD.n3109 VDD.n3107 23.1255
R19854 VDD.n3107 VDD.t48 23.1255
R19855 VDD.n3207 VDD.n3108 23.1255
R19856 VDD.n3108 VDD.t48 23.1255
R19857 VDD.n3113 VDD.n3041 23.1255
R19858 VDD.t55 VDD.n3041 23.1255
R19859 VDD.n3110 VDD.n3042 23.1255
R19860 VDD.t55 VDD.n3042 23.1255
R19861 VDD.n3124 VDD.n3123 23.1255
R19862 VDD.n3123 VDD.t48 23.1255
R19863 VDD.n3127 VDD.n3126 23.1255
R19864 VDD.n3126 VDD.t48 23.1255
R19865 VDD.n3119 VDD.n3039 23.1255
R19866 VDD.t55 VDD.n3039 23.1255
R19867 VDD.n3122 VDD.n3040 23.1255
R19868 VDD.t55 VDD.n3040 23.1255
R19869 VDD.n3210 VDD.n3012 23.1255
R19870 VDD.t48 VDD.n3012 23.1255
R19871 VDD.n3211 VDD.n3013 23.1255
R19872 VDD.t48 VDD.n3013 23.1255
R19873 VDD.n3057 VDD.n3037 23.1255
R19874 VDD.t55 VDD.n3037 23.1255
R19875 VDD.n3058 VDD.n3038 23.1255
R19876 VDD.t55 VDD.n3038 23.1255
R19877 VDD.n3079 VDD.n3077 23.1255
R19878 VDD.n3077 VDD.t48 23.1255
R19879 VDD.n3080 VDD.n3078 23.1255
R19880 VDD.n3078 VDD.t48 23.1255
R19881 VDD.n3034 VDD.n3032 23.1255
R19882 VDD.t55 VDD.n3032 23.1255
R19883 VDD.n3232 VDD.n3036 23.1255
R19884 VDD.n3232 VDD.t55 23.1255
R19885 VDD.n3027 VDD.n3025 23.1255
R19886 VDD.n3025 VDD.t48 23.1255
R19887 VDD.n3028 VDD.n3026 23.1255
R19888 VDD.n3026 VDD.t48 23.1255
R19889 VDD.n3231 VDD.n3230 23.1255
R19890 VDD.t55 VDD.n3231 23.1255
R19891 VDD.n3228 VDD.n3062 23.1255
R19892 VDD.t55 VDD.n3062 23.1255
R19893 VDD.n3361 VDD.n3359 23.1255
R19894 VDD.n3359 VDD.t135 23.1255
R19895 VDD.n3360 VDD.n3325 23.1255
R19896 VDD.n3360 VDD.t135 23.1255
R19897 VDD.n3335 VDD.n3334 23.1255
R19898 VDD.n3335 VDD.t135 23.1255
R19899 VDD.n3478 VDD.n3477 23.1255
R19900 VDD.n3477 VDD.t135 23.1255
R19901 VDD.n3329 VDD.n3314 23.1255
R19902 VDD.t92 VDD.n3314 23.1255
R19903 VDD.n3332 VDD.n3315 23.1255
R19904 VDD.t92 VDD.n3315 23.1255
R19905 VDD.n3347 VDD.n3345 23.1255
R19906 VDD.n3345 VDD.t135 23.1255
R19907 VDD.n3356 VDD.n3346 23.1255
R19908 VDD.n3346 VDD.t135 23.1255
R19909 VDD.n3351 VDD.n3312 23.1255
R19910 VDD.t92 VDD.n3312 23.1255
R19911 VDD.n3348 VDD.n3313 23.1255
R19912 VDD.t92 VDD.n3313 23.1255
R19913 VDD.n3401 VDD.n3400 23.1255
R19914 VDD.n3400 VDD.t135 23.1255
R19915 VDD.n3404 VDD.n3403 23.1255
R19916 VDD.n3403 VDD.t135 23.1255
R19917 VDD.n3396 VDD.n3310 23.1255
R19918 VDD.t92 VDD.n3310 23.1255
R19919 VDD.n3399 VDD.n3311 23.1255
R19920 VDD.t92 VDD.n3311 23.1255
R19921 VDD.n3417 VDD.n3416 23.1255
R19922 VDD.n3416 VDD.t135 23.1255
R19923 VDD.n3420 VDD.n3419 23.1255
R19924 VDD.n3419 VDD.t135 23.1255
R19925 VDD.n3412 VDD.n3308 23.1255
R19926 VDD.t92 VDD.n3308 23.1255
R19927 VDD.n3415 VDD.n3309 23.1255
R19928 VDD.t92 VDD.n3309 23.1255
R19929 VDD.n3424 VDD.n3306 23.1255
R19930 VDD.t92 VDD.n3306 23.1255
R19931 VDD.n3428 VDD.n3307 23.1255
R19932 VDD.t92 VDD.n3307 23.1255
R19933 VDD.n3440 VDD.n3439 23.1255
R19934 VDD.n3439 VDD.t135 23.1255
R19935 VDD.n3443 VDD.n3442 23.1255
R19936 VDD.n3442 VDD.t135 23.1255
R19937 VDD.n3435 VDD.n3304 23.1255
R19938 VDD.t92 VDD.n3304 23.1255
R19939 VDD.n3438 VDD.n3305 23.1255
R19940 VDD.t92 VDD.n3305 23.1255
R19941 VDD.n3456 VDD.n3455 23.1255
R19942 VDD.n3455 VDD.t135 23.1255
R19943 VDD.n3459 VDD.n3458 23.1255
R19944 VDD.n3458 VDD.t135 23.1255
R19945 VDD.n3451 VDD.n3302 23.1255
R19946 VDD.t92 VDD.n3302 23.1255
R19947 VDD.n3454 VDD.n3303 23.1255
R19948 VDD.t92 VDD.n3303 23.1255
R19949 VDD.n3368 VDD.n3366 23.1255
R19950 VDD.n3366 VDD.t135 23.1255
R19951 VDD.n3466 VDD.n3367 23.1255
R19952 VDD.n3367 VDD.t135 23.1255
R19953 VDD.n3372 VDD.n3300 23.1255
R19954 VDD.t92 VDD.n3300 23.1255
R19955 VDD.n3369 VDD.n3301 23.1255
R19956 VDD.t92 VDD.n3301 23.1255
R19957 VDD.n3383 VDD.n3382 23.1255
R19958 VDD.n3382 VDD.t135 23.1255
R19959 VDD.n3386 VDD.n3385 23.1255
R19960 VDD.n3385 VDD.t135 23.1255
R19961 VDD.n3378 VDD.n3298 23.1255
R19962 VDD.t92 VDD.n3298 23.1255
R19963 VDD.n3381 VDD.n3299 23.1255
R19964 VDD.t92 VDD.n3299 23.1255
R19965 VDD.n3469 VDD.n3271 23.1255
R19966 VDD.t135 VDD.n3271 23.1255
R19967 VDD.n3470 VDD.n3272 23.1255
R19968 VDD.t135 VDD.n3272 23.1255
R19969 VDD.n3316 VDD.n3296 23.1255
R19970 VDD.t92 VDD.n3296 23.1255
R19971 VDD.n3317 VDD.n3297 23.1255
R19972 VDD.t92 VDD.n3297 23.1255
R19973 VDD.n3338 VDD.n3336 23.1255
R19974 VDD.n3336 VDD.t135 23.1255
R19975 VDD.n3339 VDD.n3337 23.1255
R19976 VDD.n3337 VDD.t135 23.1255
R19977 VDD.n3293 VDD.n3291 23.1255
R19978 VDD.t92 VDD.n3291 23.1255
R19979 VDD.n3491 VDD.n3295 23.1255
R19980 VDD.n3491 VDD.t92 23.1255
R19981 VDD.n3286 VDD.n3284 23.1255
R19982 VDD.n3284 VDD.t135 23.1255
R19983 VDD.n3287 VDD.n3285 23.1255
R19984 VDD.n3285 VDD.t135 23.1255
R19985 VDD.n3490 VDD.n3489 23.1255
R19986 VDD.t92 VDD.n3490 23.1255
R19987 VDD.n3487 VDD.n3321 23.1255
R19988 VDD.t92 VDD.n3321 23.1255
R19989 VDD.n3620 VDD.n3618 23.1255
R19990 VDD.n3618 VDD.t24 23.1255
R19991 VDD.n3619 VDD.n3584 23.1255
R19992 VDD.n3619 VDD.t24 23.1255
R19993 VDD.n3594 VDD.n3593 23.1255
R19994 VDD.n3594 VDD.t24 23.1255
R19995 VDD.n3737 VDD.n3736 23.1255
R19996 VDD.n3736 VDD.t24 23.1255
R19997 VDD.n3588 VDD.n3573 23.1255
R19998 VDD.t14 VDD.n3573 23.1255
R19999 VDD.n3591 VDD.n3574 23.1255
R20000 VDD.t14 VDD.n3574 23.1255
R20001 VDD.n3606 VDD.n3604 23.1255
R20002 VDD.n3604 VDD.t24 23.1255
R20003 VDD.n3615 VDD.n3605 23.1255
R20004 VDD.n3605 VDD.t24 23.1255
R20005 VDD.n3610 VDD.n3571 23.1255
R20006 VDD.t14 VDD.n3571 23.1255
R20007 VDD.n3607 VDD.n3572 23.1255
R20008 VDD.t14 VDD.n3572 23.1255
R20009 VDD.n3660 VDD.n3659 23.1255
R20010 VDD.n3659 VDD.t24 23.1255
R20011 VDD.n3663 VDD.n3662 23.1255
R20012 VDD.n3662 VDD.t24 23.1255
R20013 VDD.n3655 VDD.n3569 23.1255
R20014 VDD.t14 VDD.n3569 23.1255
R20015 VDD.n3658 VDD.n3570 23.1255
R20016 VDD.t14 VDD.n3570 23.1255
R20017 VDD.n3676 VDD.n3675 23.1255
R20018 VDD.n3675 VDD.t24 23.1255
R20019 VDD.n3679 VDD.n3678 23.1255
R20020 VDD.n3678 VDD.t24 23.1255
R20021 VDD.n3671 VDD.n3567 23.1255
R20022 VDD.t14 VDD.n3567 23.1255
R20023 VDD.n3674 VDD.n3568 23.1255
R20024 VDD.t14 VDD.n3568 23.1255
R20025 VDD.n3683 VDD.n3565 23.1255
R20026 VDD.t14 VDD.n3565 23.1255
R20027 VDD.n3687 VDD.n3566 23.1255
R20028 VDD.t14 VDD.n3566 23.1255
R20029 VDD.n3699 VDD.n3698 23.1255
R20030 VDD.n3698 VDD.t24 23.1255
R20031 VDD.n3702 VDD.n3701 23.1255
R20032 VDD.n3701 VDD.t24 23.1255
R20033 VDD.n3694 VDD.n3563 23.1255
R20034 VDD.t14 VDD.n3563 23.1255
R20035 VDD.n3697 VDD.n3564 23.1255
R20036 VDD.t14 VDD.n3564 23.1255
R20037 VDD.n3715 VDD.n3714 23.1255
R20038 VDD.n3714 VDD.t24 23.1255
R20039 VDD.n3718 VDD.n3717 23.1255
R20040 VDD.n3717 VDD.t24 23.1255
R20041 VDD.n3710 VDD.n3561 23.1255
R20042 VDD.t14 VDD.n3561 23.1255
R20043 VDD.n3713 VDD.n3562 23.1255
R20044 VDD.t14 VDD.n3562 23.1255
R20045 VDD.n3627 VDD.n3625 23.1255
R20046 VDD.n3625 VDD.t24 23.1255
R20047 VDD.n3725 VDD.n3626 23.1255
R20048 VDD.n3626 VDD.t24 23.1255
R20049 VDD.n3631 VDD.n3559 23.1255
R20050 VDD.t14 VDD.n3559 23.1255
R20051 VDD.n3628 VDD.n3560 23.1255
R20052 VDD.t14 VDD.n3560 23.1255
R20053 VDD.n3642 VDD.n3641 23.1255
R20054 VDD.n3641 VDD.t24 23.1255
R20055 VDD.n3645 VDD.n3644 23.1255
R20056 VDD.n3644 VDD.t24 23.1255
R20057 VDD.n3637 VDD.n3557 23.1255
R20058 VDD.t14 VDD.n3557 23.1255
R20059 VDD.n3640 VDD.n3558 23.1255
R20060 VDD.t14 VDD.n3558 23.1255
R20061 VDD.n3728 VDD.n3530 23.1255
R20062 VDD.t24 VDD.n3530 23.1255
R20063 VDD.n3729 VDD.n3531 23.1255
R20064 VDD.t24 VDD.n3531 23.1255
R20065 VDD.n3575 VDD.n3555 23.1255
R20066 VDD.t14 VDD.n3555 23.1255
R20067 VDD.n3576 VDD.n3556 23.1255
R20068 VDD.t14 VDD.n3556 23.1255
R20069 VDD.n3597 VDD.n3595 23.1255
R20070 VDD.n3595 VDD.t24 23.1255
R20071 VDD.n3598 VDD.n3596 23.1255
R20072 VDD.n3596 VDD.t24 23.1255
R20073 VDD.n3552 VDD.n3550 23.1255
R20074 VDD.t14 VDD.n3550 23.1255
R20075 VDD.n3750 VDD.n3554 23.1255
R20076 VDD.n3750 VDD.t14 23.1255
R20077 VDD.n3545 VDD.n3543 23.1255
R20078 VDD.n3543 VDD.t24 23.1255
R20079 VDD.n3546 VDD.n3544 23.1255
R20080 VDD.n3544 VDD.t24 23.1255
R20081 VDD.n3749 VDD.n3748 23.1255
R20082 VDD.t14 VDD.n3749 23.1255
R20083 VDD.n3746 VDD.n3580 23.1255
R20084 VDD.t14 VDD.n3580 23.1255
R20085 VDD.n3879 VDD.n3877 23.1255
R20086 VDD.n3877 VDD.t199 23.1255
R20087 VDD.n3878 VDD.n3843 23.1255
R20088 VDD.n3878 VDD.t199 23.1255
R20089 VDD.n3853 VDD.n3852 23.1255
R20090 VDD.n3853 VDD.t199 23.1255
R20091 VDD.n3996 VDD.n3995 23.1255
R20092 VDD.n3995 VDD.t199 23.1255
R20093 VDD.n3847 VDD.n3832 23.1255
R20094 VDD.t116 VDD.n3832 23.1255
R20095 VDD.n3850 VDD.n3833 23.1255
R20096 VDD.t116 VDD.n3833 23.1255
R20097 VDD.n3865 VDD.n3863 23.1255
R20098 VDD.n3863 VDD.t199 23.1255
R20099 VDD.n3874 VDD.n3864 23.1255
R20100 VDD.n3864 VDD.t199 23.1255
R20101 VDD.n3869 VDD.n3830 23.1255
R20102 VDD.t116 VDD.n3830 23.1255
R20103 VDD.n3866 VDD.n3831 23.1255
R20104 VDD.t116 VDD.n3831 23.1255
R20105 VDD.n3919 VDD.n3918 23.1255
R20106 VDD.n3918 VDD.t199 23.1255
R20107 VDD.n3922 VDD.n3921 23.1255
R20108 VDD.n3921 VDD.t199 23.1255
R20109 VDD.n3914 VDD.n3828 23.1255
R20110 VDD.t116 VDD.n3828 23.1255
R20111 VDD.n3917 VDD.n3829 23.1255
R20112 VDD.t116 VDD.n3829 23.1255
R20113 VDD.n3935 VDD.n3934 23.1255
R20114 VDD.n3934 VDD.t199 23.1255
R20115 VDD.n3938 VDD.n3937 23.1255
R20116 VDD.n3937 VDD.t199 23.1255
R20117 VDD.n3930 VDD.n3826 23.1255
R20118 VDD.t116 VDD.n3826 23.1255
R20119 VDD.n3933 VDD.n3827 23.1255
R20120 VDD.t116 VDD.n3827 23.1255
R20121 VDD.n3942 VDD.n3824 23.1255
R20122 VDD.t116 VDD.n3824 23.1255
R20123 VDD.n3946 VDD.n3825 23.1255
R20124 VDD.t116 VDD.n3825 23.1255
R20125 VDD.n3958 VDD.n3957 23.1255
R20126 VDD.n3957 VDD.t199 23.1255
R20127 VDD.n3961 VDD.n3960 23.1255
R20128 VDD.n3960 VDD.t199 23.1255
R20129 VDD.n3953 VDD.n3822 23.1255
R20130 VDD.t116 VDD.n3822 23.1255
R20131 VDD.n3956 VDD.n3823 23.1255
R20132 VDD.t116 VDD.n3823 23.1255
R20133 VDD.n3974 VDD.n3973 23.1255
R20134 VDD.n3973 VDD.t199 23.1255
R20135 VDD.n3977 VDD.n3976 23.1255
R20136 VDD.n3976 VDD.t199 23.1255
R20137 VDD.n3969 VDD.n3820 23.1255
R20138 VDD.t116 VDD.n3820 23.1255
R20139 VDD.n3972 VDD.n3821 23.1255
R20140 VDD.t116 VDD.n3821 23.1255
R20141 VDD.n3886 VDD.n3884 23.1255
R20142 VDD.n3884 VDD.t199 23.1255
R20143 VDD.n3984 VDD.n3885 23.1255
R20144 VDD.n3885 VDD.t199 23.1255
R20145 VDD.n3890 VDD.n3818 23.1255
R20146 VDD.t116 VDD.n3818 23.1255
R20147 VDD.n3887 VDD.n3819 23.1255
R20148 VDD.t116 VDD.n3819 23.1255
R20149 VDD.n3901 VDD.n3900 23.1255
R20150 VDD.n3900 VDD.t199 23.1255
R20151 VDD.n3904 VDD.n3903 23.1255
R20152 VDD.n3903 VDD.t199 23.1255
R20153 VDD.n3896 VDD.n3816 23.1255
R20154 VDD.t116 VDD.n3816 23.1255
R20155 VDD.n3899 VDD.n3817 23.1255
R20156 VDD.t116 VDD.n3817 23.1255
R20157 VDD.n3987 VDD.n3789 23.1255
R20158 VDD.t199 VDD.n3789 23.1255
R20159 VDD.n3988 VDD.n3790 23.1255
R20160 VDD.t199 VDD.n3790 23.1255
R20161 VDD.n3834 VDD.n3814 23.1255
R20162 VDD.t116 VDD.n3814 23.1255
R20163 VDD.n3835 VDD.n3815 23.1255
R20164 VDD.t116 VDD.n3815 23.1255
R20165 VDD.n3856 VDD.n3854 23.1255
R20166 VDD.n3854 VDD.t199 23.1255
R20167 VDD.n3857 VDD.n3855 23.1255
R20168 VDD.n3855 VDD.t199 23.1255
R20169 VDD.n3811 VDD.n3809 23.1255
R20170 VDD.t116 VDD.n3809 23.1255
R20171 VDD.n4009 VDD.n3813 23.1255
R20172 VDD.n4009 VDD.t116 23.1255
R20173 VDD.n3804 VDD.n3802 23.1255
R20174 VDD.n3802 VDD.t199 23.1255
R20175 VDD.n3805 VDD.n3803 23.1255
R20176 VDD.n3803 VDD.t199 23.1255
R20177 VDD.n4008 VDD.n4007 23.1255
R20178 VDD.t116 VDD.n4008 23.1255
R20179 VDD.n4005 VDD.n3839 23.1255
R20180 VDD.t116 VDD.n3839 23.1255
R20181 VDD.n4138 VDD.n4136 23.1255
R20182 VDD.n4136 VDD.t8 23.1255
R20183 VDD.n4137 VDD.n4102 23.1255
R20184 VDD.n4137 VDD.t8 23.1255
R20185 VDD.n4112 VDD.n4111 23.1255
R20186 VDD.n4112 VDD.t8 23.1255
R20187 VDD.n4255 VDD.n4254 23.1255
R20188 VDD.n4254 VDD.t8 23.1255
R20189 VDD.n4106 VDD.n4091 23.1255
R20190 VDD.t6 VDD.n4091 23.1255
R20191 VDD.n4109 VDD.n4092 23.1255
R20192 VDD.t6 VDD.n4092 23.1255
R20193 VDD.n4124 VDD.n4122 23.1255
R20194 VDD.n4122 VDD.t8 23.1255
R20195 VDD.n4133 VDD.n4123 23.1255
R20196 VDD.n4123 VDD.t8 23.1255
R20197 VDD.n4128 VDD.n4089 23.1255
R20198 VDD.t6 VDD.n4089 23.1255
R20199 VDD.n4125 VDD.n4090 23.1255
R20200 VDD.t6 VDD.n4090 23.1255
R20201 VDD.n4178 VDD.n4177 23.1255
R20202 VDD.n4177 VDD.t8 23.1255
R20203 VDD.n4181 VDD.n4180 23.1255
R20204 VDD.n4180 VDD.t8 23.1255
R20205 VDD.n4173 VDD.n4087 23.1255
R20206 VDD.t6 VDD.n4087 23.1255
R20207 VDD.n4176 VDD.n4088 23.1255
R20208 VDD.t6 VDD.n4088 23.1255
R20209 VDD.n4194 VDD.n4193 23.1255
R20210 VDD.n4193 VDD.t8 23.1255
R20211 VDD.n4197 VDD.n4196 23.1255
R20212 VDD.n4196 VDD.t8 23.1255
R20213 VDD.n4189 VDD.n4085 23.1255
R20214 VDD.t6 VDD.n4085 23.1255
R20215 VDD.n4192 VDD.n4086 23.1255
R20216 VDD.t6 VDD.n4086 23.1255
R20217 VDD.n4201 VDD.n4083 23.1255
R20218 VDD.t6 VDD.n4083 23.1255
R20219 VDD.n4205 VDD.n4084 23.1255
R20220 VDD.t6 VDD.n4084 23.1255
R20221 VDD.n4217 VDD.n4216 23.1255
R20222 VDD.n4216 VDD.t8 23.1255
R20223 VDD.n4220 VDD.n4219 23.1255
R20224 VDD.n4219 VDD.t8 23.1255
R20225 VDD.n4212 VDD.n4081 23.1255
R20226 VDD.t6 VDD.n4081 23.1255
R20227 VDD.n4215 VDD.n4082 23.1255
R20228 VDD.t6 VDD.n4082 23.1255
R20229 VDD.n4233 VDD.n4232 23.1255
R20230 VDD.n4232 VDD.t8 23.1255
R20231 VDD.n4236 VDD.n4235 23.1255
R20232 VDD.n4235 VDD.t8 23.1255
R20233 VDD.n4228 VDD.n4079 23.1255
R20234 VDD.t6 VDD.n4079 23.1255
R20235 VDD.n4231 VDD.n4080 23.1255
R20236 VDD.t6 VDD.n4080 23.1255
R20237 VDD.n4145 VDD.n4143 23.1255
R20238 VDD.n4143 VDD.t8 23.1255
R20239 VDD.n4243 VDD.n4144 23.1255
R20240 VDD.n4144 VDD.t8 23.1255
R20241 VDD.n4149 VDD.n4077 23.1255
R20242 VDD.t6 VDD.n4077 23.1255
R20243 VDD.n4146 VDD.n4078 23.1255
R20244 VDD.t6 VDD.n4078 23.1255
R20245 VDD.n4160 VDD.n4159 23.1255
R20246 VDD.n4159 VDD.t8 23.1255
R20247 VDD.n4163 VDD.n4162 23.1255
R20248 VDD.n4162 VDD.t8 23.1255
R20249 VDD.n4155 VDD.n4075 23.1255
R20250 VDD.t6 VDD.n4075 23.1255
R20251 VDD.n4158 VDD.n4076 23.1255
R20252 VDD.t6 VDD.n4076 23.1255
R20253 VDD.n4246 VDD.n4048 23.1255
R20254 VDD.t8 VDD.n4048 23.1255
R20255 VDD.n4247 VDD.n4049 23.1255
R20256 VDD.t8 VDD.n4049 23.1255
R20257 VDD.n4093 VDD.n4073 23.1255
R20258 VDD.t6 VDD.n4073 23.1255
R20259 VDD.n4094 VDD.n4074 23.1255
R20260 VDD.t6 VDD.n4074 23.1255
R20261 VDD.n4115 VDD.n4113 23.1255
R20262 VDD.n4113 VDD.t8 23.1255
R20263 VDD.n4116 VDD.n4114 23.1255
R20264 VDD.n4114 VDD.t8 23.1255
R20265 VDD.n4070 VDD.n4068 23.1255
R20266 VDD.t6 VDD.n4068 23.1255
R20267 VDD.n4268 VDD.n4072 23.1255
R20268 VDD.n4268 VDD.t6 23.1255
R20269 VDD.n4063 VDD.n4061 23.1255
R20270 VDD.n4061 VDD.t8 23.1255
R20271 VDD.n4064 VDD.n4062 23.1255
R20272 VDD.n4062 VDD.t8 23.1255
R20273 VDD.n4267 VDD.n4266 23.1255
R20274 VDD.t6 VDD.n4267 23.1255
R20275 VDD.n4264 VDD.n4098 23.1255
R20276 VDD.t6 VDD.n4098 23.1255
R20277 VDD.n4397 VDD.n4395 23.1255
R20278 VDD.n4395 VDD.t76 23.1255
R20279 VDD.n4396 VDD.n4361 23.1255
R20280 VDD.n4396 VDD.t76 23.1255
R20281 VDD.n4371 VDD.n4370 23.1255
R20282 VDD.n4371 VDD.t76 23.1255
R20283 VDD.n4514 VDD.n4513 23.1255
R20284 VDD.n4513 VDD.t76 23.1255
R20285 VDD.n4365 VDD.n4350 23.1255
R20286 VDD.t175 VDD.n4350 23.1255
R20287 VDD.n4368 VDD.n4351 23.1255
R20288 VDD.t175 VDD.n4351 23.1255
R20289 VDD.n4383 VDD.n4381 23.1255
R20290 VDD.n4381 VDD.t76 23.1255
R20291 VDD.n4392 VDD.n4382 23.1255
R20292 VDD.n4382 VDD.t76 23.1255
R20293 VDD.n4387 VDD.n4348 23.1255
R20294 VDD.t175 VDD.n4348 23.1255
R20295 VDD.n4384 VDD.n4349 23.1255
R20296 VDD.t175 VDD.n4349 23.1255
R20297 VDD.n4437 VDD.n4436 23.1255
R20298 VDD.n4436 VDD.t76 23.1255
R20299 VDD.n4440 VDD.n4439 23.1255
R20300 VDD.n4439 VDD.t76 23.1255
R20301 VDD.n4432 VDD.n4346 23.1255
R20302 VDD.t175 VDD.n4346 23.1255
R20303 VDD.n4435 VDD.n4347 23.1255
R20304 VDD.t175 VDD.n4347 23.1255
R20305 VDD.n4453 VDD.n4452 23.1255
R20306 VDD.n4452 VDD.t76 23.1255
R20307 VDD.n4456 VDD.n4455 23.1255
R20308 VDD.n4455 VDD.t76 23.1255
R20309 VDD.n4448 VDD.n4344 23.1255
R20310 VDD.t175 VDD.n4344 23.1255
R20311 VDD.n4451 VDD.n4345 23.1255
R20312 VDD.t175 VDD.n4345 23.1255
R20313 VDD.n4460 VDD.n4342 23.1255
R20314 VDD.t175 VDD.n4342 23.1255
R20315 VDD.n4464 VDD.n4343 23.1255
R20316 VDD.t175 VDD.n4343 23.1255
R20317 VDD.n4476 VDD.n4475 23.1255
R20318 VDD.n4475 VDD.t76 23.1255
R20319 VDD.n4479 VDD.n4478 23.1255
R20320 VDD.n4478 VDD.t76 23.1255
R20321 VDD.n4471 VDD.n4340 23.1255
R20322 VDD.t175 VDD.n4340 23.1255
R20323 VDD.n4474 VDD.n4341 23.1255
R20324 VDD.t175 VDD.n4341 23.1255
R20325 VDD.n4492 VDD.n4491 23.1255
R20326 VDD.n4491 VDD.t76 23.1255
R20327 VDD.n4495 VDD.n4494 23.1255
R20328 VDD.n4494 VDD.t76 23.1255
R20329 VDD.n4487 VDD.n4338 23.1255
R20330 VDD.t175 VDD.n4338 23.1255
R20331 VDD.n4490 VDD.n4339 23.1255
R20332 VDD.t175 VDD.n4339 23.1255
R20333 VDD.n4404 VDD.n4402 23.1255
R20334 VDD.n4402 VDD.t76 23.1255
R20335 VDD.n4502 VDD.n4403 23.1255
R20336 VDD.n4403 VDD.t76 23.1255
R20337 VDD.n4408 VDD.n4336 23.1255
R20338 VDD.t175 VDD.n4336 23.1255
R20339 VDD.n4405 VDD.n4337 23.1255
R20340 VDD.t175 VDD.n4337 23.1255
R20341 VDD.n4419 VDD.n4418 23.1255
R20342 VDD.n4418 VDD.t76 23.1255
R20343 VDD.n4422 VDD.n4421 23.1255
R20344 VDD.n4421 VDD.t76 23.1255
R20345 VDD.n4414 VDD.n4334 23.1255
R20346 VDD.t175 VDD.n4334 23.1255
R20347 VDD.n4417 VDD.n4335 23.1255
R20348 VDD.t175 VDD.n4335 23.1255
R20349 VDD.n4505 VDD.n4307 23.1255
R20350 VDD.t76 VDD.n4307 23.1255
R20351 VDD.n4506 VDD.n4308 23.1255
R20352 VDD.t76 VDD.n4308 23.1255
R20353 VDD.n4352 VDD.n4332 23.1255
R20354 VDD.t175 VDD.n4332 23.1255
R20355 VDD.n4353 VDD.n4333 23.1255
R20356 VDD.t175 VDD.n4333 23.1255
R20357 VDD.n4374 VDD.n4372 23.1255
R20358 VDD.n4372 VDD.t76 23.1255
R20359 VDD.n4375 VDD.n4373 23.1255
R20360 VDD.n4373 VDD.t76 23.1255
R20361 VDD.n4329 VDD.n4327 23.1255
R20362 VDD.t175 VDD.n4327 23.1255
R20363 VDD.n4527 VDD.n4331 23.1255
R20364 VDD.n4527 VDD.t175 23.1255
R20365 VDD.n4323 VDD.n4321 23.1255
R20366 VDD.n4321 VDD.t76 23.1255
R20367 VDD.n4322 VDD.n4320 23.1255
R20368 VDD.n4320 VDD.t76 23.1255
R20369 VDD.n4526 VDD.n4525 23.1255
R20370 VDD.t175 VDD.n4526 23.1255
R20371 VDD.n4523 VDD.n4357 23.1255
R20372 VDD.t175 VDD.n4357 23.1255
R20373 VDD.n5022 VDD.n5021 23.1255
R20374 VDD.n5021 VDD.n5020 23.1255
R20375 VDD.n5025 VDD.n5024 23.1255
R20376 VDD.n5026 VDD.n5025 23.1255
R20377 VDD.n4559 VDD.n4557 23.1255
R20378 VDD.n5027 VDD.n4559 23.1255
R20379 VDD.n4560 VDD.n4558 23.1255
R20380 VDD.n5018 VDD.n5017 23.1255
R20381 VDD.n5019 VDD.n5018 23.1255
R20382 VDD.n5015 VDD.n5014 23.1255
R20383 VDD.n4570 VDD.n4568 23.1255
R20384 VDD.n5002 VDD.n4570 23.1255
R20385 VDD.n4571 VDD.n4569 23.1255
R20386 VDD.n5000 VDD.n4999 23.1255
R20387 VDD.n5001 VDD.n5000 23.1255
R20388 VDD.n4997 VDD.n4996 23.1255
R20389 VDD.n4981 VDD.n4980 23.1255
R20390 VDD.n4980 VDD.n4979 23.1255
R20391 VDD.n4984 VDD.n4983 23.1255
R20392 VDD.n4985 VDD.n4984 23.1255
R20393 VDD.n4578 VDD.n4576 23.1255
R20394 VDD.n4986 VDD.n4578 23.1255
R20395 VDD.n4579 VDD.n4577 23.1255
R20396 VDD.n4977 VDD.n4976 23.1255
R20397 VDD.n4978 VDD.n4977 23.1255
R20398 VDD.n4974 VDD.n4973 23.1255
R20399 VDD.n4589 VDD.n4587 23.1255
R20400 VDD.n4961 VDD.n4589 23.1255
R20401 VDD.n4590 VDD.n4588 23.1255
R20402 VDD.n4959 VDD.n4958 23.1255
R20403 VDD.n4960 VDD.n4959 23.1255
R20404 VDD.n4956 VDD.n4955 23.1255
R20405 VDD.n4940 VDD.n4939 23.1255
R20406 VDD.n4939 VDD.n4938 23.1255
R20407 VDD.n4943 VDD.n4942 23.1255
R20408 VDD.n4944 VDD.n4943 23.1255
R20409 VDD.n4597 VDD.n4595 23.1255
R20410 VDD.n4945 VDD.n4597 23.1255
R20411 VDD.n4598 VDD.n4596 23.1255
R20412 VDD.n4936 VDD.n4935 23.1255
R20413 VDD.n4937 VDD.n4936 23.1255
R20414 VDD.n4933 VDD.n4932 23.1255
R20415 VDD.n4608 VDD.n4606 23.1255
R20416 VDD.n4920 VDD.n4608 23.1255
R20417 VDD.n4609 VDD.n4607 23.1255
R20418 VDD.n4918 VDD.n4917 23.1255
R20419 VDD.n4919 VDD.n4918 23.1255
R20420 VDD.n4915 VDD.n4914 23.1255
R20421 VDD.n4899 VDD.n4898 23.1255
R20422 VDD.n4898 VDD.n4897 23.1255
R20423 VDD.n4902 VDD.n4901 23.1255
R20424 VDD.n4903 VDD.n4902 23.1255
R20425 VDD.n4616 VDD.n4614 23.1255
R20426 VDD.n4904 VDD.n4616 23.1255
R20427 VDD.n4617 VDD.n4615 23.1255
R20428 VDD.n4895 VDD.n4894 23.1255
R20429 VDD.n4896 VDD.n4895 23.1255
R20430 VDD.n4892 VDD.n4891 23.1255
R20431 VDD.n4627 VDD.n4625 23.1255
R20432 VDD.n4879 VDD.n4627 23.1255
R20433 VDD.n4628 VDD.n4626 23.1255
R20434 VDD.n4877 VDD.n4876 23.1255
R20435 VDD.n4878 VDD.n4877 23.1255
R20436 VDD.n4874 VDD.n4873 23.1255
R20437 VDD.n4858 VDD.n4857 23.1255
R20438 VDD.n4857 VDD.n4856 23.1255
R20439 VDD.n4861 VDD.n4860 23.1255
R20440 VDD.n4862 VDD.n4861 23.1255
R20441 VDD.n4635 VDD.n4633 23.1255
R20442 VDD.n4863 VDD.n4635 23.1255
R20443 VDD.n4636 VDD.n4634 23.1255
R20444 VDD.n4854 VDD.n4853 23.1255
R20445 VDD.n4855 VDD.n4854 23.1255
R20446 VDD.n4851 VDD.n4850 23.1255
R20447 VDD.n4646 VDD.n4644 23.1255
R20448 VDD.n4838 VDD.n4646 23.1255
R20449 VDD.n4647 VDD.n4645 23.1255
R20450 VDD.n4836 VDD.n4835 23.1255
R20451 VDD.n4837 VDD.n4836 23.1255
R20452 VDD.n4833 VDD.n4832 23.1255
R20453 VDD.n4817 VDD.n4816 23.1255
R20454 VDD.n4816 VDD.n4815 23.1255
R20455 VDD.n4820 VDD.n4819 23.1255
R20456 VDD.n4821 VDD.n4820 23.1255
R20457 VDD.n4654 VDD.n4652 23.1255
R20458 VDD.n4822 VDD.n4654 23.1255
R20459 VDD.n4655 VDD.n4653 23.1255
R20460 VDD.n4813 VDD.n4812 23.1255
R20461 VDD.n4814 VDD.n4813 23.1255
R20462 VDD.n4810 VDD.n4809 23.1255
R20463 VDD.n4665 VDD.n4663 23.1255
R20464 VDD.n4797 VDD.n4665 23.1255
R20465 VDD.n4666 VDD.n4664 23.1255
R20466 VDD.n4795 VDD.n4794 23.1255
R20467 VDD.n4796 VDD.n4795 23.1255
R20468 VDD.n4792 VDD.n4791 23.1255
R20469 VDD.n4776 VDD.n4775 23.1255
R20470 VDD.n4775 VDD.n4774 23.1255
R20471 VDD.n4779 VDD.n4778 23.1255
R20472 VDD.n4780 VDD.n4779 23.1255
R20473 VDD.n4673 VDD.n4671 23.1255
R20474 VDD.n4781 VDD.n4673 23.1255
R20475 VDD.n4674 VDD.n4672 23.1255
R20476 VDD.n4772 VDD.n4771 23.1255
R20477 VDD.n4773 VDD.n4772 23.1255
R20478 VDD.n4769 VDD.n4768 23.1255
R20479 VDD.n4684 VDD.n4682 23.1255
R20480 VDD.n4756 VDD.n4684 23.1255
R20481 VDD.n4685 VDD.n4683 23.1255
R20482 VDD.n4754 VDD.n4753 23.1255
R20483 VDD.n4755 VDD.n4754 23.1255
R20484 VDD.n4751 VDD.n4750 23.1255
R20485 VDD.n4735 VDD.n4734 23.1255
R20486 VDD.n4734 VDD.n4733 23.1255
R20487 VDD.n4738 VDD.n4737 23.1255
R20488 VDD.n4739 VDD.n4738 23.1255
R20489 VDD.n4692 VDD.n4690 23.1255
R20490 VDD.n4740 VDD.n4692 23.1255
R20491 VDD.n4693 VDD.n4691 23.1255
R20492 VDD.n4731 VDD.n4730 23.1255
R20493 VDD.n4732 VDD.n4731 23.1255
R20494 VDD.n4728 VDD.n4727 23.1255
R20495 VDD.n4703 VDD.n4701 23.1255
R20496 VDD.n4715 VDD.n4703 23.1255
R20497 VDD.n4704 VDD.n4702 23.1255
R20498 VDD.n4713 VDD.n4712 23.1255
R20499 VDD.n4714 VDD.n4713 23.1255
R20500 VDD.n4710 VDD.n4709 23.1255
R20501 VDD.n6064 VDD.n6060 23.1255
R20502 VDD.n6064 VDD.n6063 23.1255
R20503 VDD.n6056 VDD.n6052 23.1255
R20504 VDD.n6073 VDD.n6052 23.1255
R20505 VDD.n6077 VDD.n6051 23.1255
R20506 VDD.n6077 VDD.n6076 23.1255
R20507 VDD.n6046 VDD.n6042 23.1255
R20508 VDD.n6083 VDD.n6042 23.1255
R20509 VDD.n6087 VDD.n6041 23.1255
R20510 VDD.n6087 VDD.n6086 23.1255
R20511 VDD.n6035 VDD.n6031 23.1255
R20512 VDD.n6093 VDD.n6031 23.1255
R20513 VDD.n6097 VDD.n6030 23.1255
R20514 VDD.n6097 VDD.n6096 23.1255
R20515 VDD.n6022 VDD.n6018 23.1255
R20516 VDD.n6103 VDD.n6018 23.1255
R20517 VDD.n6107 VDD.n6017 23.1255
R20518 VDD.n6107 VDD.n6106 23.1255
R20519 VDD.n6010 VDD.n6006 23.1255
R20520 VDD.n6113 VDD.n6006 23.1255
R20521 VDD.n6116 VDD.n6115 23.1255
R20522 VDD.n6115 VDD.n6114 23.1255
R20523 VDD.n6119 VDD.n6118 23.1255
R20524 VDD.n6120 VDD.n6119 23.1255
R20525 VDD.n6124 VDD.n6002 23.1255
R20526 VDD.n6124 VDD.n6123 23.1255
R20527 VDD.n5994 VDD.n5990 23.1255
R20528 VDD.n6130 VDD.n5990 23.1255
R20529 VDD.n6134 VDD.n5989 23.1255
R20530 VDD.n6134 VDD.n6133 23.1255
R20531 VDD.n5984 VDD.n5980 23.1255
R20532 VDD.n6140 VDD.n5980 23.1255
R20533 VDD.n6144 VDD.n5979 23.1255
R20534 VDD.n6144 VDD.n6143 23.1255
R20535 VDD.n5973 VDD.n5969 23.1255
R20536 VDD.n6150 VDD.n5969 23.1255
R20537 VDD.n6154 VDD.n5968 23.1255
R20538 VDD.n6154 VDD.n6153 23.1255
R20539 VDD.n5960 VDD.n5956 23.1255
R20540 VDD.n6160 VDD.n5956 23.1255
R20541 VDD.n6164 VDD.n5955 23.1255
R20542 VDD.n6164 VDD.n6163 23.1255
R20543 VDD.n5951 VDD.n5947 23.1255
R20544 VDD.n6170 VDD.n5947 23.1255
R20545 VDD.n6172 VDD.n5945 23.1255
R20546 VDD.n6171 VDD.n5945 23.1255
R20547 VDD.n6173 VDD.n5946 23.1255
R20548 VDD.n6178 VDD.n5946 23.1255
R20549 VDD.n6198 VDD.n5936 23.1255
R20550 VDD.n6198 VDD.n6197 23.1255
R20551 VDD.n5928 VDD.n5924 23.1255
R20552 VDD.n6204 VDD.n5924 23.1255
R20553 VDD.n6208 VDD.n5923 23.1255
R20554 VDD.n6208 VDD.n6207 23.1255
R20555 VDD.n5918 VDD.n5914 23.1255
R20556 VDD.n6214 VDD.n5914 23.1255
R20557 VDD.n6218 VDD.n5913 23.1255
R20558 VDD.n6218 VDD.n6217 23.1255
R20559 VDD.n5907 VDD.n5903 23.1255
R20560 VDD.n6224 VDD.n5903 23.1255
R20561 VDD.n6228 VDD.n5902 23.1255
R20562 VDD.n6228 VDD.n6227 23.1255
R20563 VDD.n5894 VDD.n5890 23.1255
R20564 VDD.n6234 VDD.n5890 23.1255
R20565 VDD.n6238 VDD.n5889 23.1255
R20566 VDD.n6238 VDD.n6237 23.1255
R20567 VDD.n5882 VDD.n5878 23.1255
R20568 VDD.n6244 VDD.n5878 23.1255
R20569 VDD.n6247 VDD.n6246 23.1255
R20570 VDD.n6246 VDD.n6245 23.1255
R20571 VDD.n6250 VDD.n6249 23.1255
R20572 VDD.n6251 VDD.n6250 23.1255
R20573 VDD.n6255 VDD.n5874 23.1255
R20574 VDD.n6255 VDD.n6254 23.1255
R20575 VDD.n5866 VDD.n5862 23.1255
R20576 VDD.n6261 VDD.n5862 23.1255
R20577 VDD.n6265 VDD.n5861 23.1255
R20578 VDD.n6265 VDD.n6264 23.1255
R20579 VDD.n5856 VDD.n5852 23.1255
R20580 VDD.n6271 VDD.n5852 23.1255
R20581 VDD.n6275 VDD.n5851 23.1255
R20582 VDD.n6275 VDD.n6274 23.1255
R20583 VDD.n5845 VDD.n5841 23.1255
R20584 VDD.n6281 VDD.n5841 23.1255
R20585 VDD.n6285 VDD.n5840 23.1255
R20586 VDD.n6285 VDD.n6284 23.1255
R20587 VDD.n5832 VDD.n5828 23.1255
R20588 VDD.n6291 VDD.n5828 23.1255
R20589 VDD.n6295 VDD.n5827 23.1255
R20590 VDD.n6295 VDD.n6294 23.1255
R20591 VDD.n5823 VDD.n5819 23.1255
R20592 VDD.n6301 VDD.n5819 23.1255
R20593 VDD.n6303 VDD.n5817 23.1255
R20594 VDD.n6302 VDD.n5817 23.1255
R20595 VDD.n6304 VDD.n5818 23.1255
R20596 VDD.n6309 VDD.n5818 23.1255
R20597 VDD.n6329 VDD.n5808 23.1255
R20598 VDD.n6329 VDD.n6328 23.1255
R20599 VDD.n5800 VDD.n5796 23.1255
R20600 VDD.n6335 VDD.n5796 23.1255
R20601 VDD.n6339 VDD.n5795 23.1255
R20602 VDD.n6339 VDD.n6338 23.1255
R20603 VDD.n5790 VDD.n5786 23.1255
R20604 VDD.n6345 VDD.n5786 23.1255
R20605 VDD.n6349 VDD.n5785 23.1255
R20606 VDD.n6349 VDD.n6348 23.1255
R20607 VDD.n5779 VDD.n5775 23.1255
R20608 VDD.n6355 VDD.n5775 23.1255
R20609 VDD.n6359 VDD.n5774 23.1255
R20610 VDD.n6359 VDD.n6358 23.1255
R20611 VDD.n5766 VDD.n5762 23.1255
R20612 VDD.n6365 VDD.n5762 23.1255
R20613 VDD.n6369 VDD.n5761 23.1255
R20614 VDD.n6369 VDD.n6368 23.1255
R20615 VDD.n5754 VDD.n5750 23.1255
R20616 VDD.n6375 VDD.n5750 23.1255
R20617 VDD.n6378 VDD.n6377 23.1255
R20618 VDD.n6377 VDD.n6376 23.1255
R20619 VDD.n6381 VDD.n6380 23.1255
R20620 VDD.n6382 VDD.n6381 23.1255
R20621 VDD.n6386 VDD.n5746 23.1255
R20622 VDD.n6386 VDD.n6385 23.1255
R20623 VDD.n5738 VDD.n5734 23.1255
R20624 VDD.n6392 VDD.n5734 23.1255
R20625 VDD.n6396 VDD.n5733 23.1255
R20626 VDD.n6396 VDD.n6395 23.1255
R20627 VDD.n5728 VDD.n5724 23.1255
R20628 VDD.n6402 VDD.n5724 23.1255
R20629 VDD.n6406 VDD.n5723 23.1255
R20630 VDD.n6406 VDD.n6405 23.1255
R20631 VDD.n5717 VDD.n5713 23.1255
R20632 VDD.n6412 VDD.n5713 23.1255
R20633 VDD.n6416 VDD.n5712 23.1255
R20634 VDD.n6416 VDD.n6415 23.1255
R20635 VDD.n5704 VDD.n5700 23.1255
R20636 VDD.n6422 VDD.n5700 23.1255
R20637 VDD.n6426 VDD.n5699 23.1255
R20638 VDD.n6426 VDD.n6425 23.1255
R20639 VDD.n5695 VDD.n5691 23.1255
R20640 VDD.n6432 VDD.n5691 23.1255
R20641 VDD.n6434 VDD.n5689 23.1255
R20642 VDD.n6433 VDD.n5689 23.1255
R20643 VDD.n6435 VDD.n5690 23.1255
R20644 VDD.n6440 VDD.n5690 23.1255
R20645 VDD.n6460 VDD.n5680 23.1255
R20646 VDD.n6460 VDD.n6459 23.1255
R20647 VDD.n5672 VDD.n5668 23.1255
R20648 VDD.n6466 VDD.n5668 23.1255
R20649 VDD.n6470 VDD.n5667 23.1255
R20650 VDD.n6470 VDD.n6469 23.1255
R20651 VDD.n5662 VDD.n5658 23.1255
R20652 VDD.n6476 VDD.n5658 23.1255
R20653 VDD.n6480 VDD.n5657 23.1255
R20654 VDD.n6480 VDD.n6479 23.1255
R20655 VDD.n5651 VDD.n5647 23.1255
R20656 VDD.n6486 VDD.n5647 23.1255
R20657 VDD.n6490 VDD.n5646 23.1255
R20658 VDD.n6490 VDD.n6489 23.1255
R20659 VDD.n5638 VDD.n5634 23.1255
R20660 VDD.n6496 VDD.n5634 23.1255
R20661 VDD.n6500 VDD.n5633 23.1255
R20662 VDD.n6500 VDD.n6499 23.1255
R20663 VDD.n5626 VDD.n5622 23.1255
R20664 VDD.n6506 VDD.n5622 23.1255
R20665 VDD.n6509 VDD.n6508 23.1255
R20666 VDD.n6508 VDD.n6507 23.1255
R20667 VDD.n6512 VDD.n6511 23.1255
R20668 VDD.n6513 VDD.n6512 23.1255
R20669 VDD.n6517 VDD.n5618 23.1255
R20670 VDD.n6517 VDD.n6516 23.1255
R20671 VDD.n5610 VDD.n5606 23.1255
R20672 VDD.n6523 VDD.n5606 23.1255
R20673 VDD.n6527 VDD.n5605 23.1255
R20674 VDD.n6527 VDD.n6526 23.1255
R20675 VDD.n5600 VDD.n5596 23.1255
R20676 VDD.n6533 VDD.n5596 23.1255
R20677 VDD.n6537 VDD.n5595 23.1255
R20678 VDD.n6537 VDD.n6536 23.1255
R20679 VDD.n5589 VDD.n5585 23.1255
R20680 VDD.n6543 VDD.n5585 23.1255
R20681 VDD.n6547 VDD.n5584 23.1255
R20682 VDD.n6547 VDD.n6546 23.1255
R20683 VDD.n5576 VDD.n5572 23.1255
R20684 VDD.n6553 VDD.n5572 23.1255
R20685 VDD.n6557 VDD.n5571 23.1255
R20686 VDD.n6557 VDD.n6556 23.1255
R20687 VDD.n5567 VDD.n5563 23.1255
R20688 VDD.n6563 VDD.n5563 23.1255
R20689 VDD.n6565 VDD.n5561 23.1255
R20690 VDD.n6564 VDD.n5561 23.1255
R20691 VDD.n6566 VDD.n5562 23.1255
R20692 VDD.n6571 VDD.n5562 23.1255
R20693 VDD.n6591 VDD.n5552 23.1255
R20694 VDD.n6591 VDD.n6590 23.1255
R20695 VDD.n5544 VDD.n5540 23.1255
R20696 VDD.n6597 VDD.n5540 23.1255
R20697 VDD.n6601 VDD.n5539 23.1255
R20698 VDD.n6601 VDD.n6600 23.1255
R20699 VDD.n5534 VDD.n5530 23.1255
R20700 VDD.n6607 VDD.n5530 23.1255
R20701 VDD.n6611 VDD.n5529 23.1255
R20702 VDD.n6611 VDD.n6610 23.1255
R20703 VDD.n5523 VDD.n5519 23.1255
R20704 VDD.n6617 VDD.n5519 23.1255
R20705 VDD.n6621 VDD.n5518 23.1255
R20706 VDD.n6621 VDD.n6620 23.1255
R20707 VDD.n5510 VDD.n5506 23.1255
R20708 VDD.n6627 VDD.n5506 23.1255
R20709 VDD.n6631 VDD.n5505 23.1255
R20710 VDD.n6631 VDD.n6630 23.1255
R20711 VDD.n5498 VDD.n5494 23.1255
R20712 VDD.n6637 VDD.n5494 23.1255
R20713 VDD.n6640 VDD.n6639 23.1255
R20714 VDD.n6639 VDD.n6638 23.1255
R20715 VDD.n6643 VDD.n6642 23.1255
R20716 VDD.n6644 VDD.n6643 23.1255
R20717 VDD.n6648 VDD.n5490 23.1255
R20718 VDD.n6648 VDD.n6647 23.1255
R20719 VDD.n5482 VDD.n5478 23.1255
R20720 VDD.n6654 VDD.n5478 23.1255
R20721 VDD.n6658 VDD.n5477 23.1255
R20722 VDD.n6658 VDD.n6657 23.1255
R20723 VDD.n5472 VDD.n5468 23.1255
R20724 VDD.n6664 VDD.n5468 23.1255
R20725 VDD.n6668 VDD.n5467 23.1255
R20726 VDD.n6668 VDD.n6667 23.1255
R20727 VDD.n5461 VDD.n5457 23.1255
R20728 VDD.n6674 VDD.n5457 23.1255
R20729 VDD.n6678 VDD.n5456 23.1255
R20730 VDD.n6678 VDD.n6677 23.1255
R20731 VDD.n5448 VDD.n5444 23.1255
R20732 VDD.n6684 VDD.n5444 23.1255
R20733 VDD.n6688 VDD.n5443 23.1255
R20734 VDD.n6688 VDD.n6687 23.1255
R20735 VDD.n5439 VDD.n5435 23.1255
R20736 VDD.n6694 VDD.n5435 23.1255
R20737 VDD.n6696 VDD.n5433 23.1255
R20738 VDD.n6695 VDD.n5433 23.1255
R20739 VDD.n6697 VDD.n5434 23.1255
R20740 VDD.n6702 VDD.n5434 23.1255
R20741 VDD.n6722 VDD.n5424 23.1255
R20742 VDD.n6722 VDD.n6721 23.1255
R20743 VDD.n5416 VDD.n5412 23.1255
R20744 VDD.n6728 VDD.n5412 23.1255
R20745 VDD.n6732 VDD.n5411 23.1255
R20746 VDD.n6732 VDD.n6731 23.1255
R20747 VDD.n5406 VDD.n5402 23.1255
R20748 VDD.n6738 VDD.n5402 23.1255
R20749 VDD.n6742 VDD.n5401 23.1255
R20750 VDD.n6742 VDD.n6741 23.1255
R20751 VDD.n5395 VDD.n5391 23.1255
R20752 VDD.n6748 VDD.n5391 23.1255
R20753 VDD.n6752 VDD.n5390 23.1255
R20754 VDD.n6752 VDD.n6751 23.1255
R20755 VDD.n5382 VDD.n5378 23.1255
R20756 VDD.n6758 VDD.n5378 23.1255
R20757 VDD.n6762 VDD.n5377 23.1255
R20758 VDD.n6762 VDD.n6761 23.1255
R20759 VDD.n5370 VDD.n5366 23.1255
R20760 VDD.n6768 VDD.n5366 23.1255
R20761 VDD.n6771 VDD.n6770 23.1255
R20762 VDD.n6770 VDD.n6769 23.1255
R20763 VDD.n6774 VDD.n6773 23.1255
R20764 VDD.n6775 VDD.n6774 23.1255
R20765 VDD.n6779 VDD.n5362 23.1255
R20766 VDD.n6779 VDD.n6778 23.1255
R20767 VDD.n5354 VDD.n5350 23.1255
R20768 VDD.n6785 VDD.n5350 23.1255
R20769 VDD.n6789 VDD.n5349 23.1255
R20770 VDD.n6789 VDD.n6788 23.1255
R20771 VDD.n5344 VDD.n5340 23.1255
R20772 VDD.n6795 VDD.n5340 23.1255
R20773 VDD.n6799 VDD.n5339 23.1255
R20774 VDD.n6799 VDD.n6798 23.1255
R20775 VDD.n5333 VDD.n5329 23.1255
R20776 VDD.n6805 VDD.n5329 23.1255
R20777 VDD.n6809 VDD.n5328 23.1255
R20778 VDD.n6809 VDD.n6808 23.1255
R20779 VDD.n5320 VDD.n5316 23.1255
R20780 VDD.n6815 VDD.n5316 23.1255
R20781 VDD.n6819 VDD.n5315 23.1255
R20782 VDD.n6819 VDD.n6818 23.1255
R20783 VDD.n5311 VDD.n5307 23.1255
R20784 VDD.n6825 VDD.n5307 23.1255
R20785 VDD.n6827 VDD.n5305 23.1255
R20786 VDD.n6826 VDD.n5305 23.1255
R20787 VDD.n6828 VDD.n5306 23.1255
R20788 VDD.n6833 VDD.n5306 23.1255
R20789 VDD.n6853 VDD.n5296 23.1255
R20790 VDD.n6853 VDD.n6852 23.1255
R20791 VDD.n5288 VDD.n5284 23.1255
R20792 VDD.n6859 VDD.n5284 23.1255
R20793 VDD.n6863 VDD.n5283 23.1255
R20794 VDD.n6863 VDD.n6862 23.1255
R20795 VDD.n5278 VDD.n5274 23.1255
R20796 VDD.n6869 VDD.n5274 23.1255
R20797 VDD.n6873 VDD.n5273 23.1255
R20798 VDD.n6873 VDD.n6872 23.1255
R20799 VDD.n5267 VDD.n5263 23.1255
R20800 VDD.n6879 VDD.n5263 23.1255
R20801 VDD.n6883 VDD.n5262 23.1255
R20802 VDD.n6883 VDD.n6882 23.1255
R20803 VDD.n5254 VDD.n5250 23.1255
R20804 VDD.n6889 VDD.n5250 23.1255
R20805 VDD.n6893 VDD.n5249 23.1255
R20806 VDD.n6893 VDD.n6892 23.1255
R20807 VDD.n5242 VDD.n5238 23.1255
R20808 VDD.n6899 VDD.n5238 23.1255
R20809 VDD.n6902 VDD.n6901 23.1255
R20810 VDD.n6901 VDD.n6900 23.1255
R20811 VDD.n6905 VDD.n6904 23.1255
R20812 VDD.n6906 VDD.n6905 23.1255
R20813 VDD.n6910 VDD.n5234 23.1255
R20814 VDD.n6910 VDD.n6909 23.1255
R20815 VDD.n5226 VDD.n5222 23.1255
R20816 VDD.n6916 VDD.n5222 23.1255
R20817 VDD.n6920 VDD.n5221 23.1255
R20818 VDD.n6920 VDD.n6919 23.1255
R20819 VDD.n5216 VDD.n5212 23.1255
R20820 VDD.n6926 VDD.n5212 23.1255
R20821 VDD.n6930 VDD.n5211 23.1255
R20822 VDD.n6930 VDD.n6929 23.1255
R20823 VDD.n5205 VDD.n5201 23.1255
R20824 VDD.n6936 VDD.n5201 23.1255
R20825 VDD.n6940 VDD.n5200 23.1255
R20826 VDD.n6940 VDD.n6939 23.1255
R20827 VDD.n5192 VDD.n5188 23.1255
R20828 VDD.n6946 VDD.n5188 23.1255
R20829 VDD.n6950 VDD.n5187 23.1255
R20830 VDD.n6950 VDD.n6949 23.1255
R20831 VDD.n5183 VDD.n5179 23.1255
R20832 VDD.n6956 VDD.n5179 23.1255
R20833 VDD.n6958 VDD.n5177 23.1255
R20834 VDD.n6957 VDD.n5177 23.1255
R20835 VDD.n6959 VDD.n5178 23.1255
R20836 VDD.n6964 VDD.n5178 23.1255
R20837 VDD.n6984 VDD.n5168 23.1255
R20838 VDD.n6984 VDD.n6983 23.1255
R20839 VDD.n5160 VDD.n5156 23.1255
R20840 VDD.n6990 VDD.n5156 23.1255
R20841 VDD.n6994 VDD.n5155 23.1255
R20842 VDD.n6994 VDD.n6993 23.1255
R20843 VDD.n5150 VDD.n5146 23.1255
R20844 VDD.n7000 VDD.n5146 23.1255
R20845 VDD.n7004 VDD.n5145 23.1255
R20846 VDD.n7004 VDD.n7003 23.1255
R20847 VDD.n5139 VDD.n5135 23.1255
R20848 VDD.n7010 VDD.n5135 23.1255
R20849 VDD.n7014 VDD.n5134 23.1255
R20850 VDD.n7014 VDD.n7013 23.1255
R20851 VDD.n5126 VDD.n5122 23.1255
R20852 VDD.n7020 VDD.n5122 23.1255
R20853 VDD.n7024 VDD.n5121 23.1255
R20854 VDD.n7024 VDD.n7023 23.1255
R20855 VDD.n5114 VDD.n5110 23.1255
R20856 VDD.n7030 VDD.n5110 23.1255
R20857 VDD.n7033 VDD.n7032 23.1255
R20858 VDD.n7032 VDD.n7031 23.1255
R20859 VDD.n7036 VDD.n7035 23.1255
R20860 VDD.n7037 VDD.n7036 23.1255
R20861 VDD.n7041 VDD.n5106 23.1255
R20862 VDD.n7041 VDD.n7040 23.1255
R20863 VDD.n5098 VDD.n5094 23.1255
R20864 VDD.n7047 VDD.n5094 23.1255
R20865 VDD.n7051 VDD.n5093 23.1255
R20866 VDD.n7051 VDD.n7050 23.1255
R20867 VDD.n5088 VDD.n5084 23.1255
R20868 VDD.n7057 VDD.n5084 23.1255
R20869 VDD.n7061 VDD.n5083 23.1255
R20870 VDD.n7061 VDD.n7060 23.1255
R20871 VDD.n5077 VDD.n5073 23.1255
R20872 VDD.n7067 VDD.n5073 23.1255
R20873 VDD.n7071 VDD.n5072 23.1255
R20874 VDD.n7071 VDD.n7070 23.1255
R20875 VDD.n5064 VDD.n5060 23.1255
R20876 VDD.n7077 VDD.n5060 23.1255
R20877 VDD.n7081 VDD.n5059 23.1255
R20878 VDD.n7081 VDD.n7080 23.1255
R20879 VDD.n5054 VDD.n5050 23.1255
R20880 VDD.n7087 VDD.n5050 23.1255
R20881 VDD.n7091 VDD.n5049 23.1255
R20882 VDD.n7091 VDD.n7090 23.1255
R20883 VDD.n5043 VDD.n5039 23.1255
R20884 VDD.n7097 VDD.n5039 23.1255
R20885 VDD.n6075 VDD.n6074 23.1255
R20886 VDD.n6076 VDD.n6075 23.1255
R20887 VDD.n6082 VDD.n6081 23.1255
R20888 VDD.n6083 VDD.n6082 23.1255
R20889 VDD.n6085 VDD.n6084 23.1255
R20890 VDD.n6086 VDD.n6085 23.1255
R20891 VDD.n6092 VDD.n6091 23.1255
R20892 VDD.n6093 VDD.n6092 23.1255
R20893 VDD.n6095 VDD.n6094 23.1255
R20894 VDD.n6096 VDD.n6095 23.1255
R20895 VDD.n6102 VDD.n6101 23.1255
R20896 VDD.n6103 VDD.n6102 23.1255
R20897 VDD.n6105 VDD.n6104 23.1255
R20898 VDD.n6106 VDD.n6105 23.1255
R20899 VDD.n6112 VDD.n6111 23.1255
R20900 VDD.n6113 VDD.n6112 23.1255
R20901 VDD.n6122 VDD.n6121 23.1255
R20902 VDD.n6123 VDD.n6122 23.1255
R20903 VDD.n6129 VDD.n6128 23.1255
R20904 VDD.n6130 VDD.n6129 23.1255
R20905 VDD.n6132 VDD.n6131 23.1255
R20906 VDD.n6133 VDD.n6132 23.1255
R20907 VDD.n6139 VDD.n6138 23.1255
R20908 VDD.n6140 VDD.n6139 23.1255
R20909 VDD.n6142 VDD.n6141 23.1255
R20910 VDD.n6143 VDD.n6142 23.1255
R20911 VDD.n6149 VDD.n6148 23.1255
R20912 VDD.n6150 VDD.n6149 23.1255
R20913 VDD.n6152 VDD.n6151 23.1255
R20914 VDD.n6153 VDD.n6152 23.1255
R20915 VDD.n6159 VDD.n6158 23.1255
R20916 VDD.n6160 VDD.n6159 23.1255
R20917 VDD.n6162 VDD.n6161 23.1255
R20918 VDD.n6163 VDD.n6162 23.1255
R20919 VDD.n6169 VDD.n6168 23.1255
R20920 VDD.n6170 VDD.n6169 23.1255
R20921 VDD.n6181 VDD.n6179 23.1255
R20922 VDD.n6179 VDD.n6171 23.1255
R20923 VDD.n6182 VDD.n6180 23.1255
R20924 VDD.n6180 VDD.n6178 23.1255
R20925 VDD.n6176 VDD.n5940 23.1255
R20926 VDD.n6177 VDD.n6176 23.1255
R20927 VDD.n6193 VDD.n6192 23.1255
R20928 VDD.n6194 VDD.n6193 23.1255
R20929 VDD.n6196 VDD.n6195 23.1255
R20930 VDD.n6197 VDD.n6196 23.1255
R20931 VDD.n6203 VDD.n6202 23.1255
R20932 VDD.n6204 VDD.n6203 23.1255
R20933 VDD.n6206 VDD.n6205 23.1255
R20934 VDD.n6207 VDD.n6206 23.1255
R20935 VDD.n6213 VDD.n6212 23.1255
R20936 VDD.n6214 VDD.n6213 23.1255
R20937 VDD.n6216 VDD.n6215 23.1255
R20938 VDD.n6217 VDD.n6216 23.1255
R20939 VDD.n6223 VDD.n6222 23.1255
R20940 VDD.n6224 VDD.n6223 23.1255
R20941 VDD.n6226 VDD.n6225 23.1255
R20942 VDD.n6227 VDD.n6226 23.1255
R20943 VDD.n6233 VDD.n6232 23.1255
R20944 VDD.n6234 VDD.n6233 23.1255
R20945 VDD.n6236 VDD.n6235 23.1255
R20946 VDD.n6237 VDD.n6236 23.1255
R20947 VDD.n6243 VDD.n6242 23.1255
R20948 VDD.n6244 VDD.n6243 23.1255
R20949 VDD.n6253 VDD.n6252 23.1255
R20950 VDD.n6254 VDD.n6253 23.1255
R20951 VDD.n6260 VDD.n6259 23.1255
R20952 VDD.n6261 VDD.n6260 23.1255
R20953 VDD.n6263 VDD.n6262 23.1255
R20954 VDD.n6264 VDD.n6263 23.1255
R20955 VDD.n6270 VDD.n6269 23.1255
R20956 VDD.n6271 VDD.n6270 23.1255
R20957 VDD.n6273 VDD.n6272 23.1255
R20958 VDD.n6274 VDD.n6273 23.1255
R20959 VDD.n6280 VDD.n6279 23.1255
R20960 VDD.n6281 VDD.n6280 23.1255
R20961 VDD.n6283 VDD.n6282 23.1255
R20962 VDD.n6284 VDD.n6283 23.1255
R20963 VDD.n6290 VDD.n6289 23.1255
R20964 VDD.n6291 VDD.n6290 23.1255
R20965 VDD.n6293 VDD.n6292 23.1255
R20966 VDD.n6294 VDD.n6293 23.1255
R20967 VDD.n6300 VDD.n6299 23.1255
R20968 VDD.n6301 VDD.n6300 23.1255
R20969 VDD.n6312 VDD.n6310 23.1255
R20970 VDD.n6310 VDD.n6302 23.1255
R20971 VDD.n6313 VDD.n6311 23.1255
R20972 VDD.n6311 VDD.n6309 23.1255
R20973 VDD.n6307 VDD.n5812 23.1255
R20974 VDD.n6308 VDD.n6307 23.1255
R20975 VDD.n6324 VDD.n6323 23.1255
R20976 VDD.n6325 VDD.n6324 23.1255
R20977 VDD.n6327 VDD.n6326 23.1255
R20978 VDD.n6328 VDD.n6327 23.1255
R20979 VDD.n6334 VDD.n6333 23.1255
R20980 VDD.n6335 VDD.n6334 23.1255
R20981 VDD.n6337 VDD.n6336 23.1255
R20982 VDD.n6338 VDD.n6337 23.1255
R20983 VDD.n6344 VDD.n6343 23.1255
R20984 VDD.n6345 VDD.n6344 23.1255
R20985 VDD.n6347 VDD.n6346 23.1255
R20986 VDD.n6348 VDD.n6347 23.1255
R20987 VDD.n6354 VDD.n6353 23.1255
R20988 VDD.n6355 VDD.n6354 23.1255
R20989 VDD.n6357 VDD.n6356 23.1255
R20990 VDD.n6358 VDD.n6357 23.1255
R20991 VDD.n6364 VDD.n6363 23.1255
R20992 VDD.n6365 VDD.n6364 23.1255
R20993 VDD.n6367 VDD.n6366 23.1255
R20994 VDD.n6368 VDD.n6367 23.1255
R20995 VDD.n6374 VDD.n6373 23.1255
R20996 VDD.n6375 VDD.n6374 23.1255
R20997 VDD.n6384 VDD.n6383 23.1255
R20998 VDD.n6385 VDD.n6384 23.1255
R20999 VDD.n6391 VDD.n6390 23.1255
R21000 VDD.n6392 VDD.n6391 23.1255
R21001 VDD.n6394 VDD.n6393 23.1255
R21002 VDD.n6395 VDD.n6394 23.1255
R21003 VDD.n6401 VDD.n6400 23.1255
R21004 VDD.n6402 VDD.n6401 23.1255
R21005 VDD.n6404 VDD.n6403 23.1255
R21006 VDD.n6405 VDD.n6404 23.1255
R21007 VDD.n6411 VDD.n6410 23.1255
R21008 VDD.n6412 VDD.n6411 23.1255
R21009 VDD.n6414 VDD.n6413 23.1255
R21010 VDD.n6415 VDD.n6414 23.1255
R21011 VDD.n6421 VDD.n6420 23.1255
R21012 VDD.n6422 VDD.n6421 23.1255
R21013 VDD.n6424 VDD.n6423 23.1255
R21014 VDD.n6425 VDD.n6424 23.1255
R21015 VDD.n6431 VDD.n6430 23.1255
R21016 VDD.n6432 VDD.n6431 23.1255
R21017 VDD.n6443 VDD.n6441 23.1255
R21018 VDD.n6441 VDD.n6433 23.1255
R21019 VDD.n6444 VDD.n6442 23.1255
R21020 VDD.n6442 VDD.n6440 23.1255
R21021 VDD.n6438 VDD.n5684 23.1255
R21022 VDD.n6439 VDD.n6438 23.1255
R21023 VDD.n6455 VDD.n6454 23.1255
R21024 VDD.n6456 VDD.n6455 23.1255
R21025 VDD.n6458 VDD.n6457 23.1255
R21026 VDD.n6459 VDD.n6458 23.1255
R21027 VDD.n6465 VDD.n6464 23.1255
R21028 VDD.n6466 VDD.n6465 23.1255
R21029 VDD.n6468 VDD.n6467 23.1255
R21030 VDD.n6469 VDD.n6468 23.1255
R21031 VDD.n6475 VDD.n6474 23.1255
R21032 VDD.n6476 VDD.n6475 23.1255
R21033 VDD.n6478 VDD.n6477 23.1255
R21034 VDD.n6479 VDD.n6478 23.1255
R21035 VDD.n6485 VDD.n6484 23.1255
R21036 VDD.n6486 VDD.n6485 23.1255
R21037 VDD.n6488 VDD.n6487 23.1255
R21038 VDD.n6489 VDD.n6488 23.1255
R21039 VDD.n6495 VDD.n6494 23.1255
R21040 VDD.n6496 VDD.n6495 23.1255
R21041 VDD.n6498 VDD.n6497 23.1255
R21042 VDD.n6499 VDD.n6498 23.1255
R21043 VDD.n6505 VDD.n6504 23.1255
R21044 VDD.n6506 VDD.n6505 23.1255
R21045 VDD.n6515 VDD.n6514 23.1255
R21046 VDD.n6516 VDD.n6515 23.1255
R21047 VDD.n6522 VDD.n6521 23.1255
R21048 VDD.n6523 VDD.n6522 23.1255
R21049 VDD.n6525 VDD.n6524 23.1255
R21050 VDD.n6526 VDD.n6525 23.1255
R21051 VDD.n6532 VDD.n6531 23.1255
R21052 VDD.n6533 VDD.n6532 23.1255
R21053 VDD.n6535 VDD.n6534 23.1255
R21054 VDD.n6536 VDD.n6535 23.1255
R21055 VDD.n6542 VDD.n6541 23.1255
R21056 VDD.n6543 VDD.n6542 23.1255
R21057 VDD.n6545 VDD.n6544 23.1255
R21058 VDD.n6546 VDD.n6545 23.1255
R21059 VDD.n6552 VDD.n6551 23.1255
R21060 VDD.n6553 VDD.n6552 23.1255
R21061 VDD.n6555 VDD.n6554 23.1255
R21062 VDD.n6556 VDD.n6555 23.1255
R21063 VDD.n6562 VDD.n6561 23.1255
R21064 VDD.n6563 VDD.n6562 23.1255
R21065 VDD.n6574 VDD.n6572 23.1255
R21066 VDD.n6572 VDD.n6564 23.1255
R21067 VDD.n6575 VDD.n6573 23.1255
R21068 VDD.n6573 VDD.n6571 23.1255
R21069 VDD.n6569 VDD.n5556 23.1255
R21070 VDD.n6570 VDD.n6569 23.1255
R21071 VDD.n6586 VDD.n6585 23.1255
R21072 VDD.n6587 VDD.n6586 23.1255
R21073 VDD.n6589 VDD.n6588 23.1255
R21074 VDD.n6590 VDD.n6589 23.1255
R21075 VDD.n6596 VDD.n6595 23.1255
R21076 VDD.n6597 VDD.n6596 23.1255
R21077 VDD.n6599 VDD.n6598 23.1255
R21078 VDD.n6600 VDD.n6599 23.1255
R21079 VDD.n6606 VDD.n6605 23.1255
R21080 VDD.n6607 VDD.n6606 23.1255
R21081 VDD.n6609 VDD.n6608 23.1255
R21082 VDD.n6610 VDD.n6609 23.1255
R21083 VDD.n6616 VDD.n6615 23.1255
R21084 VDD.n6617 VDD.n6616 23.1255
R21085 VDD.n6619 VDD.n6618 23.1255
R21086 VDD.n6620 VDD.n6619 23.1255
R21087 VDD.n6626 VDD.n6625 23.1255
R21088 VDD.n6627 VDD.n6626 23.1255
R21089 VDD.n6629 VDD.n6628 23.1255
R21090 VDD.n6630 VDD.n6629 23.1255
R21091 VDD.n6636 VDD.n6635 23.1255
R21092 VDD.n6637 VDD.n6636 23.1255
R21093 VDD.n6646 VDD.n6645 23.1255
R21094 VDD.n6647 VDD.n6646 23.1255
R21095 VDD.n6653 VDD.n6652 23.1255
R21096 VDD.n6654 VDD.n6653 23.1255
R21097 VDD.n6656 VDD.n6655 23.1255
R21098 VDD.n6657 VDD.n6656 23.1255
R21099 VDD.n6663 VDD.n6662 23.1255
R21100 VDD.n6664 VDD.n6663 23.1255
R21101 VDD.n6666 VDD.n6665 23.1255
R21102 VDD.n6667 VDD.n6666 23.1255
R21103 VDD.n6673 VDD.n6672 23.1255
R21104 VDD.n6674 VDD.n6673 23.1255
R21105 VDD.n6676 VDD.n6675 23.1255
R21106 VDD.n6677 VDD.n6676 23.1255
R21107 VDD.n6683 VDD.n6682 23.1255
R21108 VDD.n6684 VDD.n6683 23.1255
R21109 VDD.n6686 VDD.n6685 23.1255
R21110 VDD.n6687 VDD.n6686 23.1255
R21111 VDD.n6693 VDD.n6692 23.1255
R21112 VDD.n6694 VDD.n6693 23.1255
R21113 VDD.n6705 VDD.n6703 23.1255
R21114 VDD.n6703 VDD.n6695 23.1255
R21115 VDD.n6706 VDD.n6704 23.1255
R21116 VDD.n6704 VDD.n6702 23.1255
R21117 VDD.n6700 VDD.n5428 23.1255
R21118 VDD.n6701 VDD.n6700 23.1255
R21119 VDD.n6717 VDD.n6716 23.1255
R21120 VDD.n6718 VDD.n6717 23.1255
R21121 VDD.n6720 VDD.n6719 23.1255
R21122 VDD.n6721 VDD.n6720 23.1255
R21123 VDD.n6727 VDD.n6726 23.1255
R21124 VDD.n6728 VDD.n6727 23.1255
R21125 VDD.n6730 VDD.n6729 23.1255
R21126 VDD.n6731 VDD.n6730 23.1255
R21127 VDD.n6737 VDD.n6736 23.1255
R21128 VDD.n6738 VDD.n6737 23.1255
R21129 VDD.n6740 VDD.n6739 23.1255
R21130 VDD.n6741 VDD.n6740 23.1255
R21131 VDD.n6747 VDD.n6746 23.1255
R21132 VDD.n6748 VDD.n6747 23.1255
R21133 VDD.n6750 VDD.n6749 23.1255
R21134 VDD.n6751 VDD.n6750 23.1255
R21135 VDD.n6757 VDD.n6756 23.1255
R21136 VDD.n6758 VDD.n6757 23.1255
R21137 VDD.n6760 VDD.n6759 23.1255
R21138 VDD.n6761 VDD.n6760 23.1255
R21139 VDD.n6767 VDD.n6766 23.1255
R21140 VDD.n6768 VDD.n6767 23.1255
R21141 VDD.n6777 VDD.n6776 23.1255
R21142 VDD.n6778 VDD.n6777 23.1255
R21143 VDD.n6784 VDD.n6783 23.1255
R21144 VDD.n6785 VDD.n6784 23.1255
R21145 VDD.n6787 VDD.n6786 23.1255
R21146 VDD.n6788 VDD.n6787 23.1255
R21147 VDD.n6794 VDD.n6793 23.1255
R21148 VDD.n6795 VDD.n6794 23.1255
R21149 VDD.n6797 VDD.n6796 23.1255
R21150 VDD.n6798 VDD.n6797 23.1255
R21151 VDD.n6804 VDD.n6803 23.1255
R21152 VDD.n6805 VDD.n6804 23.1255
R21153 VDD.n6807 VDD.n6806 23.1255
R21154 VDD.n6808 VDD.n6807 23.1255
R21155 VDD.n6814 VDD.n6813 23.1255
R21156 VDD.n6815 VDD.n6814 23.1255
R21157 VDD.n6817 VDD.n6816 23.1255
R21158 VDD.n6818 VDD.n6817 23.1255
R21159 VDD.n6824 VDD.n6823 23.1255
R21160 VDD.n6825 VDD.n6824 23.1255
R21161 VDD.n6836 VDD.n6834 23.1255
R21162 VDD.n6834 VDD.n6826 23.1255
R21163 VDD.n6837 VDD.n6835 23.1255
R21164 VDD.n6835 VDD.n6833 23.1255
R21165 VDD.n6831 VDD.n5300 23.1255
R21166 VDD.n6832 VDD.n6831 23.1255
R21167 VDD.n6848 VDD.n6847 23.1255
R21168 VDD.n6849 VDD.n6848 23.1255
R21169 VDD.n6851 VDD.n6850 23.1255
R21170 VDD.n6852 VDD.n6851 23.1255
R21171 VDD.n6858 VDD.n6857 23.1255
R21172 VDD.n6859 VDD.n6858 23.1255
R21173 VDD.n6861 VDD.n6860 23.1255
R21174 VDD.n6862 VDD.n6861 23.1255
R21175 VDD.n6868 VDD.n6867 23.1255
R21176 VDD.n6869 VDD.n6868 23.1255
R21177 VDD.n6871 VDD.n6870 23.1255
R21178 VDD.n6872 VDD.n6871 23.1255
R21179 VDD.n6878 VDD.n6877 23.1255
R21180 VDD.n6879 VDD.n6878 23.1255
R21181 VDD.n6881 VDD.n6880 23.1255
R21182 VDD.n6882 VDD.n6881 23.1255
R21183 VDD.n6888 VDD.n6887 23.1255
R21184 VDD.n6889 VDD.n6888 23.1255
R21185 VDD.n6891 VDD.n6890 23.1255
R21186 VDD.n6892 VDD.n6891 23.1255
R21187 VDD.n6898 VDD.n6897 23.1255
R21188 VDD.n6899 VDD.n6898 23.1255
R21189 VDD.n6908 VDD.n6907 23.1255
R21190 VDD.n6909 VDD.n6908 23.1255
R21191 VDD.n6915 VDD.n6914 23.1255
R21192 VDD.n6916 VDD.n6915 23.1255
R21193 VDD.n6918 VDD.n6917 23.1255
R21194 VDD.n6919 VDD.n6918 23.1255
R21195 VDD.n6925 VDD.n6924 23.1255
R21196 VDD.n6926 VDD.n6925 23.1255
R21197 VDD.n6928 VDD.n6927 23.1255
R21198 VDD.n6929 VDD.n6928 23.1255
R21199 VDD.n6935 VDD.n6934 23.1255
R21200 VDD.n6936 VDD.n6935 23.1255
R21201 VDD.n6938 VDD.n6937 23.1255
R21202 VDD.n6939 VDD.n6938 23.1255
R21203 VDD.n6945 VDD.n6944 23.1255
R21204 VDD.n6946 VDD.n6945 23.1255
R21205 VDD.n6948 VDD.n6947 23.1255
R21206 VDD.n6949 VDD.n6948 23.1255
R21207 VDD.n6955 VDD.n6954 23.1255
R21208 VDD.n6956 VDD.n6955 23.1255
R21209 VDD.n6967 VDD.n6965 23.1255
R21210 VDD.n6965 VDD.n6957 23.1255
R21211 VDD.n6968 VDD.n6966 23.1255
R21212 VDD.n6966 VDD.n6964 23.1255
R21213 VDD.n6962 VDD.n5172 23.1255
R21214 VDD.n6963 VDD.n6962 23.1255
R21215 VDD.n6979 VDD.n6978 23.1255
R21216 VDD.n6980 VDD.n6979 23.1255
R21217 VDD.n6982 VDD.n6981 23.1255
R21218 VDD.n6983 VDD.n6982 23.1255
R21219 VDD.n6989 VDD.n6988 23.1255
R21220 VDD.n6990 VDD.n6989 23.1255
R21221 VDD.n6992 VDD.n6991 23.1255
R21222 VDD.n6993 VDD.n6992 23.1255
R21223 VDD.n6999 VDD.n6998 23.1255
R21224 VDD.n7000 VDD.n6999 23.1255
R21225 VDD.n7002 VDD.n7001 23.1255
R21226 VDD.n7003 VDD.n7002 23.1255
R21227 VDD.n7009 VDD.n7008 23.1255
R21228 VDD.n7010 VDD.n7009 23.1255
R21229 VDD.n7012 VDD.n7011 23.1255
R21230 VDD.n7013 VDD.n7012 23.1255
R21231 VDD.n7019 VDD.n7018 23.1255
R21232 VDD.n7020 VDD.n7019 23.1255
R21233 VDD.n7022 VDD.n7021 23.1255
R21234 VDD.n7023 VDD.n7022 23.1255
R21235 VDD.n7029 VDD.n7028 23.1255
R21236 VDD.n7030 VDD.n7029 23.1255
R21237 VDD.n7039 VDD.n7038 23.1255
R21238 VDD.n7040 VDD.n7039 23.1255
R21239 VDD.n7046 VDD.n7045 23.1255
R21240 VDD.n7047 VDD.n7046 23.1255
R21241 VDD.n7049 VDD.n7048 23.1255
R21242 VDD.n7050 VDD.n7049 23.1255
R21243 VDD.n7056 VDD.n7055 23.1255
R21244 VDD.n7057 VDD.n7056 23.1255
R21245 VDD.n7059 VDD.n7058 23.1255
R21246 VDD.n7060 VDD.n7059 23.1255
R21247 VDD.n7066 VDD.n7065 23.1255
R21248 VDD.n7067 VDD.n7066 23.1255
R21249 VDD.n7069 VDD.n7068 23.1255
R21250 VDD.n7070 VDD.n7069 23.1255
R21251 VDD.n7076 VDD.n7075 23.1255
R21252 VDD.n7077 VDD.n7076 23.1255
R21253 VDD.n7079 VDD.n7078 23.1255
R21254 VDD.n7080 VDD.n7079 23.1255
R21255 VDD.n7086 VDD.n7085 23.1255
R21256 VDD.n7087 VDD.n7086 23.1255
R21257 VDD.n7089 VDD.n7088 23.1255
R21258 VDD.n7090 VDD.n7089 23.1255
R21259 VDD.n7096 VDD.n7095 23.1255
R21260 VDD.n7097 VDD.n7096 23.1255
R21261 VDD.n7098 VDD.n5035 23.1255
R21262 VDD.n7099 VDD.n7098 23.1255
R21263 VDD.n7102 VDD.n7101 23.1255
R21264 VDD.n6072 VDD.n6071 23.1255
R21265 VDD.n6073 VDD.n6072 23.1255
R21266 VDD.n6062 VDD.n6061 23.1255
R21267 VDD.n6063 VDD.n6062 23.1255
R21268 VDD.n7121 VDD.n7120 23.1255
R21269 VDD.n7122 VDD.n7121 23.1255
R21270 VDD.n7118 VDD.n7117 23.1255
R21271 VDD.n7117 VDD.n7116 23.1255
R21272 VDD.n7114 VDD.n7113 23.1255
R21273 VDD.n7115 VDD.n7114 23.1255
R21274 VDD.n7111 VDD.n7110 23.1255
R21275 VDD.n7125 VDD.n7124 23.1255
R21276 VDD.n7124 VDD.n7123 23.1255
R21277 VDD.n139 VDD.n135 23.1255
R21278 VDD.n7142 VDD.n7141 23.1255
R21279 VDD.n7143 VDD.n7142 23.1255
R21280 VDD.n7139 VDD.n7138 23.1255
R21281 VDD.n7138 VDD.n7137 23.1255
R21282 VDD.n7135 VDD.n7134 23.1255
R21283 VDD.n7136 VDD.n7135 23.1255
R21284 VDD.n7132 VDD.n7131 23.1255
R21285 VDD.n7146 VDD.n7145 23.1255
R21286 VDD.n7145 VDD.n7144 23.1255
R21287 VDD.n120 VDD.n116 23.1255
R21288 VDD.n7163 VDD.n7162 23.1255
R21289 VDD.n7164 VDD.n7163 23.1255
R21290 VDD.n7160 VDD.n7159 23.1255
R21291 VDD.n7159 VDD.n7158 23.1255
R21292 VDD.n7156 VDD.n7155 23.1255
R21293 VDD.n7157 VDD.n7156 23.1255
R21294 VDD.n7153 VDD.n7152 23.1255
R21295 VDD.n7167 VDD.n7166 23.1255
R21296 VDD.n7166 VDD.n7165 23.1255
R21297 VDD.n101 VDD.n97 23.1255
R21298 VDD.n7184 VDD.n7183 23.1255
R21299 VDD.n7185 VDD.n7184 23.1255
R21300 VDD.n7181 VDD.n7180 23.1255
R21301 VDD.n7180 VDD.n7179 23.1255
R21302 VDD.n7177 VDD.n7176 23.1255
R21303 VDD.n7178 VDD.n7177 23.1255
R21304 VDD.n7174 VDD.n7173 23.1255
R21305 VDD.n7188 VDD.n7187 23.1255
R21306 VDD.n7187 VDD.n7186 23.1255
R21307 VDD.n82 VDD.n78 23.1255
R21308 VDD.n7205 VDD.n7204 23.1255
R21309 VDD.n7206 VDD.n7205 23.1255
R21310 VDD.n7202 VDD.n7201 23.1255
R21311 VDD.n7201 VDD.n7200 23.1255
R21312 VDD.n7198 VDD.n7197 23.1255
R21313 VDD.n7199 VDD.n7198 23.1255
R21314 VDD.n7195 VDD.n7194 23.1255
R21315 VDD.n7209 VDD.n7208 23.1255
R21316 VDD.n7208 VDD.n7207 23.1255
R21317 VDD.n63 VDD.n59 23.1255
R21318 VDD.n7226 VDD.n7225 23.1255
R21319 VDD.n7227 VDD.n7226 23.1255
R21320 VDD.n7223 VDD.n7222 23.1255
R21321 VDD.n7222 VDD.n7221 23.1255
R21322 VDD.n7219 VDD.n7218 23.1255
R21323 VDD.n7220 VDD.n7219 23.1255
R21324 VDD.n7216 VDD.n7215 23.1255
R21325 VDD.n7230 VDD.n7229 23.1255
R21326 VDD.n7229 VDD.n7228 23.1255
R21327 VDD.n44 VDD.n40 23.1255
R21328 VDD.n7247 VDD.n7246 23.1255
R21329 VDD.n7248 VDD.n7247 23.1255
R21330 VDD.n7244 VDD.n7243 23.1255
R21331 VDD.n7243 VDD.n7242 23.1255
R21332 VDD.n7240 VDD.n7239 23.1255
R21333 VDD.n7241 VDD.n7240 23.1255
R21334 VDD.n7237 VDD.n7236 23.1255
R21335 VDD.n7251 VDD.n7250 23.1255
R21336 VDD.n7250 VDD.n7249 23.1255
R21337 VDD.n25 VDD.n21 23.1255
R21338 VDD.n7268 VDD.n7267 23.1255
R21339 VDD.n7269 VDD.n7268 23.1255
R21340 VDD.n7265 VDD.n7264 23.1255
R21341 VDD.n7264 VDD.n7263 23.1255
R21342 VDD.n7261 VDD.n7260 23.1255
R21343 VDD.n7262 VDD.n7261 23.1255
R21344 VDD.n7258 VDD.n7257 23.1255
R21345 VDD.n7272 VDD.n7271 23.1255
R21346 VDD.n7271 VDD.n7270 23.1255
R21347 VDD.n6 VDD.n2 23.1255
R21348 VDD.n2224 VDD 22.8404
R21349 VDD.n7309 VDD.n7279 21.3068
R21350 VDD.n7309 VDD.n7308 21.3068
R21351 VDD.n7277 VDD.t884 20.9643
R21352 VDD.n7286 VDD.n7275 20.9422
R21353 VDD.n7289 VDD.n7288 20.4313
R21354 VDD.n2484 VDD 20.4275
R21355 VDD.n2483 VDD 20.3024
R21356 VDD.n7276 VDD.t45 18.427
R21357 VDD.n7276 VDD.t43 18.427
R21358 VDD.n2742 VDD 17.7644
R21359 VDD.n2743 VDD 17.6357
R21360 VDD.n165 VDD.n160 15.5222
R21361 VDD.n668 VDD.n663 15.5222
R21362 VDD.n927 VDD.n922 15.5222
R21363 VDD.n1186 VDD.n1181 15.5222
R21364 VDD.n1445 VDD.n1440 15.5222
R21365 VDD.n1704 VDD.n1699 15.5222
R21366 VDD.n1963 VDD.n1958 15.5222
R21367 VDD.n2222 VDD.n2217 15.5222
R21368 VDD.n2481 VDD.n2476 15.5222
R21369 VDD.n2740 VDD.n2735 15.5222
R21370 VDD.n2999 VDD.n2994 15.5222
R21371 VDD.n3258 VDD.n3253 15.5222
R21372 VDD.n3517 VDD.n3512 15.5222
R21373 VDD.n3776 VDD.n3771 15.5222
R21374 VDD.n4035 VDD.n4030 15.5222
R21375 VDD.n4294 VDD.n4289 15.5222
R21376 VDD.n4553 VDD.n4548 15.5222
R21377 VDD.n3001 VDD 15.2264
R21378 VDD.n3002 VDD 14.8439
R21379 VDD.n7332 VDD.n7275 14.7125
R21380 VDD VDD.n7332 13.2701
R21381 VDD.n3260 VDD 12.6884
R21382 VDD.n3261 VDD 12.0521
R21383 VDD.n3519 VDD 10.1504
R21384 VDD.n3520 VDD 9.26028
R21385 VDD.n5034 VDD 9.24202
R21386 VDD.n414 VDD.n413 9.20653
R21387 VDD.n151 VDD.n150 8.357
R21388 VDD.n132 VDD.n131 8.357
R21389 VDD.n113 VDD.n112 8.357
R21390 VDD.n94 VDD.n93 8.357
R21391 VDD.n75 VDD.n74 8.357
R21392 VDD.n56 VDD.n55 8.357
R21393 VDD.n37 VDD.n36 8.357
R21394 VDD.n18 VDD.n17 8.357
R21395 VDD.n166 VDD.n165 8.24202
R21396 VDD.n4724 VDD 8.21517
R21397 VDD.n4747 VDD 8.21517
R21398 VDD.n4765 VDD 8.21517
R21399 VDD.n4788 VDD 8.21517
R21400 VDD.n4806 VDD 8.21517
R21401 VDD.n4829 VDD 8.21517
R21402 VDD.n4847 VDD 8.21517
R21403 VDD.n4870 VDD 8.21517
R21404 VDD.n4888 VDD 8.21517
R21405 VDD.n4911 VDD 8.21517
R21406 VDD.n4929 VDD 8.21517
R21407 VDD.n4952 VDD 8.21517
R21408 VDD.n4970 VDD 8.21517
R21409 VDD.n4993 VDD 8.21517
R21410 VDD.n5011 VDD 8.21517
R21411 VDD.n7106 VDD 8.17952
R21412 VDD.n409 VDD.n408 7.9105
R21413 VDD.n657 VDD.n656 7.9105
R21414 VDD.n916 VDD.n915 7.9105
R21415 VDD.n1175 VDD.n1174 7.9105
R21416 VDD.n1434 VDD.n1433 7.9105
R21417 VDD.n1693 VDD.n1692 7.9105
R21418 VDD.n1952 VDD.n1951 7.9105
R21419 VDD.n2211 VDD.n2210 7.9105
R21420 VDD.n2470 VDD.n2469 7.9105
R21421 VDD.n2729 VDD.n2728 7.9105
R21422 VDD.n2988 VDD.n2987 7.9105
R21423 VDD.n3247 VDD.n3246 7.9105
R21424 VDD.n3506 VDD.n3505 7.9105
R21425 VDD.n3765 VDD.n3764 7.9105
R21426 VDD.n4024 VDD.n4023 7.9105
R21427 VDD.n4283 VDD.n4282 7.9105
R21428 VDD.n4542 VDD.n4541 7.9105
R21429 VDD.n669 VDD.n668 7.83713
R21430 VDD.n928 VDD.n927 7.83713
R21431 VDD.n1187 VDD.n1186 7.83713
R21432 VDD.n1446 VDD.n1445 7.83713
R21433 VDD.n1705 VDD.n1704 7.83713
R21434 VDD.n1964 VDD.n1963 7.83713
R21435 VDD.n2223 VDD.n2222 7.83713
R21436 VDD.n2482 VDD.n2481 7.83713
R21437 VDD.n2741 VDD.n2740 7.83713
R21438 VDD.n3000 VDD.n2999 7.83713
R21439 VDD.n3259 VDD.n3258 7.83713
R21440 VDD.n3518 VDD.n3517 7.83713
R21441 VDD.n3777 VDD.n3776 7.83713
R21442 VDD.n4036 VDD.n4035 7.83713
R21443 VDD.n4295 VDD.n4294 7.83713
R21444 VDD.n4554 VDD.n4553 7.83713
R21445 VDD.n3778 VDD 7.61236
R21446 VDD.n396 VDD.n192 7.39606
R21447 VDD.n396 VDD.n193 7.39606
R21448 VDD.n405 VDD.n171 7.39606
R21449 VDD.n405 VDD.n173 7.39606
R21450 VDD.n291 VDD.n279 7.39606
R21451 VDD.n291 VDD.n290 7.39606
R21452 VDD.n367 VDD.n276 7.39606
R21453 VDD.n368 VDD.n367 7.39606
R21454 VDD.n364 VDD.n352 7.39606
R21455 VDD.n364 VDD.n363 7.39606
R21456 VDD.n348 VDD.n336 7.39606
R21457 VDD.n348 VDD.n347 7.39606
R21458 VDD.n325 VDD.n313 7.39606
R21459 VDD.n325 VDD.n324 7.39606
R21460 VDD.n309 VDD.n297 7.39606
R21461 VDD.n309 VDD.n308 7.39606
R21462 VDD.n257 VDD.n255 7.39606
R21463 VDD.n258 VDD.n257 7.39606
R21464 VDD.n383 VDD.n230 7.39606
R21465 VDD.n383 VDD.n382 7.39606
R21466 VDD.n388 VDD.n227 7.39606
R21467 VDD.n389 VDD.n388 7.39606
R21468 VDD.n644 VDD.n440 7.39606
R21469 VDD.n644 VDD.n441 7.39606
R21470 VDD.n653 VDD.n419 7.39606
R21471 VDD.n653 VDD.n421 7.39606
R21472 VDD.n539 VDD.n527 7.39606
R21473 VDD.n539 VDD.n538 7.39606
R21474 VDD.n615 VDD.n524 7.39606
R21475 VDD.n616 VDD.n615 7.39606
R21476 VDD.n612 VDD.n600 7.39606
R21477 VDD.n612 VDD.n611 7.39606
R21478 VDD.n596 VDD.n584 7.39606
R21479 VDD.n596 VDD.n595 7.39606
R21480 VDD.n573 VDD.n561 7.39606
R21481 VDD.n573 VDD.n572 7.39606
R21482 VDD.n557 VDD.n545 7.39606
R21483 VDD.n557 VDD.n556 7.39606
R21484 VDD.n505 VDD.n503 7.39606
R21485 VDD.n506 VDD.n505 7.39606
R21486 VDD.n631 VDD.n478 7.39606
R21487 VDD.n631 VDD.n630 7.39606
R21488 VDD.n636 VDD.n475 7.39606
R21489 VDD.n637 VDD.n636 7.39606
R21490 VDD.n903 VDD.n699 7.39606
R21491 VDD.n903 VDD.n700 7.39606
R21492 VDD.n912 VDD.n678 7.39606
R21493 VDD.n912 VDD.n680 7.39606
R21494 VDD.n798 VDD.n786 7.39606
R21495 VDD.n798 VDD.n797 7.39606
R21496 VDD.n874 VDD.n783 7.39606
R21497 VDD.n875 VDD.n874 7.39606
R21498 VDD.n871 VDD.n859 7.39606
R21499 VDD.n871 VDD.n870 7.39606
R21500 VDD.n855 VDD.n843 7.39606
R21501 VDD.n855 VDD.n854 7.39606
R21502 VDD.n832 VDD.n820 7.39606
R21503 VDD.n832 VDD.n831 7.39606
R21504 VDD.n816 VDD.n804 7.39606
R21505 VDD.n816 VDD.n815 7.39606
R21506 VDD.n764 VDD.n762 7.39606
R21507 VDD.n765 VDD.n764 7.39606
R21508 VDD.n890 VDD.n737 7.39606
R21509 VDD.n890 VDD.n889 7.39606
R21510 VDD.n895 VDD.n734 7.39606
R21511 VDD.n896 VDD.n895 7.39606
R21512 VDD.n1162 VDD.n958 7.39606
R21513 VDD.n1162 VDD.n959 7.39606
R21514 VDD.n1171 VDD.n937 7.39606
R21515 VDD.n1171 VDD.n939 7.39606
R21516 VDD.n1057 VDD.n1045 7.39606
R21517 VDD.n1057 VDD.n1056 7.39606
R21518 VDD.n1133 VDD.n1042 7.39606
R21519 VDD.n1134 VDD.n1133 7.39606
R21520 VDD.n1130 VDD.n1118 7.39606
R21521 VDD.n1130 VDD.n1129 7.39606
R21522 VDD.n1114 VDD.n1102 7.39606
R21523 VDD.n1114 VDD.n1113 7.39606
R21524 VDD.n1091 VDD.n1079 7.39606
R21525 VDD.n1091 VDD.n1090 7.39606
R21526 VDD.n1075 VDD.n1063 7.39606
R21527 VDD.n1075 VDD.n1074 7.39606
R21528 VDD.n1023 VDD.n1021 7.39606
R21529 VDD.n1024 VDD.n1023 7.39606
R21530 VDD.n1149 VDD.n996 7.39606
R21531 VDD.n1149 VDD.n1148 7.39606
R21532 VDD.n1154 VDD.n993 7.39606
R21533 VDD.n1155 VDD.n1154 7.39606
R21534 VDD.n1421 VDD.n1217 7.39606
R21535 VDD.n1421 VDD.n1218 7.39606
R21536 VDD.n1430 VDD.n1196 7.39606
R21537 VDD.n1430 VDD.n1198 7.39606
R21538 VDD.n1316 VDD.n1304 7.39606
R21539 VDD.n1316 VDD.n1315 7.39606
R21540 VDD.n1392 VDD.n1301 7.39606
R21541 VDD.n1393 VDD.n1392 7.39606
R21542 VDD.n1389 VDD.n1377 7.39606
R21543 VDD.n1389 VDD.n1388 7.39606
R21544 VDD.n1373 VDD.n1361 7.39606
R21545 VDD.n1373 VDD.n1372 7.39606
R21546 VDD.n1350 VDD.n1338 7.39606
R21547 VDD.n1350 VDD.n1349 7.39606
R21548 VDD.n1334 VDD.n1322 7.39606
R21549 VDD.n1334 VDD.n1333 7.39606
R21550 VDD.n1282 VDD.n1280 7.39606
R21551 VDD.n1283 VDD.n1282 7.39606
R21552 VDD.n1408 VDD.n1255 7.39606
R21553 VDD.n1408 VDD.n1407 7.39606
R21554 VDD.n1413 VDD.n1252 7.39606
R21555 VDD.n1414 VDD.n1413 7.39606
R21556 VDD.n1680 VDD.n1476 7.39606
R21557 VDD.n1680 VDD.n1477 7.39606
R21558 VDD.n1689 VDD.n1455 7.39606
R21559 VDD.n1689 VDD.n1457 7.39606
R21560 VDD.n1575 VDD.n1563 7.39606
R21561 VDD.n1575 VDD.n1574 7.39606
R21562 VDD.n1651 VDD.n1560 7.39606
R21563 VDD.n1652 VDD.n1651 7.39606
R21564 VDD.n1648 VDD.n1636 7.39606
R21565 VDD.n1648 VDD.n1647 7.39606
R21566 VDD.n1632 VDD.n1620 7.39606
R21567 VDD.n1632 VDD.n1631 7.39606
R21568 VDD.n1609 VDD.n1597 7.39606
R21569 VDD.n1609 VDD.n1608 7.39606
R21570 VDD.n1593 VDD.n1581 7.39606
R21571 VDD.n1593 VDD.n1592 7.39606
R21572 VDD.n1541 VDD.n1539 7.39606
R21573 VDD.n1542 VDD.n1541 7.39606
R21574 VDD.n1667 VDD.n1514 7.39606
R21575 VDD.n1667 VDD.n1666 7.39606
R21576 VDD.n1672 VDD.n1511 7.39606
R21577 VDD.n1673 VDD.n1672 7.39606
R21578 VDD.n1939 VDD.n1735 7.39606
R21579 VDD.n1939 VDD.n1736 7.39606
R21580 VDD.n1948 VDD.n1714 7.39606
R21581 VDD.n1948 VDD.n1716 7.39606
R21582 VDD.n1834 VDD.n1822 7.39606
R21583 VDD.n1834 VDD.n1833 7.39606
R21584 VDD.n1910 VDD.n1819 7.39606
R21585 VDD.n1911 VDD.n1910 7.39606
R21586 VDD.n1907 VDD.n1895 7.39606
R21587 VDD.n1907 VDD.n1906 7.39606
R21588 VDD.n1891 VDD.n1879 7.39606
R21589 VDD.n1891 VDD.n1890 7.39606
R21590 VDD.n1868 VDD.n1856 7.39606
R21591 VDD.n1868 VDD.n1867 7.39606
R21592 VDD.n1852 VDD.n1840 7.39606
R21593 VDD.n1852 VDD.n1851 7.39606
R21594 VDD.n1800 VDD.n1798 7.39606
R21595 VDD.n1801 VDD.n1800 7.39606
R21596 VDD.n1926 VDD.n1773 7.39606
R21597 VDD.n1926 VDD.n1925 7.39606
R21598 VDD.n1931 VDD.n1770 7.39606
R21599 VDD.n1932 VDD.n1931 7.39606
R21600 VDD.n2198 VDD.n1994 7.39606
R21601 VDD.n2198 VDD.n1995 7.39606
R21602 VDD.n2207 VDD.n1973 7.39606
R21603 VDD.n2207 VDD.n1975 7.39606
R21604 VDD.n2093 VDD.n2081 7.39606
R21605 VDD.n2093 VDD.n2092 7.39606
R21606 VDD.n2169 VDD.n2078 7.39606
R21607 VDD.n2170 VDD.n2169 7.39606
R21608 VDD.n2166 VDD.n2154 7.39606
R21609 VDD.n2166 VDD.n2165 7.39606
R21610 VDD.n2150 VDD.n2138 7.39606
R21611 VDD.n2150 VDD.n2149 7.39606
R21612 VDD.n2127 VDD.n2115 7.39606
R21613 VDD.n2127 VDD.n2126 7.39606
R21614 VDD.n2111 VDD.n2099 7.39606
R21615 VDD.n2111 VDD.n2110 7.39606
R21616 VDD.n2059 VDD.n2057 7.39606
R21617 VDD.n2060 VDD.n2059 7.39606
R21618 VDD.n2185 VDD.n2032 7.39606
R21619 VDD.n2185 VDD.n2184 7.39606
R21620 VDD.n2190 VDD.n2029 7.39606
R21621 VDD.n2191 VDD.n2190 7.39606
R21622 VDD.n2457 VDD.n2253 7.39606
R21623 VDD.n2457 VDD.n2254 7.39606
R21624 VDD.n2466 VDD.n2232 7.39606
R21625 VDD.n2466 VDD.n2234 7.39606
R21626 VDD.n2352 VDD.n2340 7.39606
R21627 VDD.n2352 VDD.n2351 7.39606
R21628 VDD.n2428 VDD.n2337 7.39606
R21629 VDD.n2429 VDD.n2428 7.39606
R21630 VDD.n2425 VDD.n2413 7.39606
R21631 VDD.n2425 VDD.n2424 7.39606
R21632 VDD.n2409 VDD.n2397 7.39606
R21633 VDD.n2409 VDD.n2408 7.39606
R21634 VDD.n2386 VDD.n2374 7.39606
R21635 VDD.n2386 VDD.n2385 7.39606
R21636 VDD.n2370 VDD.n2358 7.39606
R21637 VDD.n2370 VDD.n2369 7.39606
R21638 VDD.n2318 VDD.n2316 7.39606
R21639 VDD.n2319 VDD.n2318 7.39606
R21640 VDD.n2444 VDD.n2291 7.39606
R21641 VDD.n2444 VDD.n2443 7.39606
R21642 VDD.n2449 VDD.n2288 7.39606
R21643 VDD.n2450 VDD.n2449 7.39606
R21644 VDD.n2716 VDD.n2512 7.39606
R21645 VDD.n2716 VDD.n2513 7.39606
R21646 VDD.n2725 VDD.n2491 7.39606
R21647 VDD.n2725 VDD.n2493 7.39606
R21648 VDD.n2611 VDD.n2599 7.39606
R21649 VDD.n2611 VDD.n2610 7.39606
R21650 VDD.n2687 VDD.n2596 7.39606
R21651 VDD.n2688 VDD.n2687 7.39606
R21652 VDD.n2684 VDD.n2672 7.39606
R21653 VDD.n2684 VDD.n2683 7.39606
R21654 VDD.n2668 VDD.n2656 7.39606
R21655 VDD.n2668 VDD.n2667 7.39606
R21656 VDD.n2645 VDD.n2633 7.39606
R21657 VDD.n2645 VDD.n2644 7.39606
R21658 VDD.n2629 VDD.n2617 7.39606
R21659 VDD.n2629 VDD.n2628 7.39606
R21660 VDD.n2577 VDD.n2575 7.39606
R21661 VDD.n2578 VDD.n2577 7.39606
R21662 VDD.n2703 VDD.n2550 7.39606
R21663 VDD.n2703 VDD.n2702 7.39606
R21664 VDD.n2708 VDD.n2547 7.39606
R21665 VDD.n2709 VDD.n2708 7.39606
R21666 VDD.n2975 VDD.n2771 7.39606
R21667 VDD.n2975 VDD.n2772 7.39606
R21668 VDD.n2984 VDD.n2750 7.39606
R21669 VDD.n2984 VDD.n2752 7.39606
R21670 VDD.n2870 VDD.n2858 7.39606
R21671 VDD.n2870 VDD.n2869 7.39606
R21672 VDD.n2946 VDD.n2855 7.39606
R21673 VDD.n2947 VDD.n2946 7.39606
R21674 VDD.n2943 VDD.n2931 7.39606
R21675 VDD.n2943 VDD.n2942 7.39606
R21676 VDD.n2927 VDD.n2915 7.39606
R21677 VDD.n2927 VDD.n2926 7.39606
R21678 VDD.n2904 VDD.n2892 7.39606
R21679 VDD.n2904 VDD.n2903 7.39606
R21680 VDD.n2888 VDD.n2876 7.39606
R21681 VDD.n2888 VDD.n2887 7.39606
R21682 VDD.n2836 VDD.n2834 7.39606
R21683 VDD.n2837 VDD.n2836 7.39606
R21684 VDD.n2962 VDD.n2809 7.39606
R21685 VDD.n2962 VDD.n2961 7.39606
R21686 VDD.n2967 VDD.n2806 7.39606
R21687 VDD.n2968 VDD.n2967 7.39606
R21688 VDD.n3234 VDD.n3030 7.39606
R21689 VDD.n3234 VDD.n3031 7.39606
R21690 VDD.n3243 VDD.n3009 7.39606
R21691 VDD.n3243 VDD.n3011 7.39606
R21692 VDD.n3129 VDD.n3117 7.39606
R21693 VDD.n3129 VDD.n3128 7.39606
R21694 VDD.n3205 VDD.n3114 7.39606
R21695 VDD.n3206 VDD.n3205 7.39606
R21696 VDD.n3202 VDD.n3190 7.39606
R21697 VDD.n3202 VDD.n3201 7.39606
R21698 VDD.n3186 VDD.n3174 7.39606
R21699 VDD.n3186 VDD.n3185 7.39606
R21700 VDD.n3163 VDD.n3151 7.39606
R21701 VDD.n3163 VDD.n3162 7.39606
R21702 VDD.n3147 VDD.n3135 7.39606
R21703 VDD.n3147 VDD.n3146 7.39606
R21704 VDD.n3095 VDD.n3093 7.39606
R21705 VDD.n3096 VDD.n3095 7.39606
R21706 VDD.n3221 VDD.n3068 7.39606
R21707 VDD.n3221 VDD.n3220 7.39606
R21708 VDD.n3226 VDD.n3065 7.39606
R21709 VDD.n3227 VDD.n3226 7.39606
R21710 VDD.n3493 VDD.n3289 7.39606
R21711 VDD.n3493 VDD.n3290 7.39606
R21712 VDD.n3502 VDD.n3268 7.39606
R21713 VDD.n3502 VDD.n3270 7.39606
R21714 VDD.n3388 VDD.n3376 7.39606
R21715 VDD.n3388 VDD.n3387 7.39606
R21716 VDD.n3464 VDD.n3373 7.39606
R21717 VDD.n3465 VDD.n3464 7.39606
R21718 VDD.n3461 VDD.n3449 7.39606
R21719 VDD.n3461 VDD.n3460 7.39606
R21720 VDD.n3445 VDD.n3433 7.39606
R21721 VDD.n3445 VDD.n3444 7.39606
R21722 VDD.n3422 VDD.n3410 7.39606
R21723 VDD.n3422 VDD.n3421 7.39606
R21724 VDD.n3406 VDD.n3394 7.39606
R21725 VDD.n3406 VDD.n3405 7.39606
R21726 VDD.n3354 VDD.n3352 7.39606
R21727 VDD.n3355 VDD.n3354 7.39606
R21728 VDD.n3480 VDD.n3327 7.39606
R21729 VDD.n3480 VDD.n3479 7.39606
R21730 VDD.n3485 VDD.n3324 7.39606
R21731 VDD.n3486 VDD.n3485 7.39606
R21732 VDD.n3752 VDD.n3548 7.39606
R21733 VDD.n3752 VDD.n3549 7.39606
R21734 VDD.n3761 VDD.n3527 7.39606
R21735 VDD.n3761 VDD.n3529 7.39606
R21736 VDD.n3647 VDD.n3635 7.39606
R21737 VDD.n3647 VDD.n3646 7.39606
R21738 VDD.n3723 VDD.n3632 7.39606
R21739 VDD.n3724 VDD.n3723 7.39606
R21740 VDD.n3720 VDD.n3708 7.39606
R21741 VDD.n3720 VDD.n3719 7.39606
R21742 VDD.n3704 VDD.n3692 7.39606
R21743 VDD.n3704 VDD.n3703 7.39606
R21744 VDD.n3681 VDD.n3669 7.39606
R21745 VDD.n3681 VDD.n3680 7.39606
R21746 VDD.n3665 VDD.n3653 7.39606
R21747 VDD.n3665 VDD.n3664 7.39606
R21748 VDD.n3613 VDD.n3611 7.39606
R21749 VDD.n3614 VDD.n3613 7.39606
R21750 VDD.n3739 VDD.n3586 7.39606
R21751 VDD.n3739 VDD.n3738 7.39606
R21752 VDD.n3744 VDD.n3583 7.39606
R21753 VDD.n3745 VDD.n3744 7.39606
R21754 VDD.n4011 VDD.n3807 7.39606
R21755 VDD.n4011 VDD.n3808 7.39606
R21756 VDD.n4020 VDD.n3786 7.39606
R21757 VDD.n4020 VDD.n3788 7.39606
R21758 VDD.n3906 VDD.n3894 7.39606
R21759 VDD.n3906 VDD.n3905 7.39606
R21760 VDD.n3982 VDD.n3891 7.39606
R21761 VDD.n3983 VDD.n3982 7.39606
R21762 VDD.n3979 VDD.n3967 7.39606
R21763 VDD.n3979 VDD.n3978 7.39606
R21764 VDD.n3963 VDD.n3951 7.39606
R21765 VDD.n3963 VDD.n3962 7.39606
R21766 VDD.n3940 VDD.n3928 7.39606
R21767 VDD.n3940 VDD.n3939 7.39606
R21768 VDD.n3924 VDD.n3912 7.39606
R21769 VDD.n3924 VDD.n3923 7.39606
R21770 VDD.n3872 VDD.n3870 7.39606
R21771 VDD.n3873 VDD.n3872 7.39606
R21772 VDD.n3998 VDD.n3845 7.39606
R21773 VDD.n3998 VDD.n3997 7.39606
R21774 VDD.n4003 VDD.n3842 7.39606
R21775 VDD.n4004 VDD.n4003 7.39606
R21776 VDD.n4270 VDD.n4066 7.39606
R21777 VDD.n4270 VDD.n4067 7.39606
R21778 VDD.n4279 VDD.n4045 7.39606
R21779 VDD.n4279 VDD.n4047 7.39606
R21780 VDD.n4165 VDD.n4153 7.39606
R21781 VDD.n4165 VDD.n4164 7.39606
R21782 VDD.n4241 VDD.n4150 7.39606
R21783 VDD.n4242 VDD.n4241 7.39606
R21784 VDD.n4238 VDD.n4226 7.39606
R21785 VDD.n4238 VDD.n4237 7.39606
R21786 VDD.n4222 VDD.n4210 7.39606
R21787 VDD.n4222 VDD.n4221 7.39606
R21788 VDD.n4199 VDD.n4187 7.39606
R21789 VDD.n4199 VDD.n4198 7.39606
R21790 VDD.n4183 VDD.n4171 7.39606
R21791 VDD.n4183 VDD.n4182 7.39606
R21792 VDD.n4131 VDD.n4129 7.39606
R21793 VDD.n4132 VDD.n4131 7.39606
R21794 VDD.n4257 VDD.n4104 7.39606
R21795 VDD.n4257 VDD.n4256 7.39606
R21796 VDD.n4262 VDD.n4101 7.39606
R21797 VDD.n4263 VDD.n4262 7.39606
R21798 VDD.n4529 VDD.n4325 7.39606
R21799 VDD.n4529 VDD.n4326 7.39606
R21800 VDD.n4538 VDD.n4304 7.39606
R21801 VDD.n4538 VDD.n4306 7.39606
R21802 VDD.n4424 VDD.n4412 7.39606
R21803 VDD.n4424 VDD.n4423 7.39606
R21804 VDD.n4500 VDD.n4409 7.39606
R21805 VDD.n4501 VDD.n4500 7.39606
R21806 VDD.n4497 VDD.n4485 7.39606
R21807 VDD.n4497 VDD.n4496 7.39606
R21808 VDD.n4481 VDD.n4469 7.39606
R21809 VDD.n4481 VDD.n4480 7.39606
R21810 VDD.n4458 VDD.n4446 7.39606
R21811 VDD.n4458 VDD.n4457 7.39606
R21812 VDD.n4442 VDD.n4430 7.39606
R21813 VDD.n4442 VDD.n4441 7.39606
R21814 VDD.n4390 VDD.n4388 7.39606
R21815 VDD.n4391 VDD.n4390 7.39606
R21816 VDD.n4516 VDD.n4363 7.39606
R21817 VDD.n4516 VDD.n4515 7.39606
R21818 VDD.n4521 VDD.n4360 7.39606
R21819 VDD.n4522 VDD.n4521 7.39606
R21820 VDD.n7093 VDD.n5044 7.39606
R21821 VDD.n7094 VDD.n7093 7.39606
R21822 VDD.n7083 VDD.n5055 7.39606
R21823 VDD.n7084 VDD.n7083 7.39606
R21824 VDD.n7073 VDD.n5065 7.39606
R21825 VDD.n7074 VDD.n7073 7.39606
R21826 VDD.n7063 VDD.n5078 7.39606
R21827 VDD.n7064 VDD.n7063 7.39606
R21828 VDD.n7053 VDD.n5089 7.39606
R21829 VDD.n7054 VDD.n7053 7.39606
R21830 VDD.n7043 VDD.n5099 7.39606
R21831 VDD.n7044 VDD.n7043 7.39606
R21832 VDD.n7026 VDD.n5115 7.39606
R21833 VDD.n7027 VDD.n7026 7.39606
R21834 VDD.n7016 VDD.n5127 7.39606
R21835 VDD.n7017 VDD.n7016 7.39606
R21836 VDD.n7006 VDD.n5140 7.39606
R21837 VDD.n7007 VDD.n7006 7.39606
R21838 VDD.n6996 VDD.n5151 7.39606
R21839 VDD.n6997 VDD.n6996 7.39606
R21840 VDD.n6986 VDD.n5161 7.39606
R21841 VDD.n6987 VDD.n6986 7.39606
R21842 VDD.n6972 VDD.n5174 7.39606
R21843 VDD.n6972 VDD.n5176 7.39606
R21844 VDD.n6952 VDD.n5184 7.39606
R21845 VDD.n6953 VDD.n6952 7.39606
R21846 VDD.n6942 VDD.n5193 7.39606
R21847 VDD.n6943 VDD.n6942 7.39606
R21848 VDD.n6932 VDD.n5206 7.39606
R21849 VDD.n6933 VDD.n6932 7.39606
R21850 VDD.n6922 VDD.n5217 7.39606
R21851 VDD.n6923 VDD.n6922 7.39606
R21852 VDD.n6912 VDD.n5227 7.39606
R21853 VDD.n6913 VDD.n6912 7.39606
R21854 VDD.n6895 VDD.n5243 7.39606
R21855 VDD.n6896 VDD.n6895 7.39606
R21856 VDD.n6885 VDD.n5255 7.39606
R21857 VDD.n6886 VDD.n6885 7.39606
R21858 VDD.n6875 VDD.n5268 7.39606
R21859 VDD.n6876 VDD.n6875 7.39606
R21860 VDD.n6865 VDD.n5279 7.39606
R21861 VDD.n6866 VDD.n6865 7.39606
R21862 VDD.n6855 VDD.n5289 7.39606
R21863 VDD.n6856 VDD.n6855 7.39606
R21864 VDD.n6841 VDD.n5302 7.39606
R21865 VDD.n6841 VDD.n5304 7.39606
R21866 VDD.n6821 VDD.n5312 7.39606
R21867 VDD.n6822 VDD.n6821 7.39606
R21868 VDD.n6811 VDD.n5321 7.39606
R21869 VDD.n6812 VDD.n6811 7.39606
R21870 VDD.n6801 VDD.n5334 7.39606
R21871 VDD.n6802 VDD.n6801 7.39606
R21872 VDD.n6791 VDD.n5345 7.39606
R21873 VDD.n6792 VDD.n6791 7.39606
R21874 VDD.n6781 VDD.n5355 7.39606
R21875 VDD.n6782 VDD.n6781 7.39606
R21876 VDD.n6764 VDD.n5371 7.39606
R21877 VDD.n6765 VDD.n6764 7.39606
R21878 VDD.n6754 VDD.n5383 7.39606
R21879 VDD.n6755 VDD.n6754 7.39606
R21880 VDD.n6744 VDD.n5396 7.39606
R21881 VDD.n6745 VDD.n6744 7.39606
R21882 VDD.n6734 VDD.n5407 7.39606
R21883 VDD.n6735 VDD.n6734 7.39606
R21884 VDD.n6724 VDD.n5417 7.39606
R21885 VDD.n6725 VDD.n6724 7.39606
R21886 VDD.n6710 VDD.n5430 7.39606
R21887 VDD.n6710 VDD.n5432 7.39606
R21888 VDD.n6690 VDD.n5440 7.39606
R21889 VDD.n6691 VDD.n6690 7.39606
R21890 VDD.n6680 VDD.n5449 7.39606
R21891 VDD.n6681 VDD.n6680 7.39606
R21892 VDD.n6670 VDD.n5462 7.39606
R21893 VDD.n6671 VDD.n6670 7.39606
R21894 VDD.n6660 VDD.n5473 7.39606
R21895 VDD.n6661 VDD.n6660 7.39606
R21896 VDD.n6650 VDD.n5483 7.39606
R21897 VDD.n6651 VDD.n6650 7.39606
R21898 VDD.n6633 VDD.n5499 7.39606
R21899 VDD.n6634 VDD.n6633 7.39606
R21900 VDD.n6623 VDD.n5511 7.39606
R21901 VDD.n6624 VDD.n6623 7.39606
R21902 VDD.n6613 VDD.n5524 7.39606
R21903 VDD.n6614 VDD.n6613 7.39606
R21904 VDD.n6603 VDD.n5535 7.39606
R21905 VDD.n6604 VDD.n6603 7.39606
R21906 VDD.n6593 VDD.n5545 7.39606
R21907 VDD.n6594 VDD.n6593 7.39606
R21908 VDD.n6579 VDD.n5558 7.39606
R21909 VDD.n6579 VDD.n5560 7.39606
R21910 VDD.n6559 VDD.n5568 7.39606
R21911 VDD.n6560 VDD.n6559 7.39606
R21912 VDD.n6549 VDD.n5577 7.39606
R21913 VDD.n6550 VDD.n6549 7.39606
R21914 VDD.n6539 VDD.n5590 7.39606
R21915 VDD.n6540 VDD.n6539 7.39606
R21916 VDD.n6529 VDD.n5601 7.39606
R21917 VDD.n6530 VDD.n6529 7.39606
R21918 VDD.n6519 VDD.n5611 7.39606
R21919 VDD.n6520 VDD.n6519 7.39606
R21920 VDD.n6502 VDD.n5627 7.39606
R21921 VDD.n6503 VDD.n6502 7.39606
R21922 VDD.n6492 VDD.n5639 7.39606
R21923 VDD.n6493 VDD.n6492 7.39606
R21924 VDD.n6482 VDD.n5652 7.39606
R21925 VDD.n6483 VDD.n6482 7.39606
R21926 VDD.n6472 VDD.n5663 7.39606
R21927 VDD.n6473 VDD.n6472 7.39606
R21928 VDD.n6462 VDD.n5673 7.39606
R21929 VDD.n6463 VDD.n6462 7.39606
R21930 VDD.n6448 VDD.n5686 7.39606
R21931 VDD.n6448 VDD.n5688 7.39606
R21932 VDD.n6428 VDD.n5696 7.39606
R21933 VDD.n6429 VDD.n6428 7.39606
R21934 VDD.n6418 VDD.n5705 7.39606
R21935 VDD.n6419 VDD.n6418 7.39606
R21936 VDD.n6408 VDD.n5718 7.39606
R21937 VDD.n6409 VDD.n6408 7.39606
R21938 VDD.n6398 VDD.n5729 7.39606
R21939 VDD.n6399 VDD.n6398 7.39606
R21940 VDD.n6388 VDD.n5739 7.39606
R21941 VDD.n6389 VDD.n6388 7.39606
R21942 VDD.n6371 VDD.n5755 7.39606
R21943 VDD.n6372 VDD.n6371 7.39606
R21944 VDD.n6361 VDD.n5767 7.39606
R21945 VDD.n6362 VDD.n6361 7.39606
R21946 VDD.n6351 VDD.n5780 7.39606
R21947 VDD.n6352 VDD.n6351 7.39606
R21948 VDD.n6341 VDD.n5791 7.39606
R21949 VDD.n6342 VDD.n6341 7.39606
R21950 VDD.n6331 VDD.n5801 7.39606
R21951 VDD.n6332 VDD.n6331 7.39606
R21952 VDD.n6317 VDD.n5814 7.39606
R21953 VDD.n6317 VDD.n5816 7.39606
R21954 VDD.n6297 VDD.n5824 7.39606
R21955 VDD.n6298 VDD.n6297 7.39606
R21956 VDD.n6287 VDD.n5833 7.39606
R21957 VDD.n6288 VDD.n6287 7.39606
R21958 VDD.n6277 VDD.n5846 7.39606
R21959 VDD.n6278 VDD.n6277 7.39606
R21960 VDD.n6267 VDD.n5857 7.39606
R21961 VDD.n6268 VDD.n6267 7.39606
R21962 VDD.n6257 VDD.n5867 7.39606
R21963 VDD.n6258 VDD.n6257 7.39606
R21964 VDD.n6240 VDD.n5883 7.39606
R21965 VDD.n6241 VDD.n6240 7.39606
R21966 VDD.n6230 VDD.n5895 7.39606
R21967 VDD.n6231 VDD.n6230 7.39606
R21968 VDD.n6220 VDD.n5908 7.39606
R21969 VDD.n6221 VDD.n6220 7.39606
R21970 VDD.n6210 VDD.n5919 7.39606
R21971 VDD.n6211 VDD.n6210 7.39606
R21972 VDD.n6200 VDD.n5929 7.39606
R21973 VDD.n6201 VDD.n6200 7.39606
R21974 VDD.n6186 VDD.n5942 7.39606
R21975 VDD.n6186 VDD.n5944 7.39606
R21976 VDD.n6166 VDD.n5952 7.39606
R21977 VDD.n6167 VDD.n6166 7.39606
R21978 VDD.n6156 VDD.n5961 7.39606
R21979 VDD.n6157 VDD.n6156 7.39606
R21980 VDD.n6146 VDD.n5974 7.39606
R21981 VDD.n6147 VDD.n6146 7.39606
R21982 VDD.n6136 VDD.n5985 7.39606
R21983 VDD.n6137 VDD.n6136 7.39606
R21984 VDD.n6126 VDD.n5995 7.39606
R21985 VDD.n6127 VDD.n6126 7.39606
R21986 VDD.n6109 VDD.n6011 7.39606
R21987 VDD.n6110 VDD.n6109 7.39606
R21988 VDD.n6099 VDD.n6023 7.39606
R21989 VDD.n6100 VDD.n6099 7.39606
R21990 VDD.n6089 VDD.n6036 7.39606
R21991 VDD.n6090 VDD.n6089 7.39606
R21992 VDD.n6079 VDD.n6047 7.39606
R21993 VDD.n6080 VDD.n6079 7.39606
R21994 VDD.n6069 VDD.n6057 7.39606
R21995 VDD.n6070 VDD.n6069 7.39606
R21996 VDD.t796 VDD.n5030 7.31106
R21997 VDD.n5013 VDD.t332 7.31106
R21998 VDD.t269 VDD.n5005 7.31106
R21999 VDD.n4995 VDD.t468 7.31106
R22000 VDD.t583 VDD.n4989 7.31106
R22001 VDD.n4972 VDD.t585 7.31106
R22002 VDD.t703 VDD.n4964 7.31106
R22003 VDD.n4954 VDD.t888 7.31106
R22004 VDD.t598 VDD.n4948 7.31106
R22005 VDD.n4931 VDD.t549 7.31106
R22006 VDD.t732 VDD.n4923 7.31106
R22007 VDD.n4913 VDD.t31 7.31106
R22008 VDD.t891 VDD.n4907 7.31106
R22009 VDD.n4890 VDD.t526 7.31106
R22010 VDD.t454 VDD.n4882 7.31106
R22011 VDD.n4872 VDD.t59 7.31106
R22012 VDD.t594 VDD.n4866 7.31106
R22013 VDD.n4849 VDD.t596 7.31106
R22014 VDD.t368 VDD.n4841 7.31106
R22015 VDD.n4831 VDD.t553 7.31106
R22016 VDD.t296 VDD.n4825 7.31106
R22017 VDD.n4808 VDD.t645 7.31106
R22018 VDD.t794 VDD.n4800 7.31106
R22019 VDD.n4790 VDD.t87 7.31106
R22020 VDD.t422 VDD.n4784 7.31106
R22021 VDD.n4767 VDD.t725 7.31106
R22022 VDD.t878 VDD.n4759 7.31106
R22023 VDD.n4749 VDD.t747 7.31106
R22024 VDD.t842 VDD.n4743 7.31106
R22025 VDD.n4726 VDD.t869 7.31106
R22026 VDD.t571 VDD.n4718 7.31106
R22027 VDD.n4708 VDD.t340 7.31106
R22028 VDD.n7109 VDD.t915 7.31106
R22029 VDD.t773 VDD.n140 7.31106
R22030 VDD.n7130 VDD.t880 7.31106
R22031 VDD.t903 VDD.n121 7.31106
R22032 VDD.n7151 VDD.t544 7.31106
R22033 VDD.t855 VDD.n102 7.31106
R22034 VDD.n7172 VDD.t96 7.31106
R22035 VDD.t298 VDD.n83 7.31106
R22036 VDD.n7193 VDD.t402 7.31106
R22037 VDD.t714 VDD.n64 7.31106
R22038 VDD.n7214 VDD.t630 7.31106
R22039 VDD.t383 VDD.n45 7.31106
R22040 VDD.n7235 VDD.t301 7.31106
R22041 VDD.t895 VDD.n26 7.31106
R22042 VDD.n7256 VDD.t314 7.31106
R22043 VDD.t509 VDD.n7 7.31106
R22044 VDD.n3779 VDD 6.46848
R22045 VDD.n7329 VDD.n7313 6.37981
R22046 VDD.n7316 VDD.n7313 6.37981
R22047 VDD VDD.n7253 6.37007
R22048 VDD VDD.n7232 6.37007
R22049 VDD VDD.n7211 6.37007
R22050 VDD VDD.n7190 6.37007
R22051 VDD VDD.n7169 6.37007
R22052 VDD VDD.n7148 6.37007
R22053 VDD VDD.n7127 6.37007
R22054 VDD.n156 VDD 5.14622
R22055 VDD.n4037 VDD 5.07436
R22056 VDD.n399 VDD 4.82115
R22057 VDD.n296 VDD 4.82115
R22058 VDD.n293 VDD 4.82115
R22059 VDD.n647 VDD 4.82115
R22060 VDD.n544 VDD 4.82115
R22061 VDD.n541 VDD 4.82115
R22062 VDD.n906 VDD 4.82115
R22063 VDD.n803 VDD 4.82115
R22064 VDD.n800 VDD 4.82115
R22065 VDD.n1165 VDD 4.82115
R22066 VDD.n1062 VDD 4.82115
R22067 VDD.n1059 VDD 4.82115
R22068 VDD.n1424 VDD 4.82115
R22069 VDD.n1321 VDD 4.82115
R22070 VDD.n1318 VDD 4.82115
R22071 VDD.n1683 VDD 4.82115
R22072 VDD.n1580 VDD 4.82115
R22073 VDD.n1577 VDD 4.82115
R22074 VDD.n1942 VDD 4.82115
R22075 VDD.n1839 VDD 4.82115
R22076 VDD.n1836 VDD 4.82115
R22077 VDD.n2201 VDD 4.82115
R22078 VDD.n2098 VDD 4.82115
R22079 VDD.n2095 VDD 4.82115
R22080 VDD.n2460 VDD 4.82115
R22081 VDD.n2357 VDD 4.82115
R22082 VDD.n2354 VDD 4.82115
R22083 VDD.n2719 VDD 4.82115
R22084 VDD.n2616 VDD 4.82115
R22085 VDD.n2613 VDD 4.82115
R22086 VDD.n2978 VDD 4.82115
R22087 VDD.n2875 VDD 4.82115
R22088 VDD.n2872 VDD 4.82115
R22089 VDD.n3237 VDD 4.82115
R22090 VDD.n3134 VDD 4.82115
R22091 VDD.n3131 VDD 4.82115
R22092 VDD.n3496 VDD 4.82115
R22093 VDD.n3393 VDD 4.82115
R22094 VDD.n3390 VDD 4.82115
R22095 VDD.n3755 VDD 4.82115
R22096 VDD.n3652 VDD 4.82115
R22097 VDD.n3649 VDD 4.82115
R22098 VDD.n4014 VDD 4.82115
R22099 VDD.n3911 VDD 4.82115
R22100 VDD.n3908 VDD 4.82115
R22101 VDD.n4273 VDD 4.82115
R22102 VDD.n4170 VDD 4.82115
R22103 VDD.n4167 VDD 4.82115
R22104 VDD.n4532 VDD 4.82115
R22105 VDD.n4429 VDD 4.82115
R22106 VDD.n4426 VDD 4.82115
R22107 VDD.n155 VDD 4.63142
R22108 VDD.n165 VDD.n164 4.5005
R22109 VDD.n668 VDD.n667 4.5005
R22110 VDD.n927 VDD.n926 4.5005
R22111 VDD.n1186 VDD.n1185 4.5005
R22112 VDD.n1445 VDD.n1444 4.5005
R22113 VDD.n1704 VDD.n1703 4.5005
R22114 VDD.n1963 VDD.n1962 4.5005
R22115 VDD.n2222 VDD.n2221 4.5005
R22116 VDD.n2481 VDD.n2480 4.5005
R22117 VDD.n2740 VDD.n2739 4.5005
R22118 VDD.n2999 VDD.n2998 4.5005
R22119 VDD.n3258 VDD.n3257 4.5005
R22120 VDD.n3517 VDD.n3516 4.5005
R22121 VDD.n3776 VDD.n3775 4.5005
R22122 VDD.n4035 VDD.n4034 4.5005
R22123 VDD.n4294 VDD.n4293 4.5005
R22124 VDD.n4553 VDD.n4552 4.5005
R22125 VDD.n7100 VDD.t755 4.27344
R22126 VDD.n7288 VDD.t883 4.14288
R22127 VDD.n415 VDD.n414 4.12965
R22128 VDD.n169 VDD 3.97061
R22129 VDD.n413 VDD 3.7212
R22130 VDD.n4038 VDD 3.67668
R22131 VDD.n417 VDD 3.56572
R22132 VDD.n676 VDD 3.56572
R22133 VDD.n935 VDD 3.56572
R22134 VDD.n1194 VDD 3.56572
R22135 VDD.n1453 VDD 3.56572
R22136 VDD.n1712 VDD 3.56572
R22137 VDD.n1971 VDD 3.56572
R22138 VDD.n2230 VDD 3.56572
R22139 VDD.n2489 VDD 3.56572
R22140 VDD.n2748 VDD 3.56572
R22141 VDD.n3007 VDD 3.56572
R22142 VDD.n3266 VDD 3.56572
R22143 VDD.n3525 VDD 3.56572
R22144 VDD.n3784 VDD 3.56572
R22145 VDD.n4043 VDD 3.56572
R22146 VDD.n4302 VDD 3.56572
R22147 VDD.n7310 VDD.n7277 3.29941
R22148 VDD.n4707 VDD.n4700 3.15974
R22149 VDD.n6069 VDD.n6068 3.15974
R22150 VDD.n7315 VDD.n7314 3.08383
R22151 VDD.n7325 VDD.n7315 3.08383
R22152 VDD.n7106 VDD.n5034 2.85027
R22153 VDD.n155 VDD.n154 2.80327
R22154 VDD.n407 VDD 2.72902
R22155 VDD.n7331 VDD.t728 2.59419
R22156 VDD.n4296 VDD 2.53636
R22157 VDD.n655 VDD 2.438
R22158 VDD.n914 VDD 2.438
R22159 VDD.n1173 VDD 2.438
R22160 VDD.n1432 VDD 2.438
R22161 VDD.n1691 VDD 2.438
R22162 VDD.n1950 VDD 2.438
R22163 VDD.n2209 VDD 2.438
R22164 VDD.n2468 VDD 2.438
R22165 VDD.n2727 VDD 2.438
R22166 VDD.n2986 VDD 2.438
R22167 VDD.n3245 VDD 2.438
R22168 VDD.n3504 VDD 2.438
R22169 VDD.n3763 VDD 2.438
R22170 VDD.n4022 VDD 2.438
R22171 VDD.n4281 VDD 2.438
R22172 VDD.n4540 VDD 2.438
R22173 VDD.n7311 VDD 2.38637
R22174 VDD.n401 VDD.n400 2.3255
R22175 VDD.n397 VDD.n396 2.3255
R22176 VDD.n388 VDD.n387 2.3255
R22177 VDD.n384 VDD.n383 2.3255
R22178 VDD.n257 VDD.n229 2.3255
R22179 VDD.n310 VDD.n309 2.3255
R22180 VDD.n326 VDD.n325 2.3255
R22181 VDD.n333 VDD.n332 2.3255
R22182 VDD.n349 VDD.n348 2.3255
R22183 VDD.n365 VDD.n364 2.3255
R22184 VDD.n367 VDD.n366 2.3255
R22185 VDD.n292 VDD.n291 2.3255
R22186 VDD.n406 VDD.n405 2.3255
R22187 VDD.n649 VDD.n648 2.3255
R22188 VDD.n645 VDD.n644 2.3255
R22189 VDD.n636 VDD.n635 2.3255
R22190 VDD.n632 VDD.n631 2.3255
R22191 VDD.n505 VDD.n477 2.3255
R22192 VDD.n558 VDD.n557 2.3255
R22193 VDD.n574 VDD.n573 2.3255
R22194 VDD.n581 VDD.n580 2.3255
R22195 VDD.n597 VDD.n596 2.3255
R22196 VDD.n613 VDD.n612 2.3255
R22197 VDD.n615 VDD.n614 2.3255
R22198 VDD.n540 VDD.n539 2.3255
R22199 VDD.n654 VDD.n653 2.3255
R22200 VDD.n908 VDD.n907 2.3255
R22201 VDD.n904 VDD.n903 2.3255
R22202 VDD.n895 VDD.n894 2.3255
R22203 VDD.n891 VDD.n890 2.3255
R22204 VDD.n764 VDD.n736 2.3255
R22205 VDD.n817 VDD.n816 2.3255
R22206 VDD.n833 VDD.n832 2.3255
R22207 VDD.n840 VDD.n839 2.3255
R22208 VDD.n856 VDD.n855 2.3255
R22209 VDD.n872 VDD.n871 2.3255
R22210 VDD.n874 VDD.n873 2.3255
R22211 VDD.n799 VDD.n798 2.3255
R22212 VDD.n913 VDD.n912 2.3255
R22213 VDD.n1167 VDD.n1166 2.3255
R22214 VDD.n1163 VDD.n1162 2.3255
R22215 VDD.n1154 VDD.n1153 2.3255
R22216 VDD.n1150 VDD.n1149 2.3255
R22217 VDD.n1023 VDD.n995 2.3255
R22218 VDD.n1076 VDD.n1075 2.3255
R22219 VDD.n1092 VDD.n1091 2.3255
R22220 VDD.n1099 VDD.n1098 2.3255
R22221 VDD.n1115 VDD.n1114 2.3255
R22222 VDD.n1131 VDD.n1130 2.3255
R22223 VDD.n1133 VDD.n1132 2.3255
R22224 VDD.n1058 VDD.n1057 2.3255
R22225 VDD.n1172 VDD.n1171 2.3255
R22226 VDD.n1426 VDD.n1425 2.3255
R22227 VDD.n1422 VDD.n1421 2.3255
R22228 VDD.n1413 VDD.n1412 2.3255
R22229 VDD.n1409 VDD.n1408 2.3255
R22230 VDD.n1282 VDD.n1254 2.3255
R22231 VDD.n1335 VDD.n1334 2.3255
R22232 VDD.n1351 VDD.n1350 2.3255
R22233 VDD.n1358 VDD.n1357 2.3255
R22234 VDD.n1374 VDD.n1373 2.3255
R22235 VDD.n1390 VDD.n1389 2.3255
R22236 VDD.n1392 VDD.n1391 2.3255
R22237 VDD.n1317 VDD.n1316 2.3255
R22238 VDD.n1431 VDD.n1430 2.3255
R22239 VDD.n1685 VDD.n1684 2.3255
R22240 VDD.n1681 VDD.n1680 2.3255
R22241 VDD.n1672 VDD.n1671 2.3255
R22242 VDD.n1668 VDD.n1667 2.3255
R22243 VDD.n1541 VDD.n1513 2.3255
R22244 VDD.n1594 VDD.n1593 2.3255
R22245 VDD.n1610 VDD.n1609 2.3255
R22246 VDD.n1617 VDD.n1616 2.3255
R22247 VDD.n1633 VDD.n1632 2.3255
R22248 VDD.n1649 VDD.n1648 2.3255
R22249 VDD.n1651 VDD.n1650 2.3255
R22250 VDD.n1576 VDD.n1575 2.3255
R22251 VDD.n1690 VDD.n1689 2.3255
R22252 VDD.n1944 VDD.n1943 2.3255
R22253 VDD.n1940 VDD.n1939 2.3255
R22254 VDD.n1931 VDD.n1930 2.3255
R22255 VDD.n1927 VDD.n1926 2.3255
R22256 VDD.n1800 VDD.n1772 2.3255
R22257 VDD.n1853 VDD.n1852 2.3255
R22258 VDD.n1869 VDD.n1868 2.3255
R22259 VDD.n1876 VDD.n1875 2.3255
R22260 VDD.n1892 VDD.n1891 2.3255
R22261 VDD.n1908 VDD.n1907 2.3255
R22262 VDD.n1910 VDD.n1909 2.3255
R22263 VDD.n1835 VDD.n1834 2.3255
R22264 VDD.n1949 VDD.n1948 2.3255
R22265 VDD.n2203 VDD.n2202 2.3255
R22266 VDD.n2199 VDD.n2198 2.3255
R22267 VDD.n2190 VDD.n2189 2.3255
R22268 VDD.n2186 VDD.n2185 2.3255
R22269 VDD.n2059 VDD.n2031 2.3255
R22270 VDD.n2112 VDD.n2111 2.3255
R22271 VDD.n2128 VDD.n2127 2.3255
R22272 VDD.n2135 VDD.n2134 2.3255
R22273 VDD.n2151 VDD.n2150 2.3255
R22274 VDD.n2167 VDD.n2166 2.3255
R22275 VDD.n2169 VDD.n2168 2.3255
R22276 VDD.n2094 VDD.n2093 2.3255
R22277 VDD.n2208 VDD.n2207 2.3255
R22278 VDD.n2462 VDD.n2461 2.3255
R22279 VDD.n2458 VDD.n2457 2.3255
R22280 VDD.n2449 VDD.n2448 2.3255
R22281 VDD.n2445 VDD.n2444 2.3255
R22282 VDD.n2318 VDD.n2290 2.3255
R22283 VDD.n2371 VDD.n2370 2.3255
R22284 VDD.n2387 VDD.n2386 2.3255
R22285 VDD.n2394 VDD.n2393 2.3255
R22286 VDD.n2410 VDD.n2409 2.3255
R22287 VDD.n2426 VDD.n2425 2.3255
R22288 VDD.n2428 VDD.n2427 2.3255
R22289 VDD.n2353 VDD.n2352 2.3255
R22290 VDD.n2467 VDD.n2466 2.3255
R22291 VDD.n2721 VDD.n2720 2.3255
R22292 VDD.n2717 VDD.n2716 2.3255
R22293 VDD.n2708 VDD.n2707 2.3255
R22294 VDD.n2704 VDD.n2703 2.3255
R22295 VDD.n2577 VDD.n2549 2.3255
R22296 VDD.n2630 VDD.n2629 2.3255
R22297 VDD.n2646 VDD.n2645 2.3255
R22298 VDD.n2653 VDD.n2652 2.3255
R22299 VDD.n2669 VDD.n2668 2.3255
R22300 VDD.n2685 VDD.n2684 2.3255
R22301 VDD.n2687 VDD.n2686 2.3255
R22302 VDD.n2612 VDD.n2611 2.3255
R22303 VDD.n2726 VDD.n2725 2.3255
R22304 VDD.n2980 VDD.n2979 2.3255
R22305 VDD.n2976 VDD.n2975 2.3255
R22306 VDD.n2967 VDD.n2966 2.3255
R22307 VDD.n2963 VDD.n2962 2.3255
R22308 VDD.n2836 VDD.n2808 2.3255
R22309 VDD.n2889 VDD.n2888 2.3255
R22310 VDD.n2905 VDD.n2904 2.3255
R22311 VDD.n2912 VDD.n2911 2.3255
R22312 VDD.n2928 VDD.n2927 2.3255
R22313 VDD.n2944 VDD.n2943 2.3255
R22314 VDD.n2946 VDD.n2945 2.3255
R22315 VDD.n2871 VDD.n2870 2.3255
R22316 VDD.n2985 VDD.n2984 2.3255
R22317 VDD.n3239 VDD.n3238 2.3255
R22318 VDD.n3235 VDD.n3234 2.3255
R22319 VDD.n3226 VDD.n3225 2.3255
R22320 VDD.n3222 VDD.n3221 2.3255
R22321 VDD.n3095 VDD.n3067 2.3255
R22322 VDD.n3148 VDD.n3147 2.3255
R22323 VDD.n3164 VDD.n3163 2.3255
R22324 VDD.n3171 VDD.n3170 2.3255
R22325 VDD.n3187 VDD.n3186 2.3255
R22326 VDD.n3203 VDD.n3202 2.3255
R22327 VDD.n3205 VDD.n3204 2.3255
R22328 VDD.n3130 VDD.n3129 2.3255
R22329 VDD.n3244 VDD.n3243 2.3255
R22330 VDD.n3498 VDD.n3497 2.3255
R22331 VDD.n3494 VDD.n3493 2.3255
R22332 VDD.n3485 VDD.n3484 2.3255
R22333 VDD.n3481 VDD.n3480 2.3255
R22334 VDD.n3354 VDD.n3326 2.3255
R22335 VDD.n3407 VDD.n3406 2.3255
R22336 VDD.n3423 VDD.n3422 2.3255
R22337 VDD.n3430 VDD.n3429 2.3255
R22338 VDD.n3446 VDD.n3445 2.3255
R22339 VDD.n3462 VDD.n3461 2.3255
R22340 VDD.n3464 VDD.n3463 2.3255
R22341 VDD.n3389 VDD.n3388 2.3255
R22342 VDD.n3503 VDD.n3502 2.3255
R22343 VDD.n3757 VDD.n3756 2.3255
R22344 VDD.n3753 VDD.n3752 2.3255
R22345 VDD.n3744 VDD.n3743 2.3255
R22346 VDD.n3740 VDD.n3739 2.3255
R22347 VDD.n3613 VDD.n3585 2.3255
R22348 VDD.n3666 VDD.n3665 2.3255
R22349 VDD.n3682 VDD.n3681 2.3255
R22350 VDD.n3689 VDD.n3688 2.3255
R22351 VDD.n3705 VDD.n3704 2.3255
R22352 VDD.n3721 VDD.n3720 2.3255
R22353 VDD.n3723 VDD.n3722 2.3255
R22354 VDD.n3648 VDD.n3647 2.3255
R22355 VDD.n3762 VDD.n3761 2.3255
R22356 VDD.n4016 VDD.n4015 2.3255
R22357 VDD.n4012 VDD.n4011 2.3255
R22358 VDD.n4003 VDD.n4002 2.3255
R22359 VDD.n3999 VDD.n3998 2.3255
R22360 VDD.n3872 VDD.n3844 2.3255
R22361 VDD.n3925 VDD.n3924 2.3255
R22362 VDD.n3941 VDD.n3940 2.3255
R22363 VDD.n3948 VDD.n3947 2.3255
R22364 VDD.n3964 VDD.n3963 2.3255
R22365 VDD.n3980 VDD.n3979 2.3255
R22366 VDD.n3982 VDD.n3981 2.3255
R22367 VDD.n3907 VDD.n3906 2.3255
R22368 VDD.n4021 VDD.n4020 2.3255
R22369 VDD.n4275 VDD.n4274 2.3255
R22370 VDD.n4271 VDD.n4270 2.3255
R22371 VDD.n4262 VDD.n4261 2.3255
R22372 VDD.n4258 VDD.n4257 2.3255
R22373 VDD.n4131 VDD.n4103 2.3255
R22374 VDD.n4184 VDD.n4183 2.3255
R22375 VDD.n4200 VDD.n4199 2.3255
R22376 VDD.n4207 VDD.n4206 2.3255
R22377 VDD.n4223 VDD.n4222 2.3255
R22378 VDD.n4239 VDD.n4238 2.3255
R22379 VDD.n4241 VDD.n4240 2.3255
R22380 VDD.n4166 VDD.n4165 2.3255
R22381 VDD.n4280 VDD.n4279 2.3255
R22382 VDD.n4534 VDD.n4533 2.3255
R22383 VDD.n4530 VDD.n4529 2.3255
R22384 VDD.n4521 VDD.n4520 2.3255
R22385 VDD.n4517 VDD.n4516 2.3255
R22386 VDD.n4390 VDD.n4362 2.3255
R22387 VDD.n4443 VDD.n4442 2.3255
R22388 VDD.n4459 VDD.n4458 2.3255
R22389 VDD.n4466 VDD.n4465 2.3255
R22390 VDD.n4482 VDD.n4481 2.3255
R22391 VDD.n4498 VDD.n4497 2.3255
R22392 VDD.n4500 VDD.n4499 2.3255
R22393 VDD.n4425 VDD.n4424 2.3255
R22394 VDD.n4539 VDD.n4538 2.3255
R22395 VDD.n4721 VDD.n4720 2.3255
R22396 VDD.n4725 VDD.n4724 2.3255
R22397 VDD.n4722 VDD.n4696 2.3255
R22398 VDD.n4746 VDD.n4745 2.3255
R22399 VDD.n4748 VDD.n4747 2.3255
R22400 VDD.n4762 VDD.n4761 2.3255
R22401 VDD.n4766 VDD.n4765 2.3255
R22402 VDD.n4763 VDD.n4677 2.3255
R22403 VDD.n4787 VDD.n4786 2.3255
R22404 VDD.n4789 VDD.n4788 2.3255
R22405 VDD.n4803 VDD.n4802 2.3255
R22406 VDD.n4807 VDD.n4806 2.3255
R22407 VDD.n4804 VDD.n4658 2.3255
R22408 VDD.n4828 VDD.n4827 2.3255
R22409 VDD.n4830 VDD.n4829 2.3255
R22410 VDD.n4844 VDD.n4843 2.3255
R22411 VDD.n4848 VDD.n4847 2.3255
R22412 VDD.n4845 VDD.n4639 2.3255
R22413 VDD.n4869 VDD.n4868 2.3255
R22414 VDD.n4871 VDD.n4870 2.3255
R22415 VDD.n4885 VDD.n4884 2.3255
R22416 VDD.n4889 VDD.n4888 2.3255
R22417 VDD.n4886 VDD.n4620 2.3255
R22418 VDD.n4910 VDD.n4909 2.3255
R22419 VDD.n4912 VDD.n4911 2.3255
R22420 VDD.n4926 VDD.n4925 2.3255
R22421 VDD.n4930 VDD.n4929 2.3255
R22422 VDD.n4927 VDD.n4601 2.3255
R22423 VDD.n4951 VDD.n4950 2.3255
R22424 VDD.n4953 VDD.n4952 2.3255
R22425 VDD.n4967 VDD.n4966 2.3255
R22426 VDD.n4971 VDD.n4970 2.3255
R22427 VDD.n4968 VDD.n4582 2.3255
R22428 VDD.n4992 VDD.n4991 2.3255
R22429 VDD.n4994 VDD.n4993 2.3255
R22430 VDD.n5008 VDD.n5007 2.3255
R22431 VDD.n5012 VDD.n5011 2.3255
R22432 VDD.n5009 VDD.n4563 2.3255
R22433 VDD.n5033 VDD.n5032 2.3255
R22434 VDD.n6079 VDD.n6048 2.3255
R22435 VDD.n6089 VDD.n6038 2.3255
R22436 VDD.n6099 VDD.n6027 2.3255
R22437 VDD.n6109 VDD.n6014 2.3255
R22438 VDD.n6013 VDD.n6005 2.3255
R22439 VDD.n6126 VDD.n5999 2.3255
R22440 VDD.n6136 VDD.n5986 2.3255
R22441 VDD.n6146 VDD.n5976 2.3255
R22442 VDD.n6156 VDD.n5965 2.3255
R22443 VDD.n6166 VDD.n5941 2.3255
R22444 VDD.n6187 VDD.n6186 2.3255
R22445 VDD.n6191 VDD.n6190 2.3255
R22446 VDD.n6200 VDD.n5933 2.3255
R22447 VDD.n6210 VDD.n5920 2.3255
R22448 VDD.n6220 VDD.n5910 2.3255
R22449 VDD.n6230 VDD.n5899 2.3255
R22450 VDD.n6240 VDD.n5886 2.3255
R22451 VDD.n5885 VDD.n5877 2.3255
R22452 VDD.n6257 VDD.n5871 2.3255
R22453 VDD.n6267 VDD.n5858 2.3255
R22454 VDD.n6277 VDD.n5848 2.3255
R22455 VDD.n6287 VDD.n5837 2.3255
R22456 VDD.n6297 VDD.n5813 2.3255
R22457 VDD.n6318 VDD.n6317 2.3255
R22458 VDD.n6322 VDD.n6321 2.3255
R22459 VDD.n6331 VDD.n5805 2.3255
R22460 VDD.n6341 VDD.n5792 2.3255
R22461 VDD.n6351 VDD.n5782 2.3255
R22462 VDD.n6361 VDD.n5771 2.3255
R22463 VDD.n6371 VDD.n5758 2.3255
R22464 VDD.n5757 VDD.n5749 2.3255
R22465 VDD.n6388 VDD.n5743 2.3255
R22466 VDD.n6398 VDD.n5730 2.3255
R22467 VDD.n6408 VDD.n5720 2.3255
R22468 VDD.n6418 VDD.n5709 2.3255
R22469 VDD.n6428 VDD.n5685 2.3255
R22470 VDD.n6449 VDD.n6448 2.3255
R22471 VDD.n6453 VDD.n6452 2.3255
R22472 VDD.n6462 VDD.n5677 2.3255
R22473 VDD.n6472 VDD.n5664 2.3255
R22474 VDD.n6482 VDD.n5654 2.3255
R22475 VDD.n6492 VDD.n5643 2.3255
R22476 VDD.n6502 VDD.n5630 2.3255
R22477 VDD.n5629 VDD.n5621 2.3255
R22478 VDD.n6519 VDD.n5615 2.3255
R22479 VDD.n6529 VDD.n5602 2.3255
R22480 VDD.n6539 VDD.n5592 2.3255
R22481 VDD.n6549 VDD.n5581 2.3255
R22482 VDD.n6559 VDD.n5557 2.3255
R22483 VDD.n6580 VDD.n6579 2.3255
R22484 VDD.n6584 VDD.n6583 2.3255
R22485 VDD.n6593 VDD.n5549 2.3255
R22486 VDD.n6603 VDD.n5536 2.3255
R22487 VDD.n6613 VDD.n5526 2.3255
R22488 VDD.n6623 VDD.n5515 2.3255
R22489 VDD.n6633 VDD.n5502 2.3255
R22490 VDD.n5501 VDD.n5493 2.3255
R22491 VDD.n6650 VDD.n5487 2.3255
R22492 VDD.n6660 VDD.n5474 2.3255
R22493 VDD.n6670 VDD.n5464 2.3255
R22494 VDD.n6680 VDD.n5453 2.3255
R22495 VDD.n6690 VDD.n5429 2.3255
R22496 VDD.n6711 VDD.n6710 2.3255
R22497 VDD.n6715 VDD.n6714 2.3255
R22498 VDD.n6724 VDD.n5421 2.3255
R22499 VDD.n6734 VDD.n5408 2.3255
R22500 VDD.n6744 VDD.n5398 2.3255
R22501 VDD.n6754 VDD.n5387 2.3255
R22502 VDD.n6764 VDD.n5374 2.3255
R22503 VDD.n5373 VDD.n5365 2.3255
R22504 VDD.n6781 VDD.n5359 2.3255
R22505 VDD.n6791 VDD.n5346 2.3255
R22506 VDD.n6801 VDD.n5336 2.3255
R22507 VDD.n6811 VDD.n5325 2.3255
R22508 VDD.n6821 VDD.n5301 2.3255
R22509 VDD.n6842 VDD.n6841 2.3255
R22510 VDD.n6846 VDD.n6845 2.3255
R22511 VDD.n6855 VDD.n5293 2.3255
R22512 VDD.n6865 VDD.n5280 2.3255
R22513 VDD.n6875 VDD.n5270 2.3255
R22514 VDD.n6885 VDD.n5259 2.3255
R22515 VDD.n6895 VDD.n5246 2.3255
R22516 VDD.n5245 VDD.n5237 2.3255
R22517 VDD.n6912 VDD.n5231 2.3255
R22518 VDD.n6922 VDD.n5218 2.3255
R22519 VDD.n6932 VDD.n5208 2.3255
R22520 VDD.n6942 VDD.n5197 2.3255
R22521 VDD.n6952 VDD.n5173 2.3255
R22522 VDD.n6973 VDD.n6972 2.3255
R22523 VDD.n6977 VDD.n6976 2.3255
R22524 VDD.n6986 VDD.n5165 2.3255
R22525 VDD.n6996 VDD.n5152 2.3255
R22526 VDD.n7006 VDD.n5142 2.3255
R22527 VDD.n7016 VDD.n5131 2.3255
R22528 VDD.n7026 VDD.n5118 2.3255
R22529 VDD.n5117 VDD.n5109 2.3255
R22530 VDD.n7043 VDD.n5103 2.3255
R22531 VDD.n7053 VDD.n5090 2.3255
R22532 VDD.n7063 VDD.n5080 2.3255
R22533 VDD.n7073 VDD.n5069 2.3255
R22534 VDD.n7083 VDD.n5056 2.3255
R22535 VDD.n7093 VDD.n5046 2.3255
R22536 VDD.n7104 VDD.n7103 2.3255
R22537 VDD.n7274 VDD.n7273 2.3255
R22538 VDD.n13 VDD.n10 2.3255
R22539 VDD.n7255 VDD.n7254 2.3255
R22540 VDD.n7253 VDD.n7252 2.3255
R22541 VDD.n32 VDD.n29 2.3255
R22542 VDD.n7234 VDD.n7233 2.3255
R22543 VDD.n7232 VDD.n7231 2.3255
R22544 VDD.n51 VDD.n48 2.3255
R22545 VDD.n7213 VDD.n7212 2.3255
R22546 VDD.n7211 VDD.n7210 2.3255
R22547 VDD.n70 VDD.n67 2.3255
R22548 VDD.n7192 VDD.n7191 2.3255
R22549 VDD.n7190 VDD.n7189 2.3255
R22550 VDD.n89 VDD.n86 2.3255
R22551 VDD.n7171 VDD.n7170 2.3255
R22552 VDD.n7169 VDD.n7168 2.3255
R22553 VDD.n108 VDD.n105 2.3255
R22554 VDD.n7150 VDD.n7149 2.3255
R22555 VDD.n7148 VDD.n7147 2.3255
R22556 VDD.n127 VDD.n124 2.3255
R22557 VDD.n7129 VDD.n7128 2.3255
R22558 VDD.n7127 VDD.n7126 2.3255
R22559 VDD.n146 VDD.n143 2.3255
R22560 VDD.n7108 VDD.n7107 2.3255
R22561 VDD.n154 VDD 2.29175
R22562 VDD.n7333 VDD.n0 2.23613
R22563 VDD.n7321 VDD.n7320 2.05606
R22564 VDD.n7320 VDD.n7317 2.05606
R22565 VDD.n0 VDD 2.03645
R22566 VDD.n385 VDD 1.90811
R22567 VDD.n312 VDD 1.90811
R22568 VDD.n351 VDD 1.90811
R22569 VDD.n170 VDD 1.90811
R22570 VDD.n633 VDD 1.90811
R22571 VDD.n560 VDD 1.90811
R22572 VDD.n599 VDD 1.90811
R22573 VDD.n418 VDD 1.90811
R22574 VDD.n892 VDD 1.90811
R22575 VDD.n819 VDD 1.90811
R22576 VDD.n858 VDD 1.90811
R22577 VDD.n677 VDD 1.90811
R22578 VDD.n1151 VDD 1.90811
R22579 VDD.n1078 VDD 1.90811
R22580 VDD.n1117 VDD 1.90811
R22581 VDD.n936 VDD 1.90811
R22582 VDD.n1410 VDD 1.90811
R22583 VDD.n1337 VDD 1.90811
R22584 VDD.n1376 VDD 1.90811
R22585 VDD.n1195 VDD 1.90811
R22586 VDD.n1669 VDD 1.90811
R22587 VDD.n1596 VDD 1.90811
R22588 VDD.n1635 VDD 1.90811
R22589 VDD.n1454 VDD 1.90811
R22590 VDD.n1928 VDD 1.90811
R22591 VDD.n1855 VDD 1.90811
R22592 VDD.n1894 VDD 1.90811
R22593 VDD.n1713 VDD 1.90811
R22594 VDD.n2187 VDD 1.90811
R22595 VDD.n2114 VDD 1.90811
R22596 VDD.n2153 VDD 1.90811
R22597 VDD.n1972 VDD 1.90811
R22598 VDD.n2446 VDD 1.90811
R22599 VDD.n2373 VDD 1.90811
R22600 VDD.n2412 VDD 1.90811
R22601 VDD.n2231 VDD 1.90811
R22602 VDD.n2705 VDD 1.90811
R22603 VDD.n2632 VDD 1.90811
R22604 VDD.n2671 VDD 1.90811
R22605 VDD.n2490 VDD 1.90811
R22606 VDD.n2964 VDD 1.90811
R22607 VDD.n2891 VDD 1.90811
R22608 VDD.n2930 VDD 1.90811
R22609 VDD.n2749 VDD 1.90811
R22610 VDD.n3223 VDD 1.90811
R22611 VDD.n3150 VDD 1.90811
R22612 VDD.n3189 VDD 1.90811
R22613 VDD.n3008 VDD 1.90811
R22614 VDD.n3482 VDD 1.90811
R22615 VDD.n3409 VDD 1.90811
R22616 VDD.n3448 VDD 1.90811
R22617 VDD.n3267 VDD 1.90811
R22618 VDD.n3741 VDD 1.90811
R22619 VDD.n3668 VDD 1.90811
R22620 VDD.n3707 VDD 1.90811
R22621 VDD.n3526 VDD 1.90811
R22622 VDD.n4000 VDD 1.90811
R22623 VDD.n3927 VDD 1.90811
R22624 VDD.n3966 VDD 1.90811
R22625 VDD.n3785 VDD 1.90811
R22626 VDD.n4259 VDD 1.90811
R22627 VDD.n4186 VDD 1.90811
R22628 VDD.n4225 VDD 1.90811
R22629 VDD.n4044 VDD 1.90811
R22630 VDD.n4518 VDD 1.90811
R22631 VDD.n4445 VDD 1.90811
R22632 VDD.n4484 VDD 1.90811
R22633 VDD.n4303 VDD 1.90811
R22634 VDD.n4297 VDD.n4296 1.90557
R22635 VDD.n4038 VDD.n4037 1.90557
R22636 VDD.n3779 VDD.n3778 1.90557
R22637 VDD.n3520 VDD.n3519 1.90557
R22638 VDD.n3261 VDD.n3260 1.90557
R22639 VDD.n3002 VDD.n3001 1.90557
R22640 VDD.n2743 VDD.n2742 1.90557
R22641 VDD.n2484 VDD.n2483 1.90557
R22642 VDD.n2225 VDD.n2224 1.90557
R22643 VDD.n1966 VDD.n1965 1.90557
R22644 VDD.n1707 VDD.n1706 1.90557
R22645 VDD.n1448 VDD.n1447 1.90557
R22646 VDD.n1189 VDD.n1188 1.90557
R22647 VDD.n930 VDD.n929 1.90557
R22648 VDD.n671 VDD.n670 1.90557
R22649 VDD.n7311 VDD 1.71534
R22650 VDD.n384 VDD.n229 1.66898
R22651 VDD.n366 VDD.n365 1.66898
R22652 VDD.n632 VDD.n477 1.66898
R22653 VDD.n614 VDD.n613 1.66898
R22654 VDD.n891 VDD.n736 1.66898
R22655 VDD.n873 VDD.n872 1.66898
R22656 VDD.n1150 VDD.n995 1.66898
R22657 VDD.n1132 VDD.n1131 1.66898
R22658 VDD.n1409 VDD.n1254 1.66898
R22659 VDD.n1391 VDD.n1390 1.66898
R22660 VDD.n1668 VDD.n1513 1.66898
R22661 VDD.n1650 VDD.n1649 1.66898
R22662 VDD.n1927 VDD.n1772 1.66898
R22663 VDD.n1909 VDD.n1908 1.66898
R22664 VDD.n2186 VDD.n2031 1.66898
R22665 VDD.n2168 VDD.n2167 1.66898
R22666 VDD.n2445 VDD.n2290 1.66898
R22667 VDD.n2427 VDD.n2426 1.66898
R22668 VDD.n2704 VDD.n2549 1.66898
R22669 VDD.n2686 VDD.n2685 1.66898
R22670 VDD.n2963 VDD.n2808 1.66898
R22671 VDD.n2945 VDD.n2944 1.66898
R22672 VDD.n3222 VDD.n3067 1.66898
R22673 VDD.n3204 VDD.n3203 1.66898
R22674 VDD.n3481 VDD.n3326 1.66898
R22675 VDD.n3463 VDD.n3462 1.66898
R22676 VDD.n3740 VDD.n3585 1.66898
R22677 VDD.n3722 VDD.n3721 1.66898
R22678 VDD.n3999 VDD.n3844 1.66898
R22679 VDD.n3981 VDD.n3980 1.66898
R22680 VDD.n4258 VDD.n4103 1.66898
R22681 VDD.n4240 VDD.n4239 1.66898
R22682 VDD.n4517 VDD.n4362 1.66898
R22683 VDD.n4499 VDD.n4498 1.66898
R22684 VDD.n6048 VDD.n6038 1.66898
R22685 VDD.n5986 VDD.n5976 1.66898
R22686 VDD.n6187 VDD.n5941 1.66898
R22687 VDD.n5920 VDD.n5910 1.66898
R22688 VDD.n5858 VDD.n5848 1.66898
R22689 VDD.n6318 VDD.n5813 1.66898
R22690 VDD.n5792 VDD.n5782 1.66898
R22691 VDD.n5730 VDD.n5720 1.66898
R22692 VDD.n6449 VDD.n5685 1.66898
R22693 VDD.n5664 VDD.n5654 1.66898
R22694 VDD.n5602 VDD.n5592 1.66898
R22695 VDD.n6580 VDD.n5557 1.66898
R22696 VDD.n5536 VDD.n5526 1.66898
R22697 VDD.n5474 VDD.n5464 1.66898
R22698 VDD.n6711 VDD.n5429 1.66898
R22699 VDD.n5408 VDD.n5398 1.66898
R22700 VDD.n5346 VDD.n5336 1.66898
R22701 VDD.n6842 VDD.n5301 1.66898
R22702 VDD.n5280 VDD.n5270 1.66898
R22703 VDD.n5218 VDD.n5208 1.66898
R22704 VDD.n6973 VDD.n5173 1.66898
R22705 VDD.n5152 VDD.n5142 1.66898
R22706 VDD.n5090 VDD.n5080 1.66898
R22707 VDD.n5056 VDD.n5046 1.66898
R22708 VDD.n14 VDD 1.53854
R22709 VDD.n33 VDD 1.53854
R22710 VDD.n52 VDD 1.53854
R22711 VDD.n71 VDD 1.53854
R22712 VDD.n90 VDD 1.53854
R22713 VDD.n109 VDD 1.53854
R22714 VDD.n128 VDD 1.53854
R22715 VDD.n147 VDD 1.53854
R22716 VDD.n191 VDD 1.49898
R22717 VDD.n439 VDD 1.49898
R22718 VDD.n698 VDD 1.49898
R22719 VDD.n957 VDD 1.49898
R22720 VDD.n1216 VDD 1.49898
R22721 VDD.n1475 VDD 1.49898
R22722 VDD.n1734 VDD 1.49898
R22723 VDD.n1993 VDD 1.49898
R22724 VDD.n2252 VDD 1.49898
R22725 VDD.n2511 VDD 1.49898
R22726 VDD.n2770 VDD 1.49898
R22727 VDD.n3029 VDD 1.49898
R22728 VDD.n3288 VDD 1.49898
R22729 VDD.n3547 VDD 1.49898
R22730 VDD.n3806 VDD 1.49898
R22731 VDD.n4065 VDD 1.49898
R22732 VDD.n4324 VDD 1.49898
R22733 VDD.n335 VDD 1.4842
R22734 VDD.n583 VDD 1.4842
R22735 VDD.n842 VDD 1.4842
R22736 VDD.n1101 VDD 1.4842
R22737 VDD.n1360 VDD 1.4842
R22738 VDD.n1619 VDD 1.4842
R22739 VDD.n1878 VDD 1.4842
R22740 VDD.n2137 VDD 1.4842
R22741 VDD.n2396 VDD 1.4842
R22742 VDD.n2655 VDD 1.4842
R22743 VDD.n2914 VDD 1.4842
R22744 VDD.n3173 VDD 1.4842
R22745 VDD.n3432 VDD 1.4842
R22746 VDD.n3691 VDD 1.4842
R22747 VDD.n3950 VDD 1.4842
R22748 VDD.n4209 VDD 1.4842
R22749 VDD.n4468 VDD 1.4842
R22750 VDD VDD.n7310 1.45974
R22751 VDD.n13 VDD.n1 1.26409
R22752 VDD.n32 VDD.n20 1.26409
R22753 VDD.n51 VDD.n39 1.26409
R22754 VDD.n70 VDD.n58 1.26409
R22755 VDD.n89 VDD.n77 1.26409
R22756 VDD.n108 VDD.n96 1.26409
R22757 VDD.n127 VDD.n115 1.26409
R22758 VDD.n146 VDD.n134 1.26409
R22759 VDD.n7296 VDD.n7278 1.22567
R22760 VDD.n7296 VDD.n7283 1.22567
R22761 VDD.n7282 VDD.n7280 1.22567
R22762 VDD.n7295 VDD.n7282 1.22567
R22763 VDD.n7299 VDD.n7298 1.22567
R22764 VDD.n7287 VDD.n7286 1.163
R22765 VDD.n14 VDD.n13 1.1418
R22766 VDD.n33 VDD.n32 1.1418
R22767 VDD.n52 VDD.n51 1.1418
R22768 VDD.n71 VDD.n70 1.1418
R22769 VDD.n90 VDD.n89 1.1418
R22770 VDD.n109 VDD.n108 1.1418
R22771 VDD.n128 VDD.n127 1.1418
R22772 VDD.n147 VDD.n146 1.1418
R22773 VDD.n407 VDD.n406 1.11735
R22774 VDD.n664 VDD 1.09561
R22775 VDD.n660 VDD 1.09561
R22776 VDD.n923 VDD 1.09561
R22777 VDD.n919 VDD 1.09561
R22778 VDD.n1182 VDD 1.09561
R22779 VDD.n1178 VDD 1.09561
R22780 VDD.n1441 VDD 1.09561
R22781 VDD.n1437 VDD 1.09561
R22782 VDD.n1700 VDD 1.09561
R22783 VDD.n1696 VDD 1.09561
R22784 VDD.n1959 VDD 1.09561
R22785 VDD.n1955 VDD 1.09561
R22786 VDD.n2218 VDD 1.09561
R22787 VDD.n2214 VDD 1.09561
R22788 VDD.n2477 VDD 1.09561
R22789 VDD.n2473 VDD 1.09561
R22790 VDD.n2736 VDD 1.09561
R22791 VDD.n2732 VDD 1.09561
R22792 VDD.n2995 VDD 1.09561
R22793 VDD.n2991 VDD 1.09561
R22794 VDD.n3254 VDD 1.09561
R22795 VDD.n3250 VDD 1.09561
R22796 VDD.n3513 VDD 1.09561
R22797 VDD.n3509 VDD 1.09561
R22798 VDD.n3772 VDD 1.09561
R22799 VDD.n3768 VDD 1.09561
R22800 VDD.n4031 VDD 1.09561
R22801 VDD.n4027 VDD 1.09561
R22802 VDD.n4290 VDD 1.09561
R22803 VDD.n4286 VDD 1.09561
R22804 VDD.n4549 VDD 1.09561
R22805 VDD.n4545 VDD 1.09561
R22806 VDD.n7293 VDD.n7292 1.02828
R22807 VDD.n7294 VDD.n7293 1.02828
R22808 VDD.n7290 VDD.n7289 1.02828
R22809 VDD.n400 VDD 1.01137
R22810 VDD.n387 VDD 1.01137
R22811 VDD.n310 VDD 1.01137
R22812 VDD.n333 VDD 1.01137
R22813 VDD VDD.n326 1.01137
R22814 VDD.n349 VDD 1.01137
R22815 VDD VDD.n292 1.01137
R22816 VDD.n648 VDD 1.01137
R22817 VDD.n635 VDD 1.01137
R22818 VDD.n558 VDD 1.01137
R22819 VDD.n581 VDD 1.01137
R22820 VDD VDD.n574 1.01137
R22821 VDD.n597 VDD 1.01137
R22822 VDD VDD.n540 1.01137
R22823 VDD.n907 VDD 1.01137
R22824 VDD.n894 VDD 1.01137
R22825 VDD.n817 VDD 1.01137
R22826 VDD.n840 VDD 1.01137
R22827 VDD VDD.n833 1.01137
R22828 VDD.n856 VDD 1.01137
R22829 VDD VDD.n799 1.01137
R22830 VDD.n1166 VDD 1.01137
R22831 VDD.n1153 VDD 1.01137
R22832 VDD.n1076 VDD 1.01137
R22833 VDD.n1099 VDD 1.01137
R22834 VDD VDD.n1092 1.01137
R22835 VDD.n1115 VDD 1.01137
R22836 VDD VDD.n1058 1.01137
R22837 VDD.n1425 VDD 1.01137
R22838 VDD.n1412 VDD 1.01137
R22839 VDD.n1335 VDD 1.01137
R22840 VDD.n1358 VDD 1.01137
R22841 VDD VDD.n1351 1.01137
R22842 VDD.n1374 VDD 1.01137
R22843 VDD VDD.n1317 1.01137
R22844 VDD.n1684 VDD 1.01137
R22845 VDD.n1671 VDD 1.01137
R22846 VDD.n1594 VDD 1.01137
R22847 VDD.n1617 VDD 1.01137
R22848 VDD VDD.n1610 1.01137
R22849 VDD.n1633 VDD 1.01137
R22850 VDD VDD.n1576 1.01137
R22851 VDD.n1943 VDD 1.01137
R22852 VDD.n1930 VDD 1.01137
R22853 VDD.n1853 VDD 1.01137
R22854 VDD.n1876 VDD 1.01137
R22855 VDD VDD.n1869 1.01137
R22856 VDD.n1892 VDD 1.01137
R22857 VDD VDD.n1835 1.01137
R22858 VDD.n2202 VDD 1.01137
R22859 VDD.n2189 VDD 1.01137
R22860 VDD.n2112 VDD 1.01137
R22861 VDD.n2135 VDD 1.01137
R22862 VDD VDD.n2128 1.01137
R22863 VDD.n2151 VDD 1.01137
R22864 VDD VDD.n2094 1.01137
R22865 VDD.n2461 VDD 1.01137
R22866 VDD.n2448 VDD 1.01137
R22867 VDD.n2371 VDD 1.01137
R22868 VDD.n2394 VDD 1.01137
R22869 VDD VDD.n2387 1.01137
R22870 VDD.n2410 VDD 1.01137
R22871 VDD VDD.n2353 1.01137
R22872 VDD.n2720 VDD 1.01137
R22873 VDD.n2707 VDD 1.01137
R22874 VDD.n2630 VDD 1.01137
R22875 VDD.n2653 VDD 1.01137
R22876 VDD VDD.n2646 1.01137
R22877 VDD.n2669 VDD 1.01137
R22878 VDD VDD.n2612 1.01137
R22879 VDD.n2979 VDD 1.01137
R22880 VDD.n2966 VDD 1.01137
R22881 VDD.n2889 VDD 1.01137
R22882 VDD.n2912 VDD 1.01137
R22883 VDD VDD.n2905 1.01137
R22884 VDD.n2928 VDD 1.01137
R22885 VDD VDD.n2871 1.01137
R22886 VDD.n3238 VDD 1.01137
R22887 VDD.n3225 VDD 1.01137
R22888 VDD.n3148 VDD 1.01137
R22889 VDD.n3171 VDD 1.01137
R22890 VDD VDD.n3164 1.01137
R22891 VDD.n3187 VDD 1.01137
R22892 VDD VDD.n3130 1.01137
R22893 VDD.n3497 VDD 1.01137
R22894 VDD.n3484 VDD 1.01137
R22895 VDD.n3407 VDD 1.01137
R22896 VDD.n3430 VDD 1.01137
R22897 VDD VDD.n3423 1.01137
R22898 VDD.n3446 VDD 1.01137
R22899 VDD VDD.n3389 1.01137
R22900 VDD.n3756 VDD 1.01137
R22901 VDD.n3743 VDD 1.01137
R22902 VDD.n3666 VDD 1.01137
R22903 VDD.n3689 VDD 1.01137
R22904 VDD VDD.n3682 1.01137
R22905 VDD.n3705 VDD 1.01137
R22906 VDD VDD.n3648 1.01137
R22907 VDD.n4015 VDD 1.01137
R22908 VDD.n4002 VDD 1.01137
R22909 VDD.n3925 VDD 1.01137
R22910 VDD.n3948 VDD 1.01137
R22911 VDD VDD.n3941 1.01137
R22912 VDD.n3964 VDD 1.01137
R22913 VDD VDD.n3907 1.01137
R22914 VDD.n4274 VDD 1.01137
R22915 VDD.n4261 VDD 1.01137
R22916 VDD.n4184 VDD 1.01137
R22917 VDD.n4207 VDD 1.01137
R22918 VDD VDD.n4200 1.01137
R22919 VDD.n4223 VDD 1.01137
R22920 VDD VDD.n4166 1.01137
R22921 VDD.n4533 VDD 1.01137
R22922 VDD.n4520 VDD 1.01137
R22923 VDD.n4443 VDD 1.01137
R22924 VDD.n4466 VDD 1.01137
R22925 VDD VDD.n4459 1.01137
R22926 VDD.n4482 VDD 1.01137
R22927 VDD VDD.n4425 1.01137
R22928 VDD VDD.n4721 1.01137
R22929 VDD VDD.n4722 1.01137
R22930 VDD VDD.n4746 1.01137
R22931 VDD VDD.n4762 1.01137
R22932 VDD VDD.n4763 1.01137
R22933 VDD VDD.n4787 1.01137
R22934 VDD VDD.n4803 1.01137
R22935 VDD VDD.n4804 1.01137
R22936 VDD VDD.n4828 1.01137
R22937 VDD VDD.n4844 1.01137
R22938 VDD VDD.n4845 1.01137
R22939 VDD VDD.n4869 1.01137
R22940 VDD VDD.n4885 1.01137
R22941 VDD VDD.n4886 1.01137
R22942 VDD VDD.n4910 1.01137
R22943 VDD VDD.n4926 1.01137
R22944 VDD VDD.n4927 1.01137
R22945 VDD VDD.n4951 1.01137
R22946 VDD VDD.n4967 1.01137
R22947 VDD VDD.n4968 1.01137
R22948 VDD VDD.n4992 1.01137
R22949 VDD VDD.n5008 1.01137
R22950 VDD VDD.n5009 1.01137
R22951 VDD VDD.n5033 1.01137
R22952 VDD VDD.n6027 1.01137
R22953 VDD.n6014 VDD 1.01137
R22954 VDD VDD.n6013 1.01137
R22955 VDD VDD.n5999 1.01137
R22956 VDD VDD.n5965 1.01137
R22957 VDD.n6190 VDD 1.01137
R22958 VDD VDD.n5933 1.01137
R22959 VDD VDD.n5899 1.01137
R22960 VDD.n5886 VDD 1.01137
R22961 VDD VDD.n5885 1.01137
R22962 VDD VDD.n5871 1.01137
R22963 VDD VDD.n5837 1.01137
R22964 VDD.n6321 VDD 1.01137
R22965 VDD VDD.n5805 1.01137
R22966 VDD VDD.n5771 1.01137
R22967 VDD.n5758 VDD 1.01137
R22968 VDD VDD.n5757 1.01137
R22969 VDD VDD.n5743 1.01137
R22970 VDD VDD.n5709 1.01137
R22971 VDD.n6452 VDD 1.01137
R22972 VDD VDD.n5677 1.01137
R22973 VDD VDD.n5643 1.01137
R22974 VDD.n5630 VDD 1.01137
R22975 VDD VDD.n5629 1.01137
R22976 VDD VDD.n5615 1.01137
R22977 VDD VDD.n5581 1.01137
R22978 VDD.n6583 VDD 1.01137
R22979 VDD VDD.n5549 1.01137
R22980 VDD VDD.n5515 1.01137
R22981 VDD.n5502 VDD 1.01137
R22982 VDD VDD.n5501 1.01137
R22983 VDD VDD.n5487 1.01137
R22984 VDD VDD.n5453 1.01137
R22985 VDD.n6714 VDD 1.01137
R22986 VDD VDD.n5421 1.01137
R22987 VDD VDD.n5387 1.01137
R22988 VDD.n5374 VDD 1.01137
R22989 VDD VDD.n5373 1.01137
R22990 VDD VDD.n5359 1.01137
R22991 VDD VDD.n5325 1.01137
R22992 VDD.n6845 VDD 1.01137
R22993 VDD VDD.n5293 1.01137
R22994 VDD VDD.n5259 1.01137
R22995 VDD.n5246 VDD 1.01137
R22996 VDD VDD.n5245 1.01137
R22997 VDD VDD.n5231 1.01137
R22998 VDD VDD.n5197 1.01137
R22999 VDD.n6976 VDD 1.01137
R23000 VDD VDD.n5165 1.01137
R23001 VDD VDD.n5131 1.01137
R23002 VDD.n5118 VDD 1.01137
R23003 VDD VDD.n5117 1.01137
R23004 VDD VDD.n5103 1.01137
R23005 VDD VDD.n5069 1.01137
R23006 VDD.n7104 VDD 1.01137
R23007 VDD.n7254 VDD 1.01137
R23008 VDD.n7233 VDD 1.01137
R23009 VDD.n7212 VDD 1.01137
R23010 VDD.n7191 VDD 1.01137
R23011 VDD.n7170 VDD 1.01137
R23012 VDD.n7149 VDD 1.01137
R23013 VDD.n7128 VDD 1.01137
R23014 VDD.n7107 VDD 1.01137
R23015 VDD.n19 VDD 0.980969
R23016 VDD.n38 VDD 0.980969
R23017 VDD.n57 VDD 0.980969
R23018 VDD.n76 VDD 0.980969
R23019 VDD.n95 VDD 0.980969
R23020 VDD.n114 VDD 0.980969
R23021 VDD.n133 VDD 0.980969
R23022 VDD.n152 VDD 0.980969
R23023 VDD.n4297 VDD 0.884883
R23024 VDD.n666 VDD.n665 0.859196
R23025 VDD.n662 VDD.n661 0.859196
R23026 VDD.n925 VDD.n924 0.859196
R23027 VDD.n921 VDD.n920 0.859196
R23028 VDD.n1184 VDD.n1183 0.859196
R23029 VDD.n1180 VDD.n1179 0.859196
R23030 VDD.n1443 VDD.n1442 0.859196
R23031 VDD.n1439 VDD.n1438 0.859196
R23032 VDD.n1702 VDD.n1701 0.859196
R23033 VDD.n1698 VDD.n1697 0.859196
R23034 VDD.n1961 VDD.n1960 0.859196
R23035 VDD.n1957 VDD.n1956 0.859196
R23036 VDD.n2220 VDD.n2219 0.859196
R23037 VDD.n2216 VDD.n2215 0.859196
R23038 VDD.n2479 VDD.n2478 0.859196
R23039 VDD.n2475 VDD.n2474 0.859196
R23040 VDD.n2738 VDD.n2737 0.859196
R23041 VDD.n2734 VDD.n2733 0.859196
R23042 VDD.n2997 VDD.n2996 0.859196
R23043 VDD.n2993 VDD.n2992 0.859196
R23044 VDD.n3256 VDD.n3255 0.859196
R23045 VDD.n3252 VDD.n3251 0.859196
R23046 VDD.n3515 VDD.n3514 0.859196
R23047 VDD.n3511 VDD.n3510 0.859196
R23048 VDD.n3774 VDD.n3773 0.859196
R23049 VDD.n3770 VDD.n3769 0.859196
R23050 VDD.n4033 VDD.n4032 0.859196
R23051 VDD.n4029 VDD.n4028 0.859196
R23052 VDD.n4292 VDD.n4291 0.859196
R23053 VDD.n4288 VDD.n4287 0.859196
R23054 VDD.n4551 VDD.n4550 0.859196
R23055 VDD.n4547 VDD.n4546 0.859196
R23056 VDD.n4721 VDD.n4700 0.834739
R23057 VDD.n4722 VDD.n4689 0.834739
R23058 VDD.n4746 VDD.n4689 0.834739
R23059 VDD.n4747 VDD.n4681 0.834739
R23060 VDD.n4762 VDD.n4681 0.834739
R23061 VDD.n4763 VDD.n4670 0.834739
R23062 VDD.n4787 VDD.n4670 0.834739
R23063 VDD.n4788 VDD.n4662 0.834739
R23064 VDD.n4803 VDD.n4662 0.834739
R23065 VDD.n4804 VDD.n4651 0.834739
R23066 VDD.n4828 VDD.n4651 0.834739
R23067 VDD.n4829 VDD.n4643 0.834739
R23068 VDD.n4844 VDD.n4643 0.834739
R23069 VDD.n4845 VDD.n4632 0.834739
R23070 VDD.n4869 VDD.n4632 0.834739
R23071 VDD.n4870 VDD.n4624 0.834739
R23072 VDD.n4885 VDD.n4624 0.834739
R23073 VDD.n4886 VDD.n4613 0.834739
R23074 VDD.n4910 VDD.n4613 0.834739
R23075 VDD.n4911 VDD.n4605 0.834739
R23076 VDD.n4926 VDD.n4605 0.834739
R23077 VDD.n4927 VDD.n4594 0.834739
R23078 VDD.n4951 VDD.n4594 0.834739
R23079 VDD.n4952 VDD.n4586 0.834739
R23080 VDD.n4967 VDD.n4586 0.834739
R23081 VDD.n4968 VDD.n4575 0.834739
R23082 VDD.n4992 VDD.n4575 0.834739
R23083 VDD.n4993 VDD.n4567 0.834739
R23084 VDD.n5008 VDD.n4567 0.834739
R23085 VDD.n5009 VDD.n4556 0.834739
R23086 VDD.n5033 VDD.n4556 0.834739
R23087 VDD.n6068 VDD.n6048 0.834739
R23088 VDD.n6027 VDD.n6026 0.834739
R23089 VDD.n6026 VDD.n6014 0.834739
R23090 VDD.n5999 VDD.n5998 0.834739
R23091 VDD.n5998 VDD.n5986 0.834739
R23092 VDD.n5965 VDD.n5964 0.834739
R23093 VDD.n5964 VDD.n5941 0.834739
R23094 VDD.n5933 VDD.n5932 0.834739
R23095 VDD.n5932 VDD.n5920 0.834739
R23096 VDD.n5899 VDD.n5898 0.834739
R23097 VDD.n5898 VDD.n5886 0.834739
R23098 VDD.n5871 VDD.n5870 0.834739
R23099 VDD.n5870 VDD.n5858 0.834739
R23100 VDD.n5837 VDD.n5836 0.834739
R23101 VDD.n5836 VDD.n5813 0.834739
R23102 VDD.n5805 VDD.n5804 0.834739
R23103 VDD.n5804 VDD.n5792 0.834739
R23104 VDD.n5771 VDD.n5770 0.834739
R23105 VDD.n5770 VDD.n5758 0.834739
R23106 VDD.n5743 VDD.n5742 0.834739
R23107 VDD.n5742 VDD.n5730 0.834739
R23108 VDD.n5709 VDD.n5708 0.834739
R23109 VDD.n5708 VDD.n5685 0.834739
R23110 VDD.n5677 VDD.n5676 0.834739
R23111 VDD.n5676 VDD.n5664 0.834739
R23112 VDD.n5643 VDD.n5642 0.834739
R23113 VDD.n5642 VDD.n5630 0.834739
R23114 VDD.n5615 VDD.n5614 0.834739
R23115 VDD.n5614 VDD.n5602 0.834739
R23116 VDD.n5581 VDD.n5580 0.834739
R23117 VDD.n5580 VDD.n5557 0.834739
R23118 VDD.n5549 VDD.n5548 0.834739
R23119 VDD.n5548 VDD.n5536 0.834739
R23120 VDD.n5515 VDD.n5514 0.834739
R23121 VDD.n5514 VDD.n5502 0.834739
R23122 VDD.n5487 VDD.n5486 0.834739
R23123 VDD.n5486 VDD.n5474 0.834739
R23124 VDD.n5453 VDD.n5452 0.834739
R23125 VDD.n5452 VDD.n5429 0.834739
R23126 VDD.n5421 VDD.n5420 0.834739
R23127 VDD.n5420 VDD.n5408 0.834739
R23128 VDD.n5387 VDD.n5386 0.834739
R23129 VDD.n5386 VDD.n5374 0.834739
R23130 VDD.n5359 VDD.n5358 0.834739
R23131 VDD.n5358 VDD.n5346 0.834739
R23132 VDD.n5325 VDD.n5324 0.834739
R23133 VDD.n5324 VDD.n5301 0.834739
R23134 VDD.n5293 VDD.n5292 0.834739
R23135 VDD.n5292 VDD.n5280 0.834739
R23136 VDD.n5259 VDD.n5258 0.834739
R23137 VDD.n5258 VDD.n5246 0.834739
R23138 VDD.n5231 VDD.n5230 0.834739
R23139 VDD.n5230 VDD.n5218 0.834739
R23140 VDD.n5197 VDD.n5196 0.834739
R23141 VDD.n5196 VDD.n5173 0.834739
R23142 VDD.n5165 VDD.n5164 0.834739
R23143 VDD.n5164 VDD.n5152 0.834739
R23144 VDD.n5131 VDD.n5130 0.834739
R23145 VDD.n5130 VDD.n5118 0.834739
R23146 VDD.n5103 VDD.n5102 0.834739
R23147 VDD.n5102 VDD.n5090 0.834739
R23148 VDD.n5069 VDD.n5068 0.834739
R23149 VDD.n5068 VDD.n5056 0.834739
R23150 VDD.n7328 VDD.n7327 0.819084
R23151 VDD.n7327 VDD.n7326 0.819084
R23152 VDD.n4556 VDD.n4555 0.807565
R23153 VDD.n4567 VDD.n4566 0.807565
R23154 VDD.n4575 VDD.n4574 0.807565
R23155 VDD.n4586 VDD.n4585 0.807565
R23156 VDD.n4594 VDD.n4593 0.807565
R23157 VDD.n4605 VDD.n4604 0.807565
R23158 VDD.n4613 VDD.n4612 0.807565
R23159 VDD.n4624 VDD.n4623 0.807565
R23160 VDD.n4632 VDD.n4631 0.807565
R23161 VDD.n4643 VDD.n4642 0.807565
R23162 VDD.n4651 VDD.n4650 0.807565
R23163 VDD.n4662 VDD.n4661 0.807565
R23164 VDD.n4670 VDD.n4669 0.807565
R23165 VDD.n4681 VDD.n4680 0.807565
R23166 VDD.n4689 VDD.n4688 0.807565
R23167 VDD.n4700 VDD.n4699 0.807565
R23168 VDD.n6068 VDD.n6066 0.807565
R23169 VDD.n6068 VDD.n6067 0.807565
R23170 VDD.n6026 VDD.n6024 0.807565
R23171 VDD.n6026 VDD.n6025 0.807565
R23172 VDD.n5998 VDD.n5996 0.807565
R23173 VDD.n5998 VDD.n5997 0.807565
R23174 VDD.n5964 VDD.n5962 0.807565
R23175 VDD.n5964 VDD.n5963 0.807565
R23176 VDD.n5932 VDD.n5930 0.807565
R23177 VDD.n5932 VDD.n5931 0.807565
R23178 VDD.n5898 VDD.n5896 0.807565
R23179 VDD.n5898 VDD.n5897 0.807565
R23180 VDD.n5870 VDD.n5868 0.807565
R23181 VDD.n5870 VDD.n5869 0.807565
R23182 VDD.n5836 VDD.n5834 0.807565
R23183 VDD.n5836 VDD.n5835 0.807565
R23184 VDD.n5804 VDD.n5802 0.807565
R23185 VDD.n5804 VDD.n5803 0.807565
R23186 VDD.n5770 VDD.n5768 0.807565
R23187 VDD.n5770 VDD.n5769 0.807565
R23188 VDD.n5742 VDD.n5740 0.807565
R23189 VDD.n5742 VDD.n5741 0.807565
R23190 VDD.n5708 VDD.n5706 0.807565
R23191 VDD.n5708 VDD.n5707 0.807565
R23192 VDD.n5676 VDD.n5674 0.807565
R23193 VDD.n5676 VDD.n5675 0.807565
R23194 VDD.n5642 VDD.n5640 0.807565
R23195 VDD.n5642 VDD.n5641 0.807565
R23196 VDD.n5614 VDD.n5612 0.807565
R23197 VDD.n5614 VDD.n5613 0.807565
R23198 VDD.n5580 VDD.n5578 0.807565
R23199 VDD.n5580 VDD.n5579 0.807565
R23200 VDD.n5548 VDD.n5546 0.807565
R23201 VDD.n5548 VDD.n5547 0.807565
R23202 VDD.n5514 VDD.n5512 0.807565
R23203 VDD.n5514 VDD.n5513 0.807565
R23204 VDD.n5486 VDD.n5484 0.807565
R23205 VDD.n5486 VDD.n5485 0.807565
R23206 VDD.n5452 VDD.n5450 0.807565
R23207 VDD.n5452 VDD.n5451 0.807565
R23208 VDD.n5420 VDD.n5418 0.807565
R23209 VDD.n5420 VDD.n5419 0.807565
R23210 VDD.n5386 VDD.n5384 0.807565
R23211 VDD.n5386 VDD.n5385 0.807565
R23212 VDD.n5358 VDD.n5356 0.807565
R23213 VDD.n5358 VDD.n5357 0.807565
R23214 VDD.n5324 VDD.n5322 0.807565
R23215 VDD.n5324 VDD.n5323 0.807565
R23216 VDD.n5292 VDD.n5290 0.807565
R23217 VDD.n5292 VDD.n5291 0.807565
R23218 VDD.n5258 VDD.n5256 0.807565
R23219 VDD.n5258 VDD.n5257 0.807565
R23220 VDD.n5230 VDD.n5228 0.807565
R23221 VDD.n5230 VDD.n5229 0.807565
R23222 VDD.n5196 VDD.n5194 0.807565
R23223 VDD.n5196 VDD.n5195 0.807565
R23224 VDD.n5164 VDD.n5162 0.807565
R23225 VDD.n5164 VDD.n5163 0.807565
R23226 VDD.n5130 VDD.n5128 0.807565
R23227 VDD.n5130 VDD.n5129 0.807565
R23228 VDD.n5102 VDD.n5100 0.807565
R23229 VDD.n5102 VDD.n5101 0.807565
R23230 VDD.n5068 VDD.n5066 0.807565
R23231 VDD.n5068 VDD.n5067 0.807565
R23232 VDD.n7310 VDD.n7276 0.807565
R23233 VDD.n645 VDD.n417 0.783109
R23234 VDD.n904 VDD.n676 0.783109
R23235 VDD.n1163 VDD.n935 0.783109
R23236 VDD.n1422 VDD.n1194 0.783109
R23237 VDD.n1681 VDD.n1453 0.783109
R23238 VDD.n1940 VDD.n1712 0.783109
R23239 VDD.n2199 VDD.n1971 0.783109
R23240 VDD.n2458 VDD.n2230 0.783109
R23241 VDD.n2717 VDD.n2489 0.783109
R23242 VDD.n2976 VDD.n2748 0.783109
R23243 VDD.n3235 VDD.n3007 0.783109
R23244 VDD.n3494 VDD.n3266 0.783109
R23245 VDD.n3753 VDD.n3525 0.783109
R23246 VDD.n4012 VDD.n3784 0.783109
R23247 VDD.n4271 VDD.n4043 0.783109
R23248 VDD.n4530 VDD.n4302 0.783109
R23249 VDD.n7323 VDD.n7322 0.774559
R23250 VDD.n7324 VDD.n7323 0.774559
R23251 VDD.n387 VDD.n386 0.772239
R23252 VDD.n385 VDD.n384 0.772239
R23253 VDD.n311 VDD.n310 0.772239
R23254 VDD.n326 VDD.n312 0.772239
R23255 VDD.n350 VDD.n349 0.772239
R23256 VDD.n365 VDD.n351 0.772239
R23257 VDD.n292 VDD.n278 0.772239
R23258 VDD.n406 VDD.n170 0.772239
R23259 VDD.n635 VDD.n634 0.772239
R23260 VDD.n633 VDD.n632 0.772239
R23261 VDD.n559 VDD.n558 0.772239
R23262 VDD.n574 VDD.n560 0.772239
R23263 VDD.n598 VDD.n597 0.772239
R23264 VDD.n613 VDD.n599 0.772239
R23265 VDD.n540 VDD.n526 0.772239
R23266 VDD.n654 VDD.n418 0.772239
R23267 VDD.n894 VDD.n893 0.772239
R23268 VDD.n892 VDD.n891 0.772239
R23269 VDD.n818 VDD.n817 0.772239
R23270 VDD.n833 VDD.n819 0.772239
R23271 VDD.n857 VDD.n856 0.772239
R23272 VDD.n872 VDD.n858 0.772239
R23273 VDD.n799 VDD.n785 0.772239
R23274 VDD.n913 VDD.n677 0.772239
R23275 VDD.n1153 VDD.n1152 0.772239
R23276 VDD.n1151 VDD.n1150 0.772239
R23277 VDD.n1077 VDD.n1076 0.772239
R23278 VDD.n1092 VDD.n1078 0.772239
R23279 VDD.n1116 VDD.n1115 0.772239
R23280 VDD.n1131 VDD.n1117 0.772239
R23281 VDD.n1058 VDD.n1044 0.772239
R23282 VDD.n1172 VDD.n936 0.772239
R23283 VDD.n1412 VDD.n1411 0.772239
R23284 VDD.n1410 VDD.n1409 0.772239
R23285 VDD.n1336 VDD.n1335 0.772239
R23286 VDD.n1351 VDD.n1337 0.772239
R23287 VDD.n1375 VDD.n1374 0.772239
R23288 VDD.n1390 VDD.n1376 0.772239
R23289 VDD.n1317 VDD.n1303 0.772239
R23290 VDD.n1431 VDD.n1195 0.772239
R23291 VDD.n1671 VDD.n1670 0.772239
R23292 VDD.n1669 VDD.n1668 0.772239
R23293 VDD.n1595 VDD.n1594 0.772239
R23294 VDD.n1610 VDD.n1596 0.772239
R23295 VDD.n1634 VDD.n1633 0.772239
R23296 VDD.n1649 VDD.n1635 0.772239
R23297 VDD.n1576 VDD.n1562 0.772239
R23298 VDD.n1690 VDD.n1454 0.772239
R23299 VDD.n1930 VDD.n1929 0.772239
R23300 VDD.n1928 VDD.n1927 0.772239
R23301 VDD.n1854 VDD.n1853 0.772239
R23302 VDD.n1869 VDD.n1855 0.772239
R23303 VDD.n1893 VDD.n1892 0.772239
R23304 VDD.n1908 VDD.n1894 0.772239
R23305 VDD.n1835 VDD.n1821 0.772239
R23306 VDD.n1949 VDD.n1713 0.772239
R23307 VDD.n2189 VDD.n2188 0.772239
R23308 VDD.n2187 VDD.n2186 0.772239
R23309 VDD.n2113 VDD.n2112 0.772239
R23310 VDD.n2128 VDD.n2114 0.772239
R23311 VDD.n2152 VDD.n2151 0.772239
R23312 VDD.n2167 VDD.n2153 0.772239
R23313 VDD.n2094 VDD.n2080 0.772239
R23314 VDD.n2208 VDD.n1972 0.772239
R23315 VDD.n2448 VDD.n2447 0.772239
R23316 VDD.n2446 VDD.n2445 0.772239
R23317 VDD.n2372 VDD.n2371 0.772239
R23318 VDD.n2387 VDD.n2373 0.772239
R23319 VDD.n2411 VDD.n2410 0.772239
R23320 VDD.n2426 VDD.n2412 0.772239
R23321 VDD.n2353 VDD.n2339 0.772239
R23322 VDD.n2467 VDD.n2231 0.772239
R23323 VDD.n2707 VDD.n2706 0.772239
R23324 VDD.n2705 VDD.n2704 0.772239
R23325 VDD.n2631 VDD.n2630 0.772239
R23326 VDD.n2646 VDD.n2632 0.772239
R23327 VDD.n2670 VDD.n2669 0.772239
R23328 VDD.n2685 VDD.n2671 0.772239
R23329 VDD.n2612 VDD.n2598 0.772239
R23330 VDD.n2726 VDD.n2490 0.772239
R23331 VDD.n2966 VDD.n2965 0.772239
R23332 VDD.n2964 VDD.n2963 0.772239
R23333 VDD.n2890 VDD.n2889 0.772239
R23334 VDD.n2905 VDD.n2891 0.772239
R23335 VDD.n2929 VDD.n2928 0.772239
R23336 VDD.n2944 VDD.n2930 0.772239
R23337 VDD.n2871 VDD.n2857 0.772239
R23338 VDD.n2985 VDD.n2749 0.772239
R23339 VDD.n3225 VDD.n3224 0.772239
R23340 VDD.n3223 VDD.n3222 0.772239
R23341 VDD.n3149 VDD.n3148 0.772239
R23342 VDD.n3164 VDD.n3150 0.772239
R23343 VDD.n3188 VDD.n3187 0.772239
R23344 VDD.n3203 VDD.n3189 0.772239
R23345 VDD.n3130 VDD.n3116 0.772239
R23346 VDD.n3244 VDD.n3008 0.772239
R23347 VDD.n3484 VDD.n3483 0.772239
R23348 VDD.n3482 VDD.n3481 0.772239
R23349 VDD.n3408 VDD.n3407 0.772239
R23350 VDD.n3423 VDD.n3409 0.772239
R23351 VDD.n3447 VDD.n3446 0.772239
R23352 VDD.n3462 VDD.n3448 0.772239
R23353 VDD.n3389 VDD.n3375 0.772239
R23354 VDD.n3503 VDD.n3267 0.772239
R23355 VDD.n3743 VDD.n3742 0.772239
R23356 VDD.n3741 VDD.n3740 0.772239
R23357 VDD.n3667 VDD.n3666 0.772239
R23358 VDD.n3682 VDD.n3668 0.772239
R23359 VDD.n3706 VDD.n3705 0.772239
R23360 VDD.n3721 VDD.n3707 0.772239
R23361 VDD.n3648 VDD.n3634 0.772239
R23362 VDD.n3762 VDD.n3526 0.772239
R23363 VDD.n4002 VDD.n4001 0.772239
R23364 VDD.n4000 VDD.n3999 0.772239
R23365 VDD.n3926 VDD.n3925 0.772239
R23366 VDD.n3941 VDD.n3927 0.772239
R23367 VDD.n3965 VDD.n3964 0.772239
R23368 VDD.n3980 VDD.n3966 0.772239
R23369 VDD.n3907 VDD.n3893 0.772239
R23370 VDD.n4021 VDD.n3785 0.772239
R23371 VDD.n4261 VDD.n4260 0.772239
R23372 VDD.n4259 VDD.n4258 0.772239
R23373 VDD.n4185 VDD.n4184 0.772239
R23374 VDD.n4200 VDD.n4186 0.772239
R23375 VDD.n4224 VDD.n4223 0.772239
R23376 VDD.n4239 VDD.n4225 0.772239
R23377 VDD.n4166 VDD.n4152 0.772239
R23378 VDD.n4280 VDD.n4044 0.772239
R23379 VDD.n4520 VDD.n4519 0.772239
R23380 VDD.n4518 VDD.n4517 0.772239
R23381 VDD.n4444 VDD.n4443 0.772239
R23382 VDD.n4459 VDD.n4445 0.772239
R23383 VDD.n4483 VDD.n4482 0.772239
R23384 VDD.n4498 VDD.n4484 0.772239
R23385 VDD.n4425 VDD.n4411 0.772239
R23386 VDD.n4539 VDD.n4303 0.772239
R23387 VDD.n4300 VDD 0.716182
R23388 VDD.n4041 VDD 0.716182
R23389 VDD.n3782 VDD 0.716182
R23390 VDD.n3523 VDD 0.716182
R23391 VDD.n3264 VDD 0.716182
R23392 VDD.n3005 VDD 0.716182
R23393 VDD.n2746 VDD 0.716182
R23394 VDD.n2487 VDD 0.716182
R23395 VDD.n2228 VDD 0.716182
R23396 VDD.n1969 VDD 0.716182
R23397 VDD.n1710 VDD 0.716182
R23398 VDD.n1451 VDD 0.716182
R23399 VDD.n1192 VDD 0.716182
R23400 VDD.n933 VDD 0.716182
R23401 VDD.n674 VDD 0.716182
R23402 VDD.n415 VDD 0.716182
R23403 VDD.n167 VDD 0.716182
R23404 VDD.n655 VDD.n654 0.712457
R23405 VDD.n914 VDD.n913 0.712457
R23406 VDD.n1173 VDD.n1172 0.712457
R23407 VDD.n1432 VDD.n1431 0.712457
R23408 VDD.n1691 VDD.n1690 0.712457
R23409 VDD.n1950 VDD.n1949 0.712457
R23410 VDD.n2209 VDD.n2208 0.712457
R23411 VDD.n2468 VDD.n2467 0.712457
R23412 VDD.n2727 VDD.n2726 0.712457
R23413 VDD.n2986 VDD.n2985 0.712457
R23414 VDD.n3245 VDD.n3244 0.712457
R23415 VDD.n3504 VDD.n3503 0.712457
R23416 VDD.n3763 VDD.n3762 0.712457
R23417 VDD.n4022 VDD.n4021 0.712457
R23418 VDD.n4281 VDD.n4280 0.712457
R23419 VDD.n4540 VDD.n4539 0.712457
R23420 VDD.n666 VDD 0.662609
R23421 VDD.n662 VDD 0.662609
R23422 VDD.n925 VDD 0.662609
R23423 VDD.n921 VDD 0.662609
R23424 VDD.n1184 VDD 0.662609
R23425 VDD.n1180 VDD 0.662609
R23426 VDD.n1443 VDD 0.662609
R23427 VDD.n1439 VDD 0.662609
R23428 VDD.n1702 VDD 0.662609
R23429 VDD.n1698 VDD 0.662609
R23430 VDD.n1961 VDD 0.662609
R23431 VDD.n1957 VDD 0.662609
R23432 VDD.n2220 VDD 0.662609
R23433 VDD.n2216 VDD 0.662609
R23434 VDD.n2479 VDD 0.662609
R23435 VDD.n2475 VDD 0.662609
R23436 VDD.n2738 VDD 0.662609
R23437 VDD.n2734 VDD 0.662609
R23438 VDD.n2997 VDD 0.662609
R23439 VDD.n2993 VDD 0.662609
R23440 VDD.n3256 VDD 0.662609
R23441 VDD.n3252 VDD 0.662609
R23442 VDD.n3515 VDD 0.662609
R23443 VDD.n3511 VDD 0.662609
R23444 VDD.n3774 VDD 0.662609
R23445 VDD.n3770 VDD 0.662609
R23446 VDD.n4033 VDD 0.662609
R23447 VDD.n4029 VDD 0.662609
R23448 VDD.n4292 VDD 0.662609
R23449 VDD.n4288 VDD 0.662609
R23450 VDD.n4551 VDD 0.662609
R23451 VDD.n4547 VDD 0.662609
R23452 VDD.n149 VDD.n148 0.648317
R23453 VDD.n130 VDD.n129 0.648317
R23454 VDD.n111 VDD.n110 0.648317
R23455 VDD.n92 VDD.n91 0.648317
R23456 VDD.n73 VDD.n72 0.648317
R23457 VDD.n54 VDD.n53 0.648317
R23458 VDD.n35 VDD.n34 0.648317
R23459 VDD.n16 VDD.n15 0.648317
R23460 VDD.n4301 VDD 0.638917
R23461 VDD.n4042 VDD 0.638917
R23462 VDD.n3783 VDD 0.638917
R23463 VDD.n3524 VDD 0.638917
R23464 VDD.n3265 VDD 0.638917
R23465 VDD.n3006 VDD 0.638917
R23466 VDD.n2747 VDD 0.638917
R23467 VDD.n2488 VDD 0.638917
R23468 VDD.n2229 VDD 0.638917
R23469 VDD.n1970 VDD 0.638917
R23470 VDD.n1711 VDD 0.638917
R23471 VDD.n1452 VDD 0.638917
R23472 VDD.n1193 VDD 0.638917
R23473 VDD.n934 VDD 0.638917
R23474 VDD.n675 VDD 0.638917
R23475 VDD.n416 VDD 0.638917
R23476 VDD.n7310 VDD.n7309 0.6205
R23477 VDD.n4723 VDD 0.601043
R23478 VDD.n4764 VDD 0.601043
R23479 VDD.n4805 VDD 0.601043
R23480 VDD.n4846 VDD 0.601043
R23481 VDD.n4887 VDD 0.601043
R23482 VDD.n4928 VDD 0.601043
R23483 VDD.n4969 VDD 0.601043
R23484 VDD.n5010 VDD 0.601043
R23485 VDD.n6037 VDD 0.601043
R23486 VDD.n6012 VDD 0.601043
R23487 VDD.n5975 VDD 0.601043
R23488 VDD VDD.n6188 0.601043
R23489 VDD.n6189 VDD 0.601043
R23490 VDD.n5909 VDD 0.601043
R23491 VDD.n5884 VDD 0.601043
R23492 VDD.n5847 VDD 0.601043
R23493 VDD VDD.n6319 0.601043
R23494 VDD.n6320 VDD 0.601043
R23495 VDD.n5781 VDD 0.601043
R23496 VDD.n5756 VDD 0.601043
R23497 VDD.n5719 VDD 0.601043
R23498 VDD VDD.n6450 0.601043
R23499 VDD.n6451 VDD 0.601043
R23500 VDD.n5653 VDD 0.601043
R23501 VDD.n5628 VDD 0.601043
R23502 VDD.n5591 VDD 0.601043
R23503 VDD VDD.n6581 0.601043
R23504 VDD.n6582 VDD 0.601043
R23505 VDD.n5525 VDD 0.601043
R23506 VDD.n5500 VDD 0.601043
R23507 VDD.n5463 VDD 0.601043
R23508 VDD VDD.n6712 0.601043
R23509 VDD.n6713 VDD 0.601043
R23510 VDD.n5397 VDD 0.601043
R23511 VDD.n5372 VDD 0.601043
R23512 VDD.n5335 VDD 0.601043
R23513 VDD VDD.n6843 0.601043
R23514 VDD.n6844 VDD 0.601043
R23515 VDD.n5269 VDD 0.601043
R23516 VDD.n5244 VDD 0.601043
R23517 VDD.n5207 VDD 0.601043
R23518 VDD VDD.n6974 0.601043
R23519 VDD.n6975 VDD 0.601043
R23520 VDD.n5141 VDD 0.601043
R23521 VDD.n5116 VDD 0.601043
R23522 VDD.n5079 VDD 0.601043
R23523 VDD.n5045 VDD 0.601043
R23524 VDD VDD.n7105 0.601043
R23525 VDD.n149 VDD 0.592985
R23526 VDD.n130 VDD 0.592985
R23527 VDD.n111 VDD 0.592985
R23528 VDD.n92 VDD 0.592985
R23529 VDD.n73 VDD 0.592985
R23530 VDD.n54 VDD 0.592985
R23531 VDD.n35 VDD 0.592985
R23532 VDD.n16 VDD 0.592985
R23533 VDD.n4544 VDD.n4543 0.5833
R23534 VDD.n4285 VDD.n4284 0.5833
R23535 VDD.n4026 VDD.n4025 0.5833
R23536 VDD.n3767 VDD.n3766 0.5833
R23537 VDD.n3508 VDD.n3507 0.5833
R23538 VDD.n3249 VDD.n3248 0.5833
R23539 VDD.n2990 VDD.n2989 0.5833
R23540 VDD.n2731 VDD.n2730 0.5833
R23541 VDD.n2472 VDD.n2471 0.5833
R23542 VDD.n2213 VDD.n2212 0.5833
R23543 VDD.n1954 VDD.n1953 0.5833
R23544 VDD.n1695 VDD.n1694 0.5833
R23545 VDD.n1436 VDD.n1435 0.5833
R23546 VDD.n1177 VDD.n1176 0.5833
R23547 VDD.n918 VDD.n917 0.5833
R23548 VDD.n659 VDD.n658 0.5833
R23549 VDD.n168 VDD.n167 0.5833
R23550 VDD VDD.n399 0.538543
R23551 VDD VDD.n296 0.538543
R23552 VDD VDD.n335 0.538543
R23553 VDD.n293 VDD 0.538543
R23554 VDD VDD.n647 0.538543
R23555 VDD VDD.n544 0.538543
R23556 VDD VDD.n583 0.538543
R23557 VDD.n541 VDD 0.538543
R23558 VDD VDD.n906 0.538543
R23559 VDD VDD.n803 0.538543
R23560 VDD VDD.n842 0.538543
R23561 VDD.n800 VDD 0.538543
R23562 VDD VDD.n1165 0.538543
R23563 VDD VDD.n1062 0.538543
R23564 VDD VDD.n1101 0.538543
R23565 VDD.n1059 VDD 0.538543
R23566 VDD VDD.n1424 0.538543
R23567 VDD VDD.n1321 0.538543
R23568 VDD VDD.n1360 0.538543
R23569 VDD.n1318 VDD 0.538543
R23570 VDD VDD.n1683 0.538543
R23571 VDD VDD.n1580 0.538543
R23572 VDD VDD.n1619 0.538543
R23573 VDD.n1577 VDD 0.538543
R23574 VDD VDD.n1942 0.538543
R23575 VDD VDD.n1839 0.538543
R23576 VDD VDD.n1878 0.538543
R23577 VDD.n1836 VDD 0.538543
R23578 VDD VDD.n2201 0.538543
R23579 VDD VDD.n2098 0.538543
R23580 VDD VDD.n2137 0.538543
R23581 VDD.n2095 VDD 0.538543
R23582 VDD VDD.n2460 0.538543
R23583 VDD VDD.n2357 0.538543
R23584 VDD VDD.n2396 0.538543
R23585 VDD.n2354 VDD 0.538543
R23586 VDD VDD.n2719 0.538543
R23587 VDD VDD.n2616 0.538543
R23588 VDD VDD.n2655 0.538543
R23589 VDD.n2613 VDD 0.538543
R23590 VDD VDD.n2978 0.538543
R23591 VDD VDD.n2875 0.538543
R23592 VDD VDD.n2914 0.538543
R23593 VDD.n2872 VDD 0.538543
R23594 VDD VDD.n3237 0.538543
R23595 VDD VDD.n3134 0.538543
R23596 VDD VDD.n3173 0.538543
R23597 VDD.n3131 VDD 0.538543
R23598 VDD VDD.n3496 0.538543
R23599 VDD VDD.n3393 0.538543
R23600 VDD VDD.n3432 0.538543
R23601 VDD.n3390 VDD 0.538543
R23602 VDD VDD.n3755 0.538543
R23603 VDD VDD.n3652 0.538543
R23604 VDD VDD.n3691 0.538543
R23605 VDD.n3649 VDD 0.538543
R23606 VDD VDD.n4014 0.538543
R23607 VDD VDD.n3911 0.538543
R23608 VDD VDD.n3950 0.538543
R23609 VDD.n3908 VDD 0.538543
R23610 VDD VDD.n4273 0.538543
R23611 VDD VDD.n4170 0.538543
R23612 VDD VDD.n4209 0.538543
R23613 VDD.n4167 VDD 0.538543
R23614 VDD VDD.n4532 0.538543
R23615 VDD VDD.n4429 0.538543
R23616 VDD VDD.n4468 0.538543
R23617 VDD.n4426 VDD 0.538543
R23618 VDD.n4543 VDD 0.533879
R23619 VDD.n4284 VDD 0.533879
R23620 VDD.n4025 VDD 0.533879
R23621 VDD.n3766 VDD 0.533879
R23622 VDD.n3507 VDD 0.533879
R23623 VDD.n3248 VDD 0.533879
R23624 VDD.n2989 VDD 0.533879
R23625 VDD.n2730 VDD 0.533879
R23626 VDD.n2471 VDD 0.533879
R23627 VDD.n2212 VDD 0.533879
R23628 VDD.n1953 VDD 0.533879
R23629 VDD.n1694 VDD 0.533879
R23630 VDD.n1435 VDD 0.533879
R23631 VDD.n1176 VDD 0.533879
R23632 VDD.n917 VDD 0.533879
R23633 VDD.n658 VDD 0.533879
R23634 VDD.n161 VDD 0.524957
R23635 VDD.n157 VDD 0.524957
R23636 VDD.n7286 VDD.n7277 0.486913
R23637 VDD.n4724 VDD.n4723 0.410826
R23638 VDD.n4765 VDD.n4764 0.410826
R23639 VDD.n4806 VDD.n4805 0.410826
R23640 VDD.n4847 VDD.n4846 0.410826
R23641 VDD.n4888 VDD.n4887 0.410826
R23642 VDD.n4929 VDD.n4928 0.410826
R23643 VDD.n4970 VDD.n4969 0.410826
R23644 VDD.n5011 VDD.n5010 0.410826
R23645 VDD.n6038 VDD.n6037 0.410826
R23646 VDD.n6013 VDD.n6012 0.410826
R23647 VDD.n5976 VDD.n5975 0.410826
R23648 VDD.n6188 VDD.n6187 0.410826
R23649 VDD.n6190 VDD.n6189 0.410826
R23650 VDD.n5910 VDD.n5909 0.410826
R23651 VDD.n5885 VDD.n5884 0.410826
R23652 VDD.n5848 VDD.n5847 0.410826
R23653 VDD.n6319 VDD.n6318 0.410826
R23654 VDD.n6321 VDD.n6320 0.410826
R23655 VDD.n5782 VDD.n5781 0.410826
R23656 VDD.n5757 VDD.n5756 0.410826
R23657 VDD.n5720 VDD.n5719 0.410826
R23658 VDD.n6450 VDD.n6449 0.410826
R23659 VDD.n6452 VDD.n6451 0.410826
R23660 VDD.n5654 VDD.n5653 0.410826
R23661 VDD.n5629 VDD.n5628 0.410826
R23662 VDD.n5592 VDD.n5591 0.410826
R23663 VDD.n6581 VDD.n6580 0.410826
R23664 VDD.n6583 VDD.n6582 0.410826
R23665 VDD.n5526 VDD.n5525 0.410826
R23666 VDD.n5501 VDD.n5500 0.410826
R23667 VDD.n5464 VDD.n5463 0.410826
R23668 VDD.n6712 VDD.n6711 0.410826
R23669 VDD.n6714 VDD.n6713 0.410826
R23670 VDD.n5398 VDD.n5397 0.410826
R23671 VDD.n5373 VDD.n5372 0.410826
R23672 VDD.n5336 VDD.n5335 0.410826
R23673 VDD.n6843 VDD.n6842 0.410826
R23674 VDD.n6845 VDD.n6844 0.410826
R23675 VDD.n5270 VDD.n5269 0.410826
R23676 VDD.n5245 VDD.n5244 0.410826
R23677 VDD.n5208 VDD.n5207 0.410826
R23678 VDD.n6974 VDD.n6973 0.410826
R23679 VDD.n6976 VDD.n6975 0.410826
R23680 VDD.n5142 VDD.n5141 0.410826
R23681 VDD.n5117 VDD.n5116 0.410826
R23682 VDD.n5080 VDD.n5079 0.410826
R23683 VDD.n5046 VDD.n5045 0.410826
R23684 VDD.n7105 VDD.n7104 0.410826
R23685 VDD.n7274 VDD.n1 0.405391
R23686 VDD.n7253 VDD.n20 0.405391
R23687 VDD.n7232 VDD.n39 0.405391
R23688 VDD.n7211 VDD.n58 0.405391
R23689 VDD.n7190 VDD.n77 0.405391
R23690 VDD.n7169 VDD.n96 0.405391
R23691 VDD.n7148 VDD.n115 0.405391
R23692 VDD.n7127 VDD.n134 0.405391
R23693 VDD.n7319 VDD.n7312 0.397496
R23694 VDD.n7319 VDD.n7318 0.397496
R23695 VDD.n397 VDD.n169 0.378217
R23696 VDD.n7254 VDD.n19 0.353761
R23697 VDD.n7233 VDD.n38 0.353761
R23698 VDD.n7212 VDD.n57 0.353761
R23699 VDD.n7191 VDD.n76 0.353761
R23700 VDD.n7170 VDD.n95 0.353761
R23701 VDD.n7149 VDD.n114 0.353761
R23702 VDD.n7128 VDD.n133 0.353761
R23703 VDD.n7107 VDD.n152 0.353761
R23704 VDD.n400 VDD.n191 0.348326
R23705 VDD.n398 VDD.n397 0.348326
R23706 VDD.n295 VDD.n229 0.348326
R23707 VDD.n334 VDD.n333 0.348326
R23708 VDD.n366 VDD.n294 0.348326
R23709 VDD.n648 VDD.n439 0.348326
R23710 VDD.n646 VDD.n645 0.348326
R23711 VDD.n543 VDD.n477 0.348326
R23712 VDD.n582 VDD.n581 0.348326
R23713 VDD.n614 VDD.n542 0.348326
R23714 VDD.n907 VDD.n698 0.348326
R23715 VDD.n905 VDD.n904 0.348326
R23716 VDD.n802 VDD.n736 0.348326
R23717 VDD.n841 VDD.n840 0.348326
R23718 VDD.n873 VDD.n801 0.348326
R23719 VDD.n1166 VDD.n957 0.348326
R23720 VDD.n1164 VDD.n1163 0.348326
R23721 VDD.n1061 VDD.n995 0.348326
R23722 VDD.n1100 VDD.n1099 0.348326
R23723 VDD.n1132 VDD.n1060 0.348326
R23724 VDD.n1425 VDD.n1216 0.348326
R23725 VDD.n1423 VDD.n1422 0.348326
R23726 VDD.n1320 VDD.n1254 0.348326
R23727 VDD.n1359 VDD.n1358 0.348326
R23728 VDD.n1391 VDD.n1319 0.348326
R23729 VDD.n1684 VDD.n1475 0.348326
R23730 VDD.n1682 VDD.n1681 0.348326
R23731 VDD.n1579 VDD.n1513 0.348326
R23732 VDD.n1618 VDD.n1617 0.348326
R23733 VDD.n1650 VDD.n1578 0.348326
R23734 VDD.n1943 VDD.n1734 0.348326
R23735 VDD.n1941 VDD.n1940 0.348326
R23736 VDD.n1838 VDD.n1772 0.348326
R23737 VDD.n1877 VDD.n1876 0.348326
R23738 VDD.n1909 VDD.n1837 0.348326
R23739 VDD.n2202 VDD.n1993 0.348326
R23740 VDD.n2200 VDD.n2199 0.348326
R23741 VDD.n2097 VDD.n2031 0.348326
R23742 VDD.n2136 VDD.n2135 0.348326
R23743 VDD.n2168 VDD.n2096 0.348326
R23744 VDD.n2461 VDD.n2252 0.348326
R23745 VDD.n2459 VDD.n2458 0.348326
R23746 VDD.n2356 VDD.n2290 0.348326
R23747 VDD.n2395 VDD.n2394 0.348326
R23748 VDD.n2427 VDD.n2355 0.348326
R23749 VDD.n2720 VDD.n2511 0.348326
R23750 VDD.n2718 VDD.n2717 0.348326
R23751 VDD.n2615 VDD.n2549 0.348326
R23752 VDD.n2654 VDD.n2653 0.348326
R23753 VDD.n2686 VDD.n2614 0.348326
R23754 VDD.n2979 VDD.n2770 0.348326
R23755 VDD.n2977 VDD.n2976 0.348326
R23756 VDD.n2874 VDD.n2808 0.348326
R23757 VDD.n2913 VDD.n2912 0.348326
R23758 VDD.n2945 VDD.n2873 0.348326
R23759 VDD.n3238 VDD.n3029 0.348326
R23760 VDD.n3236 VDD.n3235 0.348326
R23761 VDD.n3133 VDD.n3067 0.348326
R23762 VDD.n3172 VDD.n3171 0.348326
R23763 VDD.n3204 VDD.n3132 0.348326
R23764 VDD.n3497 VDD.n3288 0.348326
R23765 VDD.n3495 VDD.n3494 0.348326
R23766 VDD.n3392 VDD.n3326 0.348326
R23767 VDD.n3431 VDD.n3430 0.348326
R23768 VDD.n3463 VDD.n3391 0.348326
R23769 VDD.n3756 VDD.n3547 0.348326
R23770 VDD.n3754 VDD.n3753 0.348326
R23771 VDD.n3651 VDD.n3585 0.348326
R23772 VDD.n3690 VDD.n3689 0.348326
R23773 VDD.n3722 VDD.n3650 0.348326
R23774 VDD.n4015 VDD.n3806 0.348326
R23775 VDD.n4013 VDD.n4012 0.348326
R23776 VDD.n3910 VDD.n3844 0.348326
R23777 VDD.n3949 VDD.n3948 0.348326
R23778 VDD.n3981 VDD.n3909 0.348326
R23779 VDD.n4274 VDD.n4065 0.348326
R23780 VDD.n4272 VDD.n4271 0.348326
R23781 VDD.n4169 VDD.n4103 0.348326
R23782 VDD.n4208 VDD.n4207 0.348326
R23783 VDD.n4240 VDD.n4168 0.348326
R23784 VDD.n4533 VDD.n4324 0.348326
R23785 VDD.n4531 VDD.n4530 0.348326
R23786 VDD.n4428 VDD.n4362 0.348326
R23787 VDD.n4467 VDD.n4466 0.348326
R23788 VDD.n4499 VDD.n4427 0.348326
R23789 VDD.n7330 VDD.n7329 0.344944
R23790 VDD.n398 VDD 0.295582
R23791 VDD.n295 VDD 0.295582
R23792 VDD.n294 VDD 0.295582
R23793 VDD.n646 VDD 0.295582
R23794 VDD.n543 VDD 0.295582
R23795 VDD.n542 VDD 0.295582
R23796 VDD.n905 VDD 0.295582
R23797 VDD.n802 VDD 0.295582
R23798 VDD.n801 VDD 0.295582
R23799 VDD.n1164 VDD 0.295582
R23800 VDD.n1061 VDD 0.295582
R23801 VDD.n1060 VDD 0.295582
R23802 VDD.n1423 VDD 0.295582
R23803 VDD.n1320 VDD 0.295582
R23804 VDD.n1319 VDD 0.295582
R23805 VDD.n1682 VDD 0.295582
R23806 VDD.n1579 VDD 0.295582
R23807 VDD.n1578 VDD 0.295582
R23808 VDD.n1941 VDD 0.295582
R23809 VDD.n1838 VDD 0.295582
R23810 VDD.n1837 VDD 0.295582
R23811 VDD.n2200 VDD 0.295582
R23812 VDD.n2097 VDD 0.295582
R23813 VDD.n2096 VDD 0.295582
R23814 VDD.n2459 VDD 0.295582
R23815 VDD.n2356 VDD 0.295582
R23816 VDD.n2355 VDD 0.295582
R23817 VDD.n2718 VDD 0.295582
R23818 VDD.n2615 VDD 0.295582
R23819 VDD.n2614 VDD 0.295582
R23820 VDD.n2977 VDD 0.295582
R23821 VDD.n2874 VDD 0.295582
R23822 VDD.n2873 VDD 0.295582
R23823 VDD.n3236 VDD 0.295582
R23824 VDD.n3133 VDD 0.295582
R23825 VDD.n3132 VDD 0.295582
R23826 VDD.n3495 VDD 0.295582
R23827 VDD.n3392 VDD 0.295582
R23828 VDD.n3391 VDD 0.295582
R23829 VDD.n3754 VDD 0.295582
R23830 VDD.n3651 VDD 0.295582
R23831 VDD.n3650 VDD 0.295582
R23832 VDD.n4013 VDD 0.295582
R23833 VDD.n3910 VDD 0.295582
R23834 VDD.n3909 VDD 0.295582
R23835 VDD.n4272 VDD 0.295582
R23836 VDD.n4169 VDD 0.295582
R23837 VDD.n4168 VDD 0.295582
R23838 VDD.n4531 VDD 0.295582
R23839 VDD.n4428 VDD 0.295582
R23840 VDD.n4427 VDD 0.295582
R23841 VDD.n163 VDD.n162 0.288543
R23842 VDD.n159 VDD.n158 0.288543
R23843 VDD.n163 VDD 0.252453
R23844 VDD.n159 VDD 0.252453
R23845 VDD.n168 VDD 0.20495
R23846 VDD.n191 VDD 0.161168
R23847 VDD.n334 VDD 0.161168
R23848 VDD.n439 VDD 0.161168
R23849 VDD.n582 VDD 0.161168
R23850 VDD.n698 VDD 0.161168
R23851 VDD.n841 VDD 0.161168
R23852 VDD.n957 VDD 0.161168
R23853 VDD.n1100 VDD 0.161168
R23854 VDD.n1216 VDD 0.161168
R23855 VDD.n1359 VDD 0.161168
R23856 VDD.n1475 VDD 0.161168
R23857 VDD.n1618 VDD 0.161168
R23858 VDD.n1734 VDD 0.161168
R23859 VDD.n1877 VDD 0.161168
R23860 VDD.n1993 VDD 0.161168
R23861 VDD.n2136 VDD 0.161168
R23862 VDD.n2252 VDD 0.161168
R23863 VDD.n2395 VDD 0.161168
R23864 VDD.n2511 VDD 0.161168
R23865 VDD.n2654 VDD 0.161168
R23866 VDD.n2770 VDD 0.161168
R23867 VDD.n2913 VDD 0.161168
R23868 VDD.n3029 VDD 0.161168
R23869 VDD.n3172 VDD 0.161168
R23870 VDD.n3288 VDD 0.161168
R23871 VDD.n3431 VDD 0.161168
R23872 VDD.n3547 VDD 0.161168
R23873 VDD.n3690 VDD 0.161168
R23874 VDD.n3806 VDD 0.161168
R23875 VDD.n3949 VDD 0.161168
R23876 VDD.n4065 VDD 0.161168
R23877 VDD.n4208 VDD 0.161168
R23878 VDD.n4324 VDD 0.161168
R23879 VDD.n4467 VDD 0.161168
R23880 VDD.n4301 VDD.n4300 0.149333
R23881 VDD.n4042 VDD.n4041 0.149333
R23882 VDD.n3783 VDD.n3782 0.149333
R23883 VDD.n3524 VDD.n3523 0.149333
R23884 VDD.n3265 VDD.n3264 0.149333
R23885 VDD.n3006 VDD.n3005 0.149333
R23886 VDD.n2747 VDD.n2746 0.149333
R23887 VDD.n2488 VDD.n2487 0.149333
R23888 VDD.n2229 VDD.n2228 0.149333
R23889 VDD.n1970 VDD.n1969 0.149333
R23890 VDD.n1711 VDD.n1710 0.149333
R23891 VDD.n1452 VDD.n1451 0.149333
R23892 VDD.n1193 VDD.n1192 0.149333
R23893 VDD.n934 VDD.n933 0.149333
R23894 VDD.n675 VDD.n674 0.149333
R23895 VDD.n416 VDD.n415 0.149333
R23896 VDD.n411 VDD.n410 0.149333
R23897 VDD.n410 VDD 0.139364
R23898 VDD.n386 VDD 0.112522
R23899 VDD.n311 VDD 0.112522
R23900 VDD.n350 VDD 0.112522
R23901 VDD.n278 VDD 0.112522
R23902 VDD.n634 VDD 0.112522
R23903 VDD.n559 VDD 0.112522
R23904 VDD.n598 VDD 0.112522
R23905 VDD.n526 VDD 0.112522
R23906 VDD.n893 VDD 0.112522
R23907 VDD.n818 VDD 0.112522
R23908 VDD.n857 VDD 0.112522
R23909 VDD.n785 VDD 0.112522
R23910 VDD.n1152 VDD 0.112522
R23911 VDD.n1077 VDD 0.112522
R23912 VDD.n1116 VDD 0.112522
R23913 VDD.n1044 VDD 0.112522
R23914 VDD.n1411 VDD 0.112522
R23915 VDD.n1336 VDD 0.112522
R23916 VDD.n1375 VDD 0.112522
R23917 VDD.n1303 VDD 0.112522
R23918 VDD.n1670 VDD 0.112522
R23919 VDD.n1595 VDD 0.112522
R23920 VDD.n1634 VDD 0.112522
R23921 VDD.n1562 VDD 0.112522
R23922 VDD.n1929 VDD 0.112522
R23923 VDD.n1854 VDD 0.112522
R23924 VDD.n1893 VDD 0.112522
R23925 VDD.n1821 VDD 0.112522
R23926 VDD.n2188 VDD 0.112522
R23927 VDD.n2113 VDD 0.112522
R23928 VDD.n2152 VDD 0.112522
R23929 VDD.n2080 VDD 0.112522
R23930 VDD.n2447 VDD 0.112522
R23931 VDD.n2372 VDD 0.112522
R23932 VDD.n2411 VDD 0.112522
R23933 VDD.n2339 VDD 0.112522
R23934 VDD.n2706 VDD 0.112522
R23935 VDD.n2631 VDD 0.112522
R23936 VDD.n2670 VDD 0.112522
R23937 VDD.n2598 VDD 0.112522
R23938 VDD.n2965 VDD 0.112522
R23939 VDD.n2890 VDD 0.112522
R23940 VDD.n2929 VDD 0.112522
R23941 VDD.n2857 VDD 0.112522
R23942 VDD.n3224 VDD 0.112522
R23943 VDD.n3149 VDD 0.112522
R23944 VDD.n3188 VDD 0.112522
R23945 VDD.n3116 VDD 0.112522
R23946 VDD.n3483 VDD 0.112522
R23947 VDD.n3408 VDD 0.112522
R23948 VDD.n3447 VDD 0.112522
R23949 VDD.n3375 VDD 0.112522
R23950 VDD.n3742 VDD 0.112522
R23951 VDD.n3667 VDD 0.112522
R23952 VDD.n3706 VDD 0.112522
R23953 VDD.n3634 VDD 0.112522
R23954 VDD.n4001 VDD 0.112522
R23955 VDD.n3926 VDD 0.112522
R23956 VDD.n3965 VDD 0.112522
R23957 VDD.n3893 VDD 0.112522
R23958 VDD.n4260 VDD 0.112522
R23959 VDD.n4185 VDD 0.112522
R23960 VDD.n4224 VDD 0.112522
R23961 VDD.n4152 VDD 0.112522
R23962 VDD.n4519 VDD 0.112522
R23963 VDD.n4444 VDD 0.112522
R23964 VDD.n4483 VDD 0.112522
R23965 VDD.n4411 VDD 0.112522
R23966 VDD.t42 VDD.n7301 0.086419
R23967 VDD.n162 VDD 0.063
R23968 VDD.n164 VDD.n161 0.063
R23969 VDD.n164 VDD.n163 0.063
R23970 VDD.n158 VDD 0.063
R23971 VDD.n160 VDD.n157 0.063
R23972 VDD.n160 VDD.n159 0.063
R23973 VDD.n408 VDD.n169 0.063
R23974 VDD.n408 VDD.n407 0.063
R23975 VDD.n412 VDD 0.063
R23976 VDD.n153 VDD 0.063
R23977 VDD.n656 VDD.n417 0.063
R23978 VDD.n656 VDD.n655 0.063
R23979 VDD.n665 VDD 0.063
R23980 VDD.n667 VDD.n664 0.063
R23981 VDD.n667 VDD.n666 0.063
R23982 VDD.n661 VDD 0.063
R23983 VDD.n663 VDD.n660 0.063
R23984 VDD.n663 VDD.n662 0.063
R23985 VDD.n672 VDD 0.063
R23986 VDD.n915 VDD.n676 0.063
R23987 VDD.n915 VDD.n914 0.063
R23988 VDD.n924 VDD 0.063
R23989 VDD.n926 VDD.n923 0.063
R23990 VDD.n926 VDD.n925 0.063
R23991 VDD.n920 VDD 0.063
R23992 VDD.n922 VDD.n919 0.063
R23993 VDD.n922 VDD.n921 0.063
R23994 VDD.n931 VDD 0.063
R23995 VDD.n1174 VDD.n935 0.063
R23996 VDD.n1174 VDD.n1173 0.063
R23997 VDD.n1183 VDD 0.063
R23998 VDD.n1185 VDD.n1182 0.063
R23999 VDD.n1185 VDD.n1184 0.063
R24000 VDD.n1179 VDD 0.063
R24001 VDD.n1181 VDD.n1178 0.063
R24002 VDD.n1181 VDD.n1180 0.063
R24003 VDD.n1190 VDD 0.063
R24004 VDD.n1433 VDD.n1194 0.063
R24005 VDD.n1433 VDD.n1432 0.063
R24006 VDD.n1442 VDD 0.063
R24007 VDD.n1444 VDD.n1441 0.063
R24008 VDD.n1444 VDD.n1443 0.063
R24009 VDD.n1438 VDD 0.063
R24010 VDD.n1440 VDD.n1437 0.063
R24011 VDD.n1440 VDD.n1439 0.063
R24012 VDD.n1449 VDD 0.063
R24013 VDD.n1692 VDD.n1453 0.063
R24014 VDD.n1692 VDD.n1691 0.063
R24015 VDD.n1701 VDD 0.063
R24016 VDD.n1703 VDD.n1700 0.063
R24017 VDD.n1703 VDD.n1702 0.063
R24018 VDD.n1697 VDD 0.063
R24019 VDD.n1699 VDD.n1696 0.063
R24020 VDD.n1699 VDD.n1698 0.063
R24021 VDD.n1708 VDD 0.063
R24022 VDD.n1951 VDD.n1712 0.063
R24023 VDD.n1951 VDD.n1950 0.063
R24024 VDD.n1960 VDD 0.063
R24025 VDD.n1962 VDD.n1959 0.063
R24026 VDD.n1962 VDD.n1961 0.063
R24027 VDD.n1956 VDD 0.063
R24028 VDD.n1958 VDD.n1955 0.063
R24029 VDD.n1958 VDD.n1957 0.063
R24030 VDD.n1967 VDD 0.063
R24031 VDD.n2210 VDD.n1971 0.063
R24032 VDD.n2210 VDD.n2209 0.063
R24033 VDD.n2219 VDD 0.063
R24034 VDD.n2221 VDD.n2218 0.063
R24035 VDD.n2221 VDD.n2220 0.063
R24036 VDD.n2215 VDD 0.063
R24037 VDD.n2217 VDD.n2214 0.063
R24038 VDD.n2217 VDD.n2216 0.063
R24039 VDD.n2226 VDD 0.063
R24040 VDD.n2469 VDD.n2230 0.063
R24041 VDD.n2469 VDD.n2468 0.063
R24042 VDD.n2478 VDD 0.063
R24043 VDD.n2480 VDD.n2477 0.063
R24044 VDD.n2480 VDD.n2479 0.063
R24045 VDD.n2474 VDD 0.063
R24046 VDD.n2476 VDD.n2473 0.063
R24047 VDD.n2476 VDD.n2475 0.063
R24048 VDD.n2485 VDD 0.063
R24049 VDD.n2728 VDD.n2489 0.063
R24050 VDD.n2728 VDD.n2727 0.063
R24051 VDD.n2737 VDD 0.063
R24052 VDD.n2739 VDD.n2736 0.063
R24053 VDD.n2739 VDD.n2738 0.063
R24054 VDD.n2733 VDD 0.063
R24055 VDD.n2735 VDD.n2732 0.063
R24056 VDD.n2735 VDD.n2734 0.063
R24057 VDD.n2744 VDD 0.063
R24058 VDD.n2987 VDD.n2748 0.063
R24059 VDD.n2987 VDD.n2986 0.063
R24060 VDD.n2996 VDD 0.063
R24061 VDD.n2998 VDD.n2995 0.063
R24062 VDD.n2998 VDD.n2997 0.063
R24063 VDD.n2992 VDD 0.063
R24064 VDD.n2994 VDD.n2991 0.063
R24065 VDD.n2994 VDD.n2993 0.063
R24066 VDD.n3003 VDD 0.063
R24067 VDD.n3246 VDD.n3007 0.063
R24068 VDD.n3246 VDD.n3245 0.063
R24069 VDD.n3255 VDD 0.063
R24070 VDD.n3257 VDD.n3254 0.063
R24071 VDD.n3257 VDD.n3256 0.063
R24072 VDD.n3251 VDD 0.063
R24073 VDD.n3253 VDD.n3250 0.063
R24074 VDD.n3253 VDD.n3252 0.063
R24075 VDD.n3262 VDD 0.063
R24076 VDD.n3505 VDD.n3266 0.063
R24077 VDD.n3505 VDD.n3504 0.063
R24078 VDD.n3514 VDD 0.063
R24079 VDD.n3516 VDD.n3513 0.063
R24080 VDD.n3516 VDD.n3515 0.063
R24081 VDD.n3510 VDD 0.063
R24082 VDD.n3512 VDD.n3509 0.063
R24083 VDD.n3512 VDD.n3511 0.063
R24084 VDD.n3521 VDD 0.063
R24085 VDD.n3764 VDD.n3525 0.063
R24086 VDD.n3764 VDD.n3763 0.063
R24087 VDD.n3773 VDD 0.063
R24088 VDD.n3775 VDD.n3772 0.063
R24089 VDD.n3775 VDD.n3774 0.063
R24090 VDD.n3769 VDD 0.063
R24091 VDD.n3771 VDD.n3768 0.063
R24092 VDD.n3771 VDD.n3770 0.063
R24093 VDD.n3780 VDD 0.063
R24094 VDD.n4023 VDD.n3784 0.063
R24095 VDD.n4023 VDD.n4022 0.063
R24096 VDD.n4032 VDD 0.063
R24097 VDD.n4034 VDD.n4031 0.063
R24098 VDD.n4034 VDD.n4033 0.063
R24099 VDD.n4028 VDD 0.063
R24100 VDD.n4030 VDD.n4027 0.063
R24101 VDD.n4030 VDD.n4029 0.063
R24102 VDD.n4039 VDD 0.063
R24103 VDD.n4282 VDD.n4043 0.063
R24104 VDD.n4282 VDD.n4281 0.063
R24105 VDD.n4291 VDD 0.063
R24106 VDD.n4293 VDD.n4290 0.063
R24107 VDD.n4293 VDD.n4292 0.063
R24108 VDD.n4287 VDD 0.063
R24109 VDD.n4289 VDD.n4286 0.063
R24110 VDD.n4289 VDD.n4288 0.063
R24111 VDD.n4298 VDD 0.063
R24112 VDD.n4541 VDD.n4302 0.063
R24113 VDD.n4541 VDD.n4540 0.063
R24114 VDD.n4550 VDD 0.063
R24115 VDD.n4552 VDD.n4549 0.063
R24116 VDD.n4552 VDD.n4551 0.063
R24117 VDD.n4546 VDD 0.063
R24118 VDD.n4548 VDD.n4545 0.063
R24119 VDD.n4548 VDD.n4547 0.063
R24120 VDD.n18 VDD.n14 0.063
R24121 VDD.n19 VDD.n18 0.063
R24122 VDD.n37 VDD.n33 0.063
R24123 VDD.n38 VDD.n37 0.063
R24124 VDD.n56 VDD.n52 0.063
R24125 VDD.n57 VDD.n56 0.063
R24126 VDD.n75 VDD.n71 0.063
R24127 VDD.n76 VDD.n75 0.063
R24128 VDD.n94 VDD.n90 0.063
R24129 VDD.n95 VDD.n94 0.063
R24130 VDD.n113 VDD.n109 0.063
R24131 VDD.n114 VDD.n113 0.063
R24132 VDD.n132 VDD.n128 0.063
R24133 VDD.n133 VDD.n132 0.063
R24134 VDD.n151 VDD.n147 0.063
R24135 VDD.n152 VDD.n151 0.063
R24136 VDD.n156 VDD.n155 0.0475
R24137 VDD.n154 VDD.n0 0.0475
R24138 VDD.n150 VDD.n149 0.024
R24139 VDD.n131 VDD.n130 0.024
R24140 VDD.n112 VDD.n111 0.024
R24141 VDD.n93 VDD.n92 0.024
R24142 VDD.n74 VDD.n73 0.024
R24143 VDD.n55 VDD.n54 0.024
R24144 VDD.n36 VDD.n35 0.024
R24145 VDD.n17 VDD.n16 0.024
R24146 VDD.n4542 VDD.n4301 0.024
R24147 VDD.n4543 VDD.n4542 0.024
R24148 VDD.n4299 VDD.n4297 0.024
R24149 VDD.n4300 VDD.n4299 0.024
R24150 VDD.n4296 VDD.n4295 0.024
R24151 VDD.n4283 VDD.n4042 0.024
R24152 VDD.n4284 VDD.n4283 0.024
R24153 VDD.n4040 VDD.n4038 0.024
R24154 VDD.n4041 VDD.n4040 0.024
R24155 VDD.n4037 VDD.n4036 0.024
R24156 VDD.n4024 VDD.n3783 0.024
R24157 VDD.n4025 VDD.n4024 0.024
R24158 VDD.n3781 VDD.n3779 0.024
R24159 VDD.n3782 VDD.n3781 0.024
R24160 VDD.n3778 VDD.n3777 0.024
R24161 VDD.n3765 VDD.n3524 0.024
R24162 VDD.n3766 VDD.n3765 0.024
R24163 VDD.n3522 VDD.n3520 0.024
R24164 VDD.n3523 VDD.n3522 0.024
R24165 VDD.n3519 VDD.n3518 0.024
R24166 VDD.n3506 VDD.n3265 0.024
R24167 VDD.n3507 VDD.n3506 0.024
R24168 VDD.n3263 VDD.n3261 0.024
R24169 VDD.n3264 VDD.n3263 0.024
R24170 VDD.n3260 VDD.n3259 0.024
R24171 VDD.n3247 VDD.n3006 0.024
R24172 VDD.n3248 VDD.n3247 0.024
R24173 VDD.n3004 VDD.n3002 0.024
R24174 VDD.n3005 VDD.n3004 0.024
R24175 VDD.n3001 VDD.n3000 0.024
R24176 VDD.n2988 VDD.n2747 0.024
R24177 VDD.n2989 VDD.n2988 0.024
R24178 VDD.n2745 VDD.n2743 0.024
R24179 VDD.n2746 VDD.n2745 0.024
R24180 VDD.n2742 VDD.n2741 0.024
R24181 VDD.n2729 VDD.n2488 0.024
R24182 VDD.n2730 VDD.n2729 0.024
R24183 VDD.n2486 VDD.n2484 0.024
R24184 VDD.n2487 VDD.n2486 0.024
R24185 VDD.n2483 VDD.n2482 0.024
R24186 VDD.n2470 VDD.n2229 0.024
R24187 VDD.n2471 VDD.n2470 0.024
R24188 VDD.n2227 VDD.n2225 0.024
R24189 VDD.n2228 VDD.n2227 0.024
R24190 VDD.n2224 VDD.n2223 0.024
R24191 VDD.n2211 VDD.n1970 0.024
R24192 VDD.n2212 VDD.n2211 0.024
R24193 VDD.n1968 VDD.n1966 0.024
R24194 VDD.n1969 VDD.n1968 0.024
R24195 VDD.n1965 VDD.n1964 0.024
R24196 VDD.n1952 VDD.n1711 0.024
R24197 VDD.n1953 VDD.n1952 0.024
R24198 VDD.n1709 VDD.n1707 0.024
R24199 VDD.n1710 VDD.n1709 0.024
R24200 VDD.n1706 VDD.n1705 0.024
R24201 VDD.n1693 VDD.n1452 0.024
R24202 VDD.n1694 VDD.n1693 0.024
R24203 VDD.n1450 VDD.n1448 0.024
R24204 VDD.n1451 VDD.n1450 0.024
R24205 VDD.n1447 VDD.n1446 0.024
R24206 VDD.n1434 VDD.n1193 0.024
R24207 VDD.n1435 VDD.n1434 0.024
R24208 VDD.n1191 VDD.n1189 0.024
R24209 VDD.n1192 VDD.n1191 0.024
R24210 VDD.n1188 VDD.n1187 0.024
R24211 VDD.n1175 VDD.n934 0.024
R24212 VDD.n1176 VDD.n1175 0.024
R24213 VDD.n932 VDD.n930 0.024
R24214 VDD.n933 VDD.n932 0.024
R24215 VDD.n929 VDD.n928 0.024
R24216 VDD.n916 VDD.n675 0.024
R24217 VDD.n917 VDD.n916 0.024
R24218 VDD.n673 VDD.n671 0.024
R24219 VDD.n674 VDD.n673 0.024
R24220 VDD.n670 VDD.n669 0.024
R24221 VDD.n657 VDD.n416 0.024
R24222 VDD.n658 VDD.n657 0.024
R24223 VDD.n409 VDD.n168 0.024
R24224 VDD.n410 VDD.n409 0.024
R24225 VDD.n167 VDD.n166 0.024
R24226 VDD VDD.n4554 0.0218636
R24227 VDD.n4554 VDD 0.0204394
R24228 VDD.n4295 VDD 0.0204394
R24229 VDD.n4036 VDD 0.0204394
R24230 VDD.n3777 VDD 0.0204394
R24231 VDD.n3518 VDD 0.0204394
R24232 VDD.n3259 VDD 0.0204394
R24233 VDD.n3000 VDD 0.0204394
R24234 VDD.n2741 VDD 0.0204394
R24235 VDD.n2482 VDD 0.0204394
R24236 VDD.n2223 VDD 0.0204394
R24237 VDD.n1964 VDD 0.0204394
R24238 VDD.n1705 VDD 0.0204394
R24239 VDD.n1446 VDD 0.0204394
R24240 VDD.n1187 VDD 0.0204394
R24241 VDD.n928 VDD 0.0204394
R24242 VDD.n669 VDD 0.0204394
R24243 VDD.n335 VDD.n334 0.0152815
R24244 VDD.n583 VDD.n582 0.0152815
R24245 VDD.n842 VDD.n841 0.0152815
R24246 VDD.n1101 VDD.n1100 0.0152815
R24247 VDD.n1360 VDD.n1359 0.0152815
R24248 VDD.n1619 VDD.n1618 0.0152815
R24249 VDD.n1878 VDD.n1877 0.0152815
R24250 VDD.n2137 VDD.n2136 0.0152815
R24251 VDD.n2396 VDD.n2395 0.0152815
R24252 VDD.n2655 VDD.n2654 0.0152815
R24253 VDD.n2914 VDD.n2913 0.0152815
R24254 VDD.n3173 VDD.n3172 0.0152815
R24255 VDD.n3432 VDD.n3431 0.0152815
R24256 VDD.n3691 VDD.n3690 0.0152815
R24257 VDD.n3950 VDD.n3949 0.0152815
R24258 VDD.n4209 VDD.n4208 0.0152815
R24259 VDD.n4468 VDD.n4467 0.0152815
R24260 VDD.n399 VDD.n398 0.00835519
R24261 VDD.n386 VDD.n385 0.00835519
R24262 VDD.n296 VDD.n295 0.00835519
R24263 VDD.n312 VDD.n311 0.00835519
R24264 VDD.n351 VDD.n350 0.00835519
R24265 VDD.n294 VDD.n293 0.00835519
R24266 VDD.n278 VDD.n170 0.00835519
R24267 VDD.n647 VDD.n646 0.00835519
R24268 VDD.n634 VDD.n633 0.00835519
R24269 VDD.n544 VDD.n543 0.00835519
R24270 VDD.n560 VDD.n559 0.00835519
R24271 VDD.n599 VDD.n598 0.00835519
R24272 VDD.n542 VDD.n541 0.00835519
R24273 VDD.n526 VDD.n418 0.00835519
R24274 VDD.n906 VDD.n905 0.00835519
R24275 VDD.n893 VDD.n892 0.00835519
R24276 VDD.n803 VDD.n802 0.00835519
R24277 VDD.n819 VDD.n818 0.00835519
R24278 VDD.n858 VDD.n857 0.00835519
R24279 VDD.n801 VDD.n800 0.00835519
R24280 VDD.n785 VDD.n677 0.00835519
R24281 VDD.n1165 VDD.n1164 0.00835519
R24282 VDD.n1152 VDD.n1151 0.00835519
R24283 VDD.n1062 VDD.n1061 0.00835519
R24284 VDD.n1078 VDD.n1077 0.00835519
R24285 VDD.n1117 VDD.n1116 0.00835519
R24286 VDD.n1060 VDD.n1059 0.00835519
R24287 VDD.n1044 VDD.n936 0.00835519
R24288 VDD.n1424 VDD.n1423 0.00835519
R24289 VDD.n1411 VDD.n1410 0.00835519
R24290 VDD.n1321 VDD.n1320 0.00835519
R24291 VDD.n1337 VDD.n1336 0.00835519
R24292 VDD.n1376 VDD.n1375 0.00835519
R24293 VDD.n1319 VDD.n1318 0.00835519
R24294 VDD.n1303 VDD.n1195 0.00835519
R24295 VDD.n1683 VDD.n1682 0.00835519
R24296 VDD.n1670 VDD.n1669 0.00835519
R24297 VDD.n1580 VDD.n1579 0.00835519
R24298 VDD.n1596 VDD.n1595 0.00835519
R24299 VDD.n1635 VDD.n1634 0.00835519
R24300 VDD.n1578 VDD.n1577 0.00835519
R24301 VDD.n1562 VDD.n1454 0.00835519
R24302 VDD.n1942 VDD.n1941 0.00835519
R24303 VDD.n1929 VDD.n1928 0.00835519
R24304 VDD.n1839 VDD.n1838 0.00835519
R24305 VDD.n1855 VDD.n1854 0.00835519
R24306 VDD.n1894 VDD.n1893 0.00835519
R24307 VDD.n1837 VDD.n1836 0.00835519
R24308 VDD.n1821 VDD.n1713 0.00835519
R24309 VDD.n2201 VDD.n2200 0.00835519
R24310 VDD.n2188 VDD.n2187 0.00835519
R24311 VDD.n2098 VDD.n2097 0.00835519
R24312 VDD.n2114 VDD.n2113 0.00835519
R24313 VDD.n2153 VDD.n2152 0.00835519
R24314 VDD.n2096 VDD.n2095 0.00835519
R24315 VDD.n2080 VDD.n1972 0.00835519
R24316 VDD.n2460 VDD.n2459 0.00835519
R24317 VDD.n2447 VDD.n2446 0.00835519
R24318 VDD.n2357 VDD.n2356 0.00835519
R24319 VDD.n2373 VDD.n2372 0.00835519
R24320 VDD.n2412 VDD.n2411 0.00835519
R24321 VDD.n2355 VDD.n2354 0.00835519
R24322 VDD.n2339 VDD.n2231 0.00835519
R24323 VDD.n2719 VDD.n2718 0.00835519
R24324 VDD.n2706 VDD.n2705 0.00835519
R24325 VDD.n2616 VDD.n2615 0.00835519
R24326 VDD.n2632 VDD.n2631 0.00835519
R24327 VDD.n2671 VDD.n2670 0.00835519
R24328 VDD.n2614 VDD.n2613 0.00835519
R24329 VDD.n2598 VDD.n2490 0.00835519
R24330 VDD.n2978 VDD.n2977 0.00835519
R24331 VDD.n2965 VDD.n2964 0.00835519
R24332 VDD.n2875 VDD.n2874 0.00835519
R24333 VDD.n2891 VDD.n2890 0.00835519
R24334 VDD.n2930 VDD.n2929 0.00835519
R24335 VDD.n2873 VDD.n2872 0.00835519
R24336 VDD.n2857 VDD.n2749 0.00835519
R24337 VDD.n3237 VDD.n3236 0.00835519
R24338 VDD.n3224 VDD.n3223 0.00835519
R24339 VDD.n3134 VDD.n3133 0.00835519
R24340 VDD.n3150 VDD.n3149 0.00835519
R24341 VDD.n3189 VDD.n3188 0.00835519
R24342 VDD.n3132 VDD.n3131 0.00835519
R24343 VDD.n3116 VDD.n3008 0.00835519
R24344 VDD.n3496 VDD.n3495 0.00835519
R24345 VDD.n3483 VDD.n3482 0.00835519
R24346 VDD.n3393 VDD.n3392 0.00835519
R24347 VDD.n3409 VDD.n3408 0.00835519
R24348 VDD.n3448 VDD.n3447 0.00835519
R24349 VDD.n3391 VDD.n3390 0.00835519
R24350 VDD.n3375 VDD.n3267 0.00835519
R24351 VDD.n3755 VDD.n3754 0.00835519
R24352 VDD.n3742 VDD.n3741 0.00835519
R24353 VDD.n3652 VDD.n3651 0.00835519
R24354 VDD.n3668 VDD.n3667 0.00835519
R24355 VDD.n3707 VDD.n3706 0.00835519
R24356 VDD.n3650 VDD.n3649 0.00835519
R24357 VDD.n3634 VDD.n3526 0.00835519
R24358 VDD.n4014 VDD.n4013 0.00835519
R24359 VDD.n4001 VDD.n4000 0.00835519
R24360 VDD.n3911 VDD.n3910 0.00835519
R24361 VDD.n3927 VDD.n3926 0.00835519
R24362 VDD.n3966 VDD.n3965 0.00835519
R24363 VDD.n3909 VDD.n3908 0.00835519
R24364 VDD.n3893 VDD.n3785 0.00835519
R24365 VDD.n4273 VDD.n4272 0.00835519
R24366 VDD.n4260 VDD.n4259 0.00835519
R24367 VDD.n4170 VDD.n4169 0.00835519
R24368 VDD.n4186 VDD.n4185 0.00835519
R24369 VDD.n4225 VDD.n4224 0.00835519
R24370 VDD.n4168 VDD.n4167 0.00835519
R24371 VDD.n4152 VDD.n4044 0.00835519
R24372 VDD.n4532 VDD.n4531 0.00835519
R24373 VDD.n4519 VDD.n4518 0.00835519
R24374 VDD.n4429 VDD.n4428 0.00835519
R24375 VDD.n4445 VDD.n4444 0.00835519
R24376 VDD.n4484 VDD.n4483 0.00835519
R24377 VDD.n4427 VDD.n4426 0.00835519
R24378 VDD.n4411 VDD.n4303 0.00835519
R24379 VDD.n148 VDD 0.00441667
R24380 VDD.n129 VDD 0.00441667
R24381 VDD.n110 VDD 0.00441667
R24382 VDD.n91 VDD 0.00441667
R24383 VDD.n72 VDD 0.00441667
R24384 VDD.n53 VDD 0.00441667
R24385 VDD.n34 VDD 0.00441667
R24386 VDD.n15 VDD 0.00441667
R24387 VDD.n4544 VDD 0.00441667
R24388 VDD.n4285 VDD 0.00441667
R24389 VDD.n4026 VDD 0.00441667
R24390 VDD.n3767 VDD 0.00441667
R24391 VDD.n3508 VDD 0.00441667
R24392 VDD.n3249 VDD 0.00441667
R24393 VDD.n2990 VDD 0.00441667
R24394 VDD.n2731 VDD 0.00441667
R24395 VDD.n2472 VDD 0.00441667
R24396 VDD.n2213 VDD 0.00441667
R24397 VDD.n1954 VDD 0.00441667
R24398 VDD.n1695 VDD 0.00441667
R24399 VDD.n1436 VDD 0.00441667
R24400 VDD.n1177 VDD 0.00441667
R24401 VDD.n918 VDD 0.00441667
R24402 VDD.n659 VDD 0.00441667
R24403 VDD.n411 VDD 0.00441667
R24404 VDD VDD.n7333 0.00441667
R24405 VDD.n148 VDD 0.00406061
R24406 VDD.n129 VDD 0.00406061
R24407 VDD.n110 VDD 0.00406061
R24408 VDD.n91 VDD 0.00406061
R24409 VDD.n72 VDD 0.00406061
R24410 VDD.n53 VDD 0.00406061
R24411 VDD.n34 VDD 0.00406061
R24412 VDD.n15 VDD 0.00406061
R24413 VDD VDD.n4544 0.00406061
R24414 VDD VDD.n4285 0.00406061
R24415 VDD VDD.n4026 0.00406061
R24416 VDD VDD.n3767 0.00406061
R24417 VDD VDD.n3508 0.00406061
R24418 VDD VDD.n3249 0.00406061
R24419 VDD VDD.n2990 0.00406061
R24420 VDD VDD.n2731 0.00406061
R24421 VDD VDD.n2472 0.00406061
R24422 VDD VDD.n2213 0.00406061
R24423 VDD VDD.n1954 0.00406061
R24424 VDD VDD.n1695 0.00406061
R24425 VDD VDD.n1436 0.00406061
R24426 VDD VDD.n1177 0.00406061
R24427 VDD VDD.n918 0.00406061
R24428 VDD VDD.n659 0.00406061
R24429 VDD VDD.n411 0.00406061
R24430 VDD.n7333 VDD 0.00406061
R24431 VDD.n7331 VDD.n7330 0.00241755
R24432 Ring_Counter_0.D_FlipFlop_15.Qbar.n4 Ring_Counter_0.D_FlipFlop_15.Qbar.t0 169.46
R24433 Ring_Counter_0.D_FlipFlop_15.Qbar.n4 Ring_Counter_0.D_FlipFlop_15.Qbar.t3 167.809
R24434 Ring_Counter_0.D_FlipFlop_15.Qbar.n3 Ring_Counter_0.D_FlipFlop_15.Qbar.t1 167.809
R24435 Ring_Counter_0.D_FlipFlop_15.Qbar.n1 Ring_Counter_0.D_FlipFlop_15.Qbar.t5 158.28
R24436 Ring_Counter_0.D_FlipFlop_15.Qbar.t5 Ring_Counter_0.D_FlipFlop_15.Qbar.n0 150.273
R24437 Ring_Counter_0.D_FlipFlop_15.Qbar.n0 Ring_Counter_0.D_FlipFlop_15.Qbar.t4 74.951
R24438 Ring_Counter_0.D_FlipFlop_15.Qbar.n6 Ring_Counter_0.D_FlipFlop_15.Qbar.t2 60.3943
R24439 Ring_Counter_0.D_FlipFlop_15.Qbar.n5 Ring_Counter_0.D_FlipFlop_15.Qbar.n4 11.4489
R24440 Ring_Counter_0.D_FlipFlop_15.Qbar.n3 Ring_Counter_0.D_FlipFlop_15.Qbar 8.5174
R24441 Ring_Counter_0.D_FlipFlop_15.Qbar.n6 Ring_Counter_0.D_FlipFlop_15.Qbar.n5 1.96917
R24442 Ring_Counter_0.D_FlipFlop_15.Qbar.n2 Ring_Counter_0.D_FlipFlop_15.Qbar.n1 0.42585
R24443 Ring_Counter_0.D_FlipFlop_15.Qbar.n1 Ring_Counter_0.D_FlipFlop_15.Qbar 0.390742
R24444 Ring_Counter_0.D_FlipFlop_15.Qbar.n5 Ring_Counter_0.D_FlipFlop_15.Qbar.n3 0.280391
R24445 Ring_Counter_0.D_FlipFlop_15.Qbar.n0 Ring_Counter_0.D_FlipFlop_15.Qbar 0.063
R24446 Ring_Counter_0.D_FlipFlop_15.Qbar Ring_Counter_0.D_FlipFlop_15.Qbar.n6 0.063
R24447 Ring_Counter_0.D_FlipFlop_15.Qbar.n2 Ring_Counter_0.D_FlipFlop_15.Qbar 0.00441667
R24448 Ring_Counter_0.D_FlipFlop_15.Qbar Ring_Counter_0.D_FlipFlop_15.Qbar.n2 0.00406061
R24449 Nand_Gate_1.A.n19 Nand_Gate_1.A.t0 169.46
R24450 Nand_Gate_1.A.n12 Nand_Gate_1.A.t7 168.391
R24451 Nand_Gate_1.A.n19 Nand_Gate_1.A.t3 167.809
R24452 Nand_Gate_1.A.n18 Nand_Gate_1.A.t1 167.809
R24453 Nand_Gate_1.A.n15 Nand_Gate_1.A.t10 158.565
R24454 Nand_Gate_1.A.t10 Nand_Gate_1.A.n14 151.594
R24455 Nand_Gate_1.A.t7 Nand_Gate_1.A.n2 150.293
R24456 Nand_Gate_1.A.n6 Nand_Gate_1.A.t8 150.273
R24457 Nand_Gate_1.A.n3 Nand_Gate_1.A.t6 150.273
R24458 Nand_Gate_1.A Nand_Gate_1.A.t9 99.8701
R24459 Nand_Gate_1.A.n5 Nand_Gate_1.A.t4 74.163
R24460 Nand_Gate_1.A.t9 Nand_Gate_1.A.n10 74.163
R24461 Nand_Gate_1.A.n14 Nand_Gate_1.A.t11 73.6304
R24462 Nand_Gate_1.A.n0 Nand_Gate_1.A.t5 73.6304
R24463 Nand_Gate_1.A.n21 Nand_Gate_1.A.t2 62.1634
R24464 Nand_Gate_1.A.n9 Nand_Gate_1.A.n8 12.6418
R24465 Nand_Gate_1.A.n20 Nand_Gate_1.A.n19 11.4489
R24466 Nand_Gate_1.A.n18 Nand_Gate_1.A.n17 8.21389
R24467 Nand_Gate_1.A.n13 Nand_Gate_1.A 1.2047
R24468 Nand_Gate_1.A.n2 Nand_Gate_1.A.n1 1.19615
R24469 Nand_Gate_1.A.n12 Nand_Gate_1.A.n11 0.922483
R24470 Nand_Gate_1.A.n5 Nand_Gate_1.A 0.851043
R24471 Nand_Gate_1.A.n10 Nand_Gate_1.A 0.851043
R24472 Nand_Gate_1.A.n7 Nand_Gate_1.A.n6 0.61463
R24473 Nand_Gate_1.A.n4 Nand_Gate_1.A.n3 0.61463
R24474 Nand_Gate_1.A.n7 Nand_Gate_1.A 0.486828
R24475 Nand_Gate_1.A.n4 Nand_Gate_1.A 0.486828
R24476 Nand_Gate_1.A.n2 Nand_Gate_1.A 0.447191
R24477 Nand_Gate_1.A.n17 Nand_Gate_1.A.n16 0.425067
R24478 Nand_Gate_1.A.n13 Nand_Gate_1.A.n12 0.399217
R24479 Nand_Gate_1.A.n17 Nand_Gate_1.A 0.39003
R24480 Nand_Gate_1.A.n20 Nand_Gate_1.A.n18 0.280391
R24481 Nand_Gate_1.A.n21 Nand_Gate_1.A.n20 0.200143
R24482 Nand_Gate_1.A.n1 Nand_Gate_1.A 0.1255
R24483 Nand_Gate_1.A.n14 Nand_Gate_1.A 0.063
R24484 Nand_Gate_1.A.n6 Nand_Gate_1.A 0.063
R24485 Nand_Gate_1.A.n8 Nand_Gate_1.A.n5 0.063
R24486 Nand_Gate_1.A.n8 Nand_Gate_1.A.n7 0.063
R24487 Nand_Gate_1.A.n3 Nand_Gate_1.A 0.063
R24488 Nand_Gate_1.A.n10 Nand_Gate_1.A.n9 0.063
R24489 Nand_Gate_1.A.n9 Nand_Gate_1.A.n4 0.063
R24490 Nand_Gate_1.A Nand_Gate_1.A.n21 0.063
R24491 Nand_Gate_1.A.n15 Nand_Gate_1.A.n13 0.024
R24492 Nand_Gate_1.A Nand_Gate_1.A.n15 0.0204394
R24493 Nand_Gate_1.A.n1 Nand_Gate_1.A.n0 0.0107679
R24494 Nand_Gate_1.A.n0 Nand_Gate_1.A 0.0107679
R24495 Nand_Gate_1.A.n11 Nand_Gate_1.A 0.00441667
R24496 Nand_Gate_1.A.n16 Nand_Gate_1.A 0.00441667
R24497 Nand_Gate_1.A.n11 Nand_Gate_1.A 0.00406061
R24498 Nand_Gate_1.A.n16 Nand_Gate_1.A 0.00406061
R24499 CDAC_v3_0.switch_6.Z.n131 CDAC_v3_0.switch_6.Z.t131 168.075
R24500 CDAC_v3_0.switch_6.Z.n131 CDAC_v3_0.switch_6.Z.t0 168.075
R24501 CDAC_v3_0.switch_6.Z.n0 CDAC_v3_0.switch_6.Z.t2 60.6851
R24502 CDAC_v3_0.switch_6.Z CDAC_v3_0.switch_6.Z.t1 60.6226
R24503 CDAC_v3_0.switch_6.Z.n129 CDAC_v3_0.switch_6.Z.n128 23.3141
R24504 CDAC_v3_0.switch_6.Z.n32 CDAC_v3_0.switch_6.Z.n16 9.88172
R24505 CDAC_v3_0.switch_6.Z.n113 CDAC_v3_0.switch_6.Z.t32 9.74547
R24506 CDAC_v3_0.switch_6.Z.n97 CDAC_v3_0.switch_6.Z.t23 9.74547
R24507 CDAC_v3_0.switch_6.Z.n81 CDAC_v3_0.switch_6.Z.t9 9.74547
R24508 CDAC_v3_0.switch_6.Z.n65 CDAC_v3_0.switch_6.Z.t87 9.74547
R24509 CDAC_v3_0.switch_6.Z.n126 CDAC_v3_0.switch_6.Z.t50 7.2858
R24510 CDAC_v3_0.switch_6.Z.n124 CDAC_v3_0.switch_6.Z.t98 7.2858
R24511 CDAC_v3_0.switch_6.Z.n122 CDAC_v3_0.switch_6.Z.t18 7.2858
R24512 CDAC_v3_0.switch_6.Z.n120 CDAC_v3_0.switch_6.Z.t84 7.2858
R24513 CDAC_v3_0.switch_6.Z.n118 CDAC_v3_0.switch_6.Z.t81 7.2858
R24514 CDAC_v3_0.switch_6.Z.n116 CDAC_v3_0.switch_6.Z.t8 7.2858
R24515 CDAC_v3_0.switch_6.Z.n114 CDAC_v3_0.switch_6.Z.t62 7.2858
R24516 CDAC_v3_0.switch_6.Z.n110 CDAC_v3_0.switch_6.Z.t42 7.2858
R24517 CDAC_v3_0.switch_6.Z.n108 CDAC_v3_0.switch_6.Z.t89 7.2858
R24518 CDAC_v3_0.switch_6.Z.n106 CDAC_v3_0.switch_6.Z.t12 7.2858
R24519 CDAC_v3_0.switch_6.Z.n104 CDAC_v3_0.switch_6.Z.t80 7.2858
R24520 CDAC_v3_0.switch_6.Z.n102 CDAC_v3_0.switch_6.Z.t71 7.2858
R24521 CDAC_v3_0.switch_6.Z.n100 CDAC_v3_0.switch_6.Z.t130 7.2858
R24522 CDAC_v3_0.switch_6.Z.n98 CDAC_v3_0.switch_6.Z.t56 7.2858
R24523 CDAC_v3_0.switch_6.Z.n94 CDAC_v3_0.switch_6.Z.t24 7.2858
R24524 CDAC_v3_0.switch_6.Z.n92 CDAC_v3_0.switch_6.Z.t76 7.2858
R24525 CDAC_v3_0.switch_6.Z.n90 CDAC_v3_0.switch_6.Z.t126 7.2858
R24526 CDAC_v3_0.switch_6.Z.n88 CDAC_v3_0.switch_6.Z.t68 7.2858
R24527 CDAC_v3_0.switch_6.Z.n86 CDAC_v3_0.switch_6.Z.t60 7.2858
R24528 CDAC_v3_0.switch_6.Z.n84 CDAC_v3_0.switch_6.Z.t112 7.2858
R24529 CDAC_v3_0.switch_6.Z.n82 CDAC_v3_0.switch_6.Z.t44 7.2858
R24530 CDAC_v3_0.switch_6.Z.n78 CDAC_v3_0.switch_6.Z.t106 7.2858
R24531 CDAC_v3_0.switch_6.Z.n76 CDAC_v3_0.switch_6.Z.t39 7.2858
R24532 CDAC_v3_0.switch_6.Z.n74 CDAC_v3_0.switch_6.Z.t79 7.2858
R24533 CDAC_v3_0.switch_6.Z.n72 CDAC_v3_0.switch_6.Z.t22 7.2858
R24534 CDAC_v3_0.switch_6.Z.n70 CDAC_v3_0.switch_6.Z.t14 7.2858
R24535 CDAC_v3_0.switch_6.Z.n68 CDAC_v3_0.switch_6.Z.t70 7.2858
R24536 CDAC_v3_0.switch_6.Z.n66 CDAC_v3_0.switch_6.Z.t123 7.2858
R24537 CDAC_v3_0.switch_6.Z.n63 CDAC_v3_0.switch_6.Z.t115 7.28556
R24538 CDAC_v3_0.switch_6.Z.n61 CDAC_v3_0.switch_6.Z.t117 7.28556
R24539 CDAC_v3_0.switch_6.Z.n59 CDAC_v3_0.switch_6.Z.t102 7.28556
R24540 CDAC_v3_0.switch_6.Z.n57 CDAC_v3_0.switch_6.Z.t105 7.28556
R24541 CDAC_v3_0.switch_6.Z.n55 CDAC_v3_0.switch_6.Z.t38 7.28556
R24542 CDAC_v3_0.switch_6.Z.n53 CDAC_v3_0.switch_6.Z.t93 7.28556
R24543 CDAC_v3_0.switch_6.Z.n51 CDAC_v3_0.switch_6.Z.t21 7.28556
R24544 CDAC_v3_0.switch_6.Z.n49 CDAC_v3_0.switch_6.Z.t101 7.28556
R24545 CDAC_v3_0.switch_6.Z.n47 CDAC_v3_0.switch_6.Z.t107 7.28556
R24546 CDAC_v3_0.switch_6.Z.n45 CDAC_v3_0.switch_6.Z.t108 7.28556
R24547 CDAC_v3_0.switch_6.Z.n43 CDAC_v3_0.switch_6.Z.t91 7.28556
R24548 CDAC_v3_0.switch_6.Z.n41 CDAC_v3_0.switch_6.Z.t96 7.28556
R24549 CDAC_v3_0.switch_6.Z.n39 CDAC_v3_0.switch_6.Z.t25 7.28556
R24550 CDAC_v3_0.switch_6.Z.n37 CDAC_v3_0.switch_6.Z.t82 7.28556
R24551 CDAC_v3_0.switch_6.Z.n35 CDAC_v3_0.switch_6.Z.t13 7.28556
R24552 CDAC_v3_0.switch_6.Z.n33 CDAC_v3_0.switch_6.Z.t90 7.28556
R24553 CDAC_v3_0.switch_6.Z.n31 CDAC_v3_0.switch_6.Z.t31 7.28556
R24554 CDAC_v3_0.switch_6.Z.n29 CDAC_v3_0.switch_6.Z.t33 7.28556
R24555 CDAC_v3_0.switch_6.Z.n27 CDAC_v3_0.switch_6.Z.t16 7.28556
R24556 CDAC_v3_0.switch_6.Z.n25 CDAC_v3_0.switch_6.Z.t19 7.28556
R24557 CDAC_v3_0.switch_6.Z.n23 CDAC_v3_0.switch_6.Z.t73 7.28556
R24558 CDAC_v3_0.switch_6.Z.n21 CDAC_v3_0.switch_6.Z.t7 7.28556
R24559 CDAC_v3_0.switch_6.Z.n19 CDAC_v3_0.switch_6.Z.t65 7.28556
R24560 CDAC_v3_0.switch_6.Z.n17 CDAC_v3_0.switch_6.Z.t15 7.28556
R24561 CDAC_v3_0.switch_6.Z.n16 CDAC_v3_0.switch_6.Z.t86 7.28556
R24562 CDAC_v3_0.switch_6.Z.n14 CDAC_v3_0.switch_6.Z.t72 7.28556
R24563 CDAC_v3_0.switch_6.Z.n12 CDAC_v3_0.switch_6.Z.t94 7.28556
R24564 CDAC_v3_0.switch_6.Z.n10 CDAC_v3_0.switch_6.Z.t119 7.28556
R24565 CDAC_v3_0.switch_6.Z.n8 CDAC_v3_0.switch_6.Z.t83 7.28556
R24566 CDAC_v3_0.switch_6.Z.n6 CDAC_v3_0.switch_6.Z.t40 7.28556
R24567 CDAC_v3_0.switch_6.Z.n4 CDAC_v3_0.switch_6.Z.t3 7.28556
R24568 CDAC_v3_0.switch_6.Z.n2 CDAC_v3_0.switch_6.Z.t88 7.28556
R24569 CDAC_v3_0.switch_6.Z.n128 CDAC_v3_0.switch_6.Z.n127 6.08323
R24570 CDAC_v3_0.switch_6.Z.n112 CDAC_v3_0.switch_6.Z.n111 6.08323
R24571 CDAC_v3_0.switch_6.Z.n96 CDAC_v3_0.switch_6.Z.n95 6.08323
R24572 CDAC_v3_0.switch_6.Z.n80 CDAC_v3_0.switch_6.Z.n79 6.08323
R24573 CDAC_v3_0.switch_6.Z.n64 CDAC_v3_0.switch_6.Z.n63 6.07666
R24574 CDAC_v3_0.switch_6.Z.n48 CDAC_v3_0.switch_6.Z.n47 6.07666
R24575 CDAC_v3_0.switch_6.Z.n32 CDAC_v3_0.switch_6.Z.n31 6.07666
R24576 CDAC_v3_0.switch_6.Z.n80 CDAC_v3_0.switch_6.Z.n64 4.09733
R24577 CDAC_v3_0.switch_6.Z.n48 CDAC_v3_0.switch_6.Z.n32 3.80593
R24578 CDAC_v3_0.switch_6.Z.n64 CDAC_v3_0.switch_6.Z.n48 3.80593
R24579 CDAC_v3_0.switch_6.Z.n96 CDAC_v3_0.switch_6.Z.n80 3.80593
R24580 CDAC_v3_0.switch_6.Z.n112 CDAC_v3_0.switch_6.Z.n96 3.80593
R24581 CDAC_v3_0.switch_6.Z.n128 CDAC_v3_0.switch_6.Z.n112 3.80593
R24582 CDAC_v3_0.switch_6.Z.n49 CDAC_v3_0.switch_6.Z.t11 2.76693
R24583 CDAC_v3_0.switch_6.Z.n33 CDAC_v3_0.switch_6.Z.t124 2.76693
R24584 CDAC_v3_0.switch_6.Z.n17 CDAC_v3_0.switch_6.Z.t46 2.76693
R24585 CDAC_v3_0.switch_6.Z.n2 CDAC_v3_0.switch_6.Z.t34 2.76693
R24586 CDAC_v3_0.switch_6.Z.n115 CDAC_v3_0.switch_6.Z.n114 2.46017
R24587 CDAC_v3_0.switch_6.Z.n117 CDAC_v3_0.switch_6.Z.n116 2.46017
R24588 CDAC_v3_0.switch_6.Z.n119 CDAC_v3_0.switch_6.Z.n118 2.46017
R24589 CDAC_v3_0.switch_6.Z.n121 CDAC_v3_0.switch_6.Z.n120 2.46017
R24590 CDAC_v3_0.switch_6.Z.n123 CDAC_v3_0.switch_6.Z.n122 2.46017
R24591 CDAC_v3_0.switch_6.Z.n125 CDAC_v3_0.switch_6.Z.n124 2.46017
R24592 CDAC_v3_0.switch_6.Z.n127 CDAC_v3_0.switch_6.Z.n126 2.46017
R24593 CDAC_v3_0.switch_6.Z.n99 CDAC_v3_0.switch_6.Z.n98 2.46017
R24594 CDAC_v3_0.switch_6.Z.n101 CDAC_v3_0.switch_6.Z.n100 2.46017
R24595 CDAC_v3_0.switch_6.Z.n103 CDAC_v3_0.switch_6.Z.n102 2.46017
R24596 CDAC_v3_0.switch_6.Z.n105 CDAC_v3_0.switch_6.Z.n104 2.46017
R24597 CDAC_v3_0.switch_6.Z.n107 CDAC_v3_0.switch_6.Z.n106 2.46017
R24598 CDAC_v3_0.switch_6.Z.n109 CDAC_v3_0.switch_6.Z.n108 2.46017
R24599 CDAC_v3_0.switch_6.Z.n111 CDAC_v3_0.switch_6.Z.n110 2.46017
R24600 CDAC_v3_0.switch_6.Z.n83 CDAC_v3_0.switch_6.Z.n82 2.46017
R24601 CDAC_v3_0.switch_6.Z.n85 CDAC_v3_0.switch_6.Z.n84 2.46017
R24602 CDAC_v3_0.switch_6.Z.n87 CDAC_v3_0.switch_6.Z.n86 2.46017
R24603 CDAC_v3_0.switch_6.Z.n89 CDAC_v3_0.switch_6.Z.n88 2.46017
R24604 CDAC_v3_0.switch_6.Z.n91 CDAC_v3_0.switch_6.Z.n90 2.46017
R24605 CDAC_v3_0.switch_6.Z.n93 CDAC_v3_0.switch_6.Z.n92 2.46017
R24606 CDAC_v3_0.switch_6.Z.n95 CDAC_v3_0.switch_6.Z.n94 2.46017
R24607 CDAC_v3_0.switch_6.Z.n67 CDAC_v3_0.switch_6.Z.n66 2.46017
R24608 CDAC_v3_0.switch_6.Z.n69 CDAC_v3_0.switch_6.Z.n68 2.46017
R24609 CDAC_v3_0.switch_6.Z.n71 CDAC_v3_0.switch_6.Z.n70 2.46017
R24610 CDAC_v3_0.switch_6.Z.n73 CDAC_v3_0.switch_6.Z.n72 2.46017
R24611 CDAC_v3_0.switch_6.Z.n75 CDAC_v3_0.switch_6.Z.n74 2.46017
R24612 CDAC_v3_0.switch_6.Z.n77 CDAC_v3_0.switch_6.Z.n76 2.46017
R24613 CDAC_v3_0.switch_6.Z.n79 CDAC_v3_0.switch_6.Z.n78 2.46017
R24614 CDAC_v3_0.switch_6.Z.n51 CDAC_v3_0.switch_6.Z.n50 2.45986
R24615 CDAC_v3_0.switch_6.Z.n53 CDAC_v3_0.switch_6.Z.n52 2.45986
R24616 CDAC_v3_0.switch_6.Z.n55 CDAC_v3_0.switch_6.Z.n54 2.45986
R24617 CDAC_v3_0.switch_6.Z.n57 CDAC_v3_0.switch_6.Z.n56 2.45986
R24618 CDAC_v3_0.switch_6.Z.n59 CDAC_v3_0.switch_6.Z.n58 2.45986
R24619 CDAC_v3_0.switch_6.Z.n61 CDAC_v3_0.switch_6.Z.n60 2.45986
R24620 CDAC_v3_0.switch_6.Z.n63 CDAC_v3_0.switch_6.Z.n62 2.45986
R24621 CDAC_v3_0.switch_6.Z.n35 CDAC_v3_0.switch_6.Z.n34 2.45986
R24622 CDAC_v3_0.switch_6.Z.n37 CDAC_v3_0.switch_6.Z.n36 2.45986
R24623 CDAC_v3_0.switch_6.Z.n39 CDAC_v3_0.switch_6.Z.n38 2.45986
R24624 CDAC_v3_0.switch_6.Z.n41 CDAC_v3_0.switch_6.Z.n40 2.45986
R24625 CDAC_v3_0.switch_6.Z.n43 CDAC_v3_0.switch_6.Z.n42 2.45986
R24626 CDAC_v3_0.switch_6.Z.n45 CDAC_v3_0.switch_6.Z.n44 2.45986
R24627 CDAC_v3_0.switch_6.Z.n47 CDAC_v3_0.switch_6.Z.n46 2.45986
R24628 CDAC_v3_0.switch_6.Z.n19 CDAC_v3_0.switch_6.Z.n18 2.45986
R24629 CDAC_v3_0.switch_6.Z.n21 CDAC_v3_0.switch_6.Z.n20 2.45986
R24630 CDAC_v3_0.switch_6.Z.n23 CDAC_v3_0.switch_6.Z.n22 2.45986
R24631 CDAC_v3_0.switch_6.Z.n25 CDAC_v3_0.switch_6.Z.n24 2.45986
R24632 CDAC_v3_0.switch_6.Z.n27 CDAC_v3_0.switch_6.Z.n26 2.45986
R24633 CDAC_v3_0.switch_6.Z.n29 CDAC_v3_0.switch_6.Z.n28 2.45986
R24634 CDAC_v3_0.switch_6.Z.n31 CDAC_v3_0.switch_6.Z.n30 2.45986
R24635 CDAC_v3_0.switch_6.Z.n4 CDAC_v3_0.switch_6.Z.n3 2.45986
R24636 CDAC_v3_0.switch_6.Z.n6 CDAC_v3_0.switch_6.Z.n5 2.45986
R24637 CDAC_v3_0.switch_6.Z.n8 CDAC_v3_0.switch_6.Z.n7 2.45986
R24638 CDAC_v3_0.switch_6.Z.n10 CDAC_v3_0.switch_6.Z.n9 2.45986
R24639 CDAC_v3_0.switch_6.Z.n12 CDAC_v3_0.switch_6.Z.n11 2.45986
R24640 CDAC_v3_0.switch_6.Z.n14 CDAC_v3_0.switch_6.Z.n13 2.45986
R24641 CDAC_v3_0.switch_6.Z.n16 CDAC_v3_0.switch_6.Z.n15 2.45986
R24642 CDAC_v3_0.switch_6.Z.n132 CDAC_v3_0.switch_6.Z.n130 1.34289
R24643 CDAC_v3_0.switch_6.Z.n114 CDAC_v3_0.switch_6.Z.n113 1.33843
R24644 CDAC_v3_0.switch_6.Z.n116 CDAC_v3_0.switch_6.Z.n115 1.33843
R24645 CDAC_v3_0.switch_6.Z.n118 CDAC_v3_0.switch_6.Z.n117 1.33843
R24646 CDAC_v3_0.switch_6.Z.n120 CDAC_v3_0.switch_6.Z.n119 1.33843
R24647 CDAC_v3_0.switch_6.Z.n122 CDAC_v3_0.switch_6.Z.n121 1.33843
R24648 CDAC_v3_0.switch_6.Z.n124 CDAC_v3_0.switch_6.Z.n123 1.33843
R24649 CDAC_v3_0.switch_6.Z.n126 CDAC_v3_0.switch_6.Z.n125 1.33843
R24650 CDAC_v3_0.switch_6.Z.n98 CDAC_v3_0.switch_6.Z.n97 1.33843
R24651 CDAC_v3_0.switch_6.Z.n100 CDAC_v3_0.switch_6.Z.n99 1.33843
R24652 CDAC_v3_0.switch_6.Z.n102 CDAC_v3_0.switch_6.Z.n101 1.33843
R24653 CDAC_v3_0.switch_6.Z.n104 CDAC_v3_0.switch_6.Z.n103 1.33843
R24654 CDAC_v3_0.switch_6.Z.n106 CDAC_v3_0.switch_6.Z.n105 1.33843
R24655 CDAC_v3_0.switch_6.Z.n108 CDAC_v3_0.switch_6.Z.n107 1.33843
R24656 CDAC_v3_0.switch_6.Z.n110 CDAC_v3_0.switch_6.Z.n109 1.33843
R24657 CDAC_v3_0.switch_6.Z.n82 CDAC_v3_0.switch_6.Z.n81 1.33843
R24658 CDAC_v3_0.switch_6.Z.n84 CDAC_v3_0.switch_6.Z.n83 1.33843
R24659 CDAC_v3_0.switch_6.Z.n86 CDAC_v3_0.switch_6.Z.n85 1.33843
R24660 CDAC_v3_0.switch_6.Z.n88 CDAC_v3_0.switch_6.Z.n87 1.33843
R24661 CDAC_v3_0.switch_6.Z.n90 CDAC_v3_0.switch_6.Z.n89 1.33843
R24662 CDAC_v3_0.switch_6.Z.n92 CDAC_v3_0.switch_6.Z.n91 1.33843
R24663 CDAC_v3_0.switch_6.Z.n94 CDAC_v3_0.switch_6.Z.n93 1.33843
R24664 CDAC_v3_0.switch_6.Z.n66 CDAC_v3_0.switch_6.Z.n65 1.33843
R24665 CDAC_v3_0.switch_6.Z.n68 CDAC_v3_0.switch_6.Z.n67 1.33843
R24666 CDAC_v3_0.switch_6.Z.n70 CDAC_v3_0.switch_6.Z.n69 1.33843
R24667 CDAC_v3_0.switch_6.Z.n72 CDAC_v3_0.switch_6.Z.n71 1.33843
R24668 CDAC_v3_0.switch_6.Z.n74 CDAC_v3_0.switch_6.Z.n73 1.33843
R24669 CDAC_v3_0.switch_6.Z.n76 CDAC_v3_0.switch_6.Z.n75 1.33843
R24670 CDAC_v3_0.switch_6.Z.n78 CDAC_v3_0.switch_6.Z.n77 1.33843
R24671 CDAC_v3_0.switch_6.Z.n50 CDAC_v3_0.switch_6.Z.n49 1.33813
R24672 CDAC_v3_0.switch_6.Z.n52 CDAC_v3_0.switch_6.Z.n51 1.33813
R24673 CDAC_v3_0.switch_6.Z.n54 CDAC_v3_0.switch_6.Z.n53 1.33813
R24674 CDAC_v3_0.switch_6.Z.n56 CDAC_v3_0.switch_6.Z.n55 1.33813
R24675 CDAC_v3_0.switch_6.Z.n58 CDAC_v3_0.switch_6.Z.n57 1.33813
R24676 CDAC_v3_0.switch_6.Z.n60 CDAC_v3_0.switch_6.Z.n59 1.33813
R24677 CDAC_v3_0.switch_6.Z.n62 CDAC_v3_0.switch_6.Z.n61 1.33813
R24678 CDAC_v3_0.switch_6.Z.n34 CDAC_v3_0.switch_6.Z.n33 1.33813
R24679 CDAC_v3_0.switch_6.Z.n36 CDAC_v3_0.switch_6.Z.n35 1.33813
R24680 CDAC_v3_0.switch_6.Z.n38 CDAC_v3_0.switch_6.Z.n37 1.33813
R24681 CDAC_v3_0.switch_6.Z.n40 CDAC_v3_0.switch_6.Z.n39 1.33813
R24682 CDAC_v3_0.switch_6.Z.n42 CDAC_v3_0.switch_6.Z.n41 1.33813
R24683 CDAC_v3_0.switch_6.Z.n44 CDAC_v3_0.switch_6.Z.n43 1.33813
R24684 CDAC_v3_0.switch_6.Z.n46 CDAC_v3_0.switch_6.Z.n45 1.33813
R24685 CDAC_v3_0.switch_6.Z.n18 CDAC_v3_0.switch_6.Z.n17 1.33813
R24686 CDAC_v3_0.switch_6.Z.n20 CDAC_v3_0.switch_6.Z.n19 1.33813
R24687 CDAC_v3_0.switch_6.Z.n22 CDAC_v3_0.switch_6.Z.n21 1.33813
R24688 CDAC_v3_0.switch_6.Z.n24 CDAC_v3_0.switch_6.Z.n23 1.33813
R24689 CDAC_v3_0.switch_6.Z.n26 CDAC_v3_0.switch_6.Z.n25 1.33813
R24690 CDAC_v3_0.switch_6.Z.n28 CDAC_v3_0.switch_6.Z.n27 1.33813
R24691 CDAC_v3_0.switch_6.Z.n30 CDAC_v3_0.switch_6.Z.n29 1.33813
R24692 CDAC_v3_0.switch_6.Z.n3 CDAC_v3_0.switch_6.Z.n2 1.33813
R24693 CDAC_v3_0.switch_6.Z.n5 CDAC_v3_0.switch_6.Z.n4 1.33813
R24694 CDAC_v3_0.switch_6.Z.n7 CDAC_v3_0.switch_6.Z.n6 1.33813
R24695 CDAC_v3_0.switch_6.Z.n9 CDAC_v3_0.switch_6.Z.n8 1.33813
R24696 CDAC_v3_0.switch_6.Z.n11 CDAC_v3_0.switch_6.Z.n10 1.33813
R24697 CDAC_v3_0.switch_6.Z.n13 CDAC_v3_0.switch_6.Z.n12 1.33813
R24698 CDAC_v3_0.switch_6.Z.n15 CDAC_v3_0.switch_6.Z.n14 1.33813
R24699 CDAC_v3_0.switch_6.Z.n130 CDAC_v3_0.switch_6.Z 0.42713
R24700 CDAC_v3_0.switch_6.Z.n113 CDAC_v3_0.switch_6.Z.t36 0.307567
R24701 CDAC_v3_0.switch_6.Z.n115 CDAC_v3_0.switch_6.Z.t78 0.307567
R24702 CDAC_v3_0.switch_6.Z.n117 CDAC_v3_0.switch_6.Z.t26 0.307567
R24703 CDAC_v3_0.switch_6.Z.n119 CDAC_v3_0.switch_6.Z.t85 0.307567
R24704 CDAC_v3_0.switch_6.Z.n121 CDAC_v3_0.switch_6.Z.t41 0.307567
R24705 CDAC_v3_0.switch_6.Z.n123 CDAC_v3_0.switch_6.Z.t37 0.307567
R24706 CDAC_v3_0.switch_6.Z.n125 CDAC_v3_0.switch_6.Z.t52 0.307567
R24707 CDAC_v3_0.switch_6.Z.n127 CDAC_v3_0.switch_6.Z.t51 0.307567
R24708 CDAC_v3_0.switch_6.Z.n97 CDAC_v3_0.switch_6.Z.t121 0.307567
R24709 CDAC_v3_0.switch_6.Z.n99 CDAC_v3_0.switch_6.Z.t47 0.307567
R24710 CDAC_v3_0.switch_6.Z.n101 CDAC_v3_0.switch_6.Z.t111 0.307567
R24711 CDAC_v3_0.switch_6.Z.n103 CDAC_v3_0.switch_6.Z.t55 0.307567
R24712 CDAC_v3_0.switch_6.Z.n105 CDAC_v3_0.switch_6.Z.t125 0.307567
R24713 CDAC_v3_0.switch_6.Z.n107 CDAC_v3_0.switch_6.Z.t122 0.307567
R24714 CDAC_v3_0.switch_6.Z.n109 CDAC_v3_0.switch_6.Z.t6 0.307567
R24715 CDAC_v3_0.switch_6.Z.n111 CDAC_v3_0.switch_6.Z.t5 0.307567
R24716 CDAC_v3_0.switch_6.Z.n81 CDAC_v3_0.switch_6.Z.t99 0.307567
R24717 CDAC_v3_0.switch_6.Z.n83 CDAC_v3_0.switch_6.Z.t20 0.307567
R24718 CDAC_v3_0.switch_6.Z.n85 CDAC_v3_0.switch_6.Z.t92 0.307567
R24719 CDAC_v3_0.switch_6.Z.n87 CDAC_v3_0.switch_6.Z.t35 0.307567
R24720 CDAC_v3_0.switch_6.Z.n89 CDAC_v3_0.switch_6.Z.t104 0.307567
R24721 CDAC_v3_0.switch_6.Z.n91 CDAC_v3_0.switch_6.Z.t100 0.307567
R24722 CDAC_v3_0.switch_6.Z.n93 CDAC_v3_0.switch_6.Z.t116 0.307567
R24723 CDAC_v3_0.switch_6.Z.n95 CDAC_v3_0.switch_6.Z.t114 0.307567
R24724 CDAC_v3_0.switch_6.Z.n65 CDAC_v3_0.switch_6.Z.t63 0.307567
R24725 CDAC_v3_0.switch_6.Z.n67 CDAC_v3_0.switch_6.Z.t109 0.307567
R24726 CDAC_v3_0.switch_6.Z.n69 CDAC_v3_0.switch_6.Z.t58 0.307567
R24727 CDAC_v3_0.switch_6.Z.n71 CDAC_v3_0.switch_6.Z.t120 0.307567
R24728 CDAC_v3_0.switch_6.Z.n73 CDAC_v3_0.switch_6.Z.t67 0.307567
R24729 CDAC_v3_0.switch_6.Z.n75 CDAC_v3_0.switch_6.Z.t64 0.307567
R24730 CDAC_v3_0.switch_6.Z.n77 CDAC_v3_0.switch_6.Z.t75 0.307567
R24731 CDAC_v3_0.switch_6.Z.n79 CDAC_v3_0.switch_6.Z.t74 0.307567
R24732 CDAC_v3_0.switch_6.Z.n50 CDAC_v3_0.switch_6.Z.t45 0.307567
R24733 CDAC_v3_0.switch_6.Z.n52 CDAC_v3_0.switch_6.Z.t113 0.307567
R24734 CDAC_v3_0.switch_6.Z.n54 CDAC_v3_0.switch_6.Z.t61 0.307567
R24735 CDAC_v3_0.switch_6.Z.n56 CDAC_v3_0.switch_6.Z.t69 0.307567
R24736 CDAC_v3_0.switch_6.Z.n58 CDAC_v3_0.switch_6.Z.t128 0.307567
R24737 CDAC_v3_0.switch_6.Z.n60 CDAC_v3_0.switch_6.Z.t77 0.307567
R24738 CDAC_v3_0.switch_6.Z.n62 CDAC_v3_0.switch_6.Z.t27 0.307567
R24739 CDAC_v3_0.switch_6.Z.n34 CDAC_v3_0.switch_6.Z.t28 0.307567
R24740 CDAC_v3_0.switch_6.Z.n36 CDAC_v3_0.switch_6.Z.t97 0.307567
R24741 CDAC_v3_0.switch_6.Z.n38 CDAC_v3_0.switch_6.Z.t49 0.307567
R24742 CDAC_v3_0.switch_6.Z.n40 CDAC_v3_0.switch_6.Z.t57 0.307567
R24743 CDAC_v3_0.switch_6.Z.n42 CDAC_v3_0.switch_6.Z.t110 0.307567
R24744 CDAC_v3_0.switch_6.Z.n44 CDAC_v3_0.switch_6.Z.t66 0.307567
R24745 CDAC_v3_0.switch_6.Z.n46 CDAC_v3_0.switch_6.Z.t10 0.307567
R24746 CDAC_v3_0.switch_6.Z.n18 CDAC_v3_0.switch_6.Z.t103 0.307567
R24747 CDAC_v3_0.switch_6.Z.n20 CDAC_v3_0.switch_6.Z.t29 0.307567
R24748 CDAC_v3_0.switch_6.Z.n22 CDAC_v3_0.switch_6.Z.t59 0.307567
R24749 CDAC_v3_0.switch_6.Z.n24 CDAC_v3_0.switch_6.Z.t54 0.307567
R24750 CDAC_v3_0.switch_6.Z.n26 CDAC_v3_0.switch_6.Z.t127 0.307567
R24751 CDAC_v3_0.switch_6.Z.n28 CDAC_v3_0.switch_6.Z.t4 0.307567
R24752 CDAC_v3_0.switch_6.Z.n30 CDAC_v3_0.switch_6.Z.t43 0.307567
R24753 CDAC_v3_0.switch_6.Z.n3 CDAC_v3_0.switch_6.Z.t95 0.307567
R24754 CDAC_v3_0.switch_6.Z.n5 CDAC_v3_0.switch_6.Z.t17 0.307567
R24755 CDAC_v3_0.switch_6.Z.n7 CDAC_v3_0.switch_6.Z.t53 0.307567
R24756 CDAC_v3_0.switch_6.Z.n9 CDAC_v3_0.switch_6.Z.t48 0.307567
R24757 CDAC_v3_0.switch_6.Z.n11 CDAC_v3_0.switch_6.Z.t118 0.307567
R24758 CDAC_v3_0.switch_6.Z.n13 CDAC_v3_0.switch_6.Z.t129 0.307567
R24759 CDAC_v3_0.switch_6.Z.n15 CDAC_v3_0.switch_6.Z.t30 0.307567
R24760 CDAC_v3_0.switch_6.Z.n1 CDAC_v3_0.switch_6.Z 0.182141
R24761 CDAC_v3_0.switch_6.Z CDAC_v3_0.switch_6.Z.n132 0.178175
R24762 CDAC_v3_0.switch_6.Z.n1 CDAC_v3_0.switch_6.Z.n0 0.128217
R24763 CDAC_v3_0.switch_6.Z.n0 CDAC_v3_0.switch_6.Z 0.1255
R24764 CDAC_v3_0.switch_6.Z.n0 CDAC_v3_0.switch_6.Z 0.063
R24765 CDAC_v3_0.switch_6.Z.n130 CDAC_v3_0.switch_6.Z.n129 0.063
R24766 CDAC_v3_0.switch_6.Z.n129 CDAC_v3_0.switch_6.Z.n1 0.063
R24767 CDAC_v3_0.switch_6.Z.n132 CDAC_v3_0.switch_6.Z.n131 0.0130546
R24768 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.t2 169.46
R24769 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout.t1 167.809
R24770 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.t0 167.809
R24771 D_FlipFlop_2.3-input-nand_2.Vout.t6 D_FlipFlop_2.3-input-nand_2.Vout.n11 167.227
R24772 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.t6 150.293
R24773 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.t4 150.273
R24774 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout.t7 73.6406
R24775 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout.t5 73.6304
R24776 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout.t3 60.3809
R24777 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout.n5 12.3891
R24778 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout.n9 11.4489
R24779 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout.n2 1.38365
R24780 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.n1 1.19615
R24781 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.n4 1.1717
R24782 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout 0.848156
R24783 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.Vout.n12 0.447191
R24784 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R24785 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout.n10 0.280391
R24786 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout 0.217464
R24787 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout 0.200143
R24788 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R24789 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R24790 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R24791 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R24792 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout.n7 0.0874565
R24793 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout.n3 0.063
R24794 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout.n6 0.063
R24795 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.Vout.n8 0.063
R24796 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R24797 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout.n0 0.0107679
R24798 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout 0.0107679
R24799 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 169.46
R24800 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 167.809
R24801 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 167.809
R24802 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 167.227
R24803 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 151.594
R24804 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 150.273
R24805 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 74.8641
R24806 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 73.6304
R24807 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 61.84
R24808 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 12.3891
R24809 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 11.4489
R24810 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R24811 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 0.280391
R24812 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 0.200143
R24813 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R24814 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R24815 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 0.149957
R24816 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.063
R24817 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 0.063
R24818 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 0.063
R24819 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 0.063
R24820 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R24821 CDAC_v3_0.switch_7.Z.n67 CDAC_v3_0.switch_7.Z.t67 168.075
R24822 CDAC_v3_0.switch_7.Z.n67 CDAC_v3_0.switch_7.Z.t0 168.075
R24823 CDAC_v3_0.switch_7.Z.n0 CDAC_v3_0.switch_7.Z.t66 60.6851
R24824 CDAC_v3_0.switch_7.Z CDAC_v3_0.switch_7.Z.t1 60.6226
R24825 CDAC_v3_0.switch_7.Z.n65 CDAC_v3_0.switch_7.Z.n64 39.6106
R24826 CDAC_v3_0.switch_7.Z.n16 CDAC_v3_0.switch_7.Z.n8 12.3546
R24827 CDAC_v3_0.switch_7.Z.n32 CDAC_v3_0.switch_7.Z.n31 8.54917
R24828 CDAC_v3_0.switch_7.Z.n24 CDAC_v3_0.switch_7.Z.n23 8.54917
R24829 CDAC_v3_0.switch_7.Z.n16 CDAC_v3_0.switch_7.Z.n15 8.54917
R24830 CDAC_v3_0.switch_7.Z.n40 CDAC_v3_0.switch_7.Z.n32 7.61607
R24831 CDAC_v3_0.switch_7.Z.n64 CDAC_v3_0.switch_7.Z.n63 6.08323
R24832 CDAC_v3_0.switch_7.Z.n56 CDAC_v3_0.switch_7.Z.n55 6.08323
R24833 CDAC_v3_0.switch_7.Z.n48 CDAC_v3_0.switch_7.Z.n47 6.08323
R24834 CDAC_v3_0.switch_7.Z.n40 CDAC_v3_0.switch_7.Z.n39 6.08323
R24835 CDAC_v3_0.switch_7.Z.n57 CDAC_v3_0.switch_7.Z.t57 4.1177
R24836 CDAC_v3_0.switch_7.Z.n49 CDAC_v3_0.switch_7.Z.t40 4.1177
R24837 CDAC_v3_0.switch_7.Z.n41 CDAC_v3_0.switch_7.Z.t28 4.1177
R24838 CDAC_v3_0.switch_7.Z.n33 CDAC_v3_0.switch_7.Z.t8 4.1177
R24839 CDAC_v3_0.switch_7.Z.n25 CDAC_v3_0.switch_7.Z.t41 4.1177
R24840 CDAC_v3_0.switch_7.Z.n17 CDAC_v3_0.switch_7.Z.t31 4.1177
R24841 CDAC_v3_0.switch_7.Z.n9 CDAC_v3_0.switch_7.Z.t2 4.1177
R24842 CDAC_v3_0.switch_7.Z.n2 CDAC_v3_0.switch_7.Z.t61 4.1177
R24843 CDAC_v3_0.switch_7.Z.n58 CDAC_v3_0.switch_7.Z.n57 3.81063
R24844 CDAC_v3_0.switch_7.Z.n59 CDAC_v3_0.switch_7.Z.n58 3.81063
R24845 CDAC_v3_0.switch_7.Z.n60 CDAC_v3_0.switch_7.Z.n59 3.81063
R24846 CDAC_v3_0.switch_7.Z.n61 CDAC_v3_0.switch_7.Z.n60 3.81063
R24847 CDAC_v3_0.switch_7.Z.n62 CDAC_v3_0.switch_7.Z.n61 3.81063
R24848 CDAC_v3_0.switch_7.Z.n63 CDAC_v3_0.switch_7.Z.n62 3.81063
R24849 CDAC_v3_0.switch_7.Z.n50 CDAC_v3_0.switch_7.Z.n49 3.81063
R24850 CDAC_v3_0.switch_7.Z.n51 CDAC_v3_0.switch_7.Z.n50 3.81063
R24851 CDAC_v3_0.switch_7.Z.n52 CDAC_v3_0.switch_7.Z.n51 3.81063
R24852 CDAC_v3_0.switch_7.Z.n53 CDAC_v3_0.switch_7.Z.n52 3.81063
R24853 CDAC_v3_0.switch_7.Z.n54 CDAC_v3_0.switch_7.Z.n53 3.81063
R24854 CDAC_v3_0.switch_7.Z.n55 CDAC_v3_0.switch_7.Z.n54 3.81063
R24855 CDAC_v3_0.switch_7.Z.n42 CDAC_v3_0.switch_7.Z.n41 3.81063
R24856 CDAC_v3_0.switch_7.Z.n43 CDAC_v3_0.switch_7.Z.n42 3.81063
R24857 CDAC_v3_0.switch_7.Z.n44 CDAC_v3_0.switch_7.Z.n43 3.81063
R24858 CDAC_v3_0.switch_7.Z.n45 CDAC_v3_0.switch_7.Z.n44 3.81063
R24859 CDAC_v3_0.switch_7.Z.n46 CDAC_v3_0.switch_7.Z.n45 3.81063
R24860 CDAC_v3_0.switch_7.Z.n47 CDAC_v3_0.switch_7.Z.n46 3.81063
R24861 CDAC_v3_0.switch_7.Z.n34 CDAC_v3_0.switch_7.Z.n33 3.81063
R24862 CDAC_v3_0.switch_7.Z.n35 CDAC_v3_0.switch_7.Z.n34 3.81063
R24863 CDAC_v3_0.switch_7.Z.n36 CDAC_v3_0.switch_7.Z.n35 3.81063
R24864 CDAC_v3_0.switch_7.Z.n37 CDAC_v3_0.switch_7.Z.n36 3.81063
R24865 CDAC_v3_0.switch_7.Z.n38 CDAC_v3_0.switch_7.Z.n37 3.81063
R24866 CDAC_v3_0.switch_7.Z.n39 CDAC_v3_0.switch_7.Z.n38 3.81063
R24867 CDAC_v3_0.switch_7.Z.n26 CDAC_v3_0.switch_7.Z.n25 3.81063
R24868 CDAC_v3_0.switch_7.Z.n27 CDAC_v3_0.switch_7.Z.n26 3.81063
R24869 CDAC_v3_0.switch_7.Z.n28 CDAC_v3_0.switch_7.Z.n27 3.81063
R24870 CDAC_v3_0.switch_7.Z.n29 CDAC_v3_0.switch_7.Z.n28 3.81063
R24871 CDAC_v3_0.switch_7.Z.n30 CDAC_v3_0.switch_7.Z.n29 3.81063
R24872 CDAC_v3_0.switch_7.Z.n31 CDAC_v3_0.switch_7.Z.n30 3.81063
R24873 CDAC_v3_0.switch_7.Z.n18 CDAC_v3_0.switch_7.Z.n17 3.81063
R24874 CDAC_v3_0.switch_7.Z.n19 CDAC_v3_0.switch_7.Z.n18 3.81063
R24875 CDAC_v3_0.switch_7.Z.n20 CDAC_v3_0.switch_7.Z.n19 3.81063
R24876 CDAC_v3_0.switch_7.Z.n21 CDAC_v3_0.switch_7.Z.n20 3.81063
R24877 CDAC_v3_0.switch_7.Z.n22 CDAC_v3_0.switch_7.Z.n21 3.81063
R24878 CDAC_v3_0.switch_7.Z.n23 CDAC_v3_0.switch_7.Z.n22 3.81063
R24879 CDAC_v3_0.switch_7.Z.n10 CDAC_v3_0.switch_7.Z.n9 3.81063
R24880 CDAC_v3_0.switch_7.Z.n11 CDAC_v3_0.switch_7.Z.n10 3.81063
R24881 CDAC_v3_0.switch_7.Z.n12 CDAC_v3_0.switch_7.Z.n11 3.81063
R24882 CDAC_v3_0.switch_7.Z.n13 CDAC_v3_0.switch_7.Z.n12 3.81063
R24883 CDAC_v3_0.switch_7.Z.n14 CDAC_v3_0.switch_7.Z.n13 3.81063
R24884 CDAC_v3_0.switch_7.Z.n15 CDAC_v3_0.switch_7.Z.n14 3.81063
R24885 CDAC_v3_0.switch_7.Z.n3 CDAC_v3_0.switch_7.Z.n2 3.81063
R24886 CDAC_v3_0.switch_7.Z.n4 CDAC_v3_0.switch_7.Z.n3 3.81063
R24887 CDAC_v3_0.switch_7.Z.n5 CDAC_v3_0.switch_7.Z.n4 3.81063
R24888 CDAC_v3_0.switch_7.Z.n6 CDAC_v3_0.switch_7.Z.n5 3.81063
R24889 CDAC_v3_0.switch_7.Z.n7 CDAC_v3_0.switch_7.Z.n6 3.81063
R24890 CDAC_v3_0.switch_7.Z.n8 CDAC_v3_0.switch_7.Z.n7 3.81063
R24891 CDAC_v3_0.switch_7.Z.n24 CDAC_v3_0.switch_7.Z.n16 3.80593
R24892 CDAC_v3_0.switch_7.Z.n32 CDAC_v3_0.switch_7.Z.n24 3.80593
R24893 CDAC_v3_0.switch_7.Z.n48 CDAC_v3_0.switch_7.Z.n40 3.80593
R24894 CDAC_v3_0.switch_7.Z.n56 CDAC_v3_0.switch_7.Z.n48 3.80593
R24895 CDAC_v3_0.switch_7.Z.n64 CDAC_v3_0.switch_7.Z.n56 3.80593
R24896 CDAC_v3_0.switch_7.Z.n68 CDAC_v3_0.switch_7.Z.n66 1.34289
R24897 CDAC_v3_0.switch_7.Z.n66 CDAC_v3_0.switch_7.Z 0.42713
R24898 CDAC_v3_0.switch_7.Z.n63 CDAC_v3_0.switch_7.Z.t49 0.307567
R24899 CDAC_v3_0.switch_7.Z.n62 CDAC_v3_0.switch_7.Z.t3 0.307567
R24900 CDAC_v3_0.switch_7.Z.n61 CDAC_v3_0.switch_7.Z.t42 0.307567
R24901 CDAC_v3_0.switch_7.Z.n60 CDAC_v3_0.switch_7.Z.t11 0.307567
R24902 CDAC_v3_0.switch_7.Z.n59 CDAC_v3_0.switch_7.Z.t14 0.307567
R24903 CDAC_v3_0.switch_7.Z.n58 CDAC_v3_0.switch_7.Z.t44 0.307567
R24904 CDAC_v3_0.switch_7.Z.n57 CDAC_v3_0.switch_7.Z.t21 0.307567
R24905 CDAC_v3_0.switch_7.Z.n55 CDAC_v3_0.switch_7.Z.t30 0.307567
R24906 CDAC_v3_0.switch_7.Z.n54 CDAC_v3_0.switch_7.Z.t45 0.307567
R24907 CDAC_v3_0.switch_7.Z.n53 CDAC_v3_0.switch_7.Z.t17 0.307567
R24908 CDAC_v3_0.switch_7.Z.n52 CDAC_v3_0.switch_7.Z.t55 0.307567
R24909 CDAC_v3_0.switch_7.Z.n51 CDAC_v3_0.switch_7.Z.t60 0.307567
R24910 CDAC_v3_0.switch_7.Z.n50 CDAC_v3_0.switch_7.Z.t24 0.307567
R24911 CDAC_v3_0.switch_7.Z.n49 CDAC_v3_0.switch_7.Z.t6 0.307567
R24912 CDAC_v3_0.switch_7.Z.n47 CDAC_v3_0.switch_7.Z.t19 0.307567
R24913 CDAC_v3_0.switch_7.Z.n46 CDAC_v3_0.switch_7.Z.t37 0.307567
R24914 CDAC_v3_0.switch_7.Z.n45 CDAC_v3_0.switch_7.Z.t9 0.307567
R24915 CDAC_v3_0.switch_7.Z.n44 CDAC_v3_0.switch_7.Z.t46 0.307567
R24916 CDAC_v3_0.switch_7.Z.n43 CDAC_v3_0.switch_7.Z.t48 0.307567
R24917 CDAC_v3_0.switch_7.Z.n42 CDAC_v3_0.switch_7.Z.t13 0.307567
R24918 CDAC_v3_0.switch_7.Z.n41 CDAC_v3_0.switch_7.Z.t54 0.307567
R24919 CDAC_v3_0.switch_7.Z.n39 CDAC_v3_0.switch_7.Z.t4 0.307567
R24920 CDAC_v3_0.switch_7.Z.n38 CDAC_v3_0.switch_7.Z.t15 0.307567
R24921 CDAC_v3_0.switch_7.Z.n37 CDAC_v3_0.switch_7.Z.t52 0.307567
R24922 CDAC_v3_0.switch_7.Z.n36 CDAC_v3_0.switch_7.Z.t26 0.307567
R24923 CDAC_v3_0.switch_7.Z.n35 CDAC_v3_0.switch_7.Z.t29 0.307567
R24924 CDAC_v3_0.switch_7.Z.n34 CDAC_v3_0.switch_7.Z.t59 0.307567
R24925 CDAC_v3_0.switch_7.Z.n33 CDAC_v3_0.switch_7.Z.t38 0.307567
R24926 CDAC_v3_0.switch_7.Z.n25 CDAC_v3_0.switch_7.Z.t43 0.307567
R24927 CDAC_v3_0.switch_7.Z.n26 CDAC_v3_0.switch_7.Z.t33 0.307567
R24928 CDAC_v3_0.switch_7.Z.n27 CDAC_v3_0.switch_7.Z.t36 0.307567
R24929 CDAC_v3_0.switch_7.Z.n28 CDAC_v3_0.switch_7.Z.t62 0.307567
R24930 CDAC_v3_0.switch_7.Z.n29 CDAC_v3_0.switch_7.Z.t27 0.307567
R24931 CDAC_v3_0.switch_7.Z.n30 CDAC_v3_0.switch_7.Z.t53 0.307567
R24932 CDAC_v3_0.switch_7.Z.n31 CDAC_v3_0.switch_7.Z.t32 0.307567
R24933 CDAC_v3_0.switch_7.Z.n17 CDAC_v3_0.switch_7.Z.t34 0.307567
R24934 CDAC_v3_0.switch_7.Z.n18 CDAC_v3_0.switch_7.Z.t23 0.307567
R24935 CDAC_v3_0.switch_7.Z.n19 CDAC_v3_0.switch_7.Z.t25 0.307567
R24936 CDAC_v3_0.switch_7.Z.n20 CDAC_v3_0.switch_7.Z.t51 0.307567
R24937 CDAC_v3_0.switch_7.Z.n21 CDAC_v3_0.switch_7.Z.t18 0.307567
R24938 CDAC_v3_0.switch_7.Z.n22 CDAC_v3_0.switch_7.Z.t47 0.307567
R24939 CDAC_v3_0.switch_7.Z.n23 CDAC_v3_0.switch_7.Z.t22 0.307567
R24940 CDAC_v3_0.switch_7.Z.n9 CDAC_v3_0.switch_7.Z.t56 0.307567
R24941 CDAC_v3_0.switch_7.Z.n10 CDAC_v3_0.switch_7.Z.t7 0.307567
R24942 CDAC_v3_0.switch_7.Z.n11 CDAC_v3_0.switch_7.Z.t12 0.307567
R24943 CDAC_v3_0.switch_7.Z.n12 CDAC_v3_0.switch_7.Z.t65 0.307567
R24944 CDAC_v3_0.switch_7.Z.n13 CDAC_v3_0.switch_7.Z.t39 0.307567
R24945 CDAC_v3_0.switch_7.Z.n14 CDAC_v3_0.switch_7.Z.t20 0.307567
R24946 CDAC_v3_0.switch_7.Z.n15 CDAC_v3_0.switch_7.Z.t5 0.307567
R24947 CDAC_v3_0.switch_7.Z.n2 CDAC_v3_0.switch_7.Z.t50 0.307567
R24948 CDAC_v3_0.switch_7.Z.n3 CDAC_v3_0.switch_7.Z.t64 0.307567
R24949 CDAC_v3_0.switch_7.Z.n4 CDAC_v3_0.switch_7.Z.t10 0.307567
R24950 CDAC_v3_0.switch_7.Z.n5 CDAC_v3_0.switch_7.Z.t58 0.307567
R24951 CDAC_v3_0.switch_7.Z.n6 CDAC_v3_0.switch_7.Z.t35 0.307567
R24952 CDAC_v3_0.switch_7.Z.n7 CDAC_v3_0.switch_7.Z.t16 0.307567
R24953 CDAC_v3_0.switch_7.Z.n8 CDAC_v3_0.switch_7.Z.t63 0.307567
R24954 CDAC_v3_0.switch_7.Z.n1 CDAC_v3_0.switch_7.Z 0.182141
R24955 CDAC_v3_0.switch_7.Z CDAC_v3_0.switch_7.Z.n68 0.178175
R24956 CDAC_v3_0.switch_7.Z.n1 CDAC_v3_0.switch_7.Z.n0 0.128217
R24957 CDAC_v3_0.switch_7.Z.n0 CDAC_v3_0.switch_7.Z 0.1255
R24958 CDAC_v3_0.switch_7.Z.n0 CDAC_v3_0.switch_7.Z 0.063
R24959 CDAC_v3_0.switch_7.Z.n66 CDAC_v3_0.switch_7.Z.n65 0.063
R24960 CDAC_v3_0.switch_7.Z.n65 CDAC_v3_0.switch_7.Z.n1 0.063
R24961 CDAC_v3_0.switch_7.Z.n68 CDAC_v3_0.switch_7.Z.n67 0.0130546
R24962 D_FlipFlop_4.CLK.n12 D_FlipFlop_4.CLK.t0 168.108
R24963 D_FlipFlop_4.CLK.t2 D_FlipFlop_4.CLK.n5 158.207
R24964 D_FlipFlop_4.CLK D_FlipFlop_4.CLK.t3 158.202
R24965 D_FlipFlop_4.CLK.n0 D_FlipFlop_4.CLK.t5 150.293
R24966 D_FlipFlop_4.CLK.t3 D_FlipFlop_4.CLK.n3 150.293
R24967 D_FlipFlop_4.CLK.n6 D_FlipFlop_4.CLK.t2 150.273
R24968 D_FlipFlop_4.CLK.n9 D_FlipFlop_4.CLK.t7 90.1131
R24969 D_FlipFlop_4.CLK.t7 D_FlipFlop_4.CLK.n8 73.6406
R24970 D_FlipFlop_4.CLK.n2 D_FlipFlop_4.CLK.t4 73.6304
R24971 D_FlipFlop_4.CLK.n1 D_FlipFlop_4.CLK.t6 73.6304
R24972 D_FlipFlop_4.CLK D_FlipFlop_4.CLK.t1 60.3072
R24973 D_FlipFlop_4.CLK.n2 D_FlipFlop_4.CLK.n1 16.332
R24974 D_FlipFlop_4.CLK.n12 D_FlipFlop_4.CLK.n11 1.62007
R24975 D_FlipFlop_4.CLK.n8 D_FlipFlop_4.CLK.n7 1.19615
R24976 D_FlipFlop_4.CLK.n1 D_FlipFlop_4.CLK.n0 1.1717
R24977 D_FlipFlop_4.CLK.n3 D_FlipFlop_4.CLK.n2 1.1717
R24978 D_FlipFlop_4.CLK D_FlipFlop_4.CLK.n12 0.484875
R24979 D_FlipFlop_4.CLK.n3 D_FlipFlop_4.CLK 0.447191
R24980 D_FlipFlop_4.CLK.n0 D_FlipFlop_4.CLK 0.436162
R24981 D_FlipFlop_4.CLK.n5 D_FlipFlop_4.CLK.n4 0.349867
R24982 D_FlipFlop_4.CLK.n5 D_FlipFlop_4.CLK 0.321667
R24983 D_FlipFlop_4.CLK.n8 D_FlipFlop_4.CLK 0.217464
R24984 D_FlipFlop_4.CLK.n2 D_FlipFlop_4.CLK 0.149957
R24985 D_FlipFlop_4.CLK.n11 D_FlipFlop_4.CLK 0.149957
R24986 D_FlipFlop_4.CLK.n7 D_FlipFlop_4.CLK 0.1255
R24987 D_FlipFlop_4.CLK.n1 D_FlipFlop_4.CLK 0.117348
R24988 D_FlipFlop_4.CLK.n10 D_FlipFlop_4.CLK 0.0903438
R24989 D_FlipFlop_4.CLK.n1 D_FlipFlop_4.CLK 0.0454219
R24990 D_FlipFlop_4.CLK.n2 D_FlipFlop_4.CLK 0.0454219
R24991 D_FlipFlop_4.CLK.n10 D_FlipFlop_4.CLK.n9 0.027881
R24992 D_FlipFlop_4.CLK.n9 D_FlipFlop_4.CLK 0.027881
R24993 D_FlipFlop_4.CLK.n7 D_FlipFlop_4.CLK.n6 0.0216397
R24994 D_FlipFlop_4.CLK.n6 D_FlipFlop_4.CLK 0.0216397
R24995 D_FlipFlop_4.CLK.n11 D_FlipFlop_4.CLK.n10 0.0180781
R24996 D_FlipFlop_4.CLK.n4 D_FlipFlop_4.CLK 0.00441667
R24997 D_FlipFlop_4.CLK.n4 D_FlipFlop_4.CLK 0.00406061
R24998 CLK.n1 CLK.t2 158.207
R24999 CLK.n148 CLK.t58 158.183
R25000 CLK.n144 CLK.t68 158.183
R25001 CLK.n139 CLK.t53 158.183
R25002 CLK.n135 CLK.t59 158.183
R25003 CLK.n130 CLK.t106 158.183
R25004 CLK.n126 CLK.t39 158.183
R25005 CLK.n121 CLK.t76 158.183
R25006 CLK.n117 CLK.t85 158.183
R25007 CLK.n112 CLK.t71 158.183
R25008 CLK.n108 CLK.t79 158.183
R25009 CLK.n103 CLK.t117 158.183
R25010 CLK.n99 CLK.t101 158.183
R25011 CLK.n94 CLK.t17 158.183
R25012 CLK.n90 CLK.t11 158.183
R25013 CLK.n85 CLK.t7 158.183
R25014 CLK.n81 CLK.t32 158.183
R25015 CLK.n77 CLK.t67 158.183
R25016 CLK.n72 CLK.t102 158.183
R25017 CLK.n68 CLK.t74 158.183
R25018 CLK.n63 CLK.t66 158.183
R25019 CLK.n59 CLK.t61 158.183
R25020 CLK.n54 CLK.t90 158.183
R25021 CLK.n50 CLK.t81 158.183
R25022 CLK.n45 CLK.t73 158.183
R25023 CLK.n41 CLK.t89 158.183
R25024 CLK.n36 CLK.t93 158.183
R25025 CLK.n32 CLK.t28 158.183
R25026 CLK.n27 CLK.t114 158.183
R25027 CLK.n23 CLK.t92 158.183
R25028 CLK.n18 CLK.t86 158.183
R25029 CLK.n14 CLK.t84 158.183
R25030 CLK.n9 CLK.t103 158.183
R25031 CLK.n5 CLK.t100 158.183
R25032 CLK.n142 CLK.t15 151.506
R25033 CLK.n133 CLK.t8 151.506
R25034 CLK.n124 CLK.t113 151.506
R25035 CLK.n115 CLK.t33 151.506
R25036 CLK.n106 CLK.t24 151.506
R25037 CLK.n97 CLK.t49 151.506
R25038 CLK.n88 CLK.t94 151.506
R25039 CLK.n79 CLK.t111 151.506
R25040 CLK.n75 CLK.t14 151.506
R25041 CLK.n66 CLK.t20 151.506
R25042 CLK.n57 CLK.t9 151.506
R25043 CLK.n48 CLK.t27 151.506
R25044 CLK.n39 CLK.t35 151.506
R25045 CLK.n30 CLK.t108 151.506
R25046 CLK.n21 CLK.t42 151.506
R25047 CLK.n12 CLK.t29 151.506
R25048 CLK.n3 CLK.t48 151.506
R25049 CLK.t68 CLK.n143 151.506
R25050 CLK.t59 CLK.n134 151.506
R25051 CLK.t39 CLK.n125 151.506
R25052 CLK.t85 CLK.n116 151.506
R25053 CLK.t79 CLK.n107 151.506
R25054 CLK.t101 CLK.n98 151.506
R25055 CLK.t11 CLK.n89 151.506
R25056 CLK.t32 CLK.n80 151.506
R25057 CLK.t67 CLK.n76 151.506
R25058 CLK.t74 CLK.n67 151.506
R25059 CLK.t61 CLK.n58 151.506
R25060 CLK.t81 CLK.n49 151.506
R25061 CLK.t89 CLK.n40 151.506
R25062 CLK.t28 CLK.n31 151.506
R25063 CLK.t92 CLK.n22 151.506
R25064 CLK.t84 CLK.n13 151.506
R25065 CLK.t100 CLK.n4 151.506
R25066 CLK.n187 CLK.t110 150.273
R25067 CLK.n182 CLK.t22 150.273
R25068 CLK.n177 CLK.t4 150.273
R25069 CLK.n173 CLK.t105 150.273
R25070 CLK.n168 CLK.t40 150.273
R25071 CLK.n163 CLK.t107 150.273
R25072 CLK.n158 CLK.t82 150.273
R25073 CLK.n154 CLK.t98 150.273
R25074 CLK.t58 CLK.n147 150.273
R25075 CLK.t53 CLK.n138 150.273
R25076 CLK.t106 CLK.n129 150.273
R25077 CLK.t76 CLK.n120 150.273
R25078 CLK.t71 CLK.n111 150.273
R25079 CLK.t117 CLK.n102 150.273
R25080 CLK.t17 CLK.n93 150.273
R25081 CLK.t7 CLK.n84 150.273
R25082 CLK.t102 CLK.n71 150.273
R25083 CLK.t66 CLK.n62 150.273
R25084 CLK.t90 CLK.n53 150.273
R25085 CLK.t73 CLK.n44 150.273
R25086 CLK.t93 CLK.n35 150.273
R25087 CLK.t114 CLK.n26 150.273
R25088 CLK.t86 CLK.n17 150.273
R25089 CLK.t103 CLK.n8 150.273
R25090 CLK.t2 CLK.n0 150.273
R25091 CLK.n147 CLK.t54 74.951
R25092 CLK.n138 CLK.t116 74.951
R25093 CLK.n129 CLK.t31 74.951
R25094 CLK.n120 CLK.t16 74.951
R25095 CLK.n111 CLK.t10 74.951
R25096 CLK.n102 CLK.t69 74.951
R25097 CLK.n93 CLK.t112 74.951
R25098 CLK.n84 CLK.t3 74.951
R25099 CLK.n71 CLK.t0 74.951
R25100 CLK.n62 CLK.t5 74.951
R25101 CLK.n53 CLK.t51 74.951
R25102 CLK.n44 CLK.t12 74.951
R25103 CLK.n35 CLK.t34 74.951
R25104 CLK.n26 CLK.t63 74.951
R25105 CLK.n17 CLK.t41 74.951
R25106 CLK.n8 CLK.t13 74.951
R25107 CLK.n0 CLK.t77 74.951
R25108 CLK.n184 CLK.t115 73.6304
R25109 CLK.n179 CLK.t37 73.6304
R25110 CLK.n174 CLK.t26 73.6304
R25111 CLK.n170 CLK.t97 73.6304
R25112 CLK.n165 CLK.t96 73.6304
R25113 CLK.n160 CLK.t19 73.6304
R25114 CLK.n155 CLK.t91 73.6304
R25115 CLK.n151 CLK.t18 73.6304
R25116 CLK.n143 CLK.t30 73.6304
R25117 CLK.n142 CLK.t52 73.6304
R25118 CLK.n134 CLK.t21 73.6304
R25119 CLK.n133 CLK.t45 73.6304
R25120 CLK.n125 CLK.t36 73.6304
R25121 CLK.n124 CLK.t55 73.6304
R25122 CLK.n116 CLK.t47 73.6304
R25123 CLK.n115 CLK.t70 73.6304
R25124 CLK.n107 CLK.t60 73.6304
R25125 CLK.n106 CLK.t83 73.6304
R25126 CLK.n98 CLK.t109 73.6304
R25127 CLK.n97 CLK.t1 73.6304
R25128 CLK.n89 CLK.t88 73.6304
R25129 CLK.n88 CLK.t104 73.6304
R25130 CLK.n80 CLK.t75 73.6304
R25131 CLK.n79 CLK.t95 73.6304
R25132 CLK.n76 CLK.t62 73.6304
R25133 CLK.n75 CLK.t87 73.6304
R25134 CLK.n67 CLK.t38 73.6304
R25135 CLK.n66 CLK.t57 73.6304
R25136 CLK.n58 CLK.t44 73.6304
R25137 CLK.n57 CLK.t65 73.6304
R25138 CLK.n49 CLK.t43 73.6304
R25139 CLK.n48 CLK.t64 73.6304
R25140 CLK.n40 CLK.t50 73.6304
R25141 CLK.n39 CLK.t72 73.6304
R25142 CLK.n31 CLK.t23 73.6304
R25143 CLK.n30 CLK.t46 73.6304
R25144 CLK.n22 CLK.t56 73.6304
R25145 CLK.n21 CLK.t78 73.6304
R25146 CLK.n13 CLK.t80 73.6304
R25147 CLK.n12 CLK.t99 73.6304
R25148 CLK.n4 CLK.t6 73.6304
R25149 CLK.n3 CLK.t25 73.6304
R25150 CLK.n7 CLK 42.3279
R25151 CLK.n6 CLK 40.6064
R25152 CLK.n16 CLK 39.5361
R25153 CLK.n15 CLK 38.0684
R25154 CLK.n25 CLK 36.7443
R25155 CLK.n24 CLK 35.5304
R25156 CLK.n34 CLK 33.9525
R25157 CLK.n33 CLK 32.9924
R25158 CLK.n43 CLK 31.1607
R25159 CLK.n42 CLK 30.4544
R25160 CLK.n52 CLK 28.3689
R25161 CLK.n178 CLK.n173 28.2614
R25162 CLK.n159 CLK.n154 28.2614
R25163 CLK.n51 CLK 27.9164
R25164 CLK.n61 CLK 25.5771
R25165 CLK.n60 CLK 25.3784
R25166 CLK.n183 CLK.n178 23.7614
R25167 CLK.n188 CLK.n183 23.7614
R25168 CLK.n164 CLK.n159 23.7614
R25169 CLK.n169 CLK.n164 23.7614
R25170 CLK.n69 CLK 22.8404
R25171 CLK.n70 CLK 22.7853
R25172 CLK.n78 CLK 20.3024
R25173 CLK.n149 CLK 19.9935
R25174 CLK.n141 CLK 17.7644
R25175 CLK.n140 CLK 17.2017
R25176 CLK.n143 CLK.n142 16.332
R25177 CLK.n134 CLK.n133 16.332
R25178 CLK.n125 CLK.n124 16.332
R25179 CLK.n116 CLK.n115 16.332
R25180 CLK.n107 CLK.n106 16.332
R25181 CLK.n98 CLK.n97 16.332
R25182 CLK.n89 CLK.n88 16.332
R25183 CLK.n80 CLK.n79 16.332
R25184 CLK.n76 CLK.n75 16.332
R25185 CLK.n67 CLK.n66 16.332
R25186 CLK.n58 CLK.n57 16.332
R25187 CLK.n49 CLK.n48 16.332
R25188 CLK.n40 CLK.n39 16.332
R25189 CLK.n31 CLK.n30 16.332
R25190 CLK.n22 CLK.n21 16.332
R25191 CLK.n13 CLK.n12 16.332
R25192 CLK.n4 CLK.n3 16.332
R25193 CLK.n132 CLK 15.2264
R25194 CLK.n131 CLK 14.4099
R25195 CLK.n123 CLK 12.6884
R25196 CLK.n189 CLK.n188 11.8429
R25197 CLK.n189 CLK.n169 11.8429
R25198 CLK.n122 CLK 11.6181
R25199 CLK.n114 CLK 10.1504
R25200 CLK.n113 CLK 8.82632
R25201 CLK.n105 CLK 7.61236
R25202 CLK.n190 CLK.n150 6.04157
R25203 CLK.n104 CLK 6.03452
R25204 CLK.n96 CLK 5.07436
R25205 CLK.n178 CLK.n177 4.5005
R25206 CLK.n183 CLK.n182 4.5005
R25207 CLK.n188 CLK.n187 4.5005
R25208 CLK.n159 CLK.n158 4.5005
R25209 CLK.n164 CLK.n163 4.5005
R25210 CLK.n169 CLK.n168 4.5005
R25211 CLK CLK.n189 3.43044
R25212 CLK.n95 CLK 3.24272
R25213 CLK.n87 CLK 2.53636
R25214 CLK.n87 CLK.n86 2.33953
R25215 CLK.n96 CLK.n95 2.33953
R25216 CLK.n105 CLK.n104 2.33953
R25217 CLK.n114 CLK.n113 2.33953
R25218 CLK.n123 CLK.n122 2.33953
R25219 CLK.n132 CLK.n131 2.33953
R25220 CLK.n141 CLK.n140 2.33953
R25221 CLK.n7 CLK.n6 2.33953
R25222 CLK.n16 CLK.n15 2.33953
R25223 CLK.n25 CLK.n24 2.33953
R25224 CLK.n34 CLK.n33 2.33953
R25225 CLK.n43 CLK.n42 2.33953
R25226 CLK.n52 CLK.n51 2.33953
R25227 CLK.n61 CLK.n60 2.33953
R25228 CLK.n70 CLK.n69 2.33953
R25229 CLK.n150 CLK.n78 2.12412
R25230 CLK.n186 CLK.n185 1.1717
R25231 CLK.n181 CLK.n180 1.1717
R25232 CLK.n176 CLK.n175 1.1717
R25233 CLK.n172 CLK.n171 1.1717
R25234 CLK.n167 CLK.n166 1.1717
R25235 CLK.n162 CLK.n161 1.1717
R25236 CLK.n157 CLK.n156 1.1717
R25237 CLK.n153 CLK.n152 1.1717
R25238 CLK.n186 CLK 0.932141
R25239 CLK.n181 CLK 0.932141
R25240 CLK.n176 CLK 0.932141
R25241 CLK.n172 CLK 0.932141
R25242 CLK.n167 CLK 0.932141
R25243 CLK.n162 CLK 0.932141
R25244 CLK.n157 CLK 0.932141
R25245 CLK.n153 CLK 0.932141
R25246 CLK.n86 CLK 0.450917
R25247 CLK.n83 CLK.n82 0.349867
R25248 CLK.n92 CLK.n91 0.349867
R25249 CLK.n101 CLK.n100 0.349867
R25250 CLK.n110 CLK.n109 0.349867
R25251 CLK.n119 CLK.n118 0.349867
R25252 CLK.n128 CLK.n127 0.349867
R25253 CLK.n137 CLK.n136 0.349867
R25254 CLK.n146 CLK.n145 0.349867
R25255 CLK.n2 CLK.n1 0.349867
R25256 CLK.n11 CLK.n10 0.349867
R25257 CLK.n20 CLK.n19 0.349867
R25258 CLK.n29 CLK.n28 0.349867
R25259 CLK.n38 CLK.n37 0.349867
R25260 CLK.n47 CLK.n46 0.349867
R25261 CLK.n56 CLK.n55 0.349867
R25262 CLK.n65 CLK.n64 0.349867
R25263 CLK.n74 CLK.n73 0.349867
R25264 CLK.n83 CLK 0.321667
R25265 CLK.n92 CLK 0.321667
R25266 CLK.n101 CLK 0.321667
R25267 CLK.n110 CLK 0.321667
R25268 CLK.n119 CLK 0.321667
R25269 CLK.n128 CLK 0.321667
R25270 CLK.n137 CLK 0.321667
R25271 CLK.n146 CLK 0.321667
R25272 CLK.n1 CLK 0.321667
R25273 CLK.n10 CLK 0.321667
R25274 CLK.n19 CLK 0.321667
R25275 CLK.n28 CLK 0.321667
R25276 CLK.n37 CLK 0.321667
R25277 CLK.n46 CLK 0.321667
R25278 CLK.n55 CLK 0.321667
R25279 CLK.n64 CLK 0.321667
R25280 CLK.n73 CLK 0.321667
R25281 CLK CLK.n149 0.192417
R25282 CLK.n143 CLK 0.149957
R25283 CLK.n134 CLK 0.149957
R25284 CLK.n125 CLK 0.149957
R25285 CLK.n116 CLK 0.149957
R25286 CLK.n107 CLK 0.149957
R25287 CLK.n98 CLK 0.149957
R25288 CLK.n89 CLK 0.149957
R25289 CLK.n80 CLK 0.149957
R25290 CLK.n76 CLK 0.149957
R25291 CLK.n67 CLK 0.149957
R25292 CLK.n58 CLK 0.149957
R25293 CLK.n49 CLK 0.149957
R25294 CLK.n40 CLK 0.149957
R25295 CLK.n31 CLK 0.149957
R25296 CLK.n22 CLK 0.149957
R25297 CLK.n13 CLK 0.149957
R25298 CLK.n4 CLK 0.149957
R25299 CLK.n185 CLK 0.1255
R25300 CLK.n180 CLK 0.1255
R25301 CLK.n175 CLK 0.1255
R25302 CLK.n171 CLK 0.1255
R25303 CLK.n166 CLK 0.1255
R25304 CLK.n161 CLK 0.1255
R25305 CLK.n156 CLK 0.1255
R25306 CLK.n152 CLK 0.1255
R25307 CLK.n142 CLK 0.117348
R25308 CLK.n133 CLK 0.117348
R25309 CLK.n124 CLK 0.117348
R25310 CLK.n115 CLK 0.117348
R25311 CLK.n106 CLK 0.117348
R25312 CLK.n97 CLK 0.117348
R25313 CLK.n88 CLK 0.117348
R25314 CLK.n79 CLK 0.117348
R25315 CLK.n75 CLK 0.117348
R25316 CLK.n66 CLK 0.117348
R25317 CLK.n57 CLK 0.117348
R25318 CLK.n48 CLK 0.117348
R25319 CLK.n39 CLK 0.117348
R25320 CLK.n30 CLK 0.117348
R25321 CLK.n21 CLK 0.117348
R25322 CLK.n12 CLK 0.117348
R25323 CLK.n3 CLK 0.117348
R25324 CLK.n187 CLK.n186 0.063
R25325 CLK.n182 CLK.n181 0.063
R25326 CLK.n177 CLK.n176 0.063
R25327 CLK.n173 CLK.n172 0.063
R25328 CLK.n168 CLK.n167 0.063
R25329 CLK.n163 CLK.n162 0.063
R25330 CLK.n158 CLK.n157 0.063
R25331 CLK.n154 CLK.n153 0.063
R25332 CLK.n147 CLK 0.063
R25333 CLK.n138 CLK 0.063
R25334 CLK.n129 CLK 0.063
R25335 CLK.n120 CLK 0.063
R25336 CLK.n111 CLK 0.063
R25337 CLK.n102 CLK 0.063
R25338 CLK.n93 CLK 0.063
R25339 CLK.n84 CLK 0.063
R25340 CLK.n71 CLK 0.063
R25341 CLK.n62 CLK 0.063
R25342 CLK.n53 CLK 0.063
R25343 CLK.n44 CLK 0.063
R25344 CLK.n35 CLK 0.063
R25345 CLK.n26 CLK 0.063
R25346 CLK.n17 CLK 0.063
R25347 CLK.n8 CLK 0.063
R25348 CLK.n0 CLK 0.063
R25349 CLK.n142 CLK 0.0454219
R25350 CLK.n143 CLK 0.0454219
R25351 CLK.n133 CLK 0.0454219
R25352 CLK.n134 CLK 0.0454219
R25353 CLK.n124 CLK 0.0454219
R25354 CLK.n125 CLK 0.0454219
R25355 CLK.n115 CLK 0.0454219
R25356 CLK.n116 CLK 0.0454219
R25357 CLK.n106 CLK 0.0454219
R25358 CLK.n107 CLK 0.0454219
R25359 CLK.n97 CLK 0.0454219
R25360 CLK.n98 CLK 0.0454219
R25361 CLK.n88 CLK 0.0454219
R25362 CLK.n89 CLK 0.0454219
R25363 CLK.n79 CLK 0.0454219
R25364 CLK.n80 CLK 0.0454219
R25365 CLK.n75 CLK 0.0454219
R25366 CLK.n76 CLK 0.0454219
R25367 CLK.n66 CLK 0.0454219
R25368 CLK.n67 CLK 0.0454219
R25369 CLK.n57 CLK 0.0454219
R25370 CLK.n58 CLK 0.0454219
R25371 CLK.n48 CLK 0.0454219
R25372 CLK.n49 CLK 0.0454219
R25373 CLK.n39 CLK 0.0454219
R25374 CLK.n40 CLK 0.0454219
R25375 CLK.n30 CLK 0.0454219
R25376 CLK.n31 CLK 0.0454219
R25377 CLK.n21 CLK 0.0454219
R25378 CLK.n22 CLK 0.0454219
R25379 CLK.n12 CLK 0.0454219
R25380 CLK.n13 CLK 0.0454219
R25381 CLK.n3 CLK 0.0454219
R25382 CLK.n4 CLK 0.0454219
R25383 CLK.n86 CLK.n85 0.024
R25384 CLK.n85 CLK.n83 0.024
R25385 CLK.n90 CLK.n87 0.024
R25386 CLK.n95 CLK.n94 0.024
R25387 CLK.n94 CLK.n92 0.024
R25388 CLK.n99 CLK.n96 0.024
R25389 CLK.n104 CLK.n103 0.024
R25390 CLK.n103 CLK.n101 0.024
R25391 CLK.n108 CLK.n105 0.024
R25392 CLK.n113 CLK.n112 0.024
R25393 CLK.n112 CLK.n110 0.024
R25394 CLK.n117 CLK.n114 0.024
R25395 CLK.n122 CLK.n121 0.024
R25396 CLK.n121 CLK.n119 0.024
R25397 CLK.n126 CLK.n123 0.024
R25398 CLK.n131 CLK.n130 0.024
R25399 CLK.n130 CLK.n128 0.024
R25400 CLK.n135 CLK.n132 0.024
R25401 CLK.n140 CLK.n139 0.024
R25402 CLK.n139 CLK.n137 0.024
R25403 CLK.n144 CLK.n141 0.024
R25404 CLK.n149 CLK.n148 0.024
R25405 CLK.n148 CLK.n146 0.024
R25406 CLK.n6 CLK.n5 0.024
R25407 CLK.n9 CLK.n7 0.024
R25408 CLK.n10 CLK.n9 0.024
R25409 CLK.n15 CLK.n14 0.024
R25410 CLK.n18 CLK.n16 0.024
R25411 CLK.n19 CLK.n18 0.024
R25412 CLK.n24 CLK.n23 0.024
R25413 CLK.n27 CLK.n25 0.024
R25414 CLK.n28 CLK.n27 0.024
R25415 CLK.n33 CLK.n32 0.024
R25416 CLK.n36 CLK.n34 0.024
R25417 CLK.n37 CLK.n36 0.024
R25418 CLK.n42 CLK.n41 0.024
R25419 CLK.n45 CLK.n43 0.024
R25420 CLK.n46 CLK.n45 0.024
R25421 CLK.n51 CLK.n50 0.024
R25422 CLK.n54 CLK.n52 0.024
R25423 CLK.n55 CLK.n54 0.024
R25424 CLK.n60 CLK.n59 0.024
R25425 CLK.n63 CLK.n61 0.024
R25426 CLK.n64 CLK.n63 0.024
R25427 CLK.n69 CLK.n68 0.024
R25428 CLK.n72 CLK.n70 0.024
R25429 CLK.n73 CLK.n72 0.024
R25430 CLK.n78 CLK.n77 0.024
R25431 CLK.n150 CLK 0.024
R25432 CLK.n81 CLK 0.0218636
R25433 CLK CLK.n81 0.0204394
R25434 CLK CLK.n90 0.0204394
R25435 CLK CLK.n99 0.0204394
R25436 CLK CLK.n108 0.0204394
R25437 CLK CLK.n117 0.0204394
R25438 CLK CLK.n126 0.0204394
R25439 CLK CLK.n135 0.0204394
R25440 CLK CLK.n144 0.0204394
R25441 CLK.n5 CLK 0.0204394
R25442 CLK.n14 CLK 0.0204394
R25443 CLK.n23 CLK 0.0204394
R25444 CLK.n32 CLK 0.0204394
R25445 CLK.n41 CLK 0.0204394
R25446 CLK.n50 CLK 0.0204394
R25447 CLK.n59 CLK 0.0204394
R25448 CLK.n68 CLK 0.0204394
R25449 CLK.n77 CLK 0.0204394
R25450 CLK.n185 CLK.n184 0.0107679
R25451 CLK.n184 CLK 0.0107679
R25452 CLK.n180 CLK.n179 0.0107679
R25453 CLK.n179 CLK 0.0107679
R25454 CLK.n175 CLK.n174 0.0107679
R25455 CLK.n174 CLK 0.0107679
R25456 CLK.n171 CLK.n170 0.0107679
R25457 CLK.n170 CLK 0.0107679
R25458 CLK.n166 CLK.n165 0.0107679
R25459 CLK.n165 CLK 0.0107679
R25460 CLK.n161 CLK.n160 0.0107679
R25461 CLK.n160 CLK 0.0107679
R25462 CLK.n156 CLK.n155 0.0107679
R25463 CLK.n155 CLK 0.0107679
R25464 CLK.n152 CLK.n151 0.0107679
R25465 CLK.n151 CLK 0.0107679
R25466 CLK.n82 CLK 0.00441667
R25467 CLK.n91 CLK 0.00441667
R25468 CLK.n100 CLK 0.00441667
R25469 CLK.n109 CLK 0.00441667
R25470 CLK.n118 CLK 0.00441667
R25471 CLK.n127 CLK 0.00441667
R25472 CLK.n136 CLK 0.00441667
R25473 CLK.n145 CLK 0.00441667
R25474 CLK.n2 CLK 0.00441667
R25475 CLK.n11 CLK 0.00441667
R25476 CLK.n20 CLK 0.00441667
R25477 CLK.n29 CLK 0.00441667
R25478 CLK.n38 CLK 0.00441667
R25479 CLK.n47 CLK 0.00441667
R25480 CLK.n56 CLK 0.00441667
R25481 CLK.n65 CLK 0.00441667
R25482 CLK.n74 CLK 0.00441667
R25483 CLK CLK.n190 0.00441667
R25484 CLK.n82 CLK 0.00406061
R25485 CLK.n91 CLK 0.00406061
R25486 CLK.n100 CLK 0.00406061
R25487 CLK.n109 CLK 0.00406061
R25488 CLK.n118 CLK 0.00406061
R25489 CLK.n127 CLK 0.00406061
R25490 CLK.n136 CLK 0.00406061
R25491 CLK.n145 CLK 0.00406061
R25492 CLK CLK.n2 0.00406061
R25493 CLK CLK.n11 0.00406061
R25494 CLK CLK.n20 0.00406061
R25495 CLK CLK.n29 0.00406061
R25496 CLK CLK.n38 0.00406061
R25497 CLK CLK.n47 0.00406061
R25498 CLK CLK.n56 0.00406061
R25499 CLK CLK.n65 0.00406061
R25500 CLK CLK.n74 0.00406061
R25501 CLK.n190 CLK 0.00406061
R25502 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 169.46
R25503 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 167.809
R25504 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 167.809
R25505 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 167.227
R25506 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 151.594
R25507 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 150.273
R25508 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 74.8641
R25509 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 73.6304
R25510 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 61.84
R25511 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 12.3891
R25512 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 11.4489
R25513 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R25514 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 0.280391
R25515 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 0.200143
R25516 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R25517 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R25518 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 0.149957
R25519 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.063
R25520 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 0.063
R25521 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 0.063
R25522 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 0.063
R25523 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R25524 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t0 169.46
R25525 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t3 167.809
R25526 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t2 167.809
R25527 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t7 167.226
R25528 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n6 150.273
R25529 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t6 150.273
R25530 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t4 74.951
R25531 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t5 73.6304
R25532 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t1 60.3943
R25533 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n4 12.3891
R25534 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n8 11.4489
R25535 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n10 1.68257
R25536 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n0 1.44615
R25537 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n2 1.2342
R25538 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 1.08448
R25539 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.932141
R25540 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n9 0.3496
R25541 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n7 0.280391
R25542 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.063
R25543 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.063
R25544 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n3 0.063
R25545 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.063
R25546 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n5 0.063
R25547 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n1 0.063
R25548 D_FlipFlop_0.CLK.n12 D_FlipFlop_0.CLK.t0 168.108
R25549 D_FlipFlop_0.CLK.t7 D_FlipFlop_0.CLK.n5 158.207
R25550 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.t2 158.202
R25551 D_FlipFlop_0.CLK.n0 D_FlipFlop_0.CLK.t4 150.293
R25552 D_FlipFlop_0.CLK.t2 D_FlipFlop_0.CLK.n3 150.293
R25553 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK.t7 150.273
R25554 D_FlipFlop_0.CLK.n9 D_FlipFlop_0.CLK.t6 90.1131
R25555 D_FlipFlop_0.CLK.t6 D_FlipFlop_0.CLK.n8 73.6406
R25556 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK.t3 73.6304
R25557 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK.t5 73.6304
R25558 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.t1 60.3072
R25559 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK.n1 16.332
R25560 D_FlipFlop_0.CLK.n12 D_FlipFlop_0.CLK.n11 1.62007
R25561 D_FlipFlop_0.CLK.n8 D_FlipFlop_0.CLK.n7 1.19615
R25562 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK.n0 1.1717
R25563 D_FlipFlop_0.CLK.n3 D_FlipFlop_0.CLK.n2 1.1717
R25564 D_FlipFlop_0.CLK D_FlipFlop_0.CLK.n12 0.484875
R25565 D_FlipFlop_0.CLK.n3 D_FlipFlop_0.CLK 0.447191
R25566 D_FlipFlop_0.CLK.n0 D_FlipFlop_0.CLK 0.436162
R25567 D_FlipFlop_0.CLK.n5 D_FlipFlop_0.CLK.n4 0.349867
R25568 D_FlipFlop_0.CLK.n5 D_FlipFlop_0.CLK 0.321667
R25569 D_FlipFlop_0.CLK.n8 D_FlipFlop_0.CLK 0.217464
R25570 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK 0.149957
R25571 D_FlipFlop_0.CLK.n11 D_FlipFlop_0.CLK 0.149957
R25572 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK 0.1255
R25573 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK 0.117348
R25574 D_FlipFlop_0.CLK.n10 D_FlipFlop_0.CLK 0.0903438
R25575 D_FlipFlop_0.CLK.n1 D_FlipFlop_0.CLK 0.0454219
R25576 D_FlipFlop_0.CLK.n2 D_FlipFlop_0.CLK 0.0454219
R25577 D_FlipFlop_0.CLK.n10 D_FlipFlop_0.CLK.n9 0.027881
R25578 D_FlipFlop_0.CLK.n9 D_FlipFlop_0.CLK 0.027881
R25579 D_FlipFlop_0.CLK.n7 D_FlipFlop_0.CLK.n6 0.0216397
R25580 D_FlipFlop_0.CLK.n6 D_FlipFlop_0.CLK 0.0216397
R25581 D_FlipFlop_0.CLK.n11 D_FlipFlop_0.CLK.n10 0.0180781
R25582 D_FlipFlop_0.CLK.n4 D_FlipFlop_0.CLK 0.00441667
R25583 D_FlipFlop_0.CLK.n4 D_FlipFlop_0.CLK 0.00406061
R25584 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 169.46
R25585 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 168.089
R25586 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 167.809
R25587 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 150.887
R25588 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 73.6304
R25589 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 60.3943
R25590 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 12.0358
R25591 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 11.4489
R25592 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 1.05069
R25593 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 0.981478
R25594 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.769522
R25595 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 0.745065
R25596 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.580578
R25597 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 0.533109
R25598 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.428234
R25599 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.063
R25600 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 0.063
R25601 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 0.063
R25602 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.063
R25603 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 0.063
R25604 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 0.063
R25605 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t2 316.762
R25606 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t0 169.195
R25607 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t5 150.887
R25608 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n2 150.273
R25609 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t3 74.951
R25610 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t4 73.6304
R25611 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t1 60.3943
R25612 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n6 12.0358
R25613 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n8 0.981478
R25614 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.769522
R25615 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n0 0.745065
R25616 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.580578
R25617 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n4 0.533109
R25618 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.428234
R25619 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.063
R25620 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.063
R25621 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n3 0.063
R25622 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n5 0.063
R25623 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.063
R25624 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n7 0.063
R25625 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n1 0.063
R25626 FFCLR.n195 FFCLR.t0 169.46
R25627 FFCLR.n195 FFCLR.t1 167.809
R25628 FFCLR.n194 FFCLR.t2 167.809
R25629 FFCLR.n178 FFCLR.t32 165.081
R25630 FFCLR.n142 FFCLR.t31 158.988
R25631 FFCLR.n120 FFCLR.t36 158.988
R25632 FFCLR.n98 FFCLR.t27 158.988
R25633 FFCLR.n76 FFCLR.t42 158.988
R25634 FFCLR.n54 FFCLR.t28 158.988
R25635 FFCLR.n32 FFCLR.t38 158.988
R25636 FFCLR.n11 FFCLR.t25 158.988
R25637 D_FlipFlop_0.nPRE FFCLR.t54 158.581
R25638 FFCLR.n191 FFCLR.t22 158.565
R25639 FFCLR.t22 FFCLR.n190 151.594
R25640 FFCLR.n150 FFCLR.t37 150.293
R25641 FFCLR.n144 FFCLR.t40 150.293
R25642 FFCLR.n128 FFCLR.t46 150.293
R25643 FFCLR.n122 FFCLR.t9 150.293
R25644 FFCLR.n106 FFCLR.t20 150.293
R25645 FFCLR.n100 FFCLR.t21 150.293
R25646 FFCLR.n84 FFCLR.t50 150.293
R25647 FFCLR.n78 FFCLR.t19 150.293
R25648 FFCLR.n62 FFCLR.t17 150.293
R25649 FFCLR.n56 FFCLR.t30 150.293
R25650 FFCLR.n40 FFCLR.t29 150.293
R25651 FFCLR.n34 FFCLR.t10 150.293
R25652 FFCLR.n19 FFCLR.t57 150.293
R25653 FFCLR.n13 FFCLR.t34 150.293
R25654 FFCLR.t54 FFCLR.n5 150.293
R25655 FFCLR.t32 FFCLR.n2 150.293
R25656 FFCLR.n182 FFCLR.t23 150.273
R25657 FFCLR.n179 FFCLR.t5 150.273
R25658 FFCLR.n172 FFCLR.t6 150.273
R25659 FFCLR.n166 FFCLR.t12 150.273
R25660 FFCLR.t31 FFCLR.n141 150.273
R25661 FFCLR.t36 FFCLR.n119 150.273
R25662 FFCLR.t27 FFCLR.n97 150.273
R25663 FFCLR.t42 FFCLR.n75 150.273
R25664 FFCLR.t28 FFCLR.n53 150.273
R25665 FFCLR.t38 FFCLR.n31 150.273
R25666 FFCLR.t25 FFCLR.n10 150.273
R25667 Ring_Counter_0.Q0 FFCLR.t41 99.8701
R25668 FFCLR.n181 FFCLR.t14 74.163
R25669 FFCLR.t41 FFCLR.n186 74.163
R25670 FFCLR.n170 FFCLR.t55 73.6406
R25671 FFCLR.n164 FFCLR.t56 73.6406
R25672 FFCLR.n139 FFCLR.t7 73.6406
R25673 FFCLR.n117 FFCLR.t48 73.6406
R25674 FFCLR.n95 FFCLR.t58 73.6406
R25675 FFCLR.n73 FFCLR.t15 73.6406
R25676 FFCLR.n51 FFCLR.t59 73.6406
R25677 FFCLR.n29 FFCLR.t18 73.6406
R25678 FFCLR.n8 FFCLR.t26 73.6406
R25679 FFCLR.n190 FFCLR.t13 73.6304
R25680 FFCLR.n152 FFCLR.t45 73.6304
R25681 FFCLR.n146 FFCLR.t8 73.6304
R25682 FFCLR.n130 FFCLR.t51 73.6304
R25683 FFCLR.n124 FFCLR.t16 73.6304
R25684 FFCLR.n108 FFCLR.t39 73.6304
R25685 FFCLR.n102 FFCLR.t47 73.6304
R25686 FFCLR.n86 FFCLR.t53 73.6304
R25687 FFCLR.n80 FFCLR.t24 73.6304
R25688 FFCLR.n64 FFCLR.t43 73.6304
R25689 FFCLR.n58 FFCLR.t52 73.6304
R25690 FFCLR.n42 FFCLR.t44 73.6304
R25691 FFCLR.n36 FFCLR.t33 73.6304
R25692 FFCLR.n21 FFCLR.t11 73.6304
R25693 FFCLR.n15 FFCLR.t49 73.6304
R25694 FFCLR.n3 FFCLR.t4 73.6304
R25695 FFCLR.n0 FFCLR.t35 73.6304
R25696 FFCLR.n197 FFCLR.t3 62.1634
R25697 FFCLR.n50 FFCLR.n28 27.1442
R25698 FFCLR.n161 FFCLR.n160 26.7393
R25699 FFCLR.n72 FFCLR.n50 23.7342
R25700 FFCLR.n94 FFCLR.n72 23.7342
R25701 FFCLR.n116 FFCLR.n94 23.7342
R25702 FFCLR.n138 FFCLR.n116 23.7342
R25703 FFCLR.n160 FFCLR.n138 23.7342
R25704 FFCLR.n176 FFCLR.n169 15.5222
R25705 FFCLR.n156 FFCLR.n149 15.5222
R25706 FFCLR.n134 FFCLR.n127 15.5222
R25707 FFCLR.n112 FFCLR.n105 15.5222
R25708 FFCLR.n90 FFCLR.n83 15.5222
R25709 FFCLR.n68 FFCLR.n61 15.5222
R25710 FFCLR.n46 FFCLR.n39 15.5222
R25711 FFCLR.n25 FFCLR.n18 15.5222
R25712 FFCLR.n185 FFCLR.n184 12.6418
R25713 FFCLR.n196 FFCLR.n195 11.4489
R25714 FFCLR.n177 FFCLR.n176 8.24202
R25715 FFCLR.n194 FFCLR.n193 8.21389
R25716 D_FlipFlop_1.nCLR FFCLR.n156 7.85707
R25717 D_FlipFlop_2.nCLR FFCLR.n134 7.85707
R25718 D_FlipFlop_3.nCLR FFCLR.n112 7.85707
R25719 D_FlipFlop_5.nCLR FFCLR.n90 7.85707
R25720 D_FlipFlop_4.nCLR FFCLR.n68 7.85707
R25721 D_FlipFlop_6.nCLR FFCLR.n46 7.85707
R25722 D_FlipFlop_7.nCLR FFCLR.n25 7.85707
R25723 FFCLR.n178 FFCLR.n177 5.81925
R25724 FFCLR.n176 FFCLR.n175 4.5005
R25725 FFCLR.n156 FFCLR.n155 4.5005
R25726 FFCLR.n134 FFCLR.n133 4.5005
R25727 FFCLR.n112 FFCLR.n111 4.5005
R25728 FFCLR.n90 FFCLR.n89 4.5005
R25729 FFCLR.n68 FFCLR.n67 4.5005
R25730 FFCLR.n46 FFCLR.n45 4.5005
R25731 FFCLR.n25 FFCLR.n24 4.5005
R25732 FFCLR.n188 FFCLR.n178 4.03482
R25733 FFCLR.n50 FFCLR.n49 3.4105
R25734 FFCLR.n72 FFCLR.n71 3.4105
R25735 FFCLR.n94 FFCLR.n93 3.4105
R25736 FFCLR.n116 FFCLR.n115 3.4105
R25737 FFCLR.n138 FFCLR.n137 3.4105
R25738 FFCLR.n160 FFCLR.n159 3.4105
R25739 Ring_Counter_0.D_FlipFlop_0.Q Ring_Counter_0.Q0 1.3729
R25740 Ring_Counter_0.D_FlipFlop_0.Q Ring_Counter_0.Q0 1.24814
R25741 FFCLR.n189 Ring_Counter_0.Q0 1.2047
R25742 FFCLR.n140 FFCLR.n139 1.19615
R25743 FFCLR.n118 FFCLR.n117 1.19615
R25744 FFCLR.n96 FFCLR.n95 1.19615
R25745 FFCLR.n74 FFCLR.n73 1.19615
R25746 FFCLR.n52 FFCLR.n51 1.19615
R25747 FFCLR.n30 FFCLR.n29 1.19615
R25748 FFCLR.n9 FFCLR.n8 1.19615
R25749 FFCLR.n5 FFCLR.n4 1.19615
R25750 FFCLR.n2 FFCLR.n1 1.19615
R25751 FFCLR.n151 D_FlipFlop_1.3-input-nand_3.A 1.09561
R25752 FFCLR.n145 D_FlipFlop_1.3-input-nand_5.A 1.09561
R25753 FFCLR.n129 D_FlipFlop_2.3-input-nand_3.A 1.09561
R25754 FFCLR.n123 D_FlipFlop_2.3-input-nand_5.A 1.09561
R25755 FFCLR.n107 D_FlipFlop_3.3-input-nand_3.A 1.09561
R25756 FFCLR.n101 D_FlipFlop_3.3-input-nand_5.A 1.09561
R25757 FFCLR.n85 D_FlipFlop_5.3-input-nand_3.A 1.09561
R25758 FFCLR.n79 D_FlipFlop_5.3-input-nand_5.A 1.09561
R25759 FFCLR.n63 D_FlipFlop_4.3-input-nand_3.A 1.09561
R25760 FFCLR.n57 D_FlipFlop_4.3-input-nand_5.A 1.09561
R25761 FFCLR.n41 D_FlipFlop_6.3-input-nand_3.A 1.09561
R25762 FFCLR.n35 D_FlipFlop_6.3-input-nand_5.A 1.09561
R25763 FFCLR.n20 D_FlipFlop_7.3-input-nand_3.A 1.09561
R25764 FFCLR.n14 D_FlipFlop_7.3-input-nand_5.A 1.09561
R25765 FFCLR.n188 FFCLR.n187 0.922483
R25766 FFCLR.n181 Ring_Counter_0.D_FlipFlop_1.Inverter_0.Vin 0.851043
R25767 FFCLR.n186 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.B 0.851043
R25768 FFCLR.n171 FFCLR.n170 0.796696
R25769 FFCLR.n165 FFCLR.n164 0.796696
R25770 FFCLR.n154 FFCLR.n153 0.796696
R25771 FFCLR.n148 FFCLR.n147 0.796696
R25772 FFCLR.n132 FFCLR.n131 0.796696
R25773 FFCLR.n126 FFCLR.n125 0.796696
R25774 FFCLR.n110 FFCLR.n109 0.796696
R25775 FFCLR.n104 FFCLR.n103 0.796696
R25776 FFCLR.n88 FFCLR.n87 0.796696
R25777 FFCLR.n82 FFCLR.n81 0.796696
R25778 FFCLR.n66 FFCLR.n65 0.796696
R25779 FFCLR.n60 FFCLR.n59 0.796696
R25780 FFCLR.n44 FFCLR.n43 0.796696
R25781 FFCLR.n38 FFCLR.n37 0.796696
R25782 FFCLR.n23 FFCLR.n22 0.796696
R25783 FFCLR.n17 FFCLR.n16 0.796696
R25784 FFCLR.n143 D_FlipFlop_1.nCLR 0.73135
R25785 FFCLR.n121 D_FlipFlop_2.nCLR 0.73135
R25786 FFCLR.n99 D_FlipFlop_3.nCLR 0.73135
R25787 FFCLR.n77 D_FlipFlop_5.nCLR 0.73135
R25788 FFCLR.n55 D_FlipFlop_4.nCLR 0.73135
R25789 FFCLR.n33 D_FlipFlop_6.nCLR 0.73135
R25790 FFCLR.n12 D_FlipFlop_7.nCLR 0.73135
R25791 FFCLR.n142 D_FlipFlop_1.nCLR 0.716182
R25792 FFCLR.n120 D_FlipFlop_2.nCLR 0.716182
R25793 FFCLR.n98 D_FlipFlop_3.nCLR 0.716182
R25794 FFCLR.n76 D_FlipFlop_5.nCLR 0.716182
R25795 FFCLR.n54 D_FlipFlop_4.nCLR 0.716182
R25796 FFCLR.n32 D_FlipFlop_6.nCLR 0.716182
R25797 FFCLR.n11 D_FlipFlop_7.nCLR 0.716182
R25798 FFCLR.n163 D_FlipFlop_0.nPRE 0.716182
R25799 FFCLR.n158 FFCLR.n157 0.675733
R25800 FFCLR.n136 FFCLR.n135 0.675733
R25801 FFCLR.n114 FFCLR.n113 0.675733
R25802 FFCLR.n92 FFCLR.n91 0.675733
R25803 FFCLR.n70 FFCLR.n69 0.675733
R25804 FFCLR.n48 FFCLR.n47 0.675733
R25805 FFCLR.n27 FFCLR.n26 0.675733
R25806 FFCLR.n154 D_FlipFlop_1.3-input-nand_3.A 0.662609
R25807 FFCLR.n148 D_FlipFlop_1.3-input-nand_5.A 0.662609
R25808 FFCLR.n132 D_FlipFlop_2.3-input-nand_3.A 0.662609
R25809 FFCLR.n126 D_FlipFlop_2.3-input-nand_5.A 0.662609
R25810 FFCLR.n110 D_FlipFlop_3.3-input-nand_3.A 0.662609
R25811 FFCLR.n104 D_FlipFlop_3.3-input-nand_5.A 0.662609
R25812 FFCLR.n88 D_FlipFlop_5.3-input-nand_3.A 0.662609
R25813 FFCLR.n82 D_FlipFlop_5.3-input-nand_5.A 0.662609
R25814 FFCLR.n66 D_FlipFlop_4.3-input-nand_3.A 0.662609
R25815 FFCLR.n60 D_FlipFlop_4.3-input-nand_5.A 0.662609
R25816 FFCLR.n44 D_FlipFlop_6.3-input-nand_3.A 0.662609
R25817 FFCLR.n38 D_FlipFlop_6.3-input-nand_5.A 0.662609
R25818 FFCLR.n23 D_FlipFlop_7.3-input-nand_3.A 0.662609
R25819 FFCLR.n17 D_FlipFlop_7.3-input-nand_5.A 0.662609
R25820 FFCLR.n158 D_FlipFlop_1.nCLR 0.617909
R25821 FFCLR.n136 D_FlipFlop_2.nCLR 0.617909
R25822 FFCLR.n114 D_FlipFlop_3.nCLR 0.617909
R25823 FFCLR.n92 D_FlipFlop_5.nCLR 0.617909
R25824 FFCLR.n70 D_FlipFlop_4.nCLR 0.617909
R25825 FFCLR.n48 D_FlipFlop_6.nCLR 0.617909
R25826 FFCLR.n27 D_FlipFlop_7.nCLR 0.617909
R25827 FFCLR.n183 FFCLR.n182 0.61463
R25828 FFCLR.n180 FFCLR.n179 0.61463
R25829 FFCLR.n171 D_FlipFlop_0.3-input-nand_2.A 0.524957
R25830 FFCLR.n165 D_FlipFlop_0.3-input-nand_4.A 0.524957
R25831 FFCLR.n163 FFCLR.n162 0.490867
R25832 FFCLR.n183 Ring_Counter_0.D_FlipFlop_1.Inverter_0.Vin 0.486828
R25833 FFCLR.n180 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.B 0.486828
R25834 FFCLR.n150 D_FlipFlop_1.3-input-nand_3.A 0.447191
R25835 FFCLR.n144 D_FlipFlop_1.3-input-nand_5.A 0.447191
R25836 FFCLR.n128 D_FlipFlop_2.3-input-nand_3.A 0.447191
R25837 FFCLR.n122 D_FlipFlop_2.3-input-nand_5.A 0.447191
R25838 FFCLR.n106 D_FlipFlop_3.3-input-nand_3.A 0.447191
R25839 FFCLR.n100 D_FlipFlop_3.3-input-nand_5.A 0.447191
R25840 FFCLR.n84 D_FlipFlop_5.3-input-nand_3.A 0.447191
R25841 FFCLR.n78 D_FlipFlop_5.3-input-nand_5.A 0.447191
R25842 FFCLR.n62 D_FlipFlop_4.3-input-nand_3.A 0.447191
R25843 FFCLR.n56 D_FlipFlop_4.3-input-nand_5.A 0.447191
R25844 FFCLR.n40 D_FlipFlop_6.3-input-nand_3.A 0.447191
R25845 FFCLR.n34 D_FlipFlop_6.3-input-nand_5.A 0.447191
R25846 FFCLR.n19 D_FlipFlop_7.3-input-nand_3.A 0.447191
R25847 FFCLR.n13 D_FlipFlop_7.3-input-nand_5.A 0.447191
R25848 FFCLR.n5 D_FlipFlop_0.3-input-nand_1.A 0.447191
R25849 FFCLR.n2 Nand_Gate_7.B 0.447191
R25850 FFCLR.n193 FFCLR.n192 0.425067
R25851 FFCLR.n189 FFCLR.n188 0.399217
R25852 FFCLR.n193 Ring_Counter_0.D_FlipFlop_0.Q 0.39003
R25853 FFCLR.n162 D_FlipFlop_0.nPRE 0.297383
R25854 FFCLR.n196 FFCLR.n194 0.280391
R25855 FFCLR.n174 D_FlipFlop_0.3-input-nand_2.A 0.252453
R25856 FFCLR.n168 D_FlipFlop_0.3-input-nand_4.A 0.252453
R25857 FFCLR.n7 FFCLR.n6 0.241767
R25858 FFCLR.n174 FFCLR.n173 0.226043
R25859 FFCLR.n168 FFCLR.n167 0.226043
R25860 FFCLR.n151 FFCLR.n150 0.226043
R25861 FFCLR.n145 FFCLR.n144 0.226043
R25862 FFCLR.n129 FFCLR.n128 0.226043
R25863 FFCLR.n123 FFCLR.n122 0.226043
R25864 FFCLR.n107 FFCLR.n106 0.226043
R25865 FFCLR.n101 FFCLR.n100 0.226043
R25866 FFCLR.n85 FFCLR.n84 0.226043
R25867 FFCLR.n79 FFCLR.n78 0.226043
R25868 FFCLR.n63 FFCLR.n62 0.226043
R25869 FFCLR.n57 FFCLR.n56 0.226043
R25870 FFCLR.n41 FFCLR.n40 0.226043
R25871 FFCLR.n35 FFCLR.n34 0.226043
R25872 FFCLR.n20 FFCLR.n19 0.226043
R25873 FFCLR.n14 FFCLR.n13 0.226043
R25874 FFCLR.n7 D_FlipFlop_0.nPRE 0.223394
R25875 FFCLR.n170 D_FlipFlop_0.3-input-nand_2.A 0.217464
R25876 FFCLR.n164 D_FlipFlop_0.3-input-nand_4.A 0.217464
R25877 FFCLR.n139 D_FlipFlop_1.3-input-nand_0.A 0.217464
R25878 FFCLR.n117 D_FlipFlop_2.3-input-nand_0.A 0.217464
R25879 FFCLR.n95 D_FlipFlop_3.3-input-nand_0.A 0.217464
R25880 FFCLR.n73 D_FlipFlop_5.3-input-nand_0.A 0.217464
R25881 FFCLR.n51 D_FlipFlop_4.3-input-nand_0.A 0.217464
R25882 FFCLR.n29 D_FlipFlop_6.3-input-nand_0.A 0.217464
R25883 FFCLR.n8 D_FlipFlop_7.3-input-nand_0.A 0.217464
R25884 FFCLR.n197 FFCLR.n196 0.200143
R25885 FFCLR.n173 D_FlipFlop_0.3-input-nand_2.A 0.1255
R25886 FFCLR.n167 D_FlipFlop_0.3-input-nand_4.A 0.1255
R25887 FFCLR.n140 D_FlipFlop_1.3-input-nand_0.A 0.1255
R25888 FFCLR.n153 D_FlipFlop_1.3-input-nand_3.A 0.1255
R25889 FFCLR.n147 D_FlipFlop_1.3-input-nand_5.A 0.1255
R25890 FFCLR.n118 D_FlipFlop_2.3-input-nand_0.A 0.1255
R25891 FFCLR.n131 D_FlipFlop_2.3-input-nand_3.A 0.1255
R25892 FFCLR.n125 D_FlipFlop_2.3-input-nand_5.A 0.1255
R25893 FFCLR.n96 D_FlipFlop_3.3-input-nand_0.A 0.1255
R25894 FFCLR.n109 D_FlipFlop_3.3-input-nand_3.A 0.1255
R25895 FFCLR.n103 D_FlipFlop_3.3-input-nand_5.A 0.1255
R25896 FFCLR.n74 D_FlipFlop_5.3-input-nand_0.A 0.1255
R25897 FFCLR.n87 D_FlipFlop_5.3-input-nand_3.A 0.1255
R25898 FFCLR.n81 D_FlipFlop_5.3-input-nand_5.A 0.1255
R25899 FFCLR.n52 D_FlipFlop_4.3-input-nand_0.A 0.1255
R25900 FFCLR.n65 D_FlipFlop_4.3-input-nand_3.A 0.1255
R25901 FFCLR.n59 D_FlipFlop_4.3-input-nand_5.A 0.1255
R25902 FFCLR.n30 D_FlipFlop_6.3-input-nand_0.A 0.1255
R25903 FFCLR.n43 D_FlipFlop_6.3-input-nand_3.A 0.1255
R25904 FFCLR.n37 D_FlipFlop_6.3-input-nand_5.A 0.1255
R25905 FFCLR.n9 D_FlipFlop_7.3-input-nand_0.A 0.1255
R25906 FFCLR.n22 D_FlipFlop_7.3-input-nand_3.A 0.1255
R25907 FFCLR.n16 D_FlipFlop_7.3-input-nand_5.A 0.1255
R25908 FFCLR.n4 D_FlipFlop_0.3-input-nand_1.A 0.1255
R25909 FFCLR.n1 Nand_Gate_7.B 0.1255
R25910 FFCLR.n190 Ring_Counter_0.D_FlipFlop_0.3-input-nand_5.C 0.063
R25911 FFCLR.n182 Ring_Counter_0.D_FlipFlop_1.Inverter_0.Vin 0.063
R25912 FFCLR.n184 FFCLR.n181 0.063
R25913 FFCLR.n184 FFCLR.n183 0.063
R25914 FFCLR.n179 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.B 0.063
R25915 FFCLR.n186 FFCLR.n185 0.063
R25916 FFCLR.n185 FFCLR.n180 0.063
R25917 FFCLR.n175 FFCLR.n171 0.063
R25918 FFCLR.n175 FFCLR.n174 0.063
R25919 FFCLR.n169 FFCLR.n165 0.063
R25920 FFCLR.n169 FFCLR.n168 0.063
R25921 FFCLR.n155 FFCLR.n151 0.063
R25922 FFCLR.n155 FFCLR.n154 0.063
R25923 FFCLR.n149 FFCLR.n145 0.063
R25924 FFCLR.n149 FFCLR.n148 0.063
R25925 FFCLR.n133 FFCLR.n129 0.063
R25926 FFCLR.n133 FFCLR.n132 0.063
R25927 FFCLR.n127 FFCLR.n123 0.063
R25928 FFCLR.n127 FFCLR.n126 0.063
R25929 FFCLR.n111 FFCLR.n107 0.063
R25930 FFCLR.n111 FFCLR.n110 0.063
R25931 FFCLR.n105 FFCLR.n101 0.063
R25932 FFCLR.n105 FFCLR.n104 0.063
R25933 FFCLR.n89 FFCLR.n85 0.063
R25934 FFCLR.n89 FFCLR.n88 0.063
R25935 FFCLR.n83 FFCLR.n79 0.063
R25936 FFCLR.n83 FFCLR.n82 0.063
R25937 FFCLR.n67 FFCLR.n63 0.063
R25938 FFCLR.n67 FFCLR.n66 0.063
R25939 FFCLR.n61 FFCLR.n57 0.063
R25940 FFCLR.n61 FFCLR.n60 0.063
R25941 FFCLR.n45 FFCLR.n41 0.063
R25942 FFCLR.n45 FFCLR.n44 0.063
R25943 FFCLR.n39 FFCLR.n35 0.063
R25944 FFCLR.n39 FFCLR.n38 0.063
R25945 FFCLR.n24 FFCLR.n20 0.063
R25946 FFCLR.n24 FFCLR.n23 0.063
R25947 FFCLR.n18 FFCLR.n14 0.063
R25948 FFCLR.n18 FFCLR.n17 0.063
R25949 Ring_Counter_0.D_FlipFlop_0.3-input-nand_4.Vout FFCLR.n197 0.063
R25950 FFCLR.n143 FFCLR.n142 0.0569
R25951 FFCLR.n121 FFCLR.n120 0.0569
R25952 FFCLR.n99 FFCLR.n98 0.0569
R25953 FFCLR.n77 FFCLR.n76 0.0569
R25954 FFCLR.n55 FFCLR.n54 0.0569
R25955 FFCLR.n33 FFCLR.n32 0.0569
R25956 FFCLR.n12 FFCLR.n11 0.0569
R25957 FFCLR.n159 FFCLR.n143 0.024
R25958 FFCLR.n159 FFCLR.n158 0.024
R25959 FFCLR.n137 FFCLR.n121 0.024
R25960 FFCLR.n137 FFCLR.n136 0.024
R25961 FFCLR.n115 FFCLR.n99 0.024
R25962 FFCLR.n115 FFCLR.n114 0.024
R25963 FFCLR.n93 FFCLR.n77 0.024
R25964 FFCLR.n93 FFCLR.n92 0.024
R25965 FFCLR.n71 FFCLR.n55 0.024
R25966 FFCLR.n71 FFCLR.n70 0.024
R25967 FFCLR.n49 FFCLR.n33 0.024
R25968 FFCLR.n49 FFCLR.n48 0.024
R25969 FFCLR.n28 FFCLR.n12 0.024
R25970 FFCLR.n28 FFCLR.n27 0.024
R25971 FFCLR.n162 FFCLR.n161 0.024
R25972 FFCLR.n161 FFCLR.n7 0.024
R25973 FFCLR.n177 FFCLR.n163 0.024
R25974 FFCLR.n191 FFCLR.n189 0.024
R25975 FFCLR.n173 FFCLR.n172 0.0216397
R25976 FFCLR.n172 D_FlipFlop_0.3-input-nand_2.A 0.0216397
R25977 FFCLR.n167 FFCLR.n166 0.0216397
R25978 FFCLR.n166 D_FlipFlop_0.3-input-nand_4.A 0.0216397
R25979 FFCLR.n141 FFCLR.n140 0.0216397
R25980 FFCLR.n141 D_FlipFlop_1.3-input-nand_0.A 0.0216397
R25981 FFCLR.n119 FFCLR.n118 0.0216397
R25982 FFCLR.n119 D_FlipFlop_2.3-input-nand_0.A 0.0216397
R25983 FFCLR.n97 FFCLR.n96 0.0216397
R25984 FFCLR.n97 D_FlipFlop_3.3-input-nand_0.A 0.0216397
R25985 FFCLR.n75 FFCLR.n74 0.0216397
R25986 FFCLR.n75 D_FlipFlop_5.3-input-nand_0.A 0.0216397
R25987 FFCLR.n53 FFCLR.n52 0.0216397
R25988 FFCLR.n53 D_FlipFlop_4.3-input-nand_0.A 0.0216397
R25989 FFCLR.n31 FFCLR.n30 0.0216397
R25990 FFCLR.n31 D_FlipFlop_6.3-input-nand_0.A 0.0216397
R25991 FFCLR.n10 FFCLR.n9 0.0216397
R25992 FFCLR.n10 D_FlipFlop_7.3-input-nand_0.A 0.0216397
R25993 Ring_Counter_0.D_FlipFlop_0.Q FFCLR.n191 0.0204394
R25994 FFCLR.n153 FFCLR.n152 0.0107679
R25995 FFCLR.n152 D_FlipFlop_1.3-input-nand_3.A 0.0107679
R25996 FFCLR.n147 FFCLR.n146 0.0107679
R25997 FFCLR.n146 D_FlipFlop_1.3-input-nand_5.A 0.0107679
R25998 FFCLR.n131 FFCLR.n130 0.0107679
R25999 FFCLR.n130 D_FlipFlop_2.3-input-nand_3.A 0.0107679
R26000 FFCLR.n125 FFCLR.n124 0.0107679
R26001 FFCLR.n124 D_FlipFlop_2.3-input-nand_5.A 0.0107679
R26002 FFCLR.n109 FFCLR.n108 0.0107679
R26003 FFCLR.n108 D_FlipFlop_3.3-input-nand_3.A 0.0107679
R26004 FFCLR.n103 FFCLR.n102 0.0107679
R26005 FFCLR.n102 D_FlipFlop_3.3-input-nand_5.A 0.0107679
R26006 FFCLR.n87 FFCLR.n86 0.0107679
R26007 FFCLR.n86 D_FlipFlop_5.3-input-nand_3.A 0.0107679
R26008 FFCLR.n81 FFCLR.n80 0.0107679
R26009 FFCLR.n80 D_FlipFlop_5.3-input-nand_5.A 0.0107679
R26010 FFCLR.n65 FFCLR.n64 0.0107679
R26011 FFCLR.n64 D_FlipFlop_4.3-input-nand_3.A 0.0107679
R26012 FFCLR.n59 FFCLR.n58 0.0107679
R26013 FFCLR.n58 D_FlipFlop_4.3-input-nand_5.A 0.0107679
R26014 FFCLR.n43 FFCLR.n42 0.0107679
R26015 FFCLR.n42 D_FlipFlop_6.3-input-nand_3.A 0.0107679
R26016 FFCLR.n37 FFCLR.n36 0.0107679
R26017 FFCLR.n36 D_FlipFlop_6.3-input-nand_5.A 0.0107679
R26018 FFCLR.n22 FFCLR.n21 0.0107679
R26019 FFCLR.n21 D_FlipFlop_7.3-input-nand_3.A 0.0107679
R26020 FFCLR.n16 FFCLR.n15 0.0107679
R26021 FFCLR.n15 D_FlipFlop_7.3-input-nand_5.A 0.0107679
R26022 FFCLR.n4 FFCLR.n3 0.0107679
R26023 FFCLR.n3 D_FlipFlop_0.3-input-nand_1.A 0.0107679
R26024 FFCLR.n1 FFCLR.n0 0.0107679
R26025 FFCLR.n0 Nand_Gate_7.B 0.0107679
R26026 FFCLR.n157 D_FlipFlop_1.nCLR 0.00441667
R26027 FFCLR.n135 D_FlipFlop_2.nCLR 0.00441667
R26028 FFCLR.n113 D_FlipFlop_3.nCLR 0.00441667
R26029 FFCLR.n91 D_FlipFlop_5.nCLR 0.00441667
R26030 FFCLR.n69 D_FlipFlop_4.nCLR 0.00441667
R26031 FFCLR.n47 D_FlipFlop_6.nCLR 0.00441667
R26032 FFCLR.n26 D_FlipFlop_7.nCLR 0.00441667
R26033 FFCLR.n6 D_FlipFlop_0.nPRE 0.00441667
R26034 FFCLR.n187 Ring_Counter_0.Q0 0.00441667
R26035 FFCLR.n192 Ring_Counter_0.D_FlipFlop_0.Q 0.00441667
R26036 FFCLR.n187 Ring_Counter_0.Q0 0.00406061
R26037 FFCLR.n157 D_FlipFlop_1.nCLR 0.00406061
R26038 FFCLR.n135 D_FlipFlop_2.nCLR 0.00406061
R26039 FFCLR.n113 D_FlipFlop_3.nCLR 0.00406061
R26040 FFCLR.n91 D_FlipFlop_5.nCLR 0.00406061
R26041 FFCLR.n69 D_FlipFlop_4.nCLR 0.00406061
R26042 FFCLR.n47 D_FlipFlop_6.nCLR 0.00406061
R26043 FFCLR.n26 D_FlipFlop_7.nCLR 0.00406061
R26044 FFCLR.n6 D_FlipFlop_0.nPRE 0.00406061
R26045 FFCLR.n192 Ring_Counter_0.D_FlipFlop_0.Q 0.00406061
R26046 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t3 316.762
R26047 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t0 169.195
R26048 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t4 150.887
R26049 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n2 150.273
R26050 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t5 74.951
R26051 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t2 73.6304
R26052 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t1 60.3943
R26053 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n6 12.0358
R26054 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n8 0.981478
R26055 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.769522
R26056 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n0 0.745065
R26057 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.580578
R26058 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n4 0.533109
R26059 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.428234
R26060 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.063
R26061 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.063
R26062 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n3 0.063
R26063 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n5 0.063
R26064 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.063
R26065 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n7 0.063
R26066 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n1 0.063
R26067 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 179.256
R26068 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 168.089
R26069 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 150.887
R26070 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 73.6304
R26071 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 60.3943
R26072 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 12.0358
R26073 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 1.05069
R26074 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 0.981478
R26075 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.769522
R26076 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 0.745065
R26077 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.580578
R26078 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 0.533109
R26079 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.428234
R26080 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.063
R26081 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 0.063
R26082 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 0.063
R26083 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.063
R26084 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 0.063
R26085 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 0.063
R26086 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 179.256
R26087 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 168.089
R26088 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 150.887
R26089 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 73.6304
R26090 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 60.3943
R26091 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 12.0358
R26092 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 1.05069
R26093 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 0.981478
R26094 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.769522
R26095 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 0.745065
R26096 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.580578
R26097 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 0.533109
R26098 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.428234
R26099 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.063
R26100 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 0.063
R26101 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 0.063
R26102 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.063
R26103 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 0.063
R26104 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 0.063
R26105 CDAC_v3_0.switch_5.Z.n0 CDAC_v3_0.switch_5.Z.t2 168.075
R26106 CDAC_v3_0.switch_5.Z.n0 CDAC_v3_0.switch_5.Z.t1 168.075
R26107 CDAC_v3_0.switch_5.Z.n36 CDAC_v3_0.switch_5.Z.t0 60.6851
R26108 CDAC_v3_0.switch_5.Z CDAC_v3_0.switch_5.Z.t3 60.6226
R26109 CDAC_v3_0.switch_5.Z.n34 CDAC_v3_0.switch_5.Z.n33 31.4952
R26110 CDAC_v3_0.switch_5.Z.n25 CDAC_v3_0.switch_5.Z.n17 15.5277
R26111 CDAC_v3_0.switch_5.Z.n17 CDAC_v3_0.switch_5.Z.n9 12.4517
R26112 CDAC_v3_0.switch_5.Z.n17 CDAC_v3_0.switch_5.Z.n16 8.6463
R26113 CDAC_v3_0.switch_5.Z.n33 CDAC_v3_0.switch_5.Z.n32 6.18037
R26114 CDAC_v3_0.switch_5.Z.n25 CDAC_v3_0.switch_5.Z.n24 6.18037
R26115 CDAC_v3_0.switch_5.Z.n26 CDAC_v3_0.switch_5.Z.t21 4.1177
R26116 CDAC_v3_0.switch_5.Z.n18 CDAC_v3_0.switch_5.Z.t16 4.1177
R26117 CDAC_v3_0.switch_5.Z.n10 CDAC_v3_0.switch_5.Z.t22 4.1177
R26118 CDAC_v3_0.switch_5.Z.n3 CDAC_v3_0.switch_5.Z.t34 4.1177
R26119 CDAC_v3_0.switch_5.Z.n32 CDAC_v3_0.switch_5.Z.n31 3.81063
R26120 CDAC_v3_0.switch_5.Z.n31 CDAC_v3_0.switch_5.Z.n30 3.81063
R26121 CDAC_v3_0.switch_5.Z.n30 CDAC_v3_0.switch_5.Z.n29 3.81063
R26122 CDAC_v3_0.switch_5.Z.n29 CDAC_v3_0.switch_5.Z.n28 3.81063
R26123 CDAC_v3_0.switch_5.Z.n28 CDAC_v3_0.switch_5.Z.n27 3.81063
R26124 CDAC_v3_0.switch_5.Z.n27 CDAC_v3_0.switch_5.Z.n26 3.81063
R26125 CDAC_v3_0.switch_5.Z.n24 CDAC_v3_0.switch_5.Z.n23 3.81063
R26126 CDAC_v3_0.switch_5.Z.n23 CDAC_v3_0.switch_5.Z.n22 3.81063
R26127 CDAC_v3_0.switch_5.Z.n22 CDAC_v3_0.switch_5.Z.n21 3.81063
R26128 CDAC_v3_0.switch_5.Z.n21 CDAC_v3_0.switch_5.Z.n20 3.81063
R26129 CDAC_v3_0.switch_5.Z.n20 CDAC_v3_0.switch_5.Z.n19 3.81063
R26130 CDAC_v3_0.switch_5.Z.n19 CDAC_v3_0.switch_5.Z.n18 3.81063
R26131 CDAC_v3_0.switch_5.Z.n16 CDAC_v3_0.switch_5.Z.n15 3.81063
R26132 CDAC_v3_0.switch_5.Z.n15 CDAC_v3_0.switch_5.Z.n14 3.81063
R26133 CDAC_v3_0.switch_5.Z.n14 CDAC_v3_0.switch_5.Z.n13 3.81063
R26134 CDAC_v3_0.switch_5.Z.n13 CDAC_v3_0.switch_5.Z.n12 3.81063
R26135 CDAC_v3_0.switch_5.Z.n12 CDAC_v3_0.switch_5.Z.n11 3.81063
R26136 CDAC_v3_0.switch_5.Z.n11 CDAC_v3_0.switch_5.Z.n10 3.81063
R26137 CDAC_v3_0.switch_5.Z.n9 CDAC_v3_0.switch_5.Z.n8 3.81063
R26138 CDAC_v3_0.switch_5.Z.n8 CDAC_v3_0.switch_5.Z.n7 3.81063
R26139 CDAC_v3_0.switch_5.Z.n7 CDAC_v3_0.switch_5.Z.n6 3.81063
R26140 CDAC_v3_0.switch_5.Z.n6 CDAC_v3_0.switch_5.Z.n5 3.81063
R26141 CDAC_v3_0.switch_5.Z.n5 CDAC_v3_0.switch_5.Z.n4 3.81063
R26142 CDAC_v3_0.switch_5.Z.n4 CDAC_v3_0.switch_5.Z.n3 3.81063
R26143 CDAC_v3_0.switch_5.Z.n33 CDAC_v3_0.switch_5.Z.n25 3.80593
R26144 CDAC_v3_0.switch_5.Z.n2 CDAC_v3_0.switch_5.Z.n1 1.34289
R26145 CDAC_v3_0.switch_5.Z.n2 CDAC_v3_0.switch_5.Z 0.42713
R26146 CDAC_v3_0.switch_5.Z.n32 CDAC_v3_0.switch_5.Z.t28 0.307567
R26147 CDAC_v3_0.switch_5.Z.n31 CDAC_v3_0.switch_5.Z.t30 0.307567
R26148 CDAC_v3_0.switch_5.Z.n30 CDAC_v3_0.switch_5.Z.t23 0.307567
R26149 CDAC_v3_0.switch_5.Z.n29 CDAC_v3_0.switch_5.Z.t24 0.307567
R26150 CDAC_v3_0.switch_5.Z.n28 CDAC_v3_0.switch_5.Z.t10 0.307567
R26151 CDAC_v3_0.switch_5.Z.n27 CDAC_v3_0.switch_5.Z.t18 0.307567
R26152 CDAC_v3_0.switch_5.Z.n26 CDAC_v3_0.switch_5.Z.t4 0.307567
R26153 CDAC_v3_0.switch_5.Z.n24 CDAC_v3_0.switch_5.Z.t26 0.307567
R26154 CDAC_v3_0.switch_5.Z.n23 CDAC_v3_0.switch_5.Z.t27 0.307567
R26155 CDAC_v3_0.switch_5.Z.n22 CDAC_v3_0.switch_5.Z.t17 0.307567
R26156 CDAC_v3_0.switch_5.Z.n21 CDAC_v3_0.switch_5.Z.t19 0.307567
R26157 CDAC_v3_0.switch_5.Z.n20 CDAC_v3_0.switch_5.Z.t6 0.307567
R26158 CDAC_v3_0.switch_5.Z.n19 CDAC_v3_0.switch_5.Z.t14 0.307567
R26159 CDAC_v3_0.switch_5.Z.n18 CDAC_v3_0.switch_5.Z.t35 0.307567
R26160 CDAC_v3_0.switch_5.Z.n10 CDAC_v3_0.switch_5.Z.t32 0.307567
R26161 CDAC_v3_0.switch_5.Z.n11 CDAC_v3_0.switch_5.Z.t13 0.307567
R26162 CDAC_v3_0.switch_5.Z.n12 CDAC_v3_0.switch_5.Z.t7 0.307567
R26163 CDAC_v3_0.switch_5.Z.n13 CDAC_v3_0.switch_5.Z.t9 0.307567
R26164 CDAC_v3_0.switch_5.Z.n14 CDAC_v3_0.switch_5.Z.t15 0.307567
R26165 CDAC_v3_0.switch_5.Z.n15 CDAC_v3_0.switch_5.Z.t11 0.307567
R26166 CDAC_v3_0.switch_5.Z.n16 CDAC_v3_0.switch_5.Z.t29 0.307567
R26167 CDAC_v3_0.switch_5.Z.n3 CDAC_v3_0.switch_5.Z.t12 0.307567
R26168 CDAC_v3_0.switch_5.Z.n4 CDAC_v3_0.switch_5.Z.t31 0.307567
R26169 CDAC_v3_0.switch_5.Z.n5 CDAC_v3_0.switch_5.Z.t8 0.307567
R26170 CDAC_v3_0.switch_5.Z.n6 CDAC_v3_0.switch_5.Z.t5 0.307567
R26171 CDAC_v3_0.switch_5.Z.n7 CDAC_v3_0.switch_5.Z.t20 0.307567
R26172 CDAC_v3_0.switch_5.Z.n8 CDAC_v3_0.switch_5.Z.t25 0.307567
R26173 CDAC_v3_0.switch_5.Z.n9 CDAC_v3_0.switch_5.Z.t33 0.307567
R26174 CDAC_v3_0.switch_5.Z.n35 CDAC_v3_0.switch_5.Z 0.182141
R26175 CDAC_v3_0.switch_5.Z.n1 CDAC_v3_0.switch_5.Z 0.178175
R26176 CDAC_v3_0.switch_5.Z.n36 CDAC_v3_0.switch_5.Z.n35 0.128217
R26177 CDAC_v3_0.switch_5.Z.n36 CDAC_v3_0.switch_5.Z 0.1255
R26178 CDAC_v3_0.switch_5.Z.n34 CDAC_v3_0.switch_5.Z.n2 0.063
R26179 CDAC_v3_0.switch_5.Z.n35 CDAC_v3_0.switch_5.Z.n34 0.063
R26180 CDAC_v3_0.switch_5.Z CDAC_v3_0.switch_5.Z.n36 0.063
R26181 CDAC_v3_0.switch_5.Z.n1 CDAC_v3_0.switch_5.Z.n0 0.0130546
R26182 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 169.46
R26183 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 167.809
R26184 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 167.809
R26185 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 167.227
R26186 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 151.594
R26187 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 150.273
R26188 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 74.8641
R26189 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 73.6304
R26190 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 61.84
R26191 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 12.3891
R26192 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 11.4489
R26193 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.38637
R26194 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 0.280391
R26195 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 0.200143
R26196 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.152844
R26197 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.149957
R26198 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 0.149957
R26199 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.063
R26200 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 0.063
R26201 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 0.063
R26202 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 0.063
R26203 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.0454219
R26204 D_FlipFlop_2.CLK.n12 D_FlipFlop_2.CLK.t0 168.108
R26205 D_FlipFlop_2.CLK.t5 D_FlipFlop_2.CLK.n5 158.207
R26206 D_FlipFlop_2.CLK D_FlipFlop_2.CLK.t6 158.202
R26207 D_FlipFlop_2.CLK.n0 D_FlipFlop_2.CLK.t4 150.293
R26208 D_FlipFlop_2.CLK.t6 D_FlipFlop_2.CLK.n3 150.293
R26209 D_FlipFlop_2.CLK.n6 D_FlipFlop_2.CLK.t5 150.273
R26210 D_FlipFlop_2.CLK.n9 D_FlipFlop_2.CLK.t3 90.1131
R26211 D_FlipFlop_2.CLK.t3 D_FlipFlop_2.CLK.n8 73.6406
R26212 D_FlipFlop_2.CLK.n2 D_FlipFlop_2.CLK.t2 73.6304
R26213 D_FlipFlop_2.CLK.n1 D_FlipFlop_2.CLK.t7 73.6304
R26214 D_FlipFlop_2.CLK D_FlipFlop_2.CLK.t1 60.3072
R26215 D_FlipFlop_2.CLK.n2 D_FlipFlop_2.CLK.n1 16.332
R26216 D_FlipFlop_2.CLK.n12 D_FlipFlop_2.CLK.n11 1.62007
R26217 D_FlipFlop_2.CLK.n8 D_FlipFlop_2.CLK.n7 1.19615
R26218 D_FlipFlop_2.CLK.n1 D_FlipFlop_2.CLK.n0 1.1717
R26219 D_FlipFlop_2.CLK.n3 D_FlipFlop_2.CLK.n2 1.1717
R26220 D_FlipFlop_2.CLK D_FlipFlop_2.CLK.n12 0.484875
R26221 D_FlipFlop_2.CLK.n3 D_FlipFlop_2.CLK 0.447191
R26222 D_FlipFlop_2.CLK.n0 D_FlipFlop_2.CLK 0.436162
R26223 D_FlipFlop_2.CLK.n5 D_FlipFlop_2.CLK.n4 0.349867
R26224 D_FlipFlop_2.CLK.n5 D_FlipFlop_2.CLK 0.321667
R26225 D_FlipFlop_2.CLK.n8 D_FlipFlop_2.CLK 0.217464
R26226 D_FlipFlop_2.CLK.n2 D_FlipFlop_2.CLK 0.149957
R26227 D_FlipFlop_2.CLK.n11 D_FlipFlop_2.CLK 0.149957
R26228 D_FlipFlop_2.CLK.n7 D_FlipFlop_2.CLK 0.1255
R26229 D_FlipFlop_2.CLK.n1 D_FlipFlop_2.CLK 0.117348
R26230 D_FlipFlop_2.CLK.n10 D_FlipFlop_2.CLK 0.0903438
R26231 D_FlipFlop_2.CLK.n1 D_FlipFlop_2.CLK 0.0454219
R26232 D_FlipFlop_2.CLK.n2 D_FlipFlop_2.CLK 0.0454219
R26233 D_FlipFlop_2.CLK.n10 D_FlipFlop_2.CLK.n9 0.027881
R26234 D_FlipFlop_2.CLK.n9 D_FlipFlop_2.CLK 0.027881
R26235 D_FlipFlop_2.CLK.n7 D_FlipFlop_2.CLK.n6 0.0216397
R26236 D_FlipFlop_2.CLK.n6 D_FlipFlop_2.CLK 0.0216397
R26237 D_FlipFlop_2.CLK.n11 D_FlipFlop_2.CLK.n10 0.0180781
R26238 D_FlipFlop_2.CLK.n4 D_FlipFlop_2.CLK 0.00441667
R26239 D_FlipFlop_2.CLK.n4 D_FlipFlop_2.CLK 0.00406061
R26240 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t0 169.46
R26241 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t1 167.809
R26242 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t3 167.809
R26243 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t5 167.226
R26244 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n6 150.273
R26245 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t6 150.273
R26246 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t4 74.951
R26247 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t7 73.6304
R26248 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t2 60.3943
R26249 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n4 12.3891
R26250 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n8 11.4489
R26251 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n10 1.68257
R26252 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n0 1.44615
R26253 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n2 1.2342
R26254 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 1.08448
R26255 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.932141
R26256 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n9 0.3496
R26257 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n7 0.280391
R26258 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.063
R26259 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.063
R26260 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n3 0.063
R26261 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.063
R26262 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n5 0.063
R26263 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n1 0.063
R26264 a_51632_31172.n0 a_51632_31172.t3 1302.5
R26265 a_51632_31172.n0 a_51632_31172.t1 1301.07
R26266 a_51632_31172.t0 a_51632_31172.n1 30.7707
R26267 a_51632_31172.n1 a_51632_31172.t2 18.2748
R26268 a_51632_31172.n1 a_51632_31172.n0 0.340816
R26269 Nand_Gate_6.A.n19 Nand_Gate_6.A.t3 169.46
R26270 Nand_Gate_6.A.n19 Nand_Gate_6.A.t2 167.809
R26271 Nand_Gate_6.A.n18 Nand_Gate_6.A.t0 167.809
R26272 Nand_Gate_6.A.n12 Nand_Gate_6.A.t10 167.268
R26273 Nand_Gate_6.A.n15 Nand_Gate_6.A.t5 158.565
R26274 Nand_Gate_6.A.t5 Nand_Gate_6.A.n14 151.594
R26275 Nand_Gate_6.A.t10 Nand_Gate_6.A.n2 150.293
R26276 Nand_Gate_6.A.n6 Nand_Gate_6.A.t11 150.273
R26277 Nand_Gate_6.A.n3 Nand_Gate_6.A.t9 150.273
R26278 Nand_Gate_6.A Nand_Gate_6.A.t8 99.8701
R26279 Nand_Gate_6.A.n5 Nand_Gate_6.A.t4 74.163
R26280 Nand_Gate_6.A.t8 Nand_Gate_6.A.n10 74.163
R26281 Nand_Gate_6.A.n14 Nand_Gate_6.A.t7 73.6304
R26282 Nand_Gate_6.A.n0 Nand_Gate_6.A.t6 73.6304
R26283 Nand_Gate_6.A.n21 Nand_Gate_6.A.t1 62.1634
R26284 Nand_Gate_6.A.n9 Nand_Gate_6.A.n8 12.6418
R26285 Nand_Gate_6.A.n20 Nand_Gate_6.A.n19 11.4489
R26286 Nand_Gate_6.A.n18 Nand_Gate_6.A.n17 8.21389
R26287 Nand_Gate_6.A.n13 Nand_Gate_6.A 1.2047
R26288 Nand_Gate_6.A.n2 Nand_Gate_6.A.n1 1.19615
R26289 Nand_Gate_6.A.n12 Nand_Gate_6.A.n11 0.922483
R26290 Nand_Gate_6.A.n5 Nand_Gate_6.A 0.851043
R26291 Nand_Gate_6.A.n10 Nand_Gate_6.A 0.851043
R26292 Nand_Gate_6.A.n7 Nand_Gate_6.A.n6 0.61463
R26293 Nand_Gate_6.A.n4 Nand_Gate_6.A.n3 0.61463
R26294 Nand_Gate_6.A.n7 Nand_Gate_6.A 0.486828
R26295 Nand_Gate_6.A.n4 Nand_Gate_6.A 0.486828
R26296 Nand_Gate_6.A.n2 Nand_Gate_6.A 0.447191
R26297 Nand_Gate_6.A.n17 Nand_Gate_6.A.n16 0.425067
R26298 Nand_Gate_6.A.n13 Nand_Gate_6.A.n12 0.399217
R26299 Nand_Gate_6.A.n17 Nand_Gate_6.A 0.39003
R26300 Nand_Gate_6.A.n20 Nand_Gate_6.A.n18 0.280391
R26301 Nand_Gate_6.A.n21 Nand_Gate_6.A.n20 0.200143
R26302 Nand_Gate_6.A.n1 Nand_Gate_6.A 0.1255
R26303 Nand_Gate_6.A.n14 Nand_Gate_6.A 0.063
R26304 Nand_Gate_6.A.n6 Nand_Gate_6.A 0.063
R26305 Nand_Gate_6.A.n8 Nand_Gate_6.A.n5 0.063
R26306 Nand_Gate_6.A.n8 Nand_Gate_6.A.n7 0.063
R26307 Nand_Gate_6.A.n3 Nand_Gate_6.A 0.063
R26308 Nand_Gate_6.A.n10 Nand_Gate_6.A.n9 0.063
R26309 Nand_Gate_6.A.n9 Nand_Gate_6.A.n4 0.063
R26310 Nand_Gate_6.A Nand_Gate_6.A.n21 0.063
R26311 Nand_Gate_6.A.n15 Nand_Gate_6.A.n13 0.024
R26312 Nand_Gate_6.A Nand_Gate_6.A.n15 0.0204394
R26313 Nand_Gate_6.A.n1 Nand_Gate_6.A.n0 0.0107679
R26314 Nand_Gate_6.A.n0 Nand_Gate_6.A 0.0107679
R26315 Nand_Gate_6.A.n11 Nand_Gate_6.A 0.00441667
R26316 Nand_Gate_6.A.n16 Nand_Gate_6.A 0.00441667
R26317 Nand_Gate_6.A.n11 Nand_Gate_6.A 0.00406061
R26318 Nand_Gate_6.A.n16 Nand_Gate_6.A 0.00406061
R26319 D_FlipFlop_6.CLK.n12 D_FlipFlop_6.CLK.t0 168.108
R26320 D_FlipFlop_6.CLK.t7 D_FlipFlop_6.CLK.n5 158.207
R26321 D_FlipFlop_6.CLK D_FlipFlop_6.CLK.t2 158.202
R26322 D_FlipFlop_6.CLK.n0 D_FlipFlop_6.CLK.t5 150.293
R26323 D_FlipFlop_6.CLK.t2 D_FlipFlop_6.CLK.n3 150.293
R26324 D_FlipFlop_6.CLK.n6 D_FlipFlop_6.CLK.t7 150.273
R26325 D_FlipFlop_6.CLK.n9 D_FlipFlop_6.CLK.t4 90.1131
R26326 D_FlipFlop_6.CLK.t4 D_FlipFlop_6.CLK.n8 73.6406
R26327 D_FlipFlop_6.CLK.n2 D_FlipFlop_6.CLK.t6 73.6304
R26328 D_FlipFlop_6.CLK.n1 D_FlipFlop_6.CLK.t3 73.6304
R26329 D_FlipFlop_6.CLK D_FlipFlop_6.CLK.t1 60.3072
R26330 D_FlipFlop_6.CLK.n2 D_FlipFlop_6.CLK.n1 16.332
R26331 D_FlipFlop_6.CLK.n12 D_FlipFlop_6.CLK.n11 1.62007
R26332 D_FlipFlop_6.CLK.n8 D_FlipFlop_6.CLK.n7 1.19615
R26333 D_FlipFlop_6.CLK.n1 D_FlipFlop_6.CLK.n0 1.1717
R26334 D_FlipFlop_6.CLK.n3 D_FlipFlop_6.CLK.n2 1.1717
R26335 D_FlipFlop_6.CLK D_FlipFlop_6.CLK.n12 0.484875
R26336 D_FlipFlop_6.CLK.n3 D_FlipFlop_6.CLK 0.447191
R26337 D_FlipFlop_6.CLK.n0 D_FlipFlop_6.CLK 0.436162
R26338 D_FlipFlop_6.CLK.n5 D_FlipFlop_6.CLK.n4 0.349867
R26339 D_FlipFlop_6.CLK.n5 D_FlipFlop_6.CLK 0.321667
R26340 D_FlipFlop_6.CLK.n8 D_FlipFlop_6.CLK 0.217464
R26341 D_FlipFlop_6.CLK.n2 D_FlipFlop_6.CLK 0.149957
R26342 D_FlipFlop_6.CLK.n11 D_FlipFlop_6.CLK 0.149957
R26343 D_FlipFlop_6.CLK.n7 D_FlipFlop_6.CLK 0.1255
R26344 D_FlipFlop_6.CLK.n1 D_FlipFlop_6.CLK 0.117348
R26345 D_FlipFlop_6.CLK.n10 D_FlipFlop_6.CLK 0.0903438
R26346 D_FlipFlop_6.CLK.n1 D_FlipFlop_6.CLK 0.0454219
R26347 D_FlipFlop_6.CLK.n2 D_FlipFlop_6.CLK 0.0454219
R26348 D_FlipFlop_6.CLK.n10 D_FlipFlop_6.CLK.n9 0.027881
R26349 D_FlipFlop_6.CLK.n9 D_FlipFlop_6.CLK 0.027881
R26350 D_FlipFlop_6.CLK.n7 D_FlipFlop_6.CLK.n6 0.0216397
R26351 D_FlipFlop_6.CLK.n6 D_FlipFlop_6.CLK 0.0216397
R26352 D_FlipFlop_6.CLK.n11 D_FlipFlop_6.CLK.n10 0.0180781
R26353 D_FlipFlop_6.CLK.n4 D_FlipFlop_6.CLK 0.00441667
R26354 D_FlipFlop_6.CLK.n4 D_FlipFlop_6.CLK 0.00406061
R26355 D_FlipFlop_7.D.t18 D_FlipFlop_7.D.n129 180.444
R26356 D_FlipFlop_7.D.n118 D_FlipFlop_7.D.t8 150.273
R26357 D_FlipFlop_7.D.n104 D_FlipFlop_7.D.t16 150.273
R26358 D_FlipFlop_7.D.n99 D_FlipFlop_7.D.t21 150.273
R26359 D_FlipFlop_7.D.n88 D_FlipFlop_7.D.t35 150.273
R26360 D_FlipFlop_7.D.n83 D_FlipFlop_7.D.t27 150.273
R26361 D_FlipFlop_7.D.n72 D_FlipFlop_7.D.t4 150.273
R26362 D_FlipFlop_7.D.n67 D_FlipFlop_7.D.t3 150.273
R26363 D_FlipFlop_7.D.n56 D_FlipFlop_7.D.t12 150.273
R26364 D_FlipFlop_7.D.n51 D_FlipFlop_7.D.t20 150.273
R26365 D_FlipFlop_7.D.n40 D_FlipFlop_7.D.t14 150.273
R26366 D_FlipFlop_7.D.n35 D_FlipFlop_7.D.t33 150.273
R26367 D_FlipFlop_7.D.n24 D_FlipFlop_7.D.t22 150.273
R26368 D_FlipFlop_7.D.n19 D_FlipFlop_7.D.t28 150.273
R26369 D_FlipFlop_7.D.n9 D_FlipFlop_7.D.t15 150.273
R26370 D_FlipFlop_7.D.n4 D_FlipFlop_7.D.t10 150.273
R26371 D_FlipFlop_7.D.n130 D_FlipFlop_7.D.t18 150.273
R26372 D_FlipFlop_7.D.n116 D_FlipFlop_7.D.t26 73.6406
R26373 D_FlipFlop_7.D.n97 D_FlipFlop_7.D.t7 73.6406
R26374 D_FlipFlop_7.D.n102 D_FlipFlop_7.D.t34 73.6406
R26375 D_FlipFlop_7.D.n81 D_FlipFlop_7.D.t13 73.6406
R26376 D_FlipFlop_7.D.n86 D_FlipFlop_7.D.t19 73.6406
R26377 D_FlipFlop_7.D.n65 D_FlipFlop_7.D.t32 73.6406
R26378 D_FlipFlop_7.D.n70 D_FlipFlop_7.D.t25 73.6406
R26379 D_FlipFlop_7.D.n49 D_FlipFlop_7.D.t6 73.6406
R26380 D_FlipFlop_7.D.n54 D_FlipFlop_7.D.t17 73.6406
R26381 D_FlipFlop_7.D.n33 D_FlipFlop_7.D.t24 73.6406
R26382 D_FlipFlop_7.D.n38 D_FlipFlop_7.D.t31 73.6406
R26383 D_FlipFlop_7.D.n17 D_FlipFlop_7.D.t5 73.6406
R26384 D_FlipFlop_7.D.n22 D_FlipFlop_7.D.t11 73.6406
R26385 D_FlipFlop_7.D.n2 D_FlipFlop_7.D.t30 73.6406
R26386 D_FlipFlop_7.D.n7 D_FlipFlop_7.D.t23 73.6406
R26387 D_FlipFlop_7.D.n0 D_FlipFlop_7.D.t9 73.6406
R26388 D_FlipFlop_7.D.n128 D_FlipFlop_7.D.t0 28.4497
R26389 D_FlipFlop_7.D.n32 D_FlipFlop_7.D.n16 28.2614
R26390 D_FlipFlop_7.D.n113 D_FlipFlop_7.D.n112 28.2614
R26391 D_FlipFlop_7.D.n129 D_FlipFlop_7.D.t1 25.7849
R26392 D_FlipFlop_7.D.n48 D_FlipFlop_7.D.n32 23.7614
R26393 D_FlipFlop_7.D.n64 D_FlipFlop_7.D.n48 23.7614
R26394 D_FlipFlop_7.D.n80 D_FlipFlop_7.D.n64 23.7614
R26395 D_FlipFlop_7.D.n96 D_FlipFlop_7.D.n80 23.7614
R26396 D_FlipFlop_7.D.n112 D_FlipFlop_7.D.n96 23.7614
R26397 D_FlipFlop_7.D.n122 D_FlipFlop_7.D.n121 12.6418
R26398 D_FlipFlop_7.D.n108 D_FlipFlop_7.D.n107 12.6418
R26399 D_FlipFlop_7.D.n92 D_FlipFlop_7.D.n91 12.6418
R26400 D_FlipFlop_7.D.n76 D_FlipFlop_7.D.n75 12.6418
R26401 D_FlipFlop_7.D.n60 D_FlipFlop_7.D.n59 12.6418
R26402 D_FlipFlop_7.D.n44 D_FlipFlop_7.D.n43 12.6418
R26403 D_FlipFlop_7.D.n28 D_FlipFlop_7.D.n27 12.6418
R26404 D_FlipFlop_7.D.n13 D_FlipFlop_7.D.n12 12.6418
R26405 D_FlipFlop_7.D.n129 D_FlipFlop_7.D.n128 7.83398
R26406 D_FlipFlop_7.D.n32 D_FlipFlop_7.D.n31 4.5005
R26407 D_FlipFlop_7.D.n48 D_FlipFlop_7.D.n47 4.5005
R26408 D_FlipFlop_7.D.n64 D_FlipFlop_7.D.n63 4.5005
R26409 D_FlipFlop_7.D.n80 D_FlipFlop_7.D.n79 4.5005
R26410 D_FlipFlop_7.D.n96 D_FlipFlop_7.D.n95 4.5005
R26411 D_FlipFlop_7.D.n112 D_FlipFlop_7.D.n111 4.5005
R26412 D_FlipFlop_7.D.n128 D_FlipFlop_7.D.n127 3.8456
R26413 D_FlipFlop_7.D.n125 D_FlipFlop_7.D.t29 1.13717
R26414 D_FlipFlop_7.D.n98 D_FlipFlop_1.Inverter_0.Vin 1.10104
R26415 D_FlipFlop_7.D.n82 D_FlipFlop_2.Inverter_0.Vin 1.10104
R26416 D_FlipFlop_7.D.n66 D_FlipFlop_3.Inverter_0.Vin 1.10104
R26417 D_FlipFlop_7.D.n50 D_FlipFlop_5.Inverter_0.Vin 1.10104
R26418 D_FlipFlop_7.D.n34 D_FlipFlop_4.Inverter_0.Vin 1.10104
R26419 D_FlipFlop_7.D.n18 D_FlipFlop_6.Inverter_0.Vin 1.10104
R26420 D_FlipFlop_7.D.n3 D_FlipFlop_7.Inverter_0.Vin 1.10104
R26421 D_FlipFlop_7.D.n1 D_FlipFlop_0.Inverter_0.Vin 1.10104
R26422 D_FlipFlop_7.D.n117 D_FlipFlop_0.3-input-nand_0.B 0.851043
R26423 D_FlipFlop_7.D.n103 D_FlipFlop_1.3-input-nand_0.B 0.851043
R26424 D_FlipFlop_7.D.n109 D_FlipFlop_1.Inverter_0.Vin 0.851043
R26425 D_FlipFlop_7.D.n87 D_FlipFlop_2.3-input-nand_0.B 0.851043
R26426 D_FlipFlop_7.D.n93 D_FlipFlop_2.Inverter_0.Vin 0.851043
R26427 D_FlipFlop_7.D.n71 D_FlipFlop_3.3-input-nand_0.B 0.851043
R26428 D_FlipFlop_7.D.n77 D_FlipFlop_3.Inverter_0.Vin 0.851043
R26429 D_FlipFlop_7.D.n55 D_FlipFlop_5.3-input-nand_0.B 0.851043
R26430 D_FlipFlop_7.D.n61 D_FlipFlop_5.Inverter_0.Vin 0.851043
R26431 D_FlipFlop_7.D.n39 D_FlipFlop_4.3-input-nand_0.B 0.851043
R26432 D_FlipFlop_7.D.n45 D_FlipFlop_4.Inverter_0.Vin 0.851043
R26433 D_FlipFlop_7.D.n23 D_FlipFlop_6.3-input-nand_0.B 0.851043
R26434 D_FlipFlop_7.D.n29 D_FlipFlop_6.Inverter_0.Vin 0.851043
R26435 D_FlipFlop_7.D.n8 D_FlipFlop_7.3-input-nand_0.B 0.851043
R26436 D_FlipFlop_7.D.n14 D_FlipFlop_7.Inverter_0.Vin 0.851043
R26437 D_FlipFlop_7.D.n115 D_FlipFlop_0.Inverter_0.Vin 0.851043
R26438 D_FlipFlop_7.D.n110 D_FlipFlop_1.Inverter_0.Vin 0.666516
R26439 D_FlipFlop_7.D.n94 D_FlipFlop_2.Inverter_0.Vin 0.666516
R26440 D_FlipFlop_7.D.n78 D_FlipFlop_3.Inverter_0.Vin 0.666516
R26441 D_FlipFlop_7.D.n62 D_FlipFlop_5.Inverter_0.Vin 0.666516
R26442 D_FlipFlop_7.D.n46 D_FlipFlop_4.Inverter_0.Vin 0.666516
R26443 D_FlipFlop_7.D.n30 D_FlipFlop_6.Inverter_0.Vin 0.666516
R26444 D_FlipFlop_7.D.n15 D_FlipFlop_7.Inverter_0.Vin 0.666516
R26445 D_FlipFlop_7.D.n114 D_FlipFlop_0.Inverter_0.Vin 0.666516
R26446 D_FlipFlop_7.D.n120 D_FlipFlop_7.D.n119 0.55213
R26447 D_FlipFlop_7.D.n106 D_FlipFlop_7.D.n105 0.55213
R26448 D_FlipFlop_7.D.n101 D_FlipFlop_7.D.n100 0.55213
R26449 D_FlipFlop_7.D.n90 D_FlipFlop_7.D.n89 0.55213
R26450 D_FlipFlop_7.D.n85 D_FlipFlop_7.D.n84 0.55213
R26451 D_FlipFlop_7.D.n74 D_FlipFlop_7.D.n73 0.55213
R26452 D_FlipFlop_7.D.n69 D_FlipFlop_7.D.n68 0.55213
R26453 D_FlipFlop_7.D.n58 D_FlipFlop_7.D.n57 0.55213
R26454 D_FlipFlop_7.D.n53 D_FlipFlop_7.D.n52 0.55213
R26455 D_FlipFlop_7.D.n42 D_FlipFlop_7.D.n41 0.55213
R26456 D_FlipFlop_7.D.n37 D_FlipFlop_7.D.n36 0.55213
R26457 D_FlipFlop_7.D.n26 D_FlipFlop_7.D.n25 0.55213
R26458 D_FlipFlop_7.D.n21 D_FlipFlop_7.D.n20 0.55213
R26459 D_FlipFlop_7.D.n11 D_FlipFlop_7.D.n10 0.55213
R26460 D_FlipFlop_7.D.n6 D_FlipFlop_7.D.n5 0.55213
R26461 D_FlipFlop_7.D.n124 D_FlipFlop_7.D.n123 0.55213
R26462 D_FlipFlop_7.D.n120 D_FlipFlop_0.3-input-nand_0.B 0.486828
R26463 D_FlipFlop_7.D.n106 D_FlipFlop_1.3-input-nand_0.B 0.486828
R26464 D_FlipFlop_7.D.n101 D_FlipFlop_1.Inverter_0.Vin 0.486828
R26465 D_FlipFlop_7.D.n90 D_FlipFlop_2.3-input-nand_0.B 0.486828
R26466 D_FlipFlop_7.D.n85 D_FlipFlop_2.Inverter_0.Vin 0.486828
R26467 D_FlipFlop_7.D.n74 D_FlipFlop_3.3-input-nand_0.B 0.486828
R26468 D_FlipFlop_7.D.n69 D_FlipFlop_3.Inverter_0.Vin 0.486828
R26469 D_FlipFlop_7.D.n58 D_FlipFlop_5.3-input-nand_0.B 0.486828
R26470 D_FlipFlop_7.D.n53 D_FlipFlop_5.Inverter_0.Vin 0.486828
R26471 D_FlipFlop_7.D.n42 D_FlipFlop_4.3-input-nand_0.B 0.486828
R26472 D_FlipFlop_7.D.n37 D_FlipFlop_4.Inverter_0.Vin 0.486828
R26473 D_FlipFlop_7.D.n26 D_FlipFlop_6.3-input-nand_0.B 0.486828
R26474 D_FlipFlop_7.D.n21 D_FlipFlop_6.Inverter_0.Vin 0.486828
R26475 D_FlipFlop_7.D.n11 D_FlipFlop_7.3-input-nand_0.B 0.486828
R26476 D_FlipFlop_7.D.n6 D_FlipFlop_7.Inverter_0.Vin 0.486828
R26477 D_FlipFlop_7.D.n123 D_FlipFlop_0.Inverter_0.Vin 0.486828
R26478 D_FlipFlop_7.D.n117 D_FlipFlop_7.D.n116 0.470609
R26479 D_FlipFlop_7.D.n103 D_FlipFlop_7.D.n102 0.470609
R26480 D_FlipFlop_7.D.n87 D_FlipFlop_7.D.n86 0.470609
R26481 D_FlipFlop_7.D.n71 D_FlipFlop_7.D.n70 0.470609
R26482 D_FlipFlop_7.D.n55 D_FlipFlop_7.D.n54 0.470609
R26483 D_FlipFlop_7.D.n39 D_FlipFlop_7.D.n38 0.470609
R26484 D_FlipFlop_7.D.n23 D_FlipFlop_7.D.n22 0.470609
R26485 D_FlipFlop_7.D.n8 D_FlipFlop_7.D.n7 0.470609
R26486 D_FlipFlop_7.D.n127 D_FlipFlop_7.D.t2 0.465687
R26487 D_FlipFlop_7.D.n127 D_FlipFlop_7.D.n126 0.386019
R26488 D_FlipFlop_7.D.n98 D_FlipFlop_7.D.n97 0.220609
R26489 D_FlipFlop_7.D.n82 D_FlipFlop_7.D.n81 0.220609
R26490 D_FlipFlop_7.D.n66 D_FlipFlop_7.D.n65 0.220609
R26491 D_FlipFlop_7.D.n50 D_FlipFlop_7.D.n49 0.220609
R26492 D_FlipFlop_7.D.n34 D_FlipFlop_7.D.n33 0.220609
R26493 D_FlipFlop_7.D.n18 D_FlipFlop_7.D.n17 0.220609
R26494 D_FlipFlop_7.D.n3 D_FlipFlop_7.D.n2 0.220609
R26495 D_FlipFlop_7.D.n1 D_FlipFlop_7.D.n0 0.220609
R26496 D_FlipFlop_7.D.n116 D_FlipFlop_0.3-input-nand_0.B 0.217464
R26497 D_FlipFlop_7.D.n97 D_FlipFlop_1.Inverter_0.Vin 0.217464
R26498 D_FlipFlop_7.D.n102 D_FlipFlop_1.3-input-nand_0.B 0.217464
R26499 D_FlipFlop_7.D.n81 D_FlipFlop_2.Inverter_0.Vin 0.217464
R26500 D_FlipFlop_7.D.n86 D_FlipFlop_2.3-input-nand_0.B 0.217464
R26501 D_FlipFlop_7.D.n65 D_FlipFlop_3.Inverter_0.Vin 0.217464
R26502 D_FlipFlop_7.D.n70 D_FlipFlop_3.3-input-nand_0.B 0.217464
R26503 D_FlipFlop_7.D.n49 D_FlipFlop_5.Inverter_0.Vin 0.217464
R26504 D_FlipFlop_7.D.n54 D_FlipFlop_5.3-input-nand_0.B 0.217464
R26505 D_FlipFlop_7.D.n33 D_FlipFlop_4.Inverter_0.Vin 0.217464
R26506 D_FlipFlop_7.D.n38 D_FlipFlop_4.3-input-nand_0.B 0.217464
R26507 D_FlipFlop_7.D.n17 D_FlipFlop_6.Inverter_0.Vin 0.217464
R26508 D_FlipFlop_7.D.n22 D_FlipFlop_6.3-input-nand_0.B 0.217464
R26509 D_FlipFlop_7.D.n2 D_FlipFlop_7.Inverter_0.Vin 0.217464
R26510 D_FlipFlop_7.D.n7 D_FlipFlop_7.3-input-nand_0.B 0.217464
R26511 D_FlipFlop_7.D.n0 D_FlipFlop_0.Inverter_0.Vin 0.217464
R26512 D_FlipFlop_7.D.n119 D_FlipFlop_0.3-input-nand_0.B 0.1255
R26513 D_FlipFlop_7.D.n105 D_FlipFlop_1.3-input-nand_0.B 0.1255
R26514 D_FlipFlop_7.D.n100 D_FlipFlop_1.Inverter_0.Vin 0.1255
R26515 D_FlipFlop_7.D.n89 D_FlipFlop_2.3-input-nand_0.B 0.1255
R26516 D_FlipFlop_7.D.n84 D_FlipFlop_2.Inverter_0.Vin 0.1255
R26517 D_FlipFlop_7.D.n73 D_FlipFlop_3.3-input-nand_0.B 0.1255
R26518 D_FlipFlop_7.D.n68 D_FlipFlop_3.Inverter_0.Vin 0.1255
R26519 D_FlipFlop_7.D.n57 D_FlipFlop_5.3-input-nand_0.B 0.1255
R26520 D_FlipFlop_7.D.n52 D_FlipFlop_5.Inverter_0.Vin 0.1255
R26521 D_FlipFlop_7.D.n41 D_FlipFlop_4.3-input-nand_0.B 0.1255
R26522 D_FlipFlop_7.D.n36 D_FlipFlop_4.Inverter_0.Vin 0.1255
R26523 D_FlipFlop_7.D.n25 D_FlipFlop_6.3-input-nand_0.B 0.1255
R26524 D_FlipFlop_7.D.n20 D_FlipFlop_6.Inverter_0.Vin 0.1255
R26525 D_FlipFlop_7.D.n10 D_FlipFlop_7.3-input-nand_0.B 0.1255
R26526 D_FlipFlop_7.D.n5 D_FlipFlop_7.Inverter_0.Vin 0.1255
R26527 D_FlipFlop_7.D.n124 D_FlipFlop_0.Inverter_0.Vin 0.1255
R26528 D_FlipFlop_7.D.n110 D_FlipFlop_7.D.n109 0.076587
R26529 D_FlipFlop_7.D.n94 D_FlipFlop_7.D.n93 0.076587
R26530 D_FlipFlop_7.D.n78 D_FlipFlop_7.D.n77 0.076587
R26531 D_FlipFlop_7.D.n62 D_FlipFlop_7.D.n61 0.076587
R26532 D_FlipFlop_7.D.n46 D_FlipFlop_7.D.n45 0.076587
R26533 D_FlipFlop_7.D.n30 D_FlipFlop_7.D.n29 0.076587
R26534 D_FlipFlop_7.D.n15 D_FlipFlop_7.D.n14 0.076587
R26535 D_FlipFlop_7.D.n115 D_FlipFlop_7.D.n114 0.076587
R26536 D_FlipFlop_7.D.n121 D_FlipFlop_7.D.n117 0.063
R26537 D_FlipFlop_7.D.n121 D_FlipFlop_7.D.n120 0.063
R26538 D_FlipFlop_7.D.n107 D_FlipFlop_7.D.n103 0.063
R26539 D_FlipFlop_7.D.n107 D_FlipFlop_7.D.n106 0.063
R26540 D_FlipFlop_7.D.n109 D_FlipFlop_7.D.n108 0.063
R26541 D_FlipFlop_7.D.n108 D_FlipFlop_7.D.n101 0.063
R26542 D_FlipFlop_7.D.n111 D_FlipFlop_7.D.n98 0.063
R26543 D_FlipFlop_7.D.n111 D_FlipFlop_7.D.n110 0.063
R26544 D_FlipFlop_7.D.n91 D_FlipFlop_7.D.n87 0.063
R26545 D_FlipFlop_7.D.n91 D_FlipFlop_7.D.n90 0.063
R26546 D_FlipFlop_7.D.n93 D_FlipFlop_7.D.n92 0.063
R26547 D_FlipFlop_7.D.n92 D_FlipFlop_7.D.n85 0.063
R26548 D_FlipFlop_7.D.n95 D_FlipFlop_7.D.n82 0.063
R26549 D_FlipFlop_7.D.n95 D_FlipFlop_7.D.n94 0.063
R26550 D_FlipFlop_7.D.n75 D_FlipFlop_7.D.n71 0.063
R26551 D_FlipFlop_7.D.n75 D_FlipFlop_7.D.n74 0.063
R26552 D_FlipFlop_7.D.n77 D_FlipFlop_7.D.n76 0.063
R26553 D_FlipFlop_7.D.n76 D_FlipFlop_7.D.n69 0.063
R26554 D_FlipFlop_7.D.n79 D_FlipFlop_7.D.n66 0.063
R26555 D_FlipFlop_7.D.n79 D_FlipFlop_7.D.n78 0.063
R26556 D_FlipFlop_7.D.n59 D_FlipFlop_7.D.n55 0.063
R26557 D_FlipFlop_7.D.n59 D_FlipFlop_7.D.n58 0.063
R26558 D_FlipFlop_7.D.n61 D_FlipFlop_7.D.n60 0.063
R26559 D_FlipFlop_7.D.n60 D_FlipFlop_7.D.n53 0.063
R26560 D_FlipFlop_7.D.n63 D_FlipFlop_7.D.n50 0.063
R26561 D_FlipFlop_7.D.n63 D_FlipFlop_7.D.n62 0.063
R26562 D_FlipFlop_7.D.n43 D_FlipFlop_7.D.n39 0.063
R26563 D_FlipFlop_7.D.n43 D_FlipFlop_7.D.n42 0.063
R26564 D_FlipFlop_7.D.n45 D_FlipFlop_7.D.n44 0.063
R26565 D_FlipFlop_7.D.n44 D_FlipFlop_7.D.n37 0.063
R26566 D_FlipFlop_7.D.n47 D_FlipFlop_7.D.n34 0.063
R26567 D_FlipFlop_7.D.n47 D_FlipFlop_7.D.n46 0.063
R26568 D_FlipFlop_7.D.n27 D_FlipFlop_7.D.n23 0.063
R26569 D_FlipFlop_7.D.n27 D_FlipFlop_7.D.n26 0.063
R26570 D_FlipFlop_7.D.n29 D_FlipFlop_7.D.n28 0.063
R26571 D_FlipFlop_7.D.n28 D_FlipFlop_7.D.n21 0.063
R26572 D_FlipFlop_7.D.n31 D_FlipFlop_7.D.n18 0.063
R26573 D_FlipFlop_7.D.n31 D_FlipFlop_7.D.n30 0.063
R26574 D_FlipFlop_7.D.n12 D_FlipFlop_7.D.n8 0.063
R26575 D_FlipFlop_7.D.n12 D_FlipFlop_7.D.n11 0.063
R26576 D_FlipFlop_7.D.n14 D_FlipFlop_7.D.n13 0.063
R26577 D_FlipFlop_7.D.n13 D_FlipFlop_7.D.n6 0.063
R26578 D_FlipFlop_7.D.n16 D_FlipFlop_7.D.n3 0.063
R26579 D_FlipFlop_7.D.n16 D_FlipFlop_7.D.n15 0.063
R26580 D_FlipFlop_7.D.n113 D_FlipFlop_7.D.n1 0.063
R26581 D_FlipFlop_7.D.n114 D_FlipFlop_7.D.n113 0.063
R26582 D_FlipFlop_7.D.n122 D_FlipFlop_7.D.n115 0.063
R26583 D_FlipFlop_7.D.n123 D_FlipFlop_7.D.n122 0.063
R26584 D_FlipFlop_7.D.n126 Comparator_0.Vout 0.0620344
R26585 D_FlipFlop_7.D.n126 D_FlipFlop_7.D.n125 0.0413995
R26586 D_FlipFlop_7.D.n119 D_FlipFlop_7.D.n118 0.0216397
R26587 D_FlipFlop_7.D.n118 D_FlipFlop_0.3-input-nand_0.B 0.0216397
R26588 D_FlipFlop_7.D.n105 D_FlipFlop_7.D.n104 0.0216397
R26589 D_FlipFlop_7.D.n104 D_FlipFlop_1.3-input-nand_0.B 0.0216397
R26590 D_FlipFlop_7.D.n100 D_FlipFlop_7.D.n99 0.0216397
R26591 D_FlipFlop_7.D.n99 D_FlipFlop_1.Inverter_0.Vin 0.0216397
R26592 D_FlipFlop_7.D.n89 D_FlipFlop_7.D.n88 0.0216397
R26593 D_FlipFlop_7.D.n88 D_FlipFlop_2.3-input-nand_0.B 0.0216397
R26594 D_FlipFlop_7.D.n84 D_FlipFlop_7.D.n83 0.0216397
R26595 D_FlipFlop_7.D.n83 D_FlipFlop_2.Inverter_0.Vin 0.0216397
R26596 D_FlipFlop_7.D.n73 D_FlipFlop_7.D.n72 0.0216397
R26597 D_FlipFlop_7.D.n72 D_FlipFlop_3.3-input-nand_0.B 0.0216397
R26598 D_FlipFlop_7.D.n68 D_FlipFlop_7.D.n67 0.0216397
R26599 D_FlipFlop_7.D.n67 D_FlipFlop_3.Inverter_0.Vin 0.0216397
R26600 D_FlipFlop_7.D.n57 D_FlipFlop_7.D.n56 0.0216397
R26601 D_FlipFlop_7.D.n56 D_FlipFlop_5.3-input-nand_0.B 0.0216397
R26602 D_FlipFlop_7.D.n52 D_FlipFlop_7.D.n51 0.0216397
R26603 D_FlipFlop_7.D.n51 D_FlipFlop_5.Inverter_0.Vin 0.0216397
R26604 D_FlipFlop_7.D.n41 D_FlipFlop_7.D.n40 0.0216397
R26605 D_FlipFlop_7.D.n40 D_FlipFlop_4.3-input-nand_0.B 0.0216397
R26606 D_FlipFlop_7.D.n36 D_FlipFlop_7.D.n35 0.0216397
R26607 D_FlipFlop_7.D.n35 D_FlipFlop_4.Inverter_0.Vin 0.0216397
R26608 D_FlipFlop_7.D.n25 D_FlipFlop_7.D.n24 0.0216397
R26609 D_FlipFlop_7.D.n24 D_FlipFlop_6.3-input-nand_0.B 0.0216397
R26610 D_FlipFlop_7.D.n20 D_FlipFlop_7.D.n19 0.0216397
R26611 D_FlipFlop_7.D.n19 D_FlipFlop_6.Inverter_0.Vin 0.0216397
R26612 D_FlipFlop_7.D.n10 D_FlipFlop_7.D.n9 0.0216397
R26613 D_FlipFlop_7.D.n9 D_FlipFlop_7.3-input-nand_0.B 0.0216397
R26614 D_FlipFlop_7.D.n5 D_FlipFlop_7.D.n4 0.0216397
R26615 D_FlipFlop_7.D.n4 D_FlipFlop_7.Inverter_0.Vin 0.0216397
R26616 D_FlipFlop_7.D.n130 D_FlipFlop_7.D.n124 0.0216397
R26617 D_FlipFlop_0.Inverter_0.Vin D_FlipFlop_7.D.n130 0.0216397
R26618 D_FlipFlop_7.D.n125 Comparator_0.Vout 0.0131087
R26619 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t4 316.762
R26620 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t0 169.195
R26621 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t3 150.887
R26622 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n2 150.273
R26623 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t5 74.951
R26624 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t2 73.6304
R26625 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t1 60.3943
R26626 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n6 12.0358
R26627 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n8 0.981478
R26628 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.769522
R26629 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n0 0.745065
R26630 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.580578
R26631 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n4 0.533109
R26632 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.428234
R26633 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.063
R26634 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.063
R26635 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n3 0.063
R26636 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n5 0.063
R26637 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.063
R26638 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n7 0.063
R26639 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n1 0.063
R26640 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 179.256
R26641 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 168.089
R26642 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 150.887
R26643 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 73.6304
R26644 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 60.3943
R26645 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 12.0358
R26646 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 1.05069
R26647 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 0.981478
R26648 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.769522
R26649 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 0.745065
R26650 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.580578
R26651 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 0.533109
R26652 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.428234
R26653 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.063
R26654 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 0.063
R26655 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 0.063
R26656 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.063
R26657 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 0.063
R26658 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 0.063
R26659 D_FlipFlop_3.nPRE.n39 D_FlipFlop_3.nPRE.t1 169.46
R26660 D_FlipFlop_3.nPRE.n38 D_FlipFlop_3.nPRE.t2 167.809
R26661 D_FlipFlop_3.nPRE.n39 D_FlipFlop_3.nPRE.t0 167.809
R26662 D_FlipFlop_3.nPRE.n22 D_FlipFlop_3.nPRE.t16 161.88
R26663 D_FlipFlop_3.nPRE D_FlipFlop_3.nPRE.t12 158.581
R26664 D_FlipFlop_3.nPRE.n35 D_FlipFlop_3.nPRE.t5 158.565
R26665 D_FlipFlop_3.nPRE.t5 D_FlipFlop_3.nPRE.n34 151.594
R26666 D_FlipFlop_3.nPRE.t16 D_FlipFlop_3.nPRE.n21 150.293
R26667 D_FlipFlop_3.nPRE.t12 D_FlipFlop_3.nPRE.n2 150.293
R26668 D_FlipFlop_3.nPRE.n26 D_FlipFlop_3.nPRE.t4 150.273
R26669 D_FlipFlop_3.nPRE.n23 D_FlipFlop_3.nPRE.t15 150.273
R26670 D_FlipFlop_3.nPRE.n13 D_FlipFlop_3.nPRE.t9 150.273
R26671 D_FlipFlop_3.nPRE.n7 D_FlipFlop_3.nPRE.t10 150.273
R26672 D_FlipFlop_3.nPRE D_FlipFlop_3.nPRE.t14 99.8701
R26673 D_FlipFlop_3.nPRE.n25 D_FlipFlop_3.nPRE.t7 74.163
R26674 D_FlipFlop_3.nPRE.t14 D_FlipFlop_3.nPRE.n30 74.163
R26675 D_FlipFlop_3.nPRE.n11 D_FlipFlop_3.nPRE.t6 73.6406
R26676 D_FlipFlop_3.nPRE.n5 D_FlipFlop_3.nPRE.t8 73.6406
R26677 D_FlipFlop_3.nPRE.n34 D_FlipFlop_3.nPRE.t11 73.6304
R26678 D_FlipFlop_3.nPRE.n19 D_FlipFlop_3.nPRE.t17 73.6304
R26679 D_FlipFlop_3.nPRE.n0 D_FlipFlop_3.nPRE.t13 73.6304
R26680 D_FlipFlop_3.nPRE.n41 D_FlipFlop_3.nPRE.t3 62.1634
R26681 D_FlipFlop_3.nPRE.n17 D_FlipFlop_3.nPRE.n10 15.5222
R26682 D_FlipFlop_3.nPRE.n29 D_FlipFlop_3.nPRE.n28 12.6418
R26683 D_FlipFlop_3.nPRE.n40 D_FlipFlop_3.nPRE.n39 11.4489
R26684 D_FlipFlop_3.nPRE.n22 D_FlipFlop_3.nPRE.n18 9.02465
R26685 D_FlipFlop_3.nPRE.n18 D_FlipFlop_3.nPRE.n17 8.24202
R26686 D_FlipFlop_3.nPRE.n38 D_FlipFlop_3.nPRE.n37 8.21389
R26687 D_FlipFlop_3.nPRE.n32 D_FlipFlop_3.nPRE.n22 4.66462
R26688 D_FlipFlop_3.nPRE.n17 D_FlipFlop_3.nPRE.n16 4.5005
R26689 D_FlipFlop_3.nPRE.n33 D_FlipFlop_3.nPRE 1.2047
R26690 D_FlipFlop_3.nPRE.n21 D_FlipFlop_3.nPRE.n20 1.19615
R26691 D_FlipFlop_3.nPRE.n2 D_FlipFlop_3.nPRE.n1 1.19615
R26692 D_FlipFlop_3.nPRE.n32 D_FlipFlop_3.nPRE.n31 0.922483
R26693 D_FlipFlop_3.nPRE.n25 D_FlipFlop_3.nPRE 0.851043
R26694 D_FlipFlop_3.nPRE.n30 D_FlipFlop_3.nPRE 0.851043
R26695 D_FlipFlop_3.nPRE.n12 D_FlipFlop_3.nPRE.n11 0.796696
R26696 D_FlipFlop_3.nPRE.n6 D_FlipFlop_3.nPRE.n5 0.796696
R26697 D_FlipFlop_3.nPRE.n4 D_FlipFlop_3.nPRE.n3 0.783833
R26698 D_FlipFlop_3.nPRE.n4 D_FlipFlop_3.nPRE 0.716182
R26699 D_FlipFlop_3.nPRE.n27 D_FlipFlop_3.nPRE.n26 0.61463
R26700 D_FlipFlop_3.nPRE.n24 D_FlipFlop_3.nPRE.n23 0.61463
R26701 D_FlipFlop_3.nPRE.n12 D_FlipFlop_3.nPRE 0.524957
R26702 D_FlipFlop_3.nPRE.n6 D_FlipFlop_3.nPRE 0.524957
R26703 D_FlipFlop_3.nPRE.n27 D_FlipFlop_3.nPRE 0.486828
R26704 D_FlipFlop_3.nPRE.n24 D_FlipFlop_3.nPRE 0.486828
R26705 D_FlipFlop_3.nPRE.n21 D_FlipFlop_3.nPRE 0.447191
R26706 D_FlipFlop_3.nPRE.n2 D_FlipFlop_3.nPRE 0.447191
R26707 D_FlipFlop_3.nPRE.n37 D_FlipFlop_3.nPRE.n36 0.425067
R26708 D_FlipFlop_3.nPRE.n33 D_FlipFlop_3.nPRE.n32 0.399217
R26709 D_FlipFlop_3.nPRE.n37 D_FlipFlop_3.nPRE 0.39003
R26710 D_FlipFlop_3.nPRE.n40 D_FlipFlop_3.nPRE.n38 0.280391
R26711 D_FlipFlop_3.nPRE.n15 D_FlipFlop_3.nPRE 0.252453
R26712 D_FlipFlop_3.nPRE.n9 D_FlipFlop_3.nPRE 0.252453
R26713 D_FlipFlop_3.nPRE.n15 D_FlipFlop_3.nPRE.n14 0.226043
R26714 D_FlipFlop_3.nPRE.n9 D_FlipFlop_3.nPRE.n8 0.226043
R26715 D_FlipFlop_3.nPRE.n11 D_FlipFlop_3.nPRE 0.217464
R26716 D_FlipFlop_3.nPRE.n5 D_FlipFlop_3.nPRE 0.217464
R26717 D_FlipFlop_3.nPRE.n41 D_FlipFlop_3.nPRE.n40 0.200143
R26718 D_FlipFlop_3.nPRE.n20 D_FlipFlop_3.nPRE 0.1255
R26719 D_FlipFlop_3.nPRE.n14 D_FlipFlop_3.nPRE 0.1255
R26720 D_FlipFlop_3.nPRE.n8 D_FlipFlop_3.nPRE 0.1255
R26721 D_FlipFlop_3.nPRE.n1 D_FlipFlop_3.nPRE 0.1255
R26722 D_FlipFlop_3.nPRE.n34 D_FlipFlop_3.nPRE 0.063
R26723 D_FlipFlop_3.nPRE.n26 D_FlipFlop_3.nPRE 0.063
R26724 D_FlipFlop_3.nPRE.n28 D_FlipFlop_3.nPRE.n25 0.063
R26725 D_FlipFlop_3.nPRE.n28 D_FlipFlop_3.nPRE.n27 0.063
R26726 D_FlipFlop_3.nPRE.n23 D_FlipFlop_3.nPRE 0.063
R26727 D_FlipFlop_3.nPRE.n30 D_FlipFlop_3.nPRE.n29 0.063
R26728 D_FlipFlop_3.nPRE.n29 D_FlipFlop_3.nPRE.n24 0.063
R26729 D_FlipFlop_3.nPRE.n16 D_FlipFlop_3.nPRE.n12 0.063
R26730 D_FlipFlop_3.nPRE.n16 D_FlipFlop_3.nPRE.n15 0.063
R26731 D_FlipFlop_3.nPRE.n10 D_FlipFlop_3.nPRE.n6 0.063
R26732 D_FlipFlop_3.nPRE.n10 D_FlipFlop_3.nPRE.n9 0.063
R26733 D_FlipFlop_3.nPRE D_FlipFlop_3.nPRE.n41 0.063
R26734 D_FlipFlop_3.nPRE.n18 D_FlipFlop_3.nPRE.n4 0.024
R26735 D_FlipFlop_3.nPRE.n35 D_FlipFlop_3.nPRE.n33 0.024
R26736 D_FlipFlop_3.nPRE.n14 D_FlipFlop_3.nPRE.n13 0.0216397
R26737 D_FlipFlop_3.nPRE.n13 D_FlipFlop_3.nPRE 0.0216397
R26738 D_FlipFlop_3.nPRE.n8 D_FlipFlop_3.nPRE.n7 0.0216397
R26739 D_FlipFlop_3.nPRE.n7 D_FlipFlop_3.nPRE 0.0216397
R26740 D_FlipFlop_3.nPRE D_FlipFlop_3.nPRE.n35 0.0204394
R26741 D_FlipFlop_3.nPRE.n20 D_FlipFlop_3.nPRE.n19 0.0107679
R26742 D_FlipFlop_3.nPRE.n19 D_FlipFlop_3.nPRE 0.0107679
R26743 D_FlipFlop_3.nPRE.n1 D_FlipFlop_3.nPRE.n0 0.0107679
R26744 D_FlipFlop_3.nPRE.n0 D_FlipFlop_3.nPRE 0.0107679
R26745 D_FlipFlop_3.nPRE.n3 D_FlipFlop_3.nPRE 0.00441667
R26746 D_FlipFlop_3.nPRE.n31 D_FlipFlop_3.nPRE 0.00441667
R26747 D_FlipFlop_3.nPRE.n36 D_FlipFlop_3.nPRE 0.00441667
R26748 D_FlipFlop_3.nPRE.n31 D_FlipFlop_3.nPRE 0.00406061
R26749 D_FlipFlop_3.nPRE.n3 D_FlipFlop_3.nPRE 0.00406061
R26750 D_FlipFlop_3.nPRE.n36 D_FlipFlop_3.nPRE 0.00406061
R26751 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 169.46
R26752 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 167.809
R26753 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 167.809
R26754 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 167.227
R26755 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 151.594
R26756 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 150.273
R26757 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 74.8641
R26758 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 73.6304
R26759 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 61.84
R26760 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 12.3891
R26761 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 11.4489
R26762 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 0.38637
R26763 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 0.280391
R26764 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 0.200143
R26765 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.152844
R26766 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.149957
R26767 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 0.149957
R26768 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.063
R26769 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.063
R26770 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 0.063
R26771 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 0.063
R26772 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.0454219
R26773 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t1 169.46
R26774 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t2 167.809
R26775 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t0 167.809
R26776 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n9 167.226
R26777 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t5 150.273
R26778 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t7 150.273
R26779 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t4 74.951
R26780 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t6 73.6304
R26781 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t3 60.3943
R26782 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n4 12.3891
R26783 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n7 11.4489
R26784 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 1.68257
R26785 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n0 1.44615
R26786 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n2 1.2342
R26787 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 1.08448
R26788 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.932141
R26789 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n6 0.3496
R26790 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n8 0.280391
R26791 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.063
R26792 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n3 0.063
R26793 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.063
R26794 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n5 0.063
R26795 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n1 0.063
R26796 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n10 0.063
R26797 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 169.46
R26798 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 167.809
R26799 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 167.809
R26800 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 167.227
R26801 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 151.594
R26802 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 150.273
R26803 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 74.8641
R26804 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 73.6304
R26805 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 61.84
R26806 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 12.3891
R26807 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 11.4489
R26808 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 0.38637
R26809 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 0.280391
R26810 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 0.200143
R26811 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.152844
R26812 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.149957
R26813 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 0.149957
R26814 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.063
R26815 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.063
R26816 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 0.063
R26817 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 0.063
R26818 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.0454219
R26819 D_FlipFlop_5.CLK.n12 D_FlipFlop_5.CLK.t0 168.108
R26820 D_FlipFlop_5.CLK.t3 D_FlipFlop_5.CLK.n5 158.207
R26821 D_FlipFlop_5.CLK D_FlipFlop_5.CLK.t4 158.202
R26822 D_FlipFlop_5.CLK.n0 D_FlipFlop_5.CLK.t5 150.293
R26823 D_FlipFlop_5.CLK.t4 D_FlipFlop_5.CLK.n3 150.293
R26824 D_FlipFlop_5.CLK.n6 D_FlipFlop_5.CLK.t3 150.273
R26825 D_FlipFlop_5.CLK.n9 D_FlipFlop_5.CLK.t2 90.1131
R26826 D_FlipFlop_5.CLK.t2 D_FlipFlop_5.CLK.n8 73.6406
R26827 D_FlipFlop_5.CLK.n2 D_FlipFlop_5.CLK.t6 73.6304
R26828 D_FlipFlop_5.CLK.n1 D_FlipFlop_5.CLK.t7 73.6304
R26829 D_FlipFlop_5.CLK D_FlipFlop_5.CLK.t1 60.3072
R26830 D_FlipFlop_5.CLK.n2 D_FlipFlop_5.CLK.n1 16.332
R26831 D_FlipFlop_5.CLK.n12 D_FlipFlop_5.CLK.n11 1.62007
R26832 D_FlipFlop_5.CLK.n8 D_FlipFlop_5.CLK.n7 1.19615
R26833 D_FlipFlop_5.CLK.n1 D_FlipFlop_5.CLK.n0 1.1717
R26834 D_FlipFlop_5.CLK.n3 D_FlipFlop_5.CLK.n2 1.1717
R26835 D_FlipFlop_5.CLK D_FlipFlop_5.CLK.n12 0.484875
R26836 D_FlipFlop_5.CLK.n3 D_FlipFlop_5.CLK 0.447191
R26837 D_FlipFlop_5.CLK.n0 D_FlipFlop_5.CLK 0.436162
R26838 D_FlipFlop_5.CLK.n5 D_FlipFlop_5.CLK.n4 0.349867
R26839 D_FlipFlop_5.CLK.n5 D_FlipFlop_5.CLK 0.321667
R26840 D_FlipFlop_5.CLK.n8 D_FlipFlop_5.CLK 0.217464
R26841 D_FlipFlop_5.CLK.n2 D_FlipFlop_5.CLK 0.149957
R26842 D_FlipFlop_5.CLK.n11 D_FlipFlop_5.CLK 0.149957
R26843 D_FlipFlop_5.CLK.n7 D_FlipFlop_5.CLK 0.1255
R26844 D_FlipFlop_5.CLK.n1 D_FlipFlop_5.CLK 0.117348
R26845 D_FlipFlop_5.CLK.n10 D_FlipFlop_5.CLK 0.0903438
R26846 D_FlipFlop_5.CLK.n1 D_FlipFlop_5.CLK 0.0454219
R26847 D_FlipFlop_5.CLK.n2 D_FlipFlop_5.CLK 0.0454219
R26848 D_FlipFlop_5.CLK.n10 D_FlipFlop_5.CLK.n9 0.027881
R26849 D_FlipFlop_5.CLK.n9 D_FlipFlop_5.CLK 0.027881
R26850 D_FlipFlop_5.CLK.n7 D_FlipFlop_5.CLK.n6 0.0216397
R26851 D_FlipFlop_5.CLK.n6 D_FlipFlop_5.CLK 0.0216397
R26852 D_FlipFlop_5.CLK.n11 D_FlipFlop_5.CLK.n10 0.0180781
R26853 D_FlipFlop_5.CLK.n4 D_FlipFlop_5.CLK 0.00441667
R26854 D_FlipFlop_5.CLK.n4 D_FlipFlop_5.CLK 0.00406061
R26855 D_FlipFlop_2.nPRE.n39 D_FlipFlop_2.nPRE.t3 169.46
R26856 D_FlipFlop_2.nPRE.n39 D_FlipFlop_2.nPRE.t2 167.809
R26857 D_FlipFlop_2.nPRE.n38 D_FlipFlop_2.nPRE.t0 167.809
R26858 D_FlipFlop_2.nPRE.n22 D_FlipFlop_2.nPRE.t17 162.52
R26859 D_FlipFlop_2.nPRE D_FlipFlop_2.nPRE.t14 158.581
R26860 D_FlipFlop_2.nPRE.n35 D_FlipFlop_2.nPRE.t7 158.565
R26861 D_FlipFlop_2.nPRE.t7 D_FlipFlop_2.nPRE.n34 151.594
R26862 D_FlipFlop_2.nPRE.t14 D_FlipFlop_2.nPRE.n5 150.293
R26863 D_FlipFlop_2.nPRE.t17 D_FlipFlop_2.nPRE.n2 150.293
R26864 D_FlipFlop_2.nPRE.n26 D_FlipFlop_2.nPRE.t5 150.273
R26865 D_FlipFlop_2.nPRE.n23 D_FlipFlop_2.nPRE.t16 150.273
R26866 D_FlipFlop_2.nPRE.n16 D_FlipFlop_2.nPRE.t15 150.273
R26867 D_FlipFlop_2.nPRE.n10 D_FlipFlop_2.nPRE.t4 150.273
R26868 D_FlipFlop_2.nPRE D_FlipFlop_2.nPRE.t12 99.8701
R26869 D_FlipFlop_2.nPRE.n25 D_FlipFlop_2.nPRE.t6 74.163
R26870 D_FlipFlop_2.nPRE.t12 D_FlipFlop_2.nPRE.n30 74.163
R26871 D_FlipFlop_2.nPRE.n14 D_FlipFlop_2.nPRE.t8 73.6406
R26872 D_FlipFlop_2.nPRE.n8 D_FlipFlop_2.nPRE.t11 73.6406
R26873 D_FlipFlop_2.nPRE.n34 D_FlipFlop_2.nPRE.t10 73.6304
R26874 D_FlipFlop_2.nPRE.n3 D_FlipFlop_2.nPRE.t9 73.6304
R26875 D_FlipFlop_2.nPRE.n0 D_FlipFlop_2.nPRE.t13 73.6304
R26876 D_FlipFlop_2.nPRE.n41 D_FlipFlop_2.nPRE.t1 62.1634
R26877 D_FlipFlop_2.nPRE.n20 D_FlipFlop_2.nPRE.n13 15.5222
R26878 D_FlipFlop_2.nPRE.n29 D_FlipFlop_2.nPRE.n28 12.6418
R26879 D_FlipFlop_2.nPRE.n40 D_FlipFlop_2.nPRE.n39 11.4489
R26880 D_FlipFlop_2.nPRE.n22 D_FlipFlop_2.nPRE.n21 8.37918
R26881 D_FlipFlop_2.nPRE.n21 D_FlipFlop_2.nPRE.n20 8.24202
R26882 D_FlipFlop_2.nPRE.n38 D_FlipFlop_2.nPRE.n37 8.21389
R26883 D_FlipFlop_2.nPRE.n20 D_FlipFlop_2.nPRE.n19 4.5005
R26884 D_FlipFlop_2.nPRE.n32 D_FlipFlop_2.nPRE.n22 4.03482
R26885 D_FlipFlop_2.nPRE.n33 D_FlipFlop_2.nPRE 1.2047
R26886 D_FlipFlop_2.nPRE.n5 D_FlipFlop_2.nPRE.n4 1.19615
R26887 D_FlipFlop_2.nPRE.n2 D_FlipFlop_2.nPRE.n1 1.19615
R26888 D_FlipFlop_2.nPRE.n32 D_FlipFlop_2.nPRE.n31 0.922483
R26889 D_FlipFlop_2.nPRE.n25 D_FlipFlop_2.nPRE 0.851043
R26890 D_FlipFlop_2.nPRE.n30 D_FlipFlop_2.nPRE 0.851043
R26891 D_FlipFlop_2.nPRE.n15 D_FlipFlop_2.nPRE.n14 0.796696
R26892 D_FlipFlop_2.nPRE.n9 D_FlipFlop_2.nPRE.n8 0.796696
R26893 D_FlipFlop_2.nPRE.n7 D_FlipFlop_2.nPRE.n6 0.783833
R26894 D_FlipFlop_2.nPRE.n7 D_FlipFlop_2.nPRE 0.716182
R26895 D_FlipFlop_2.nPRE.n27 D_FlipFlop_2.nPRE.n26 0.61463
R26896 D_FlipFlop_2.nPRE.n24 D_FlipFlop_2.nPRE.n23 0.61463
R26897 D_FlipFlop_2.nPRE.n15 D_FlipFlop_2.nPRE 0.524957
R26898 D_FlipFlop_2.nPRE.n9 D_FlipFlop_2.nPRE 0.524957
R26899 D_FlipFlop_2.nPRE.n27 D_FlipFlop_2.nPRE 0.486828
R26900 D_FlipFlop_2.nPRE.n24 D_FlipFlop_2.nPRE 0.486828
R26901 D_FlipFlop_2.nPRE.n5 D_FlipFlop_2.nPRE 0.447191
R26902 D_FlipFlop_2.nPRE.n2 D_FlipFlop_2.nPRE 0.447191
R26903 D_FlipFlop_2.nPRE.n37 D_FlipFlop_2.nPRE.n36 0.425067
R26904 D_FlipFlop_2.nPRE.n33 D_FlipFlop_2.nPRE.n32 0.399217
R26905 D_FlipFlop_2.nPRE.n37 D_FlipFlop_2.nPRE 0.39003
R26906 D_FlipFlop_2.nPRE.n40 D_FlipFlop_2.nPRE.n38 0.280391
R26907 D_FlipFlop_2.nPRE.n18 D_FlipFlop_2.nPRE 0.252453
R26908 D_FlipFlop_2.nPRE.n12 D_FlipFlop_2.nPRE 0.252453
R26909 D_FlipFlop_2.nPRE.n18 D_FlipFlop_2.nPRE.n17 0.226043
R26910 D_FlipFlop_2.nPRE.n12 D_FlipFlop_2.nPRE.n11 0.226043
R26911 D_FlipFlop_2.nPRE.n14 D_FlipFlop_2.nPRE 0.217464
R26912 D_FlipFlop_2.nPRE.n8 D_FlipFlop_2.nPRE 0.217464
R26913 D_FlipFlop_2.nPRE.n41 D_FlipFlop_2.nPRE.n40 0.200143
R26914 D_FlipFlop_2.nPRE.n17 D_FlipFlop_2.nPRE 0.1255
R26915 D_FlipFlop_2.nPRE.n11 D_FlipFlop_2.nPRE 0.1255
R26916 D_FlipFlop_2.nPRE.n4 D_FlipFlop_2.nPRE 0.1255
R26917 D_FlipFlop_2.nPRE.n1 D_FlipFlop_2.nPRE 0.1255
R26918 D_FlipFlop_2.nPRE.n34 D_FlipFlop_2.nPRE 0.063
R26919 D_FlipFlop_2.nPRE.n26 D_FlipFlop_2.nPRE 0.063
R26920 D_FlipFlop_2.nPRE.n28 D_FlipFlop_2.nPRE.n25 0.063
R26921 D_FlipFlop_2.nPRE.n28 D_FlipFlop_2.nPRE.n27 0.063
R26922 D_FlipFlop_2.nPRE.n23 D_FlipFlop_2.nPRE 0.063
R26923 D_FlipFlop_2.nPRE.n30 D_FlipFlop_2.nPRE.n29 0.063
R26924 D_FlipFlop_2.nPRE.n29 D_FlipFlop_2.nPRE.n24 0.063
R26925 D_FlipFlop_2.nPRE.n19 D_FlipFlop_2.nPRE.n15 0.063
R26926 D_FlipFlop_2.nPRE.n19 D_FlipFlop_2.nPRE.n18 0.063
R26927 D_FlipFlop_2.nPRE.n13 D_FlipFlop_2.nPRE.n9 0.063
R26928 D_FlipFlop_2.nPRE.n13 D_FlipFlop_2.nPRE.n12 0.063
R26929 D_FlipFlop_2.nPRE D_FlipFlop_2.nPRE.n41 0.063
R26930 D_FlipFlop_2.nPRE.n21 D_FlipFlop_2.nPRE.n7 0.024
R26931 D_FlipFlop_2.nPRE.n35 D_FlipFlop_2.nPRE.n33 0.024
R26932 D_FlipFlop_2.nPRE.n17 D_FlipFlop_2.nPRE.n16 0.0216397
R26933 D_FlipFlop_2.nPRE.n16 D_FlipFlop_2.nPRE 0.0216397
R26934 D_FlipFlop_2.nPRE.n11 D_FlipFlop_2.nPRE.n10 0.0216397
R26935 D_FlipFlop_2.nPRE.n10 D_FlipFlop_2.nPRE 0.0216397
R26936 D_FlipFlop_2.nPRE D_FlipFlop_2.nPRE.n35 0.0204394
R26937 D_FlipFlop_2.nPRE.n4 D_FlipFlop_2.nPRE.n3 0.0107679
R26938 D_FlipFlop_2.nPRE.n3 D_FlipFlop_2.nPRE 0.0107679
R26939 D_FlipFlop_2.nPRE.n1 D_FlipFlop_2.nPRE.n0 0.0107679
R26940 D_FlipFlop_2.nPRE.n0 D_FlipFlop_2.nPRE 0.0107679
R26941 D_FlipFlop_2.nPRE.n6 D_FlipFlop_2.nPRE 0.00441667
R26942 D_FlipFlop_2.nPRE.n31 D_FlipFlop_2.nPRE 0.00441667
R26943 D_FlipFlop_2.nPRE.n36 D_FlipFlop_2.nPRE 0.00441667
R26944 D_FlipFlop_2.nPRE.n31 D_FlipFlop_2.nPRE 0.00406061
R26945 D_FlipFlop_2.nPRE.n6 D_FlipFlop_2.nPRE 0.00406061
R26946 D_FlipFlop_2.nPRE.n36 D_FlipFlop_2.nPRE 0.00406061
R26947 CDAC_v3_0.switch_3.Z.n11 CDAC_v3_0.switch_3.Z.t11 168.075
R26948 CDAC_v3_0.switch_3.Z.n11 CDAC_v3_0.switch_3.Z.t0 168.075
R26949 CDAC_v3_0.switch_3.Z.n0 CDAC_v3_0.switch_3.Z.t10 60.6851
R26950 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_3.Z.t1 60.6226
R26951 CDAC_v3_0.switch_3.Z.n9 CDAC_v3_0.switch_3.Z.n8 43.6322
R26952 CDAC_v3_0.switch_3.Z.n8 CDAC_v3_0.switch_3.Z.n4 23.4184
R26953 CDAC_v3_0.switch_3.Z.n5 CDAC_v3_0.switch_3.Z.t8 7.92783
R26954 CDAC_v3_0.switch_3.Z.n2 CDAC_v3_0.switch_3.Z.t3 7.92783
R26955 CDAC_v3_0.switch_3.Z.n7 CDAC_v3_0.switch_3.Z.n6 7.62077
R26956 CDAC_v3_0.switch_3.Z.n6 CDAC_v3_0.switch_3.Z.n5 7.62077
R26957 CDAC_v3_0.switch_3.Z.n4 CDAC_v3_0.switch_3.Z.n3 7.62077
R26958 CDAC_v3_0.switch_3.Z.n3 CDAC_v3_0.switch_3.Z.n2 7.62077
R26959 CDAC_v3_0.switch_3.Z.n8 CDAC_v3_0.switch_3.Z.n7 6.83837
R26960 CDAC_v3_0.switch_3.Z.n12 CDAC_v3_0.switch_3.Z.n10 1.34289
R26961 CDAC_v3_0.switch_3.Z.n10 CDAC_v3_0.switch_3.Z 0.42713
R26962 CDAC_v3_0.switch_3.Z.n5 CDAC_v3_0.switch_3.Z.t9 0.307567
R26963 CDAC_v3_0.switch_3.Z.n6 CDAC_v3_0.switch_3.Z.t4 0.307567
R26964 CDAC_v3_0.switch_3.Z.n7 CDAC_v3_0.switch_3.Z.t5 0.307567
R26965 CDAC_v3_0.switch_3.Z.n4 CDAC_v3_0.switch_3.Z.t7 0.307567
R26966 CDAC_v3_0.switch_3.Z.n3 CDAC_v3_0.switch_3.Z.t6 0.307567
R26967 CDAC_v3_0.switch_3.Z.n2 CDAC_v3_0.switch_3.Z.t2 0.307567
R26968 CDAC_v3_0.switch_3.Z.n1 CDAC_v3_0.switch_3.Z 0.182141
R26969 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_3.Z.n12 0.178175
R26970 CDAC_v3_0.switch_3.Z.n1 CDAC_v3_0.switch_3.Z.n0 0.128217
R26971 CDAC_v3_0.switch_3.Z.n0 CDAC_v3_0.switch_3.Z 0.1255
R26972 CDAC_v3_0.switch_3.Z.n0 CDAC_v3_0.switch_3.Z 0.063
R26973 CDAC_v3_0.switch_3.Z.n10 CDAC_v3_0.switch_3.Z.n9 0.063
R26974 CDAC_v3_0.switch_3.Z.n9 CDAC_v3_0.switch_3.Z.n1 0.063
R26975 CDAC_v3_0.switch_3.Z.n12 CDAC_v3_0.switch_3.Z.n11 0.0130546
R26976 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t4 316.762
R26977 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t0 169.195
R26978 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t3 150.887
R26979 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n2 150.273
R26980 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t2 74.951
R26981 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t5 73.6304
R26982 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t1 60.3943
R26983 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n6 12.0358
R26984 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n8 0.981478
R26985 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.769522
R26986 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n0 0.745065
R26987 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.580578
R26988 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n4 0.533109
R26989 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.428234
R26990 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.063
R26991 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.063
R26992 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n3 0.063
R26993 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n5 0.063
R26994 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.063
R26995 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n7 0.063
R26996 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n1 0.063
R26997 D_FlipFlop_4.nPRE.n39 D_FlipFlop_4.nPRE.t2 169.46
R26998 D_FlipFlop_4.nPRE.n39 D_FlipFlop_4.nPRE.t1 167.809
R26999 D_FlipFlop_4.nPRE.n38 D_FlipFlop_4.nPRE.t3 167.809
R27000 D_FlipFlop_4.nPRE.n22 D_FlipFlop_4.nPRE.t16 161.88
R27001 D_FlipFlop_4.nPRE D_FlipFlop_4.nPRE.t12 158.581
R27002 D_FlipFlop_4.nPRE.n35 D_FlipFlop_4.nPRE.t4 158.565
R27003 D_FlipFlop_4.nPRE.t4 D_FlipFlop_4.nPRE.n34 151.594
R27004 D_FlipFlop_4.nPRE.t16 D_FlipFlop_4.nPRE.n21 150.293
R27005 D_FlipFlop_4.nPRE.t12 D_FlipFlop_4.nPRE.n2 150.293
R27006 D_FlipFlop_4.nPRE.n26 D_FlipFlop_4.nPRE.t11 150.273
R27007 D_FlipFlop_4.nPRE.n23 D_FlipFlop_4.nPRE.t6 150.273
R27008 D_FlipFlop_4.nPRE.n13 D_FlipFlop_4.nPRE.t7 150.273
R27009 D_FlipFlop_4.nPRE.n7 D_FlipFlop_4.nPRE.t13 150.273
R27010 D_FlipFlop_4.nPRE D_FlipFlop_4.nPRE.t15 99.8701
R27011 D_FlipFlop_4.nPRE.n25 D_FlipFlop_4.nPRE.t10 74.163
R27012 D_FlipFlop_4.nPRE.t15 D_FlipFlop_4.nPRE.n30 74.163
R27013 D_FlipFlop_4.nPRE.n11 D_FlipFlop_4.nPRE.t5 73.6406
R27014 D_FlipFlop_4.nPRE.n5 D_FlipFlop_4.nPRE.t8 73.6406
R27015 D_FlipFlop_4.nPRE.n34 D_FlipFlop_4.nPRE.t9 73.6304
R27016 D_FlipFlop_4.nPRE.n19 D_FlipFlop_4.nPRE.t17 73.6304
R27017 D_FlipFlop_4.nPRE.n0 D_FlipFlop_4.nPRE.t14 73.6304
R27018 D_FlipFlop_4.nPRE.n41 D_FlipFlop_4.nPRE.t0 62.1634
R27019 D_FlipFlop_4.nPRE.n17 D_FlipFlop_4.nPRE.n10 15.5222
R27020 D_FlipFlop_4.nPRE.n29 D_FlipFlop_4.nPRE.n28 12.6418
R27021 D_FlipFlop_4.nPRE.n40 D_FlipFlop_4.nPRE.n39 11.4489
R27022 D_FlipFlop_4.nPRE.n22 D_FlipFlop_4.nPRE.n18 9.02465
R27023 D_FlipFlop_4.nPRE.n18 D_FlipFlop_4.nPRE.n17 8.24202
R27024 D_FlipFlop_4.nPRE.n38 D_FlipFlop_4.nPRE.n37 8.21389
R27025 D_FlipFlop_4.nPRE.n32 D_FlipFlop_4.nPRE.n22 7.22455
R27026 D_FlipFlop_4.nPRE.n17 D_FlipFlop_4.nPRE.n16 4.5005
R27027 D_FlipFlop_4.nPRE.n33 D_FlipFlop_4.nPRE 1.2047
R27028 D_FlipFlop_4.nPRE.n21 D_FlipFlop_4.nPRE.n20 1.19615
R27029 D_FlipFlop_4.nPRE.n2 D_FlipFlop_4.nPRE.n1 1.19615
R27030 D_FlipFlop_4.nPRE.n32 D_FlipFlop_4.nPRE.n31 0.922483
R27031 D_FlipFlop_4.nPRE.n25 D_FlipFlop_4.nPRE 0.851043
R27032 D_FlipFlop_4.nPRE.n30 D_FlipFlop_4.nPRE 0.851043
R27033 D_FlipFlop_4.nPRE.n12 D_FlipFlop_4.nPRE.n11 0.796696
R27034 D_FlipFlop_4.nPRE.n6 D_FlipFlop_4.nPRE.n5 0.796696
R27035 D_FlipFlop_4.nPRE.n4 D_FlipFlop_4.nPRE.n3 0.783833
R27036 D_FlipFlop_4.nPRE.n4 D_FlipFlop_4.nPRE 0.716182
R27037 D_FlipFlop_4.nPRE.n27 D_FlipFlop_4.nPRE.n26 0.61463
R27038 D_FlipFlop_4.nPRE.n24 D_FlipFlop_4.nPRE.n23 0.61463
R27039 D_FlipFlop_4.nPRE.n12 D_FlipFlop_4.nPRE 0.524957
R27040 D_FlipFlop_4.nPRE.n6 D_FlipFlop_4.nPRE 0.524957
R27041 D_FlipFlop_4.nPRE.n27 D_FlipFlop_4.nPRE 0.486828
R27042 D_FlipFlop_4.nPRE.n24 D_FlipFlop_4.nPRE 0.486828
R27043 D_FlipFlop_4.nPRE.n21 D_FlipFlop_4.nPRE 0.447191
R27044 D_FlipFlop_4.nPRE.n2 D_FlipFlop_4.nPRE 0.447191
R27045 D_FlipFlop_4.nPRE.n37 D_FlipFlop_4.nPRE.n36 0.425067
R27046 D_FlipFlop_4.nPRE.n33 D_FlipFlop_4.nPRE.n32 0.399217
R27047 D_FlipFlop_4.nPRE.n37 D_FlipFlop_4.nPRE 0.39003
R27048 D_FlipFlop_4.nPRE.n40 D_FlipFlop_4.nPRE.n38 0.280391
R27049 D_FlipFlop_4.nPRE.n15 D_FlipFlop_4.nPRE 0.252453
R27050 D_FlipFlop_4.nPRE.n9 D_FlipFlop_4.nPRE 0.252453
R27051 D_FlipFlop_4.nPRE.n15 D_FlipFlop_4.nPRE.n14 0.226043
R27052 D_FlipFlop_4.nPRE.n9 D_FlipFlop_4.nPRE.n8 0.226043
R27053 D_FlipFlop_4.nPRE.n11 D_FlipFlop_4.nPRE 0.217464
R27054 D_FlipFlop_4.nPRE.n5 D_FlipFlop_4.nPRE 0.217464
R27055 D_FlipFlop_4.nPRE.n41 D_FlipFlop_4.nPRE.n40 0.200143
R27056 D_FlipFlop_4.nPRE.n20 D_FlipFlop_4.nPRE 0.1255
R27057 D_FlipFlop_4.nPRE.n14 D_FlipFlop_4.nPRE 0.1255
R27058 D_FlipFlop_4.nPRE.n8 D_FlipFlop_4.nPRE 0.1255
R27059 D_FlipFlop_4.nPRE.n1 D_FlipFlop_4.nPRE 0.1255
R27060 D_FlipFlop_4.nPRE.n34 D_FlipFlop_4.nPRE 0.063
R27061 D_FlipFlop_4.nPRE.n26 D_FlipFlop_4.nPRE 0.063
R27062 D_FlipFlop_4.nPRE.n28 D_FlipFlop_4.nPRE.n25 0.063
R27063 D_FlipFlop_4.nPRE.n28 D_FlipFlop_4.nPRE.n27 0.063
R27064 D_FlipFlop_4.nPRE.n23 D_FlipFlop_4.nPRE 0.063
R27065 D_FlipFlop_4.nPRE.n30 D_FlipFlop_4.nPRE.n29 0.063
R27066 D_FlipFlop_4.nPRE.n29 D_FlipFlop_4.nPRE.n24 0.063
R27067 D_FlipFlop_4.nPRE.n16 D_FlipFlop_4.nPRE.n12 0.063
R27068 D_FlipFlop_4.nPRE.n16 D_FlipFlop_4.nPRE.n15 0.063
R27069 D_FlipFlop_4.nPRE.n10 D_FlipFlop_4.nPRE.n6 0.063
R27070 D_FlipFlop_4.nPRE.n10 D_FlipFlop_4.nPRE.n9 0.063
R27071 D_FlipFlop_4.nPRE D_FlipFlop_4.nPRE.n41 0.063
R27072 D_FlipFlop_4.nPRE.n18 D_FlipFlop_4.nPRE.n4 0.024
R27073 D_FlipFlop_4.nPRE.n35 D_FlipFlop_4.nPRE.n33 0.024
R27074 D_FlipFlop_4.nPRE.n14 D_FlipFlop_4.nPRE.n13 0.0216397
R27075 D_FlipFlop_4.nPRE.n13 D_FlipFlop_4.nPRE 0.0216397
R27076 D_FlipFlop_4.nPRE.n8 D_FlipFlop_4.nPRE.n7 0.0216397
R27077 D_FlipFlop_4.nPRE.n7 D_FlipFlop_4.nPRE 0.0216397
R27078 D_FlipFlop_4.nPRE D_FlipFlop_4.nPRE.n35 0.0204394
R27079 D_FlipFlop_4.nPRE.n20 D_FlipFlop_4.nPRE.n19 0.0107679
R27080 D_FlipFlop_4.nPRE.n19 D_FlipFlop_4.nPRE 0.0107679
R27081 D_FlipFlop_4.nPRE.n1 D_FlipFlop_4.nPRE.n0 0.0107679
R27082 D_FlipFlop_4.nPRE.n0 D_FlipFlop_4.nPRE 0.0107679
R27083 D_FlipFlop_4.nPRE.n3 D_FlipFlop_4.nPRE 0.00441667
R27084 D_FlipFlop_4.nPRE.n31 D_FlipFlop_4.nPRE 0.00441667
R27085 D_FlipFlop_4.nPRE.n36 D_FlipFlop_4.nPRE 0.00441667
R27086 D_FlipFlop_4.nPRE.n31 D_FlipFlop_4.nPRE 0.00406061
R27087 D_FlipFlop_4.nPRE.n3 D_FlipFlop_4.nPRE 0.00406061
R27088 D_FlipFlop_4.nPRE.n36 D_FlipFlop_4.nPRE 0.00406061
R27089 Ring_Counter_0.D_FlipFlop_10.Qbar.n4 Ring_Counter_0.D_FlipFlop_10.Qbar.t1 169.46
R27090 Ring_Counter_0.D_FlipFlop_10.Qbar.n3 Ring_Counter_0.D_FlipFlop_10.Qbar.t2 167.809
R27091 Ring_Counter_0.D_FlipFlop_10.Qbar.n4 Ring_Counter_0.D_FlipFlop_10.Qbar.t0 167.809
R27092 Ring_Counter_0.D_FlipFlop_10.Qbar.n1 Ring_Counter_0.D_FlipFlop_10.Qbar.t5 158.28
R27093 Ring_Counter_0.D_FlipFlop_10.Qbar.t5 Ring_Counter_0.D_FlipFlop_10.Qbar.n0 150.273
R27094 Ring_Counter_0.D_FlipFlop_10.Qbar.n0 Ring_Counter_0.D_FlipFlop_10.Qbar.t4 74.951
R27095 Ring_Counter_0.D_FlipFlop_10.Qbar.n6 Ring_Counter_0.D_FlipFlop_10.Qbar.t3 60.3943
R27096 Ring_Counter_0.D_FlipFlop_10.Qbar.n5 Ring_Counter_0.D_FlipFlop_10.Qbar.n4 11.4489
R27097 Ring_Counter_0.D_FlipFlop_10.Qbar.n3 Ring_Counter_0.D_FlipFlop_10.Qbar 8.5174
R27098 Ring_Counter_0.D_FlipFlop_10.Qbar.n6 Ring_Counter_0.D_FlipFlop_10.Qbar.n5 1.96917
R27099 Ring_Counter_0.D_FlipFlop_10.Qbar.n2 Ring_Counter_0.D_FlipFlop_10.Qbar.n1 0.42585
R27100 Ring_Counter_0.D_FlipFlop_10.Qbar.n1 Ring_Counter_0.D_FlipFlop_10.Qbar 0.390742
R27101 Ring_Counter_0.D_FlipFlop_10.Qbar.n5 Ring_Counter_0.D_FlipFlop_10.Qbar.n3 0.280391
R27102 Ring_Counter_0.D_FlipFlop_10.Qbar.n0 Ring_Counter_0.D_FlipFlop_10.Qbar 0.063
R27103 Ring_Counter_0.D_FlipFlop_10.Qbar Ring_Counter_0.D_FlipFlop_10.Qbar.n6 0.063
R27104 Ring_Counter_0.D_FlipFlop_10.Qbar.n2 Ring_Counter_0.D_FlipFlop_10.Qbar 0.00441667
R27105 Ring_Counter_0.D_FlipFlop_10.Qbar Ring_Counter_0.D_FlipFlop_10.Qbar.n2 0.00406061
R27106 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t3 169.46
R27107 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t1 168.089
R27108 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n7 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t0 167.809
R27109 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t5 150.273
R27110 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t4 74.163
R27111 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t2 61.1389
R27112 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n4 12.0358
R27113 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n8 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n7 11.4489
R27114 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n0 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 1.08746
R27115 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n1 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.851043
R27116 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n9 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n6 0.851043
R27117 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.65675
R27118 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n2 0.61463
R27119 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n3 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.486828
R27120 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n9 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n8 0.200143
R27121 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n2 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.063
R27122 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n1 0.063
R27123 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n4 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n3 0.063
R27124 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n5 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n0 0.063
R27125 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n6 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n5 0.063
R27126 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n9 0.063
R27127 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t1 169.46
R27128 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R27129 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t0 167.809
R27130 D_FlipFlop_2.3-input-nand_2.C.t5 D_FlipFlop_2.3-input-nand_2.C.n13 167.226
R27131 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C.t4 150.273
R27132 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.t5 150.273
R27133 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C.t7 73.6406
R27134 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C.t6 73.6304
R27135 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.C.t3 60.3943
R27136 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C.n7 12.3891
R27137 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.n11 11.4489
R27138 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C 1.68257
R27139 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C.n2 1.38365
R27140 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C.n0 1.19615
R27141 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C.n5 1.1717
R27142 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C 1.08448
R27143 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C 0.932141
R27144 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C 0.720633
R27145 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.n12 0.280391
R27146 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C 0.217464
R27147 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27148 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27149 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C 0.1255
R27150 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C.n9 0.0874565
R27151 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C.n6 0.063
R27152 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C 0.063
R27153 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C.n8 0.063
R27154 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C.n3 0.063
R27155 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.n10 0.0435206
R27156 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.n1 0.0216397
R27157 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.C.n14 0.0216397
R27158 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C.n4 0.0107679
R27159 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C 0.0107679
R27160 D_FlipFlop_7.nPRE.n39 D_FlipFlop_7.nPRE.t2 169.46
R27161 D_FlipFlop_7.nPRE.n39 D_FlipFlop_7.nPRE.t1 167.809
R27162 D_FlipFlop_7.nPRE.n38 D_FlipFlop_7.nPRE.t3 167.809
R27163 D_FlipFlop_7.nPRE.n22 D_FlipFlop_7.nPRE.t6 161.88
R27164 D_FlipFlop_7.nPRE D_FlipFlop_7.nPRE.t10 158.581
R27165 D_FlipFlop_7.nPRE.n35 D_FlipFlop_7.nPRE.t7 158.565
R27166 D_FlipFlop_7.nPRE.t7 D_FlipFlop_7.nPRE.n34 151.594
R27167 D_FlipFlop_7.nPRE.t6 D_FlipFlop_7.nPRE.n21 150.293
R27168 D_FlipFlop_7.nPRE.t10 D_FlipFlop_7.nPRE.n2 150.293
R27169 D_FlipFlop_7.nPRE.n26 D_FlipFlop_7.nPRE.t13 150.273
R27170 D_FlipFlop_7.nPRE.n23 D_FlipFlop_7.nPRE.t8 150.273
R27171 D_FlipFlop_7.nPRE.n13 D_FlipFlop_7.nPRE.t15 150.273
R27172 D_FlipFlop_7.nPRE.n7 D_FlipFlop_7.nPRE.t12 150.273
R27173 D_FlipFlop_7.nPRE D_FlipFlop_7.nPRE.t9 99.8701
R27174 D_FlipFlop_7.nPRE.n25 D_FlipFlop_7.nPRE.t16 74.163
R27175 D_FlipFlop_7.nPRE.t9 D_FlipFlop_7.nPRE.n30 74.163
R27176 D_FlipFlop_7.nPRE.n11 D_FlipFlop_7.nPRE.t11 73.6406
R27177 D_FlipFlop_7.nPRE.n5 D_FlipFlop_7.nPRE.t5 73.6406
R27178 D_FlipFlop_7.nPRE.n34 D_FlipFlop_7.nPRE.t17 73.6304
R27179 D_FlipFlop_7.nPRE.n19 D_FlipFlop_7.nPRE.t14 73.6304
R27180 D_FlipFlop_7.nPRE.n0 D_FlipFlop_7.nPRE.t4 73.6304
R27181 D_FlipFlop_7.nPRE.n41 D_FlipFlop_7.nPRE.t0 62.1634
R27182 D_FlipFlop_7.nPRE.n17 D_FlipFlop_7.nPRE.n10 15.5222
R27183 D_FlipFlop_7.nPRE.n29 D_FlipFlop_7.nPRE.n28 12.6418
R27184 D_FlipFlop_7.nPRE.n40 D_FlipFlop_7.nPRE.n39 11.4489
R27185 D_FlipFlop_7.nPRE.n32 D_FlipFlop_7.nPRE.n22 9.78448
R27186 D_FlipFlop_7.nPRE.n22 D_FlipFlop_7.nPRE.n18 9.02465
R27187 D_FlipFlop_7.nPRE.n18 D_FlipFlop_7.nPRE.n17 8.24202
R27188 D_FlipFlop_7.nPRE.n38 D_FlipFlop_7.nPRE.n37 8.21389
R27189 D_FlipFlop_7.nPRE.n17 D_FlipFlop_7.nPRE.n16 4.5005
R27190 D_FlipFlop_7.nPRE.n33 D_FlipFlop_7.nPRE 1.2047
R27191 D_FlipFlop_7.nPRE.n21 D_FlipFlop_7.nPRE.n20 1.19615
R27192 D_FlipFlop_7.nPRE.n2 D_FlipFlop_7.nPRE.n1 1.19615
R27193 D_FlipFlop_7.nPRE.n32 D_FlipFlop_7.nPRE.n31 0.922483
R27194 D_FlipFlop_7.nPRE.n25 D_FlipFlop_7.nPRE 0.851043
R27195 D_FlipFlop_7.nPRE.n30 D_FlipFlop_7.nPRE 0.851043
R27196 D_FlipFlop_7.nPRE.n12 D_FlipFlop_7.nPRE.n11 0.796696
R27197 D_FlipFlop_7.nPRE.n6 D_FlipFlop_7.nPRE.n5 0.796696
R27198 D_FlipFlop_7.nPRE.n4 D_FlipFlop_7.nPRE.n3 0.783833
R27199 D_FlipFlop_7.nPRE.n4 D_FlipFlop_7.nPRE 0.716182
R27200 D_FlipFlop_7.nPRE.n27 D_FlipFlop_7.nPRE.n26 0.61463
R27201 D_FlipFlop_7.nPRE.n24 D_FlipFlop_7.nPRE.n23 0.61463
R27202 D_FlipFlop_7.nPRE.n12 D_FlipFlop_7.nPRE 0.524957
R27203 D_FlipFlop_7.nPRE.n6 D_FlipFlop_7.nPRE 0.524957
R27204 D_FlipFlop_7.nPRE.n27 D_FlipFlop_7.nPRE 0.486828
R27205 D_FlipFlop_7.nPRE.n24 D_FlipFlop_7.nPRE 0.486828
R27206 D_FlipFlop_7.nPRE.n21 D_FlipFlop_7.nPRE 0.447191
R27207 D_FlipFlop_7.nPRE.n2 D_FlipFlop_7.nPRE 0.447191
R27208 D_FlipFlop_7.nPRE.n37 D_FlipFlop_7.nPRE.n36 0.425067
R27209 D_FlipFlop_7.nPRE.n33 D_FlipFlop_7.nPRE.n32 0.399217
R27210 D_FlipFlop_7.nPRE.n37 D_FlipFlop_7.nPRE 0.39003
R27211 D_FlipFlop_7.nPRE.n40 D_FlipFlop_7.nPRE.n38 0.280391
R27212 D_FlipFlop_7.nPRE.n15 D_FlipFlop_7.nPRE 0.252453
R27213 D_FlipFlop_7.nPRE.n9 D_FlipFlop_7.nPRE 0.252453
R27214 D_FlipFlop_7.nPRE.n15 D_FlipFlop_7.nPRE.n14 0.226043
R27215 D_FlipFlop_7.nPRE.n9 D_FlipFlop_7.nPRE.n8 0.226043
R27216 D_FlipFlop_7.nPRE.n11 D_FlipFlop_7.nPRE 0.217464
R27217 D_FlipFlop_7.nPRE.n5 D_FlipFlop_7.nPRE 0.217464
R27218 D_FlipFlop_7.nPRE.n41 D_FlipFlop_7.nPRE.n40 0.200143
R27219 D_FlipFlop_7.nPRE.n20 D_FlipFlop_7.nPRE 0.1255
R27220 D_FlipFlop_7.nPRE.n14 D_FlipFlop_7.nPRE 0.1255
R27221 D_FlipFlop_7.nPRE.n8 D_FlipFlop_7.nPRE 0.1255
R27222 D_FlipFlop_7.nPRE.n1 D_FlipFlop_7.nPRE 0.1255
R27223 D_FlipFlop_7.nPRE.n34 D_FlipFlop_7.nPRE 0.063
R27224 D_FlipFlop_7.nPRE.n26 D_FlipFlop_7.nPRE 0.063
R27225 D_FlipFlop_7.nPRE.n28 D_FlipFlop_7.nPRE.n25 0.063
R27226 D_FlipFlop_7.nPRE.n28 D_FlipFlop_7.nPRE.n27 0.063
R27227 D_FlipFlop_7.nPRE.n23 D_FlipFlop_7.nPRE 0.063
R27228 D_FlipFlop_7.nPRE.n30 D_FlipFlop_7.nPRE.n29 0.063
R27229 D_FlipFlop_7.nPRE.n29 D_FlipFlop_7.nPRE.n24 0.063
R27230 D_FlipFlop_7.nPRE.n16 D_FlipFlop_7.nPRE.n12 0.063
R27231 D_FlipFlop_7.nPRE.n16 D_FlipFlop_7.nPRE.n15 0.063
R27232 D_FlipFlop_7.nPRE.n10 D_FlipFlop_7.nPRE.n6 0.063
R27233 D_FlipFlop_7.nPRE.n10 D_FlipFlop_7.nPRE.n9 0.063
R27234 D_FlipFlop_7.nPRE D_FlipFlop_7.nPRE.n41 0.063
R27235 D_FlipFlop_7.nPRE.n18 D_FlipFlop_7.nPRE.n4 0.024
R27236 D_FlipFlop_7.nPRE.n35 D_FlipFlop_7.nPRE.n33 0.024
R27237 D_FlipFlop_7.nPRE.n14 D_FlipFlop_7.nPRE.n13 0.0216397
R27238 D_FlipFlop_7.nPRE.n13 D_FlipFlop_7.nPRE 0.0216397
R27239 D_FlipFlop_7.nPRE.n8 D_FlipFlop_7.nPRE.n7 0.0216397
R27240 D_FlipFlop_7.nPRE.n7 D_FlipFlop_7.nPRE 0.0216397
R27241 D_FlipFlop_7.nPRE D_FlipFlop_7.nPRE.n35 0.0204394
R27242 D_FlipFlop_7.nPRE.n20 D_FlipFlop_7.nPRE.n19 0.0107679
R27243 D_FlipFlop_7.nPRE.n19 D_FlipFlop_7.nPRE 0.0107679
R27244 D_FlipFlop_7.nPRE.n1 D_FlipFlop_7.nPRE.n0 0.0107679
R27245 D_FlipFlop_7.nPRE.n0 D_FlipFlop_7.nPRE 0.0107679
R27246 D_FlipFlop_7.nPRE.n3 D_FlipFlop_7.nPRE 0.00441667
R27247 D_FlipFlop_7.nPRE.n31 D_FlipFlop_7.nPRE 0.00441667
R27248 D_FlipFlop_7.nPRE.n36 D_FlipFlop_7.nPRE 0.00441667
R27249 D_FlipFlop_7.nPRE.n31 D_FlipFlop_7.nPRE 0.00406061
R27250 D_FlipFlop_7.nPRE.n3 D_FlipFlop_7.nPRE 0.00406061
R27251 D_FlipFlop_7.nPRE.n36 D_FlipFlop_7.nPRE 0.00406061
R27252 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t2 316.762
R27253 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t0 169.195
R27254 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t4 150.887
R27255 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n2 150.273
R27256 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t3 74.951
R27257 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t5 73.6304
R27258 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t1 60.3943
R27259 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n6 12.0358
R27260 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n8 0.981478
R27261 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.769522
R27262 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n0 0.745065
R27263 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.580578
R27264 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n4 0.533109
R27265 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.428234
R27266 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.063
R27267 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.063
R27268 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n3 0.063
R27269 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n5 0.063
R27270 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.063
R27271 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n7 0.063
R27272 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n1 0.063
R27273 Nand_Gate_3.A.n19 Nand_Gate_3.A.t3 169.46
R27274 Nand_Gate_3.A.n12 Nand_Gate_3.A.t9 168.548
R27275 Nand_Gate_3.A.n18 Nand_Gate_3.A.t1 167.809
R27276 Nand_Gate_3.A.n19 Nand_Gate_3.A.t0 167.809
R27277 Nand_Gate_3.A.n15 Nand_Gate_3.A.t6 158.565
R27278 Nand_Gate_3.A.t6 Nand_Gate_3.A.n14 151.594
R27279 Nand_Gate_3.A.t9 Nand_Gate_3.A.n2 150.293
R27280 Nand_Gate_3.A.n6 Nand_Gate_3.A.t7 150.273
R27281 Nand_Gate_3.A.n3 Nand_Gate_3.A.t4 150.273
R27282 Nand_Gate_3.A Nand_Gate_3.A.t11 99.8701
R27283 Nand_Gate_3.A.n5 Nand_Gate_3.A.t5 74.163
R27284 Nand_Gate_3.A.t11 Nand_Gate_3.A.n10 74.163
R27285 Nand_Gate_3.A.n14 Nand_Gate_3.A.t8 73.6304
R27286 Nand_Gate_3.A.n0 Nand_Gate_3.A.t10 73.6304
R27287 Nand_Gate_3.A.n21 Nand_Gate_3.A.t2 62.1634
R27288 Nand_Gate_3.A.n9 Nand_Gate_3.A.n8 12.6418
R27289 Nand_Gate_3.A.n20 Nand_Gate_3.A.n19 11.4489
R27290 Nand_Gate_3.A.n18 Nand_Gate_3.A.n17 8.21389
R27291 Nand_Gate_3.A.n13 Nand_Gate_3.A 1.2047
R27292 Nand_Gate_3.A.n2 Nand_Gate_3.A.n1 1.19615
R27293 Nand_Gate_3.A.n12 Nand_Gate_3.A.n11 0.922483
R27294 Nand_Gate_3.A.n5 Nand_Gate_3.A 0.851043
R27295 Nand_Gate_3.A.n10 Nand_Gate_3.A 0.851043
R27296 Nand_Gate_3.A.n7 Nand_Gate_3.A.n6 0.61463
R27297 Nand_Gate_3.A.n4 Nand_Gate_3.A.n3 0.61463
R27298 Nand_Gate_3.A.n7 Nand_Gate_3.A 0.486828
R27299 Nand_Gate_3.A.n4 Nand_Gate_3.A 0.486828
R27300 Nand_Gate_3.A.n2 Nand_Gate_3.A 0.447191
R27301 Nand_Gate_3.A.n17 Nand_Gate_3.A.n16 0.425067
R27302 Nand_Gate_3.A.n13 Nand_Gate_3.A.n12 0.399217
R27303 Nand_Gate_3.A.n17 Nand_Gate_3.A 0.39003
R27304 Nand_Gate_3.A.n20 Nand_Gate_3.A.n18 0.280391
R27305 Nand_Gate_3.A.n21 Nand_Gate_3.A.n20 0.200143
R27306 Nand_Gate_3.A.n1 Nand_Gate_3.A 0.1255
R27307 Nand_Gate_3.A.n14 Nand_Gate_3.A 0.063
R27308 Nand_Gate_3.A.n6 Nand_Gate_3.A 0.063
R27309 Nand_Gate_3.A.n8 Nand_Gate_3.A.n5 0.063
R27310 Nand_Gate_3.A.n8 Nand_Gate_3.A.n7 0.063
R27311 Nand_Gate_3.A.n3 Nand_Gate_3.A 0.063
R27312 Nand_Gate_3.A.n10 Nand_Gate_3.A.n9 0.063
R27313 Nand_Gate_3.A.n9 Nand_Gate_3.A.n4 0.063
R27314 Nand_Gate_3.A Nand_Gate_3.A.n21 0.063
R27315 Nand_Gate_3.A.n15 Nand_Gate_3.A.n13 0.024
R27316 Nand_Gate_3.A Nand_Gate_3.A.n15 0.0204394
R27317 Nand_Gate_3.A.n1 Nand_Gate_3.A.n0 0.0107679
R27318 Nand_Gate_3.A.n0 Nand_Gate_3.A 0.0107679
R27319 Nand_Gate_3.A.n11 Nand_Gate_3.A 0.00441667
R27320 Nand_Gate_3.A.n16 Nand_Gate_3.A 0.00441667
R27321 Nand_Gate_3.A.n11 Nand_Gate_3.A 0.00406061
R27322 Nand_Gate_3.A.n16 Nand_Gate_3.A 0.00406061
R27323 D_FlipFlop_1.nPRE.n39 D_FlipFlop_1.nPRE.t2 169.46
R27324 D_FlipFlop_1.nPRE.n39 D_FlipFlop_1.nPRE.t3 167.809
R27325 D_FlipFlop_1.nPRE.n38 D_FlipFlop_1.nPRE.t0 167.809
R27326 D_FlipFlop_1.nPRE.n22 D_FlipFlop_1.nPRE.t16 163.8
R27327 D_FlipFlop_1.nPRE D_FlipFlop_1.nPRE.t12 158.581
R27328 D_FlipFlop_1.nPRE.n35 D_FlipFlop_1.nPRE.t7 158.565
R27329 D_FlipFlop_1.nPRE.t7 D_FlipFlop_1.nPRE.n34 151.594
R27330 D_FlipFlop_1.nPRE.t12 D_FlipFlop_1.nPRE.n5 150.293
R27331 D_FlipFlop_1.nPRE.t16 D_FlipFlop_1.nPRE.n2 150.293
R27332 D_FlipFlop_1.nPRE.n26 D_FlipFlop_1.nPRE.t8 150.273
R27333 D_FlipFlop_1.nPRE.n23 D_FlipFlop_1.nPRE.t6 150.273
R27334 D_FlipFlop_1.nPRE.n16 D_FlipFlop_1.nPRE.t13 150.273
R27335 D_FlipFlop_1.nPRE.n10 D_FlipFlop_1.nPRE.t14 150.273
R27336 D_FlipFlop_1.nPRE D_FlipFlop_1.nPRE.t4 99.8701
R27337 D_FlipFlop_1.nPRE.n25 D_FlipFlop_1.nPRE.t11 74.163
R27338 D_FlipFlop_1.nPRE.t4 D_FlipFlop_1.nPRE.n30 74.163
R27339 D_FlipFlop_1.nPRE.n14 D_FlipFlop_1.nPRE.t5 73.6406
R27340 D_FlipFlop_1.nPRE.n8 D_FlipFlop_1.nPRE.t9 73.6406
R27341 D_FlipFlop_1.nPRE.n34 D_FlipFlop_1.nPRE.t10 73.6304
R27342 D_FlipFlop_1.nPRE.n3 D_FlipFlop_1.nPRE.t15 73.6304
R27343 D_FlipFlop_1.nPRE.n0 D_FlipFlop_1.nPRE.t17 73.6304
R27344 D_FlipFlop_1.nPRE.n41 D_FlipFlop_1.nPRE.t1 62.1634
R27345 D_FlipFlop_1.nPRE.n20 D_FlipFlop_1.nPRE.n13 15.5222
R27346 D_FlipFlop_1.nPRE.n29 D_FlipFlop_1.nPRE.n28 12.6418
R27347 D_FlipFlop_1.nPRE.n40 D_FlipFlop_1.nPRE.n39 11.4489
R27348 D_FlipFlop_1.nPRE.n21 D_FlipFlop_1.nPRE.n20 8.24202
R27349 D_FlipFlop_1.nPRE.n38 D_FlipFlop_1.nPRE.n37 8.21389
R27350 D_FlipFlop_1.nPRE.n22 D_FlipFlop_1.nPRE.n21 7.09922
R27351 D_FlipFlop_1.nPRE.n20 D_FlipFlop_1.nPRE.n19 4.5005
R27352 D_FlipFlop_1.nPRE.n32 D_FlipFlop_1.nPRE.n22 4.03482
R27353 D_FlipFlop_1.nPRE.n33 D_FlipFlop_1.nPRE 1.2047
R27354 D_FlipFlop_1.nPRE.n5 D_FlipFlop_1.nPRE.n4 1.19615
R27355 D_FlipFlop_1.nPRE.n2 D_FlipFlop_1.nPRE.n1 1.19615
R27356 D_FlipFlop_1.nPRE.n32 D_FlipFlop_1.nPRE.n31 0.922483
R27357 D_FlipFlop_1.nPRE.n25 D_FlipFlop_1.nPRE 0.851043
R27358 D_FlipFlop_1.nPRE.n30 D_FlipFlop_1.nPRE 0.851043
R27359 D_FlipFlop_1.nPRE.n15 D_FlipFlop_1.nPRE.n14 0.796696
R27360 D_FlipFlop_1.nPRE.n9 D_FlipFlop_1.nPRE.n8 0.796696
R27361 D_FlipFlop_1.nPRE.n7 D_FlipFlop_1.nPRE.n6 0.783833
R27362 D_FlipFlop_1.nPRE.n7 D_FlipFlop_1.nPRE 0.716182
R27363 D_FlipFlop_1.nPRE.n27 D_FlipFlop_1.nPRE.n26 0.61463
R27364 D_FlipFlop_1.nPRE.n24 D_FlipFlop_1.nPRE.n23 0.61463
R27365 D_FlipFlop_1.nPRE.n15 D_FlipFlop_1.nPRE 0.524957
R27366 D_FlipFlop_1.nPRE.n9 D_FlipFlop_1.nPRE 0.524957
R27367 D_FlipFlop_1.nPRE.n27 D_FlipFlop_1.nPRE 0.486828
R27368 D_FlipFlop_1.nPRE.n24 D_FlipFlop_1.nPRE 0.486828
R27369 D_FlipFlop_1.nPRE.n5 D_FlipFlop_1.nPRE 0.447191
R27370 D_FlipFlop_1.nPRE.n2 D_FlipFlop_1.nPRE 0.447191
R27371 D_FlipFlop_1.nPRE.n37 D_FlipFlop_1.nPRE.n36 0.425067
R27372 D_FlipFlop_1.nPRE.n33 D_FlipFlop_1.nPRE.n32 0.399217
R27373 D_FlipFlop_1.nPRE.n37 D_FlipFlop_1.nPRE 0.39003
R27374 D_FlipFlop_1.nPRE.n40 D_FlipFlop_1.nPRE.n38 0.280391
R27375 D_FlipFlop_1.nPRE.n18 D_FlipFlop_1.nPRE 0.252453
R27376 D_FlipFlop_1.nPRE.n12 D_FlipFlop_1.nPRE 0.252453
R27377 D_FlipFlop_1.nPRE.n18 D_FlipFlop_1.nPRE.n17 0.226043
R27378 D_FlipFlop_1.nPRE.n12 D_FlipFlop_1.nPRE.n11 0.226043
R27379 D_FlipFlop_1.nPRE.n14 D_FlipFlop_1.nPRE 0.217464
R27380 D_FlipFlop_1.nPRE.n8 D_FlipFlop_1.nPRE 0.217464
R27381 D_FlipFlop_1.nPRE.n41 D_FlipFlop_1.nPRE.n40 0.200143
R27382 D_FlipFlop_1.nPRE.n17 D_FlipFlop_1.nPRE 0.1255
R27383 D_FlipFlop_1.nPRE.n11 D_FlipFlop_1.nPRE 0.1255
R27384 D_FlipFlop_1.nPRE.n4 D_FlipFlop_1.nPRE 0.1255
R27385 D_FlipFlop_1.nPRE.n1 D_FlipFlop_1.nPRE 0.1255
R27386 D_FlipFlop_1.nPRE.n34 D_FlipFlop_1.nPRE 0.063
R27387 D_FlipFlop_1.nPRE.n26 D_FlipFlop_1.nPRE 0.063
R27388 D_FlipFlop_1.nPRE.n28 D_FlipFlop_1.nPRE.n25 0.063
R27389 D_FlipFlop_1.nPRE.n28 D_FlipFlop_1.nPRE.n27 0.063
R27390 D_FlipFlop_1.nPRE.n23 D_FlipFlop_1.nPRE 0.063
R27391 D_FlipFlop_1.nPRE.n30 D_FlipFlop_1.nPRE.n29 0.063
R27392 D_FlipFlop_1.nPRE.n29 D_FlipFlop_1.nPRE.n24 0.063
R27393 D_FlipFlop_1.nPRE.n19 D_FlipFlop_1.nPRE.n15 0.063
R27394 D_FlipFlop_1.nPRE.n19 D_FlipFlop_1.nPRE.n18 0.063
R27395 D_FlipFlop_1.nPRE.n13 D_FlipFlop_1.nPRE.n9 0.063
R27396 D_FlipFlop_1.nPRE.n13 D_FlipFlop_1.nPRE.n12 0.063
R27397 D_FlipFlop_1.nPRE D_FlipFlop_1.nPRE.n41 0.063
R27398 D_FlipFlop_1.nPRE.n21 D_FlipFlop_1.nPRE.n7 0.024
R27399 D_FlipFlop_1.nPRE.n35 D_FlipFlop_1.nPRE.n33 0.024
R27400 D_FlipFlop_1.nPRE.n17 D_FlipFlop_1.nPRE.n16 0.0216397
R27401 D_FlipFlop_1.nPRE.n16 D_FlipFlop_1.nPRE 0.0216397
R27402 D_FlipFlop_1.nPRE.n11 D_FlipFlop_1.nPRE.n10 0.0216397
R27403 D_FlipFlop_1.nPRE.n10 D_FlipFlop_1.nPRE 0.0216397
R27404 D_FlipFlop_1.nPRE D_FlipFlop_1.nPRE.n35 0.0204394
R27405 D_FlipFlop_1.nPRE.n4 D_FlipFlop_1.nPRE.n3 0.0107679
R27406 D_FlipFlop_1.nPRE.n3 D_FlipFlop_1.nPRE 0.0107679
R27407 D_FlipFlop_1.nPRE.n1 D_FlipFlop_1.nPRE.n0 0.0107679
R27408 D_FlipFlop_1.nPRE.n0 D_FlipFlop_1.nPRE 0.0107679
R27409 D_FlipFlop_1.nPRE.n6 D_FlipFlop_1.nPRE 0.00441667
R27410 D_FlipFlop_1.nPRE.n31 D_FlipFlop_1.nPRE 0.00441667
R27411 D_FlipFlop_1.nPRE.n36 D_FlipFlop_1.nPRE 0.00441667
R27412 D_FlipFlop_1.nPRE.n31 D_FlipFlop_1.nPRE 0.00406061
R27413 D_FlipFlop_1.nPRE.n6 D_FlipFlop_1.nPRE 0.00406061
R27414 D_FlipFlop_1.nPRE.n36 D_FlipFlop_1.nPRE 0.00406061
R27415 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t2 169.46
R27416 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t3 167.809
R27417 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t1 167.809
R27418 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t7 167.226
R27419 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t6 150.273
R27420 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n0 150.273
R27421 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t4 74.951
R27422 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t5 73.6304
R27423 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t0 60.3943
R27424 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n7 12.3891
R27425 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n2 11.4489
R27426 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 1.68257
R27427 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n9 1.44615
R27428 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n5 1.2342
R27429 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 1.08448
R27430 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.932141
R27431 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n3 0.3496
R27432 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n1 0.280391
R27433 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.063
R27434 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n6 0.063
R27435 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.063
R27436 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n4 0.063
R27437 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n8 0.063
R27438 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n10 0.063
R27439 D_FlipFlop_7.CLK.n12 D_FlipFlop_7.CLK.t0 168.108
R27440 D_FlipFlop_7.CLK.t3 D_FlipFlop_7.CLK.n5 158.207
R27441 D_FlipFlop_7.CLK D_FlipFlop_7.CLK.t4 158.202
R27442 D_FlipFlop_7.CLK.n0 D_FlipFlop_7.CLK.t7 150.293
R27443 D_FlipFlop_7.CLK.t4 D_FlipFlop_7.CLK.n3 150.293
R27444 D_FlipFlop_7.CLK.n6 D_FlipFlop_7.CLK.t3 150.273
R27445 D_FlipFlop_7.CLK.n9 D_FlipFlop_7.CLK.t6 90.1131
R27446 D_FlipFlop_7.CLK.t6 D_FlipFlop_7.CLK.n8 73.6406
R27447 D_FlipFlop_7.CLK.n2 D_FlipFlop_7.CLK.t5 73.6304
R27448 D_FlipFlop_7.CLK.n1 D_FlipFlop_7.CLK.t2 73.6304
R27449 D_FlipFlop_7.CLK D_FlipFlop_7.CLK.t1 60.3072
R27450 D_FlipFlop_7.CLK.n2 D_FlipFlop_7.CLK.n1 16.332
R27451 D_FlipFlop_7.CLK.n12 D_FlipFlop_7.CLK.n11 1.62007
R27452 D_FlipFlop_7.CLK.n8 D_FlipFlop_7.CLK.n7 1.19615
R27453 D_FlipFlop_7.CLK.n1 D_FlipFlop_7.CLK.n0 1.1717
R27454 D_FlipFlop_7.CLK.n3 D_FlipFlop_7.CLK.n2 1.1717
R27455 D_FlipFlop_7.CLK D_FlipFlop_7.CLK.n12 0.484875
R27456 D_FlipFlop_7.CLK.n3 D_FlipFlop_7.CLK 0.447191
R27457 D_FlipFlop_7.CLK.n0 D_FlipFlop_7.CLK 0.436162
R27458 D_FlipFlop_7.CLK.n5 D_FlipFlop_7.CLK.n4 0.349867
R27459 D_FlipFlop_7.CLK.n5 D_FlipFlop_7.CLK 0.321667
R27460 D_FlipFlop_7.CLK.n8 D_FlipFlop_7.CLK 0.217464
R27461 D_FlipFlop_7.CLK.n2 D_FlipFlop_7.CLK 0.149957
R27462 D_FlipFlop_7.CLK.n11 D_FlipFlop_7.CLK 0.149957
R27463 D_FlipFlop_7.CLK.n7 D_FlipFlop_7.CLK 0.1255
R27464 D_FlipFlop_7.CLK.n1 D_FlipFlop_7.CLK 0.117348
R27465 D_FlipFlop_7.CLK.n10 D_FlipFlop_7.CLK 0.0903438
R27466 D_FlipFlop_7.CLK.n1 D_FlipFlop_7.CLK 0.0454219
R27467 D_FlipFlop_7.CLK.n2 D_FlipFlop_7.CLK 0.0454219
R27468 D_FlipFlop_7.CLK.n10 D_FlipFlop_7.CLK.n9 0.027881
R27469 D_FlipFlop_7.CLK.n9 D_FlipFlop_7.CLK 0.027881
R27470 D_FlipFlop_7.CLK.n7 D_FlipFlop_7.CLK.n6 0.0216397
R27471 D_FlipFlop_7.CLK.n6 D_FlipFlop_7.CLK 0.0216397
R27472 D_FlipFlop_7.CLK.n11 D_FlipFlop_7.CLK.n10 0.0180781
R27473 D_FlipFlop_7.CLK.n4 D_FlipFlop_7.CLK 0.00441667
R27474 D_FlipFlop_7.CLK.n4 D_FlipFlop_7.CLK 0.00406061
R27475 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 169.46
R27476 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 168.089
R27477 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 167.809
R27478 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 150.887
R27479 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 73.6304
R27480 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 60.3943
R27481 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 12.0358
R27482 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 11.4489
R27483 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 1.05069
R27484 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 0.981478
R27485 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.769522
R27486 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 0.745065
R27487 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.580578
R27488 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 0.533109
R27489 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.428234
R27490 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.063
R27491 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 0.063
R27492 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 0.063
R27493 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.063
R27494 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 0.063
R27495 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 0.063
R27496 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t1 169.46
R27497 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t2 167.809
R27498 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t0 167.809
R27499 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t5 167.226
R27500 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n6 150.273
R27501 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t6 150.273
R27502 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t7 74.951
R27503 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t4 73.6304
R27504 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t3 60.3943
R27505 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n4 12.3891
R27506 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n8 11.4489
R27507 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n10 1.68257
R27508 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n0 1.44615
R27509 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n2 1.2342
R27510 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 1.08448
R27511 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.932141
R27512 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n9 0.3496
R27513 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n7 0.280391
R27514 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.063
R27515 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.063
R27516 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n3 0.063
R27517 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.063
R27518 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n5 0.063
R27519 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n1 0.063
R27520 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t0 169.46
R27521 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R27522 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t3 167.809
R27523 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t4 167.226
R27524 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n6 150.273
R27525 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t7 150.273
R27526 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t5 74.951
R27527 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t6 73.6304
R27528 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t1 60.3943
R27529 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n4 12.3891
R27530 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n8 11.4489
R27531 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n10 1.68257
R27532 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n0 1.44615
R27533 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n2 1.2342
R27534 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 1.08448
R27535 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.932141
R27536 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n9 0.3496
R27537 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n7 0.280391
R27538 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.063
R27539 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.063
R27540 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n3 0.063
R27541 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.063
R27542 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n5 0.063
R27543 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n1 0.063
R27544 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 169.46
R27545 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 167.809
R27546 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 167.809
R27547 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 167.227
R27548 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 151.594
R27549 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 150.273
R27550 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 74.8641
R27551 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 73.6304
R27552 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 61.84
R27553 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 12.3891
R27554 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 11.4489
R27555 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R27556 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 0.280391
R27557 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 0.200143
R27558 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R27559 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R27560 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 0.149957
R27561 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.063
R27562 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 0.063
R27563 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 0.063
R27564 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 0.063
R27565 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R27566 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 169.46
R27567 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 167.809
R27568 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 167.809
R27569 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 167.227
R27570 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 151.594
R27571 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 150.273
R27572 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 74.8641
R27573 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 73.6304
R27574 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 61.84
R27575 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 12.3891
R27576 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 11.4489
R27577 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.38637
R27578 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 0.280391
R27579 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 0.200143
R27580 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.152844
R27581 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.149957
R27582 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 0.149957
R27583 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.063
R27584 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 0.063
R27585 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 0.063
R27586 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 0.063
R27587 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.0454219
R27588 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t2 169.46
R27589 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t3 167.809
R27590 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.t0 167.809
R27591 D_FlipFlop_0.3-input-nand_2.Vout.t4 D_FlipFlop_0.3-input-nand_2.Vout.n11 167.227
R27592 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.t4 150.293
R27593 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.t6 150.273
R27594 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout.t7 73.6406
R27595 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout.t5 73.6304
R27596 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout.t1 60.3809
R27597 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n5 12.3891
R27598 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout.n9 11.4489
R27599 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout.n2 1.38365
R27600 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.n1 1.19615
R27601 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.n4 1.1717
R27602 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout 0.848156
R27603 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.Vout.n12 0.447191
R27604 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout 0.38637
R27605 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.n10 0.280391
R27606 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout 0.217464
R27607 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout 0.200143
R27608 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout 0.152844
R27609 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.149957
R27610 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R27611 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R27612 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout.n7 0.0874565
R27613 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n3 0.063
R27614 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout.n6 0.063
R27615 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.Vout.n8 0.063
R27616 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.0454219
R27617 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout.n0 0.0107679
R27618 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout 0.0107679
R27619 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 169.46
R27620 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 168.089
R27621 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 167.809
R27622 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 150.887
R27623 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 73.6304
R27624 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 60.3943
R27625 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 12.0358
R27626 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 11.4489
R27627 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 1.05069
R27628 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 0.981478
R27629 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.769522
R27630 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 0.745065
R27631 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.580578
R27632 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 0.533109
R27633 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.428234
R27634 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.063
R27635 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 0.063
R27636 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 0.063
R27637 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.063
R27638 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 0.063
R27639 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 0.063
R27640 Q6.n2 Q6.t2 169.46
R27641 Q6.n4 Q6.t0 167.809
R27642 Q6.n2 Q6.t3 167.809
R27643 Q6.n10 Q6.t4 158.565
R27644 Q6.n14 Q6.t8 150.543
R27645 Q6.n12 Q6.t9 150.543
R27646 Q6.t4 Q6.n9 150.293
R27647 Q6.n14 Q6.t5 74.4613
R27648 Q6.n12 Q6.t7 74.4613
R27649 Q6.n7 Q6.t6 73.6304
R27650 Q6.n0 Q6.t1 60.3809
R27651 Q6 Q6.n16 12.6656
R27652 Q6.n17 Q6.n11 12.3631
R27653 Q6.n3 Q6.n2 11.4489
R27654 Q6.n11 Q6 11.2399
R27655 Q6.n5 Q6.n4 8.21389
R27656 Q6.n11 Q6.n10 4.8158
R27657 Q6.n1 Q6.n0 1.64452
R27658 Q6.n9 Q6.n8 1.19615
R27659 Q6.n13 Q6 0.984196
R27660 Q6.n0 Q6 0.848156
R27661 Q6.n15 Q6.n14 0.747783
R27662 Q6.n13 Q6.n12 0.747783
R27663 Q6.n15 Q6 0.582531
R27664 Q6.n9 Q6 0.447191
R27665 Q6.n6 Q6.n5 0.425067
R27666 Q6.n5 Q6 0.39003
R27667 Q6.n4 Q6.n3 0.280391
R27668 Q6.n3 Q6 0.200143
R27669 Q6.n8 Q6 0.1255
R27670 Q6.n1 Q6 0.1255
R27671 Q6.n14 Q6 0.063
R27672 Q6.n16 Q6.n13 0.063
R27673 Q6.n16 Q6.n15 0.063
R27674 Q6 Q6.n1 0.063
R27675 Q6.n10 Q6 0.0204394
R27676 Q6.n8 Q6.n7 0.0107679
R27677 Q6.n7 Q6 0.0107679
R27678 Q6.n6 Q6 0.00441667
R27679 Q6 Q6.n6 0.00406061
R27680 Q6.n17 Q6 0.00128333
R27681 Q6.n17 Q6 0.00121212
R27682 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 179.256
R27683 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 168.089
R27684 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 150.887
R27685 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 73.6304
R27686 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 60.3943
R27687 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 12.0358
R27688 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 1.05069
R27689 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 0.981478
R27690 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.769522
R27691 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 0.745065
R27692 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.580578
R27693 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 0.533109
R27694 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.428234
R27695 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.063
R27696 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 0.063
R27697 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 0.063
R27698 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.063
R27699 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 0.063
R27700 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 0.063
R27701 Ring_Counter_0.D_FlipFlop_3.Qbar.n4 Ring_Counter_0.D_FlipFlop_3.Qbar.t0 169.46
R27702 Ring_Counter_0.D_FlipFlop_3.Qbar.n4 Ring_Counter_0.D_FlipFlop_3.Qbar.t2 167.809
R27703 Ring_Counter_0.D_FlipFlop_3.Qbar.n3 Ring_Counter_0.D_FlipFlop_3.Qbar.t3 167.809
R27704 Ring_Counter_0.D_FlipFlop_3.Qbar.n1 Ring_Counter_0.D_FlipFlop_3.Qbar.t4 158.28
R27705 Ring_Counter_0.D_FlipFlop_3.Qbar.t4 Ring_Counter_0.D_FlipFlop_3.Qbar.n0 150.273
R27706 Ring_Counter_0.D_FlipFlop_3.Qbar.n0 Ring_Counter_0.D_FlipFlop_3.Qbar.t5 74.951
R27707 Ring_Counter_0.D_FlipFlop_3.Qbar.n6 Ring_Counter_0.D_FlipFlop_3.Qbar.t1 60.3943
R27708 Ring_Counter_0.D_FlipFlop_3.Qbar.n5 Ring_Counter_0.D_FlipFlop_3.Qbar.n4 11.4489
R27709 Ring_Counter_0.D_FlipFlop_3.Qbar.n3 Ring_Counter_0.D_FlipFlop_3.Qbar 8.5174
R27710 Ring_Counter_0.D_FlipFlop_3.Qbar.n6 Ring_Counter_0.D_FlipFlop_3.Qbar.n5 1.96917
R27711 Ring_Counter_0.D_FlipFlop_3.Qbar.n2 Ring_Counter_0.D_FlipFlop_3.Qbar.n1 0.42585
R27712 Ring_Counter_0.D_FlipFlop_3.Qbar.n1 Ring_Counter_0.D_FlipFlop_3.Qbar 0.390742
R27713 Ring_Counter_0.D_FlipFlop_3.Qbar.n5 Ring_Counter_0.D_FlipFlop_3.Qbar.n3 0.280391
R27714 Ring_Counter_0.D_FlipFlop_3.Qbar.n0 Ring_Counter_0.D_FlipFlop_3.Qbar 0.063
R27715 Ring_Counter_0.D_FlipFlop_3.Qbar Ring_Counter_0.D_FlipFlop_3.Qbar.n6 0.063
R27716 Ring_Counter_0.D_FlipFlop_3.Qbar.n2 Ring_Counter_0.D_FlipFlop_3.Qbar 0.00441667
R27717 Ring_Counter_0.D_FlipFlop_3.Qbar Ring_Counter_0.D_FlipFlop_3.Qbar.n2 0.00406061
R27718 Q5.n2 Q5.t0 169.46
R27719 Q5.n4 Q5.t2 167.809
R27720 Q5.n2 Q5.t1 167.809
R27721 Q5.n10 Q5.t7 158.565
R27722 Q5.n14 Q5.t9 150.543
R27723 Q5.n12 Q5.t6 150.543
R27724 Q5.t7 Q5.n9 150.293
R27725 Q5.n14 Q5.t5 74.4613
R27726 Q5.n12 Q5.t4 74.4613
R27727 Q5.n7 Q5.t8 73.6304
R27728 Q5.n0 Q5.t3 60.3809
R27729 Q5 Q5.n16 12.5653
R27730 Q5.n3 Q5.n2 11.4489
R27731 Q5.n17 Q5.n11 8.58897
R27732 Q5.n5 Q5.n4 8.21389
R27733 Q5.n11 Q5 7.80891
R27734 Q5.n11 Q5.n10 4.91607
R27735 Q5.n1 Q5.n0 1.64452
R27736 Q5.n9 Q5.n8 1.19615
R27737 Q5.n13 Q5 0.984196
R27738 Q5.n0 Q5 0.848156
R27739 Q5.n15 Q5.n14 0.747783
R27740 Q5.n13 Q5.n12 0.747783
R27741 Q5.n15 Q5 0.582531
R27742 Q5.n9 Q5 0.447191
R27743 Q5.n6 Q5.n5 0.425067
R27744 Q5.n5 Q5 0.39003
R27745 Q5.n4 Q5.n3 0.280391
R27746 Q5.n3 Q5 0.200143
R27747 Q5.n8 Q5 0.1255
R27748 Q5.n1 Q5 0.1255
R27749 Q5.n14 Q5 0.063
R27750 Q5.n16 Q5.n13 0.063
R27751 Q5.n16 Q5.n15 0.063
R27752 Q5 Q5.n1 0.063
R27753 Q5.n10 Q5 0.0204394
R27754 Q5.n8 Q5.n7 0.0107679
R27755 Q5.n7 Q5 0.0107679
R27756 Q5.n6 Q5 0.00441667
R27757 Q5 Q5.n6 0.00406061
R27758 Q5.n17 Q5 0.00128333
R27759 Q5.n17 Q5 0.00121212
R27760 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 169.46
R27761 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 167.809
R27762 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 167.809
R27763 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 167.227
R27764 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 151.594
R27765 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 150.273
R27766 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 74.8641
R27767 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6304
R27768 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 61.84
R27769 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 12.3891
R27770 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 11.4489
R27771 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 0.38637
R27772 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 0.280391
R27773 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 0.200143
R27774 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R27775 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R27776 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 0.149957
R27777 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.063
R27778 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.063
R27779 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 0.063
R27780 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 0.063
R27781 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R27782 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t0 169.46
R27783 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t3 167.809
R27784 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t1 167.809
R27785 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t4 167.226
R27786 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n6 150.273
R27787 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t7 150.273
R27788 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t5 74.951
R27789 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t6 73.6304
R27790 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t2 60.3943
R27791 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n4 12.3891
R27792 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n8 11.4489
R27793 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n10 1.68257
R27794 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n0 1.44615
R27795 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n2 1.2342
R27796 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 1.08448
R27797 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.932141
R27798 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n9 0.3496
R27799 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n7 0.280391
R27800 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.063
R27801 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.063
R27802 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n3 0.063
R27803 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.063
R27804 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n5 0.063
R27805 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n1 0.063
R27806 D_FlipFlop_3.CLK.n12 D_FlipFlop_3.CLK.t0 168.108
R27807 D_FlipFlop_3.CLK.t3 D_FlipFlop_3.CLK.n5 158.207
R27808 D_FlipFlop_3.CLK D_FlipFlop_3.CLK.t4 158.202
R27809 D_FlipFlop_3.CLK.n0 D_FlipFlop_3.CLK.t2 150.293
R27810 D_FlipFlop_3.CLK.t4 D_FlipFlop_3.CLK.n3 150.293
R27811 D_FlipFlop_3.CLK.n6 D_FlipFlop_3.CLK.t3 150.273
R27812 D_FlipFlop_3.CLK.n9 D_FlipFlop_3.CLK.t7 90.1131
R27813 D_FlipFlop_3.CLK.t7 D_FlipFlop_3.CLK.n8 73.6406
R27814 D_FlipFlop_3.CLK.n2 D_FlipFlop_3.CLK.t5 73.6304
R27815 D_FlipFlop_3.CLK.n1 D_FlipFlop_3.CLK.t6 73.6304
R27816 D_FlipFlop_3.CLK D_FlipFlop_3.CLK.t1 60.3072
R27817 D_FlipFlop_3.CLK.n2 D_FlipFlop_3.CLK.n1 16.332
R27818 D_FlipFlop_3.CLK.n12 D_FlipFlop_3.CLK.n11 1.62007
R27819 D_FlipFlop_3.CLK.n8 D_FlipFlop_3.CLK.n7 1.19615
R27820 D_FlipFlop_3.CLK.n1 D_FlipFlop_3.CLK.n0 1.1717
R27821 D_FlipFlop_3.CLK.n3 D_FlipFlop_3.CLK.n2 1.1717
R27822 D_FlipFlop_3.CLK D_FlipFlop_3.CLK.n12 0.484875
R27823 D_FlipFlop_3.CLK.n3 D_FlipFlop_3.CLK 0.447191
R27824 D_FlipFlop_3.CLK.n0 D_FlipFlop_3.CLK 0.436162
R27825 D_FlipFlop_3.CLK.n5 D_FlipFlop_3.CLK.n4 0.349867
R27826 D_FlipFlop_3.CLK.n5 D_FlipFlop_3.CLK 0.321667
R27827 D_FlipFlop_3.CLK.n8 D_FlipFlop_3.CLK 0.217464
R27828 D_FlipFlop_3.CLK.n2 D_FlipFlop_3.CLK 0.149957
R27829 D_FlipFlop_3.CLK.n11 D_FlipFlop_3.CLK 0.149957
R27830 D_FlipFlop_3.CLK.n7 D_FlipFlop_3.CLK 0.1255
R27831 D_FlipFlop_3.CLK.n1 D_FlipFlop_3.CLK 0.117348
R27832 D_FlipFlop_3.CLK.n10 D_FlipFlop_3.CLK 0.0903438
R27833 D_FlipFlop_3.CLK.n1 D_FlipFlop_3.CLK 0.0454219
R27834 D_FlipFlop_3.CLK.n2 D_FlipFlop_3.CLK 0.0454219
R27835 D_FlipFlop_3.CLK.n10 D_FlipFlop_3.CLK.n9 0.027881
R27836 D_FlipFlop_3.CLK.n9 D_FlipFlop_3.CLK 0.027881
R27837 D_FlipFlop_3.CLK.n7 D_FlipFlop_3.CLK.n6 0.0216397
R27838 D_FlipFlop_3.CLK.n6 D_FlipFlop_3.CLK 0.0216397
R27839 D_FlipFlop_3.CLK.n11 D_FlipFlop_3.CLK.n10 0.0180781
R27840 D_FlipFlop_3.CLK.n4 D_FlipFlop_3.CLK 0.00441667
R27841 D_FlipFlop_3.CLK.n4 D_FlipFlop_3.CLK 0.00406061
R27842 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t0 169.46
R27843 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t2 167.809
R27844 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t1 167.809
R27845 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t4 167.226
R27846 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n6 150.273
R27847 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t5 150.273
R27848 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t7 74.951
R27849 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t6 73.6304
R27850 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t3 60.3943
R27851 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n4 12.3891
R27852 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n8 11.4489
R27853 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n10 1.68257
R27854 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n0 1.44615
R27855 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n2 1.2342
R27856 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 1.08448
R27857 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.932141
R27858 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n9 0.3496
R27859 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n7 0.280391
R27860 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.063
R27861 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.063
R27862 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n3 0.063
R27863 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.063
R27864 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n5 0.063
R27865 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n1 0.063
R27866 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 169.46
R27867 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 167.809
R27868 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 167.809
R27869 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 167.227
R27870 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 151.594
R27871 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 150.273
R27872 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 74.8641
R27873 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 73.6304
R27874 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 61.84
R27875 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 12.3891
R27876 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 11.4489
R27877 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R27878 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 0.280391
R27879 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 0.200143
R27880 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R27881 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R27882 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 0.149957
R27883 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.063
R27884 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 0.063
R27885 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 0.063
R27886 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 0.063
R27887 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R27888 Q7.n2 Q7.t2 169.46
R27889 Q7.n4 Q7.t0 167.809
R27890 Q7.n2 Q7.t3 167.809
R27891 Q7.n10 Q7.t4 158.565
R27892 Q7.n14 Q7.t5 150.543
R27893 Q7.n12 Q7.t9 150.543
R27894 Q7.t4 Q7.n9 150.293
R27895 Q7.n14 Q7.t6 74.4613
R27896 Q7.n12 Q7.t7 74.4613
R27897 Q7.n7 Q7.t8 73.6304
R27898 Q7.n0 Q7.t1 60.3809
R27899 Q7.n17 Q7.n11 16.1372
R27900 Q7.n11 Q7 14.6709
R27901 Q7 Q7.n16 12.7658
R27902 Q7.n3 Q7.n2 11.4489
R27903 Q7.n5 Q7.n4 8.21389
R27904 Q7.n11 Q7.n10 4.71553
R27905 Q7.n1 Q7.n0 1.64452
R27906 Q7.n9 Q7.n8 1.19615
R27907 Q7.n13 Q7 0.984196
R27908 Q7.n0 Q7 0.848156
R27909 Q7.n15 Q7.n14 0.747783
R27910 Q7.n13 Q7.n12 0.747783
R27911 Q7.n15 Q7 0.582531
R27912 Q7.n9 Q7 0.447191
R27913 Q7.n6 Q7.n5 0.425067
R27914 Q7.n5 Q7 0.39003
R27915 Q7.n4 Q7.n3 0.280391
R27916 Q7.n3 Q7 0.200143
R27917 Q7.n8 Q7 0.1255
R27918 Q7.n1 Q7 0.1255
R27919 Q7.n14 Q7 0.063
R27920 Q7.n16 Q7.n13 0.063
R27921 Q7.n16 Q7.n15 0.063
R27922 Q7 Q7.n1 0.063
R27923 Q7.n10 Q7 0.0204394
R27924 Q7.n8 Q7.n7 0.0107679
R27925 Q7.n7 Q7 0.0107679
R27926 Q7.n6 Q7 0.00441667
R27927 Q7 Q7.n6 0.00406061
R27928 Q7.n17 Q7 0.00128333
R27929 Q7.n17 Q7 0.00121212
R27930 D_FlipFlop_6.nPRE.n39 D_FlipFlop_6.nPRE.t3 169.46
R27931 D_FlipFlop_6.nPRE.n38 D_FlipFlop_6.nPRE.t1 167.809
R27932 D_FlipFlop_6.nPRE.n39 D_FlipFlop_6.nPRE.t0 167.809
R27933 D_FlipFlop_6.nPRE.n22 D_FlipFlop_6.nPRE.t9 161.98
R27934 D_FlipFlop_6.nPRE D_FlipFlop_6.nPRE.t14 158.581
R27935 D_FlipFlop_6.nPRE.n35 D_FlipFlop_6.nPRE.t8 158.565
R27936 D_FlipFlop_6.nPRE.t8 D_FlipFlop_6.nPRE.n34 151.594
R27937 D_FlipFlop_6.nPRE.t9 D_FlipFlop_6.nPRE.n21 150.293
R27938 D_FlipFlop_6.nPRE.t14 D_FlipFlop_6.nPRE.n2 150.293
R27939 D_FlipFlop_6.nPRE.n26 D_FlipFlop_6.nPRE.t4 150.273
R27940 D_FlipFlop_6.nPRE.n23 D_FlipFlop_6.nPRE.t15 150.273
R27941 D_FlipFlop_6.nPRE.n13 D_FlipFlop_6.nPRE.t11 150.273
R27942 D_FlipFlop_6.nPRE.n7 D_FlipFlop_6.nPRE.t5 150.273
R27943 D_FlipFlop_6.nPRE D_FlipFlop_6.nPRE.t13 99.8701
R27944 D_FlipFlop_6.nPRE.n25 D_FlipFlop_6.nPRE.t7 74.163
R27945 D_FlipFlop_6.nPRE.t13 D_FlipFlop_6.nPRE.n30 74.163
R27946 D_FlipFlop_6.nPRE.n11 D_FlipFlop_6.nPRE.t6 73.6406
R27947 D_FlipFlop_6.nPRE.n5 D_FlipFlop_6.nPRE.t17 73.6406
R27948 D_FlipFlop_6.nPRE.n34 D_FlipFlop_6.nPRE.t12 73.6304
R27949 D_FlipFlop_6.nPRE.n19 D_FlipFlop_6.nPRE.t10 73.6304
R27950 D_FlipFlop_6.nPRE.n0 D_FlipFlop_6.nPRE.t16 73.6304
R27951 D_FlipFlop_6.nPRE.n41 D_FlipFlop_6.nPRE.t2 62.1634
R27952 D_FlipFlop_6.nPRE.n17 D_FlipFlop_6.nPRE.n10 15.5222
R27953 D_FlipFlop_6.nPRE.n29 D_FlipFlop_6.nPRE.n28 12.6418
R27954 D_FlipFlop_6.nPRE.n40 D_FlipFlop_6.nPRE.n39 11.4489
R27955 D_FlipFlop_6.nPRE.n22 D_FlipFlop_6.nPRE.n18 9.12492
R27956 D_FlipFlop_6.nPRE.n32 D_FlipFlop_6.nPRE.n22 8.40425
R27957 D_FlipFlop_6.nPRE.n18 D_FlipFlop_6.nPRE.n17 8.24202
R27958 D_FlipFlop_6.nPRE.n38 D_FlipFlop_6.nPRE.n37 8.21389
R27959 D_FlipFlop_6.nPRE.n17 D_FlipFlop_6.nPRE.n16 4.5005
R27960 D_FlipFlop_6.nPRE.n33 D_FlipFlop_6.nPRE 1.2047
R27961 D_FlipFlop_6.nPRE.n21 D_FlipFlop_6.nPRE.n20 1.19615
R27962 D_FlipFlop_6.nPRE.n2 D_FlipFlop_6.nPRE.n1 1.19615
R27963 D_FlipFlop_6.nPRE.n32 D_FlipFlop_6.nPRE.n31 0.922483
R27964 D_FlipFlop_6.nPRE.n25 D_FlipFlop_6.nPRE 0.851043
R27965 D_FlipFlop_6.nPRE.n30 D_FlipFlop_6.nPRE 0.851043
R27966 D_FlipFlop_6.nPRE.n12 D_FlipFlop_6.nPRE.n11 0.796696
R27967 D_FlipFlop_6.nPRE.n6 D_FlipFlop_6.nPRE.n5 0.796696
R27968 D_FlipFlop_6.nPRE.n4 D_FlipFlop_6.nPRE.n3 0.783833
R27969 D_FlipFlop_6.nPRE.n4 D_FlipFlop_6.nPRE 0.716182
R27970 D_FlipFlop_6.nPRE.n27 D_FlipFlop_6.nPRE.n26 0.61463
R27971 D_FlipFlop_6.nPRE.n24 D_FlipFlop_6.nPRE.n23 0.61463
R27972 D_FlipFlop_6.nPRE.n12 D_FlipFlop_6.nPRE 0.524957
R27973 D_FlipFlop_6.nPRE.n6 D_FlipFlop_6.nPRE 0.524957
R27974 D_FlipFlop_6.nPRE.n27 D_FlipFlop_6.nPRE 0.486828
R27975 D_FlipFlop_6.nPRE.n24 D_FlipFlop_6.nPRE 0.486828
R27976 D_FlipFlop_6.nPRE.n21 D_FlipFlop_6.nPRE 0.447191
R27977 D_FlipFlop_6.nPRE.n2 D_FlipFlop_6.nPRE 0.447191
R27978 D_FlipFlop_6.nPRE.n37 D_FlipFlop_6.nPRE.n36 0.425067
R27979 D_FlipFlop_6.nPRE.n33 D_FlipFlop_6.nPRE.n32 0.399217
R27980 D_FlipFlop_6.nPRE.n37 D_FlipFlop_6.nPRE 0.39003
R27981 D_FlipFlop_6.nPRE.n40 D_FlipFlop_6.nPRE.n38 0.280391
R27982 D_FlipFlop_6.nPRE.n15 D_FlipFlop_6.nPRE 0.252453
R27983 D_FlipFlop_6.nPRE.n9 D_FlipFlop_6.nPRE 0.252453
R27984 D_FlipFlop_6.nPRE.n15 D_FlipFlop_6.nPRE.n14 0.226043
R27985 D_FlipFlop_6.nPRE.n9 D_FlipFlop_6.nPRE.n8 0.226043
R27986 D_FlipFlop_6.nPRE.n11 D_FlipFlop_6.nPRE 0.217464
R27987 D_FlipFlop_6.nPRE.n5 D_FlipFlop_6.nPRE 0.217464
R27988 D_FlipFlop_6.nPRE.n41 D_FlipFlop_6.nPRE.n40 0.200143
R27989 D_FlipFlop_6.nPRE.n20 D_FlipFlop_6.nPRE 0.1255
R27990 D_FlipFlop_6.nPRE.n14 D_FlipFlop_6.nPRE 0.1255
R27991 D_FlipFlop_6.nPRE.n8 D_FlipFlop_6.nPRE 0.1255
R27992 D_FlipFlop_6.nPRE.n1 D_FlipFlop_6.nPRE 0.1255
R27993 D_FlipFlop_6.nPRE.n34 D_FlipFlop_6.nPRE 0.063
R27994 D_FlipFlop_6.nPRE.n26 D_FlipFlop_6.nPRE 0.063
R27995 D_FlipFlop_6.nPRE.n28 D_FlipFlop_6.nPRE.n25 0.063
R27996 D_FlipFlop_6.nPRE.n28 D_FlipFlop_6.nPRE.n27 0.063
R27997 D_FlipFlop_6.nPRE.n23 D_FlipFlop_6.nPRE 0.063
R27998 D_FlipFlop_6.nPRE.n30 D_FlipFlop_6.nPRE.n29 0.063
R27999 D_FlipFlop_6.nPRE.n29 D_FlipFlop_6.nPRE.n24 0.063
R28000 D_FlipFlop_6.nPRE.n16 D_FlipFlop_6.nPRE.n12 0.063
R28001 D_FlipFlop_6.nPRE.n16 D_FlipFlop_6.nPRE.n15 0.063
R28002 D_FlipFlop_6.nPRE.n10 D_FlipFlop_6.nPRE.n6 0.063
R28003 D_FlipFlop_6.nPRE.n10 D_FlipFlop_6.nPRE.n9 0.063
R28004 D_FlipFlop_6.nPRE D_FlipFlop_6.nPRE.n41 0.063
R28005 D_FlipFlop_6.nPRE.n18 D_FlipFlop_6.nPRE.n4 0.024
R28006 D_FlipFlop_6.nPRE.n35 D_FlipFlop_6.nPRE.n33 0.024
R28007 D_FlipFlop_6.nPRE.n14 D_FlipFlop_6.nPRE.n13 0.0216397
R28008 D_FlipFlop_6.nPRE.n13 D_FlipFlop_6.nPRE 0.0216397
R28009 D_FlipFlop_6.nPRE.n8 D_FlipFlop_6.nPRE.n7 0.0216397
R28010 D_FlipFlop_6.nPRE.n7 D_FlipFlop_6.nPRE 0.0216397
R28011 D_FlipFlop_6.nPRE D_FlipFlop_6.nPRE.n35 0.0204394
R28012 D_FlipFlop_6.nPRE.n20 D_FlipFlop_6.nPRE.n19 0.0107679
R28013 D_FlipFlop_6.nPRE.n19 D_FlipFlop_6.nPRE 0.0107679
R28014 D_FlipFlop_6.nPRE.n1 D_FlipFlop_6.nPRE.n0 0.0107679
R28015 D_FlipFlop_6.nPRE.n0 D_FlipFlop_6.nPRE 0.0107679
R28016 D_FlipFlop_6.nPRE.n3 D_FlipFlop_6.nPRE 0.00441667
R28017 D_FlipFlop_6.nPRE.n31 D_FlipFlop_6.nPRE 0.00441667
R28018 D_FlipFlop_6.nPRE.n36 D_FlipFlop_6.nPRE 0.00441667
R28019 D_FlipFlop_6.nPRE.n31 D_FlipFlop_6.nPRE 0.00406061
R28020 D_FlipFlop_6.nPRE.n3 D_FlipFlop_6.nPRE 0.00406061
R28021 D_FlipFlop_6.nPRE.n36 D_FlipFlop_6.nPRE 0.00406061
R28022 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.t1 169.46
R28023 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C.t2 167.809
R28024 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.t0 167.809
R28025 D_FlipFlop_0.3-input-nand_2.C.t4 D_FlipFlop_0.3-input-nand_2.C.n13 167.226
R28026 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C.t5 150.273
R28027 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.t4 150.273
R28028 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C.t7 73.6406
R28029 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C.t6 73.6304
R28030 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_2.C.t3 60.3943
R28031 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C.n7 12.3891
R28032 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n11 11.4489
R28033 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C 1.68257
R28034 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C.n2 1.38365
R28035 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C.n0 1.19615
R28036 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C.n5 1.1717
R28037 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C 1.08448
R28038 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C 0.932141
R28039 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C 0.720633
R28040 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C.n12 0.280391
R28041 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C 0.217464
R28042 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C 0.1255
R28043 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C 0.1255
R28044 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C 0.1255
R28045 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C.n9 0.0874565
R28046 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C.n6 0.063
R28047 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C 0.063
R28048 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C.n8 0.063
R28049 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C.n3 0.063
R28050 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n10 0.0435206
R28051 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.n1 0.0216397
R28052 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_2.C.n14 0.0216397
R28053 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C.n4 0.0107679
R28054 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C 0.0107679
R28055 Nand_Gate_0.A.n19 Nand_Gate_0.A.t2 169.46
R28056 Nand_Gate_0.A.n19 Nand_Gate_0.A.t3 167.809
R28057 Nand_Gate_0.A.n18 Nand_Gate_0.A.t0 167.809
R28058 Nand_Gate_0.A.n12 Nand_Gate_0.A.t7 167.111
R28059 Nand_Gate_0.A.n15 Nand_Gate_0.A.t5 158.565
R28060 Nand_Gate_0.A.t5 Nand_Gate_0.A.n14 151.594
R28061 Nand_Gate_0.A.t7 Nand_Gate_0.A.n2 150.293
R28062 Nand_Gate_0.A.n6 Nand_Gate_0.A.t9 150.273
R28063 Nand_Gate_0.A.n3 Nand_Gate_0.A.t6 150.273
R28064 Nand_Gate_0.A Nand_Gate_0.A.t4 99.8701
R28065 Nand_Gate_0.A.n5 Nand_Gate_0.A.t11 74.163
R28066 Nand_Gate_0.A.t4 Nand_Gate_0.A.n10 74.163
R28067 Nand_Gate_0.A.n14 Nand_Gate_0.A.t10 73.6304
R28068 Nand_Gate_0.A.n0 Nand_Gate_0.A.t8 73.6304
R28069 Nand_Gate_0.A.n21 Nand_Gate_0.A.t1 62.1634
R28070 Nand_Gate_0.A.n9 Nand_Gate_0.A.n8 12.6418
R28071 Nand_Gate_0.A.n20 Nand_Gate_0.A.n19 11.4489
R28072 Nand_Gate_0.A.n18 Nand_Gate_0.A.n17 8.21389
R28073 Nand_Gate_0.A.n13 Nand_Gate_0.A 1.2047
R28074 Nand_Gate_0.A.n2 Nand_Gate_0.A.n1 1.19615
R28075 Nand_Gate_0.A.n12 Nand_Gate_0.A.n11 0.922483
R28076 Nand_Gate_0.A.n5 Nand_Gate_0.A 0.851043
R28077 Nand_Gate_0.A.n10 Nand_Gate_0.A 0.851043
R28078 Nand_Gate_0.A.n7 Nand_Gate_0.A.n6 0.61463
R28079 Nand_Gate_0.A.n4 Nand_Gate_0.A.n3 0.61463
R28080 Nand_Gate_0.A.n7 Nand_Gate_0.A 0.486828
R28081 Nand_Gate_0.A.n4 Nand_Gate_0.A 0.486828
R28082 Nand_Gate_0.A.n2 Nand_Gate_0.A 0.447191
R28083 Nand_Gate_0.A.n17 Nand_Gate_0.A.n16 0.425067
R28084 Nand_Gate_0.A.n13 Nand_Gate_0.A.n12 0.399217
R28085 Nand_Gate_0.A.n17 Nand_Gate_0.A 0.39003
R28086 Nand_Gate_0.A.n20 Nand_Gate_0.A.n18 0.280391
R28087 Nand_Gate_0.A.n21 Nand_Gate_0.A.n20 0.200143
R28088 Nand_Gate_0.A.n1 Nand_Gate_0.A 0.1255
R28089 Nand_Gate_0.A.n14 Nand_Gate_0.A 0.063
R28090 Nand_Gate_0.A.n6 Nand_Gate_0.A 0.063
R28091 Nand_Gate_0.A.n8 Nand_Gate_0.A.n5 0.063
R28092 Nand_Gate_0.A.n8 Nand_Gate_0.A.n7 0.063
R28093 Nand_Gate_0.A.n3 Nand_Gate_0.A 0.063
R28094 Nand_Gate_0.A.n10 Nand_Gate_0.A.n9 0.063
R28095 Nand_Gate_0.A.n9 Nand_Gate_0.A.n4 0.063
R28096 Nand_Gate_0.A Nand_Gate_0.A.n21 0.063
R28097 Nand_Gate_0.A.n15 Nand_Gate_0.A.n13 0.024
R28098 Nand_Gate_0.A Nand_Gate_0.A.n15 0.0204394
R28099 Nand_Gate_0.A.n1 Nand_Gate_0.A.n0 0.0107679
R28100 Nand_Gate_0.A.n0 Nand_Gate_0.A 0.0107679
R28101 Nand_Gate_0.A.n11 Nand_Gate_0.A 0.00441667
R28102 Nand_Gate_0.A.n16 Nand_Gate_0.A 0.00441667
R28103 Nand_Gate_0.A.n11 Nand_Gate_0.A 0.00406061
R28104 Nand_Gate_0.A.n16 Nand_Gate_0.A 0.00406061
R28105 Vin Vin.t0 467.404
R28106 a_50502_29172.n0 a_50502_29172.t2 1546.57
R28107 a_50502_29172.n1 a_50502_29172.t1 27.7124
R28108 a_50502_29172.t0 a_50502_29172.n1 21.1744
R28109 a_50502_29172.n0 a_50502_29172.t3 11.1233
R28110 a_50502_29172.n1 a_50502_29172.n0 5.89691
R28111 a_51773_21431.n0 a_51773_21431.t1 25.9955
R28112 a_51773_21431.n0 a_51773_21431.t2 14.4333
R28113 a_51773_21431.t0 a_51773_21431.n0 14.4333
R28114 Vbias.n17 Vbias.n16 93853.1
R28115 Vbias.n43 Vbias.n16 93853.1
R28116 Vbias.n43 Vbias.n14 93853.1
R28117 Vbias.n19 Vbias.n16 41816.1
R28118 Vbias.n58 Vbias.n8 7992.36
R28119 Vbias.n58 Vbias.n9 7992.36
R28120 Vbias.n23 Vbias.n9 7992.36
R28121 Vbias.n23 Vbias.n8 7992.36
R28122 Vbias.n35 Vbias.n20 7992.36
R28123 Vbias.n35 Vbias.n21 7992.36
R28124 Vbias.n40 Vbias.n21 7992.36
R28125 Vbias.n40 Vbias.n20 7992.36
R28126 Vbias.n65 Vbias.n5 6345.81
R28127 Vbias.n65 Vbias.n6 6345.81
R28128 Vbias.n61 Vbias.n6 6345.81
R28129 Vbias.n61 Vbias.n5 6345.81
R28130 Vbias.n33 Vbias.n28 6345.81
R28131 Vbias.n28 Vbias.n25 6345.81
R28132 Vbias.n26 Vbias.n25 6345.81
R28133 Vbias.n33 Vbias.n26 6345.81
R28134 Vbias.n44 Vbias.n15 6098.07
R28135 Vbias.n15 Vbias.n13 6098.07
R28136 Vbias.n45 Vbias.n44 5912.48
R28137 Vbias.n45 Vbias.n13 5912.48
R28138 Vbias.n70 Vbias.n4 4699.26
R28139 Vbias.n67 Vbias.n2 4699.26
R28140 Vbias.n67 Vbias.n4 4699.26
R28141 Vbias.n37 Vbias.n36 918.212
R28142 Vbias.n57 Vbias.n10 918.212
R28143 Vbias.n11 Vbias.n10 918.212
R28144 Vbias.n39 Vbias.n37 918.212
R28145 Vbias.n57 Vbias.n56 861.144
R28146 Vbias.n39 Vbias.n38 861.144
R28147 Vbias.n36 Vbias.n12 819.201
R28148 Vbias.n55 Vbias.n11 819.201
R28149 Vbias.n64 Vbias.n7 729.976
R28150 Vbias.n64 Vbias.n63 729.976
R28151 Vbias.n63 Vbias.n62 729.976
R28152 Vbias.n62 Vbias.n7 729.976
R28153 Vbias.n32 Vbias.n31 729.976
R28154 Vbias.n31 Vbias.n30 729.976
R28155 Vbias.n30 Vbias.n29 729.976
R28156 Vbias.n32 Vbias.n29 729.976
R28157 Vbias.n71 Vbias.n3 541.741
R28158 Vbias.n3 Vbias.n1 541.741
R28159 Vbias.n72 Vbias.n71 484.675
R28160 Vbias.n72 Vbias.n1 484.675
R28161 Vbias.n42 Vbias.n41 296.86
R28162 Vbias.n18 Vbias.n17 190.803
R28163 Vbias.n42 Vbias.n19 186.645
R28164 Vbias.n68 Vbias.n66 164.214
R28165 Vbias.n37 Vbias.n20 117.001
R28166 Vbias.n20 Vbias.t2 117.001
R28167 Vbias.n38 Vbias.n21 117.001
R28168 Vbias.n21 Vbias.t2 117.001
R28169 Vbias.n4 Vbias.n3 117.001
R28170 Vbias.t7 Vbias.n4 117.001
R28171 Vbias.n72 Vbias.n2 117.001
R28172 Vbias.n10 Vbias.n8 117.001
R28173 Vbias.n8 Vbias.t5 117.001
R28174 Vbias.n56 Vbias.n9 117.001
R28175 Vbias.n9 Vbias.t5 117.001
R28176 Vbias.n33 Vbias.n32 117.001
R28177 Vbias.t9 Vbias.n33 117.001
R28178 Vbias.n30 Vbias.n25 117.001
R28179 Vbias.t9 Vbias.n25 117.001
R28180 Vbias.n7 Vbias.n5 117.001
R28181 Vbias.n5 Vbias.t0 117.001
R28182 Vbias.n63 Vbias.n6 117.001
R28183 Vbias.n6 Vbias.t0 117.001
R28184 Vbias.n69 Vbias.n2 112.052
R28185 Vbias.n70 Vbias.n69 86.728
R28186 Vbias.n41 Vbias.t2 72.8308
R28187 Vbias.n66 Vbias.t0 72.8308
R28188 Vbias.t7 Vbias.n68 72.8308
R28189 Vbias.n34 Vbias.n22 71.4462
R28190 Vbias.n60 Vbias.n59 71.4462
R28191 Vbias.n27 Vbias.n24 41.5387
R28192 Vbias.n16 Vbias.n15 32.5005
R28193 Vbias.n45 Vbias.n14 32.5005
R28194 Vbias.n18 Vbias.n14 32.4237
R28195 Vbias.t9 Vbias.n24 31.2926
R28196 Vbias.n27 Vbias.t5 31.2926
R28197 Vbias.n67 Vbias.n1 17.7278
R28198 Vbias.n68 Vbias.n67 17.7278
R28199 Vbias.n71 Vbias.n70 17.7278
R28200 Vbias.n38 Vbias.n12 17.443
R28201 Vbias.n56 Vbias.n55 17.443
R28202 Vbias.n48 Vbias.t8 16.8637
R28203 Vbias.n50 Vbias.t3 14.4765
R28204 Vbias.n49 Vbias.t6 14.02
R28205 Vbias.n29 Vbias.n26 12.4473
R28206 Vbias.n26 Vbias.n22 12.4473
R28207 Vbias.n31 Vbias.n28 12.4473
R28208 Vbias.n28 Vbias.n27 12.4473
R28209 Vbias.n62 Vbias.n61 12.4473
R28210 Vbias.n61 Vbias.n60 12.4473
R28211 Vbias.n65 Vbias.n64 12.4473
R28212 Vbias.n66 Vbias.n65 12.4473
R28213 Vbias.n53 Vbias.n50 11.6088
R28214 Vbias.n47 Vbias.t1 9.73694
R28215 Vbias.n40 Vbias.n39 9.43598
R28216 Vbias.n41 Vbias.n40 9.43598
R28217 Vbias.n36 Vbias.n35 9.43598
R28218 Vbias.n35 Vbias.n34 9.43598
R28219 Vbias.n23 Vbias.n11 9.43598
R28220 Vbias.n24 Vbias.n23 9.43598
R28221 Vbias.n58 Vbias.n57 9.43598
R28222 Vbias.n59 Vbias.n58 9.43598
R28223 Vbias.n47 Vbias.n0 8.19877
R28224 Vbias.n46 Vbias.n45 6.82745
R28225 Vbias.n52 Vbias 3.91652
R28226 Vbias.n54 Vbias.n12 3.91345
R28227 Vbias.n55 Vbias.n54 3.91345
R28228 Vbias.n48 Vbias.n47 3.4105
R28229 Vbias.n19 Vbias.t4 3.30535
R28230 Vbias.n51 Vbias 2.76137
R28231 Vbias.n52 Vbias.n51 2.688
R28232 Vbias.n69 Vbias.t7 2.16029
R28233 Vbias.n73 Vbias.n72 1.8605
R28234 Vbias Vbias.n74 1.85988
R28235 Vbias.n74 Vbias.n73 1.69615
R28236 Vbias.n49 Vbias.n48 1.57387
R28237 Vbias.n22 Vbias.t2 1.38511
R28238 Vbias.n34 Vbias.t9 1.38511
R28239 Vbias.n60 Vbias.t5 1.38511
R28240 Vbias.n59 Vbias.t0 1.38511
R28241 Vbias.n44 Vbias.n43 1.28905
R28242 Vbias.n43 Vbias.n42 1.28905
R28243 Vbias.n17 Vbias.n13 1.28905
R28244 Vbias.n50 Vbias.n49 1.16354
R28245 Vbias.n73 Vbias 0.891804
R28246 Vbias.n54 Vbias.n53 0.664786
R28247 Vbias.t4 Vbias.n18 0.0670719
R28248 Vbias.n53 Vbias.n52 0.063
R28249 Vbias.n51 Vbias.n0 0.063
R28250 Vbias.n74 Vbias.n0 0.063
R28251 Vbias.n53 Vbias 0.0512812
R28252 Vbias.n46 Vbias 0.0168043
R28253 Vbias Vbias.n46 0.0122188
R28254 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t3 316.762
R28255 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t0 169.195
R28256 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t4 150.887
R28257 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n2 150.273
R28258 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t2 74.951
R28259 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t5 73.6304
R28260 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t1 60.3943
R28261 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n6 12.0358
R28262 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n8 0.981478
R28263 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.769522
R28264 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n0 0.745065
R28265 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.580578
R28266 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n4 0.533109
R28267 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.428234
R28268 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.063
R28269 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.063
R28270 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n3 0.063
R28271 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n5 0.063
R28272 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.063
R28273 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n7 0.063
R28274 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n1 0.063
R28275 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t3 316.762
R28276 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t0 169.195
R28277 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t4 150.887
R28278 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n2 150.273
R28279 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t5 74.951
R28280 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t2 73.6304
R28281 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t1 60.3943
R28282 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n6 12.0358
R28283 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n8 0.981478
R28284 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.769522
R28285 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n0 0.745065
R28286 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.580578
R28287 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n4 0.533109
R28288 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.428234
R28289 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.063
R28290 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.063
R28291 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n3 0.063
R28292 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n5 0.063
R28293 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.063
R28294 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n7 0.063
R28295 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n1 0.063
R28296 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 179.256
R28297 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 168.089
R28298 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 150.887
R28299 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 73.6304
R28300 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 60.3943
R28301 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 12.0358
R28302 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 1.05069
R28303 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 0.981478
R28304 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.769522
R28305 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 0.745065
R28306 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.580578
R28307 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 0.533109
R28308 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.428234
R28309 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.063
R28310 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 0.063
R28311 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 0.063
R28312 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.063
R28313 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 0.063
R28314 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 0.063
R28315 Ring_Counter_0.D_FlipFlop_14.Qbar.n4 Ring_Counter_0.D_FlipFlop_14.Qbar.t0 169.46
R28316 Ring_Counter_0.D_FlipFlop_14.Qbar.n4 Ring_Counter_0.D_FlipFlop_14.Qbar.t3 167.809
R28317 Ring_Counter_0.D_FlipFlop_14.Qbar.n3 Ring_Counter_0.D_FlipFlop_14.Qbar.t1 167.809
R28318 Ring_Counter_0.D_FlipFlop_14.Qbar.n1 Ring_Counter_0.D_FlipFlop_14.Qbar.t4 158.28
R28319 Ring_Counter_0.D_FlipFlop_14.Qbar.t4 Ring_Counter_0.D_FlipFlop_14.Qbar.n0 150.273
R28320 Ring_Counter_0.D_FlipFlop_14.Qbar.n0 Ring_Counter_0.D_FlipFlop_14.Qbar.t5 74.951
R28321 Ring_Counter_0.D_FlipFlop_14.Qbar.n6 Ring_Counter_0.D_FlipFlop_14.Qbar.t2 60.3943
R28322 Ring_Counter_0.D_FlipFlop_14.Qbar.n5 Ring_Counter_0.D_FlipFlop_14.Qbar.n4 11.4489
R28323 Ring_Counter_0.D_FlipFlop_14.Qbar.n3 Ring_Counter_0.D_FlipFlop_14.Qbar 8.5174
R28324 Ring_Counter_0.D_FlipFlop_14.Qbar.n6 Ring_Counter_0.D_FlipFlop_14.Qbar.n5 1.96917
R28325 Ring_Counter_0.D_FlipFlop_14.Qbar.n2 Ring_Counter_0.D_FlipFlop_14.Qbar.n1 0.42585
R28326 Ring_Counter_0.D_FlipFlop_14.Qbar.n1 Ring_Counter_0.D_FlipFlop_14.Qbar 0.390742
R28327 Ring_Counter_0.D_FlipFlop_14.Qbar.n5 Ring_Counter_0.D_FlipFlop_14.Qbar.n3 0.280391
R28328 Ring_Counter_0.D_FlipFlop_14.Qbar.n0 Ring_Counter_0.D_FlipFlop_14.Qbar 0.063
R28329 Ring_Counter_0.D_FlipFlop_14.Qbar Ring_Counter_0.D_FlipFlop_14.Qbar.n6 0.063
R28330 Ring_Counter_0.D_FlipFlop_14.Qbar.n2 Ring_Counter_0.D_FlipFlop_14.Qbar 0.00441667
R28331 Ring_Counter_0.D_FlipFlop_14.Qbar Ring_Counter_0.D_FlipFlop_14.Qbar.n2 0.00406061
R28332 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t0 169.46
R28333 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t1 167.809
R28334 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t2 167.809
R28335 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t6 167.226
R28336 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n6 150.273
R28337 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t5 150.273
R28338 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t7 74.951
R28339 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t4 73.6304
R28340 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t3 60.3943
R28341 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n4 12.3891
R28342 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n8 11.4489
R28343 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n10 1.68257
R28344 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n0 1.44615
R28345 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n2 1.2342
R28346 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 1.08448
R28347 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.932141
R28348 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n9 0.3496
R28349 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n7 0.280391
R28350 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.063
R28351 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.063
R28352 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n3 0.063
R28353 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.063
R28354 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n5 0.063
R28355 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n1 0.063
R28356 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t2 316.762
R28357 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t0 169.195
R28358 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t3 150.887
R28359 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n2 150.273
R28360 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t4 74.951
R28361 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t5 73.6304
R28362 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t1 60.3943
R28363 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n6 12.0358
R28364 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n8 0.981478
R28365 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.769522
R28366 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n0 0.745065
R28367 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.580578
R28368 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n4 0.533109
R28369 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.428234
R28370 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.063
R28371 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.063
R28372 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n3 0.063
R28373 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n5 0.063
R28374 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.063
R28375 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n7 0.063
R28376 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n1 0.063
R28377 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 179.256
R28378 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 168.089
R28379 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 150.887
R28380 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 73.6304
R28381 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 60.3943
R28382 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 12.0358
R28383 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 1.05069
R28384 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.981478
R28385 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.769522
R28386 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 0.745065
R28387 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.580578
R28388 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 0.533109
R28389 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.428234
R28390 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.063
R28391 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 0.063
R28392 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 0.063
R28393 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 0.063
R28394 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 0.063
R28395 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 0.063
R28396 D_FlipFlop_1.CLK.n12 D_FlipFlop_1.CLK.t0 168.108
R28397 D_FlipFlop_1.CLK.t2 D_FlipFlop_1.CLK.n5 158.207
R28398 D_FlipFlop_1.CLK D_FlipFlop_1.CLK.t3 158.202
R28399 D_FlipFlop_1.CLK.n0 D_FlipFlop_1.CLK.t5 150.293
R28400 D_FlipFlop_1.CLK.t3 D_FlipFlop_1.CLK.n3 150.293
R28401 D_FlipFlop_1.CLK.n6 D_FlipFlop_1.CLK.t2 150.273
R28402 D_FlipFlop_1.CLK.n9 D_FlipFlop_1.CLK.t4 90.1131
R28403 D_FlipFlop_1.CLK.t4 D_FlipFlop_1.CLK.n8 73.6406
R28404 D_FlipFlop_1.CLK.n2 D_FlipFlop_1.CLK.t6 73.6304
R28405 D_FlipFlop_1.CLK.n1 D_FlipFlop_1.CLK.t7 73.6304
R28406 D_FlipFlop_1.CLK D_FlipFlop_1.CLK.t1 60.3072
R28407 D_FlipFlop_1.CLK.n2 D_FlipFlop_1.CLK.n1 16.332
R28408 D_FlipFlop_1.CLK.n12 D_FlipFlop_1.CLK.n11 1.62007
R28409 D_FlipFlop_1.CLK.n8 D_FlipFlop_1.CLK.n7 1.19615
R28410 D_FlipFlop_1.CLK.n1 D_FlipFlop_1.CLK.n0 1.1717
R28411 D_FlipFlop_1.CLK.n3 D_FlipFlop_1.CLK.n2 1.1717
R28412 D_FlipFlop_1.CLK D_FlipFlop_1.CLK.n12 0.484875
R28413 D_FlipFlop_1.CLK.n3 D_FlipFlop_1.CLK 0.447191
R28414 D_FlipFlop_1.CLK.n0 D_FlipFlop_1.CLK 0.436162
R28415 D_FlipFlop_1.CLK.n5 D_FlipFlop_1.CLK.n4 0.349867
R28416 D_FlipFlop_1.CLK.n5 D_FlipFlop_1.CLK 0.321667
R28417 D_FlipFlop_1.CLK.n8 D_FlipFlop_1.CLK 0.217464
R28418 D_FlipFlop_1.CLK.n2 D_FlipFlop_1.CLK 0.149957
R28419 D_FlipFlop_1.CLK.n11 D_FlipFlop_1.CLK 0.149957
R28420 D_FlipFlop_1.CLK.n7 D_FlipFlop_1.CLK 0.1255
R28421 D_FlipFlop_1.CLK.n1 D_FlipFlop_1.CLK 0.117348
R28422 D_FlipFlop_1.CLK.n10 D_FlipFlop_1.CLK 0.0903438
R28423 D_FlipFlop_1.CLK.n1 D_FlipFlop_1.CLK 0.0454219
R28424 D_FlipFlop_1.CLK.n2 D_FlipFlop_1.CLK 0.0454219
R28425 D_FlipFlop_1.CLK.n10 D_FlipFlop_1.CLK.n9 0.027881
R28426 D_FlipFlop_1.CLK.n9 D_FlipFlop_1.CLK 0.027881
R28427 D_FlipFlop_1.CLK.n7 D_FlipFlop_1.CLK.n6 0.0216397
R28428 D_FlipFlop_1.CLK.n6 D_FlipFlop_1.CLK 0.0216397
R28429 D_FlipFlop_1.CLK.n11 D_FlipFlop_1.CLK.n10 0.0180781
R28430 D_FlipFlop_1.CLK.n4 D_FlipFlop_1.CLK 0.00441667
R28431 D_FlipFlop_1.CLK.n4 D_FlipFlop_1.CLK 0.00406061
R28432 D_FlipFlop_5.nPRE.n39 D_FlipFlop_5.nPRE.t2 169.46
R28433 D_FlipFlop_5.nPRE.n39 D_FlipFlop_5.nPRE.t3 167.809
R28434 D_FlipFlop_5.nPRE.n38 D_FlipFlop_5.nPRE.t1 167.809
R28435 D_FlipFlop_5.nPRE.n22 D_FlipFlop_5.nPRE.t15 161.88
R28436 D_FlipFlop_5.nPRE D_FlipFlop_5.nPRE.t10 158.581
R28437 D_FlipFlop_5.nPRE.n35 D_FlipFlop_5.nPRE.t4 158.565
R28438 D_FlipFlop_5.nPRE.t4 D_FlipFlop_5.nPRE.n34 151.594
R28439 D_FlipFlop_5.nPRE.t15 D_FlipFlop_5.nPRE.n21 150.293
R28440 D_FlipFlop_5.nPRE.t10 D_FlipFlop_5.nPRE.n2 150.293
R28441 D_FlipFlop_5.nPRE.n26 D_FlipFlop_5.nPRE.t16 150.273
R28442 D_FlipFlop_5.nPRE.n23 D_FlipFlop_5.nPRE.t11 150.273
R28443 D_FlipFlop_5.nPRE.n13 D_FlipFlop_5.nPRE.t12 150.273
R28444 D_FlipFlop_5.nPRE.n7 D_FlipFlop_5.nPRE.t6 150.273
R28445 D_FlipFlop_5.nPRE D_FlipFlop_5.nPRE.t17 99.8701
R28446 D_FlipFlop_5.nPRE.n25 D_FlipFlop_5.nPRE.t8 74.163
R28447 D_FlipFlop_5.nPRE.t17 D_FlipFlop_5.nPRE.n30 74.163
R28448 D_FlipFlop_5.nPRE.n11 D_FlipFlop_5.nPRE.t7 73.6406
R28449 D_FlipFlop_5.nPRE.n5 D_FlipFlop_5.nPRE.t14 73.6406
R28450 D_FlipFlop_5.nPRE.n34 D_FlipFlop_5.nPRE.t9 73.6304
R28451 D_FlipFlop_5.nPRE.n19 D_FlipFlop_5.nPRE.t5 73.6304
R28452 D_FlipFlop_5.nPRE.n0 D_FlipFlop_5.nPRE.t13 73.6304
R28453 D_FlipFlop_5.nPRE.n41 D_FlipFlop_5.nPRE.t0 62.1634
R28454 D_FlipFlop_5.nPRE.n17 D_FlipFlop_5.nPRE.n10 15.5222
R28455 D_FlipFlop_5.nPRE.n29 D_FlipFlop_5.nPRE.n28 12.6418
R28456 D_FlipFlop_5.nPRE.n40 D_FlipFlop_5.nPRE.n39 11.4489
R28457 D_FlipFlop_5.nPRE.n22 D_FlipFlop_5.nPRE.n18 9.02465
R28458 D_FlipFlop_5.nPRE.n18 D_FlipFlop_5.nPRE.n17 8.24202
R28459 D_FlipFlop_5.nPRE.n38 D_FlipFlop_5.nPRE.n37 8.21389
R28460 D_FlipFlop_5.nPRE.n32 D_FlipFlop_5.nPRE.n22 5.94458
R28461 D_FlipFlop_5.nPRE.n17 D_FlipFlop_5.nPRE.n16 4.5005
R28462 D_FlipFlop_5.nPRE.n33 D_FlipFlop_5.nPRE 1.2047
R28463 D_FlipFlop_5.nPRE.n21 D_FlipFlop_5.nPRE.n20 1.19615
R28464 D_FlipFlop_5.nPRE.n2 D_FlipFlop_5.nPRE.n1 1.19615
R28465 D_FlipFlop_5.nPRE.n32 D_FlipFlop_5.nPRE.n31 0.922483
R28466 D_FlipFlop_5.nPRE.n25 D_FlipFlop_5.nPRE 0.851043
R28467 D_FlipFlop_5.nPRE.n30 D_FlipFlop_5.nPRE 0.851043
R28468 D_FlipFlop_5.nPRE.n12 D_FlipFlop_5.nPRE.n11 0.796696
R28469 D_FlipFlop_5.nPRE.n6 D_FlipFlop_5.nPRE.n5 0.796696
R28470 D_FlipFlop_5.nPRE.n4 D_FlipFlop_5.nPRE.n3 0.783833
R28471 D_FlipFlop_5.nPRE.n4 D_FlipFlop_5.nPRE 0.716182
R28472 D_FlipFlop_5.nPRE.n27 D_FlipFlop_5.nPRE.n26 0.61463
R28473 D_FlipFlop_5.nPRE.n24 D_FlipFlop_5.nPRE.n23 0.61463
R28474 D_FlipFlop_5.nPRE.n12 D_FlipFlop_5.nPRE 0.524957
R28475 D_FlipFlop_5.nPRE.n6 D_FlipFlop_5.nPRE 0.524957
R28476 D_FlipFlop_5.nPRE.n27 D_FlipFlop_5.nPRE 0.486828
R28477 D_FlipFlop_5.nPRE.n24 D_FlipFlop_5.nPRE 0.486828
R28478 D_FlipFlop_5.nPRE.n21 D_FlipFlop_5.nPRE 0.447191
R28479 D_FlipFlop_5.nPRE.n2 D_FlipFlop_5.nPRE 0.447191
R28480 D_FlipFlop_5.nPRE.n37 D_FlipFlop_5.nPRE.n36 0.425067
R28481 D_FlipFlop_5.nPRE.n33 D_FlipFlop_5.nPRE.n32 0.399217
R28482 D_FlipFlop_5.nPRE.n37 D_FlipFlop_5.nPRE 0.39003
R28483 D_FlipFlop_5.nPRE.n40 D_FlipFlop_5.nPRE.n38 0.280391
R28484 D_FlipFlop_5.nPRE.n15 D_FlipFlop_5.nPRE 0.252453
R28485 D_FlipFlop_5.nPRE.n9 D_FlipFlop_5.nPRE 0.252453
R28486 D_FlipFlop_5.nPRE.n15 D_FlipFlop_5.nPRE.n14 0.226043
R28487 D_FlipFlop_5.nPRE.n9 D_FlipFlop_5.nPRE.n8 0.226043
R28488 D_FlipFlop_5.nPRE.n11 D_FlipFlop_5.nPRE 0.217464
R28489 D_FlipFlop_5.nPRE.n5 D_FlipFlop_5.nPRE 0.217464
R28490 D_FlipFlop_5.nPRE.n41 D_FlipFlop_5.nPRE.n40 0.200143
R28491 D_FlipFlop_5.nPRE.n20 D_FlipFlop_5.nPRE 0.1255
R28492 D_FlipFlop_5.nPRE.n14 D_FlipFlop_5.nPRE 0.1255
R28493 D_FlipFlop_5.nPRE.n8 D_FlipFlop_5.nPRE 0.1255
R28494 D_FlipFlop_5.nPRE.n1 D_FlipFlop_5.nPRE 0.1255
R28495 D_FlipFlop_5.nPRE.n34 D_FlipFlop_5.nPRE 0.063
R28496 D_FlipFlop_5.nPRE.n26 D_FlipFlop_5.nPRE 0.063
R28497 D_FlipFlop_5.nPRE.n28 D_FlipFlop_5.nPRE.n25 0.063
R28498 D_FlipFlop_5.nPRE.n28 D_FlipFlop_5.nPRE.n27 0.063
R28499 D_FlipFlop_5.nPRE.n23 D_FlipFlop_5.nPRE 0.063
R28500 D_FlipFlop_5.nPRE.n30 D_FlipFlop_5.nPRE.n29 0.063
R28501 D_FlipFlop_5.nPRE.n29 D_FlipFlop_5.nPRE.n24 0.063
R28502 D_FlipFlop_5.nPRE.n16 D_FlipFlop_5.nPRE.n12 0.063
R28503 D_FlipFlop_5.nPRE.n16 D_FlipFlop_5.nPRE.n15 0.063
R28504 D_FlipFlop_5.nPRE.n10 D_FlipFlop_5.nPRE.n6 0.063
R28505 D_FlipFlop_5.nPRE.n10 D_FlipFlop_5.nPRE.n9 0.063
R28506 D_FlipFlop_5.nPRE D_FlipFlop_5.nPRE.n41 0.063
R28507 D_FlipFlop_5.nPRE.n18 D_FlipFlop_5.nPRE.n4 0.024
R28508 D_FlipFlop_5.nPRE.n35 D_FlipFlop_5.nPRE.n33 0.024
R28509 D_FlipFlop_5.nPRE.n14 D_FlipFlop_5.nPRE.n13 0.0216397
R28510 D_FlipFlop_5.nPRE.n13 D_FlipFlop_5.nPRE 0.0216397
R28511 D_FlipFlop_5.nPRE.n8 D_FlipFlop_5.nPRE.n7 0.0216397
R28512 D_FlipFlop_5.nPRE.n7 D_FlipFlop_5.nPRE 0.0216397
R28513 D_FlipFlop_5.nPRE D_FlipFlop_5.nPRE.n35 0.0204394
R28514 D_FlipFlop_5.nPRE.n20 D_FlipFlop_5.nPRE.n19 0.0107679
R28515 D_FlipFlop_5.nPRE.n19 D_FlipFlop_5.nPRE 0.0107679
R28516 D_FlipFlop_5.nPRE.n1 D_FlipFlop_5.nPRE.n0 0.0107679
R28517 D_FlipFlop_5.nPRE.n0 D_FlipFlop_5.nPRE 0.0107679
R28518 D_FlipFlop_5.nPRE.n3 D_FlipFlop_5.nPRE 0.00441667
R28519 D_FlipFlop_5.nPRE.n31 D_FlipFlop_5.nPRE 0.00441667
R28520 D_FlipFlop_5.nPRE.n36 D_FlipFlop_5.nPRE 0.00441667
R28521 D_FlipFlop_5.nPRE.n31 D_FlipFlop_5.nPRE 0.00406061
R28522 D_FlipFlop_5.nPRE.n3 D_FlipFlop_5.nPRE 0.00406061
R28523 D_FlipFlop_5.nPRE.n36 D_FlipFlop_5.nPRE 0.00406061
R28524 Ring_Counter_0.D_FlipFlop_8.Qbar.n4 Ring_Counter_0.D_FlipFlop_8.Qbar.t0 169.46
R28525 Ring_Counter_0.D_FlipFlop_8.Qbar.n4 Ring_Counter_0.D_FlipFlop_8.Qbar.t3 167.809
R28526 Ring_Counter_0.D_FlipFlop_8.Qbar.n3 Ring_Counter_0.D_FlipFlop_8.Qbar.t1 167.809
R28527 Ring_Counter_0.D_FlipFlop_8.Qbar.n1 Ring_Counter_0.D_FlipFlop_8.Qbar.t5 158.28
R28528 Ring_Counter_0.D_FlipFlop_8.Qbar.t5 Ring_Counter_0.D_FlipFlop_8.Qbar.n0 150.273
R28529 Ring_Counter_0.D_FlipFlop_8.Qbar.n0 Ring_Counter_0.D_FlipFlop_8.Qbar.t4 74.951
R28530 Ring_Counter_0.D_FlipFlop_8.Qbar.n6 Ring_Counter_0.D_FlipFlop_8.Qbar.t2 60.3943
R28531 Ring_Counter_0.D_FlipFlop_8.Qbar.n5 Ring_Counter_0.D_FlipFlop_8.Qbar.n4 11.4489
R28532 Ring_Counter_0.D_FlipFlop_8.Qbar.n3 Ring_Counter_0.D_FlipFlop_8.Qbar 8.5174
R28533 Ring_Counter_0.D_FlipFlop_8.Qbar.n6 Ring_Counter_0.D_FlipFlop_8.Qbar.n5 1.96917
R28534 Ring_Counter_0.D_FlipFlop_8.Qbar.n2 Ring_Counter_0.D_FlipFlop_8.Qbar.n1 0.42585
R28535 Ring_Counter_0.D_FlipFlop_8.Qbar.n1 Ring_Counter_0.D_FlipFlop_8.Qbar 0.390742
R28536 Ring_Counter_0.D_FlipFlop_8.Qbar.n5 Ring_Counter_0.D_FlipFlop_8.Qbar.n3 0.280391
R28537 Ring_Counter_0.D_FlipFlop_8.Qbar.n0 Ring_Counter_0.D_FlipFlop_8.Qbar 0.063
R28538 Ring_Counter_0.D_FlipFlop_8.Qbar Ring_Counter_0.D_FlipFlop_8.Qbar.n6 0.063
R28539 Ring_Counter_0.D_FlipFlop_8.Qbar.n2 Ring_Counter_0.D_FlipFlop_8.Qbar 0.00441667
R28540 Ring_Counter_0.D_FlipFlop_8.Qbar Ring_Counter_0.D_FlipFlop_8.Qbar.n2 0.00406061
R28541 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 169.46
R28542 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 167.809
R28543 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 167.809
R28544 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 167.227
R28545 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 151.594
R28546 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 150.273
R28547 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 74.8641
R28548 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 73.6304
R28549 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 61.84
R28550 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 12.3891
R28551 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 11.4489
R28552 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R28553 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 0.280391
R28554 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 0.200143
R28555 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R28556 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R28557 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 0.149957
R28558 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.063
R28559 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 0.063
R28560 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 0.063
R28561 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 0.063
R28562 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R28563 Q1.n8 Q1.t2 169.46
R28564 Q1.n10 Q1.t0 167.809
R28565 Q1.n8 Q1.t3 167.809
R28566 Q1.n16 Q1.t5 158.565
R28567 Q1.n2 Q1.t9 150.543
R28568 Q1.n0 Q1.t8 150.543
R28569 Q1.t5 Q1.n15 150.293
R28570 Q1.n2 Q1.t4 74.4613
R28571 Q1.n0 Q1.t6 74.4613
R28572 Q1.n13 Q1.t7 73.6304
R28573 Q1.n6 Q1.t1 60.3809
R28574 Q1.n5 Q1.n4 12.1649
R28575 Q1.n9 Q1.n8 11.4489
R28576 Q1.n11 Q1.n10 8.21389
R28577 Q1.n17 Q1.n5 6.40503
R28578 Q1.n5 Q1 5.82352
R28579 Q1 Q1.n16 5.31642
R28580 Q1.n7 Q1.n6 1.64452
R28581 Q1.n15 Q1.n14 1.19615
R28582 Q1.n1 Q1 0.984196
R28583 Q1.n6 Q1 0.848156
R28584 Q1.n3 Q1.n2 0.747783
R28585 Q1.n1 Q1.n0 0.747783
R28586 Q1.n3 Q1 0.582531
R28587 Q1.n15 Q1 0.447191
R28588 Q1.n12 Q1.n11 0.425067
R28589 Q1.n11 Q1 0.39003
R28590 Q1.n10 Q1.n9 0.280391
R28591 Q1.n9 Q1 0.200143
R28592 Q1.n14 Q1 0.1255
R28593 Q1.n7 Q1 0.1255
R28594 Q1 Q1.n7 0.063
R28595 Q1.n2 Q1 0.063
R28596 Q1.n4 Q1.n1 0.063
R28597 Q1.n4 Q1.n3 0.063
R28598 Q1.n16 Q1 0.0204394
R28599 Q1.n14 Q1.n13 0.0107679
R28600 Q1.n13 Q1 0.0107679
R28601 Q1.n12 Q1 0.00441667
R28602 Q1 Q1.n12 0.00406061
R28603 Q1.n17 Q1 0.00128333
R28604 Q1.n17 Q1 0.00121212
R28605 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 169.46
R28606 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 168.089
R28607 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 167.809
R28608 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 150.887
R28609 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 73.6304
R28610 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 60.3943
R28611 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 12.0358
R28612 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 11.4489
R28613 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 1.05069
R28614 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 0.981478
R28615 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.769522
R28616 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 0.745065
R28617 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.580578
R28618 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 0.533109
R28619 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.428234
R28620 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.063
R28621 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 0.063
R28622 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 0.063
R28623 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.063
R28624 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 0.063
R28625 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 0.063
R28626 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.t3 169.46
R28627 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.t2 167.809
R28628 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.t0 167.809
R28629 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.t4 167.226
R28630 D_FlipFlop_4.3-input-nand_2.C.t4 D_FlipFlop_4.3-input-nand_2.C.n10 150.273
R28631 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C.t5 150.273
R28632 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C.t6 73.6406
R28633 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C.t7 73.6304
R28634 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_2.C.t1 60.3943
R28635 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C.n5 12.3891
R28636 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C.n12 11.4489
R28637 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C 1.68257
R28638 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C.n0 1.38365
R28639 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C.n8 1.19615
R28640 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C.n3 1.1717
R28641 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C 1.08448
R28642 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C 0.932141
R28643 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_2.C.n14 0.720633
R28644 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C.n11 0.280391
R28645 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C 0.217464
R28646 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C 0.1255
R28647 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C 0.1255
R28648 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C 0.1255
R28649 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.n7 0.0874565
R28650 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C.n4 0.063
R28651 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C 0.063
R28652 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C.n6 0.063
R28653 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C.n1 0.063
R28654 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.n13 0.0435206
R28655 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C.n9 0.0216397
R28656 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C 0.0216397
R28657 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C.n2 0.0107679
R28658 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C 0.0107679
R28659 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t2 169.46
R28660 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t3 167.809
R28661 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.t0 167.809
R28662 D_FlipFlop_4.3-input-nand_2.Vout.t4 D_FlipFlop_4.3-input-nand_2.Vout.n11 167.227
R28663 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.t4 150.293
R28664 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.t7 150.273
R28665 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout.t5 73.6406
R28666 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6304
R28667 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout.t1 60.3809
R28668 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n5 12.3891
R28669 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout.n9 11.4489
R28670 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout.n2 1.38365
R28671 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.n1 1.19615
R28672 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.n4 1.1717
R28673 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout 0.848156
R28674 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.Vout.n12 0.447191
R28675 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout 0.38637
R28676 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.n10 0.280391
R28677 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout 0.217464
R28678 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout 0.200143
R28679 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R28680 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R28681 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R28682 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R28683 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout.n7 0.0874565
R28684 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n3 0.063
R28685 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout.n6 0.063
R28686 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.Vout.n8 0.063
R28687 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R28688 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout.n0 0.0107679
R28689 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout 0.0107679
R28690 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 169.46
R28691 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 167.809
R28692 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 167.809
R28693 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 167.227
R28694 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 151.594
R28695 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 150.273
R28696 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 74.8641
R28697 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 73.6304
R28698 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 61.84
R28699 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 12.3891
R28700 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 11.4489
R28701 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.38637
R28702 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 0.280391
R28703 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 0.200143
R28704 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.152844
R28705 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.149957
R28706 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 0.149957
R28707 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.063
R28708 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 0.063
R28709 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 0.063
R28710 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 0.063
R28711 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.0454219
R28712 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t0 169.46
R28713 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t3 167.809
R28714 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t2 167.809
R28715 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t5 167.226
R28716 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n6 150.273
R28717 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t7 150.273
R28718 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t6 74.951
R28719 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t4 73.6304
R28720 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t1 60.3943
R28721 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n4 12.3891
R28722 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n8 11.4489
R28723 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n10 1.68257
R28724 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n0 1.44615
R28725 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n2 1.2342
R28726 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 1.08448
R28727 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.932141
R28728 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n9 0.3496
R28729 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n7 0.280391
R28730 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.063
R28731 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.063
R28732 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n3 0.063
R28733 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.063
R28734 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n5 0.063
R28735 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n1 0.063
R28736 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t3 316.762
R28737 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t0 169.195
R28738 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t4 150.887
R28739 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n2 150.273
R28740 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t5 74.951
R28741 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t2 73.6304
R28742 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t1 60.3943
R28743 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n6 12.0358
R28744 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n8 0.981478
R28745 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.769522
R28746 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n0 0.745065
R28747 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.580578
R28748 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n4 0.533109
R28749 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.428234
R28750 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.063
R28751 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.063
R28752 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n3 0.063
R28753 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n5 0.063
R28754 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.063
R28755 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n7 0.063
R28756 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n1 0.063
R28757 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 179.256
R28758 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 168.089
R28759 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 150.887
R28760 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 73.6304
R28761 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 60.3943
R28762 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 12.0358
R28763 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 1.05069
R28764 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 0.981478
R28765 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.769522
R28766 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 0.745065
R28767 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.580578
R28768 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 0.533109
R28769 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.428234
R28770 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.063
R28771 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 0.063
R28772 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 0.063
R28773 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.063
R28774 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 0.063
R28775 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 0.063
R28776 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.t3 169.46
R28777 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout.t2 167.809
R28778 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.t0 167.809
R28779 D_FlipFlop_6.3-input-nand_2.Vout.t5 D_FlipFlop_6.3-input-nand_2.Vout.n11 167.227
R28780 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.t5 150.293
R28781 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.t4 150.273
R28782 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout.t6 73.6406
R28783 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout.t7 73.6304
R28784 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout.t1 60.3809
R28785 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout.n5 12.3891
R28786 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout.n9 11.4489
R28787 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout.n2 1.38365
R28788 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.n1 1.19615
R28789 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.n4 1.1717
R28790 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout 0.848156
R28791 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.Vout.n12 0.447191
R28792 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R28793 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout.n10 0.280391
R28794 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout 0.217464
R28795 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout 0.200143
R28796 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R28797 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R28798 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R28799 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R28800 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout.n7 0.0874565
R28801 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout.n3 0.063
R28802 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout.n6 0.063
R28803 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.Vout.n8 0.063
R28804 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R28805 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout.n0 0.0107679
R28806 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout 0.0107679
R28807 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 169.46
R28808 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 167.809
R28809 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 167.809
R28810 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 167.227
R28811 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 151.594
R28812 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 150.273
R28813 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 74.8641
R28814 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 73.6304
R28815 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 61.84
R28816 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 12.3891
R28817 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 11.4489
R28818 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.38637
R28819 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 0.280391
R28820 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 0.200143
R28821 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.152844
R28822 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.149957
R28823 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 0.149957
R28824 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.063
R28825 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 0.063
R28826 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 0.063
R28827 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 0.063
R28828 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.0454219
R28829 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 169.46
R28830 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 167.809
R28831 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 167.809
R28832 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 167.227
R28833 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 151.594
R28834 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 150.273
R28835 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 74.8641
R28836 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 73.6304
R28837 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 61.84
R28838 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 12.3891
R28839 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 11.4489
R28840 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 0.38637
R28841 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 0.280391
R28842 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 0.200143
R28843 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.152844
R28844 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.149957
R28845 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 0.149957
R28846 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.063
R28847 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.063
R28848 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 0.063
R28849 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 0.063
R28850 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.0454219
R28851 CDAC_v3_0.switch_0.Z.n0 CDAC_v3_0.switch_0.Z.t4 168.075
R28852 CDAC_v3_0.switch_0.Z.n0 CDAC_v3_0.switch_0.Z.t1 168.075
R28853 CDAC_v3_0.switch_0.Z.n4 CDAC_v3_0.switch_0.Z.n3 69.4722
R28854 CDAC_v3_0.switch_0.Z.n6 CDAC_v3_0.switch_0.Z.t0 60.6851
R28855 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_0.Z.t5 60.6226
R28856 CDAC_v3_0.switch_0.Z.n3 CDAC_v3_0.switch_0.Z.t3 21.3216
R28857 CDAC_v3_0.switch_0.Z.n2 CDAC_v3_0.switch_0.Z.n1 1.34289
R28858 CDAC_v3_0.switch_0.Z.n2 CDAC_v3_0.switch_0.Z 0.42713
R28859 CDAC_v3_0.switch_0.Z.n3 CDAC_v3_0.switch_0.Z.t2 0.307567
R28860 CDAC_v3_0.switch_0.Z.n5 CDAC_v3_0.switch_0.Z 0.182141
R28861 CDAC_v3_0.switch_0.Z.n1 CDAC_v3_0.switch_0.Z 0.178175
R28862 CDAC_v3_0.switch_0.Z.n6 CDAC_v3_0.switch_0.Z.n5 0.128217
R28863 CDAC_v3_0.switch_0.Z.n6 CDAC_v3_0.switch_0.Z 0.1255
R28864 CDAC_v3_0.switch_0.Z.n4 CDAC_v3_0.switch_0.Z.n2 0.063
R28865 CDAC_v3_0.switch_0.Z.n5 CDAC_v3_0.switch_0.Z.n4 0.063
R28866 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_0.Z.n6 0.063
R28867 CDAC_v3_0.switch_0.Z.n1 CDAC_v3_0.switch_0.Z.n0 0.0130546
R28868 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 179.256
R28869 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 168.089
R28870 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 150.887
R28871 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 73.6304
R28872 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 60.3943
R28873 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 12.0358
R28874 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 1.05069
R28875 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 0.981478
R28876 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.769522
R28877 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 0.745065
R28878 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.580578
R28879 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 0.533109
R28880 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.428234
R28881 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.063
R28882 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 0.063
R28883 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 0.063
R28884 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.063
R28885 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 0.063
R28886 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 0.063
R28887 CDAC_v3_0.switch_2.Z.n7 CDAC_v3_0.switch_2.Z.t7 168.075
R28888 CDAC_v3_0.switch_2.Z.n7 CDAC_v3_0.switch_2.Z.t0 168.075
R28889 CDAC_v3_0.switch_2.Z.n0 CDAC_v3_0.switch_2.Z.t6 60.6851
R28890 CDAC_v3_0.switch_2.Z CDAC_v3_0.switch_2.Z.t1 60.6226
R28891 CDAC_v3_0.switch_2.Z.n5 CDAC_v3_0.switch_2.Z.n4 49.1102
R28892 CDAC_v3_0.switch_2.Z.n3 CDAC_v3_0.switch_2.Z.n2 16.5787
R28893 CDAC_v3_0.switch_2.Z.n2 CDAC_v3_0.switch_2.Z.t2 13.7008
R28894 CDAC_v3_0.switch_2.Z.n3 CDAC_v3_0.switch_2.Z.t4 7.43126
R28895 CDAC_v3_0.switch_2.Z.n4 CDAC_v3_0.switch_2.Z.n3 6.26999
R28896 CDAC_v3_0.switch_2.Z.n8 CDAC_v3_0.switch_2.Z.n6 1.34289
R28897 CDAC_v3_0.switch_2.Z.n6 CDAC_v3_0.switch_2.Z 0.42713
R28898 CDAC_v3_0.switch_2.Z.n2 CDAC_v3_0.switch_2.Z.t5 0.307567
R28899 CDAC_v3_0.switch_2.Z.n4 CDAC_v3_0.switch_2.Z.t3 0.307567
R28900 CDAC_v3_0.switch_2.Z.n1 CDAC_v3_0.switch_2.Z 0.182141
R28901 CDAC_v3_0.switch_2.Z CDAC_v3_0.switch_2.Z.n8 0.178175
R28902 CDAC_v3_0.switch_2.Z.n1 CDAC_v3_0.switch_2.Z.n0 0.128217
R28903 CDAC_v3_0.switch_2.Z.n0 CDAC_v3_0.switch_2.Z 0.1255
R28904 CDAC_v3_0.switch_2.Z.n0 CDAC_v3_0.switch_2.Z 0.063
R28905 CDAC_v3_0.switch_2.Z.n6 CDAC_v3_0.switch_2.Z.n5 0.063
R28906 CDAC_v3_0.switch_2.Z.n5 CDAC_v3_0.switch_2.Z.n1 0.063
R28907 CDAC_v3_0.switch_2.Z.n8 CDAC_v3_0.switch_2.Z.n7 0.0130546
R28908 Nand_Gate_2.A.n19 Nand_Gate_2.A.t3 169.46
R28909 Nand_Gate_2.A.n18 Nand_Gate_2.A.t2 167.809
R28910 Nand_Gate_2.A.n19 Nand_Gate_2.A.t0 167.809
R28911 Nand_Gate_2.A.n12 Nand_Gate_2.A.t10 159.107
R28912 Nand_Gate_2.A.n15 Nand_Gate_2.A.t9 158.565
R28913 Nand_Gate_2.A.t9 Nand_Gate_2.A.n14 151.594
R28914 Nand_Gate_2.A.t10 Nand_Gate_2.A.n2 150.293
R28915 Nand_Gate_2.A.n6 Nand_Gate_2.A.t4 150.273
R28916 Nand_Gate_2.A.n3 Nand_Gate_2.A.t8 150.273
R28917 Nand_Gate_2.A Nand_Gate_2.A.t7 99.8701
R28918 Nand_Gate_2.A.n5 Nand_Gate_2.A.t5 74.163
R28919 Nand_Gate_2.A.t7 Nand_Gate_2.A.n10 74.163
R28920 Nand_Gate_2.A.n14 Nand_Gate_2.A.t6 73.6304
R28921 Nand_Gate_2.A.n0 Nand_Gate_2.A.t11 73.6304
R28922 Nand_Gate_2.A.n21 Nand_Gate_2.A.t1 62.1634
R28923 Nand_Gate_2.A.n9 Nand_Gate_2.A.n8 12.6418
R28924 Nand_Gate_2.A.n20 Nand_Gate_2.A.n19 11.4489
R28925 Nand_Gate_2.A.n18 Nand_Gate_2.A.n17 8.21389
R28926 Nand_Gate_2.A.n13 Nand_Gate_2.A 1.2047
R28927 Nand_Gate_2.A.n2 Nand_Gate_2.A.n1 1.19615
R28928 Nand_Gate_2.A.n12 Nand_Gate_2.A.n11 1.00082
R28929 Nand_Gate_2.A.n5 Nand_Gate_2.A 0.851043
R28930 Nand_Gate_2.A.n10 Nand_Gate_2.A 0.851043
R28931 Nand_Gate_2.A.n7 Nand_Gate_2.A.n6 0.61463
R28932 Nand_Gate_2.A.n4 Nand_Gate_2.A.n3 0.61463
R28933 Nand_Gate_2.A.n7 Nand_Gate_2.A 0.486828
R28934 Nand_Gate_2.A.n4 Nand_Gate_2.A 0.486828
R28935 Nand_Gate_2.A.n2 Nand_Gate_2.A 0.447191
R28936 Nand_Gate_2.A.n17 Nand_Gate_2.A.n16 0.425067
R28937 Nand_Gate_2.A.n17 Nand_Gate_2.A 0.39003
R28938 Nand_Gate_2.A.n13 Nand_Gate_2.A.n12 0.320883
R28939 Nand_Gate_2.A.n20 Nand_Gate_2.A.n18 0.280391
R28940 Nand_Gate_2.A.n21 Nand_Gate_2.A.n20 0.200143
R28941 Nand_Gate_2.A.n1 Nand_Gate_2.A 0.1255
R28942 Nand_Gate_2.A.n14 Nand_Gate_2.A 0.063
R28943 Nand_Gate_2.A.n6 Nand_Gate_2.A 0.063
R28944 Nand_Gate_2.A.n8 Nand_Gate_2.A.n5 0.063
R28945 Nand_Gate_2.A.n8 Nand_Gate_2.A.n7 0.063
R28946 Nand_Gate_2.A.n3 Nand_Gate_2.A 0.063
R28947 Nand_Gate_2.A.n10 Nand_Gate_2.A.n9 0.063
R28948 Nand_Gate_2.A.n9 Nand_Gate_2.A.n4 0.063
R28949 Nand_Gate_2.A Nand_Gate_2.A.n21 0.063
R28950 Nand_Gate_2.A.n15 Nand_Gate_2.A.n13 0.024
R28951 Nand_Gate_2.A Nand_Gate_2.A.n15 0.0204394
R28952 Nand_Gate_2.A.n1 Nand_Gate_2.A.n0 0.0107679
R28953 Nand_Gate_2.A.n0 Nand_Gate_2.A 0.0107679
R28954 Nand_Gate_2.A.n11 Nand_Gate_2.A 0.00441667
R28955 Nand_Gate_2.A.n16 Nand_Gate_2.A 0.00441667
R28956 Nand_Gate_2.A.n11 Nand_Gate_2.A 0.00406061
R28957 Nand_Gate_2.A.n16 Nand_Gate_2.A 0.00406061
R28958 Ring_Counter_0.D_FlipFlop_5.Qbar.n4 Ring_Counter_0.D_FlipFlop_5.Qbar.t3 169.46
R28959 Ring_Counter_0.D_FlipFlop_5.Qbar.n4 Ring_Counter_0.D_FlipFlop_5.Qbar.t1 167.809
R28960 Ring_Counter_0.D_FlipFlop_5.Qbar.n3 Ring_Counter_0.D_FlipFlop_5.Qbar.t2 167.809
R28961 Ring_Counter_0.D_FlipFlop_5.Qbar.n1 Ring_Counter_0.D_FlipFlop_5.Qbar.t4 158.28
R28962 Ring_Counter_0.D_FlipFlop_5.Qbar.t4 Ring_Counter_0.D_FlipFlop_5.Qbar.n0 150.273
R28963 Ring_Counter_0.D_FlipFlop_5.Qbar.n0 Ring_Counter_0.D_FlipFlop_5.Qbar.t5 74.951
R28964 Ring_Counter_0.D_FlipFlop_5.Qbar.n6 Ring_Counter_0.D_FlipFlop_5.Qbar.t0 60.3943
R28965 Ring_Counter_0.D_FlipFlop_5.Qbar.n5 Ring_Counter_0.D_FlipFlop_5.Qbar.n4 11.4489
R28966 Ring_Counter_0.D_FlipFlop_5.Qbar.n3 Ring_Counter_0.D_FlipFlop_5.Qbar 8.5174
R28967 Ring_Counter_0.D_FlipFlop_5.Qbar.n6 Ring_Counter_0.D_FlipFlop_5.Qbar.n5 1.96917
R28968 Ring_Counter_0.D_FlipFlop_5.Qbar.n2 Ring_Counter_0.D_FlipFlop_5.Qbar.n1 0.42585
R28969 Ring_Counter_0.D_FlipFlop_5.Qbar.n1 Ring_Counter_0.D_FlipFlop_5.Qbar 0.390742
R28970 Ring_Counter_0.D_FlipFlop_5.Qbar.n5 Ring_Counter_0.D_FlipFlop_5.Qbar.n3 0.280391
R28971 Ring_Counter_0.D_FlipFlop_5.Qbar.n0 Ring_Counter_0.D_FlipFlop_5.Qbar 0.063
R28972 Ring_Counter_0.D_FlipFlop_5.Qbar Ring_Counter_0.D_FlipFlop_5.Qbar.n6 0.063
R28973 Ring_Counter_0.D_FlipFlop_5.Qbar.n2 Ring_Counter_0.D_FlipFlop_5.Qbar 0.00441667
R28974 Ring_Counter_0.D_FlipFlop_5.Qbar Ring_Counter_0.D_FlipFlop_5.Qbar.n2 0.00406061
R28975 Nand_Gate_4.A.n12 Nand_Gate_4.A.t6 169.827
R28976 Nand_Gate_4.A.n19 Nand_Gate_4.A.t3 169.46
R28977 Nand_Gate_4.A.n18 Nand_Gate_4.A.t1 167.809
R28978 Nand_Gate_4.A.n19 Nand_Gate_4.A.t0 167.809
R28979 Nand_Gate_4.A.n15 Nand_Gate_4.A.t4 158.565
R28980 Nand_Gate_4.A.t4 Nand_Gate_4.A.n14 151.594
R28981 Nand_Gate_4.A.t6 Nand_Gate_4.A.n2 150.293
R28982 Nand_Gate_4.A.n6 Nand_Gate_4.A.t5 150.273
R28983 Nand_Gate_4.A.n3 Nand_Gate_4.A.t10 150.273
R28984 Nand_Gate_4.A Nand_Gate_4.A.t11 99.8701
R28985 Nand_Gate_4.A.n5 Nand_Gate_4.A.t9 74.163
R28986 Nand_Gate_4.A.t11 Nand_Gate_4.A.n10 74.163
R28987 Nand_Gate_4.A.n14 Nand_Gate_4.A.t8 73.6304
R28988 Nand_Gate_4.A.n0 Nand_Gate_4.A.t7 73.6304
R28989 Nand_Gate_4.A.n21 Nand_Gate_4.A.t2 62.1634
R28990 Nand_Gate_4.A.n9 Nand_Gate_4.A.n8 12.6418
R28991 Nand_Gate_4.A.n20 Nand_Gate_4.A.n19 11.4489
R28992 Nand_Gate_4.A.n18 Nand_Gate_4.A.n17 8.21389
R28993 Nand_Gate_4.A.n13 Nand_Gate_4.A 1.2047
R28994 Nand_Gate_4.A.n2 Nand_Gate_4.A.n1 1.19615
R28995 Nand_Gate_4.A.n12 Nand_Gate_4.A.n11 0.922483
R28996 Nand_Gate_4.A.n5 Nand_Gate_4.A 0.851043
R28997 Nand_Gate_4.A.n10 Nand_Gate_4.A 0.851043
R28998 Nand_Gate_4.A.n7 Nand_Gate_4.A.n6 0.61463
R28999 Nand_Gate_4.A.n4 Nand_Gate_4.A.n3 0.61463
R29000 Nand_Gate_4.A.n7 Nand_Gate_4.A 0.486828
R29001 Nand_Gate_4.A.n4 Nand_Gate_4.A 0.486828
R29002 Nand_Gate_4.A.n2 Nand_Gate_4.A 0.447191
R29003 Nand_Gate_4.A.n17 Nand_Gate_4.A.n16 0.425067
R29004 Nand_Gate_4.A.n13 Nand_Gate_4.A.n12 0.399217
R29005 Nand_Gate_4.A.n17 Nand_Gate_4.A 0.39003
R29006 Nand_Gate_4.A.n20 Nand_Gate_4.A.n18 0.280391
R29007 Nand_Gate_4.A.n21 Nand_Gate_4.A.n20 0.200143
R29008 Nand_Gate_4.A.n1 Nand_Gate_4.A 0.1255
R29009 Nand_Gate_4.A.n14 Nand_Gate_4.A 0.063
R29010 Nand_Gate_4.A.n6 Nand_Gate_4.A 0.063
R29011 Nand_Gate_4.A.n8 Nand_Gate_4.A.n5 0.063
R29012 Nand_Gate_4.A.n8 Nand_Gate_4.A.n7 0.063
R29013 Nand_Gate_4.A.n3 Nand_Gate_4.A 0.063
R29014 Nand_Gate_4.A.n10 Nand_Gate_4.A.n9 0.063
R29015 Nand_Gate_4.A.n9 Nand_Gate_4.A.n4 0.063
R29016 Nand_Gate_4.A Nand_Gate_4.A.n21 0.063
R29017 Nand_Gate_4.A.n15 Nand_Gate_4.A.n13 0.024
R29018 Nand_Gate_4.A Nand_Gate_4.A.n15 0.0204394
R29019 Nand_Gate_4.A.n1 Nand_Gate_4.A.n0 0.0107679
R29020 Nand_Gate_4.A.n0 Nand_Gate_4.A 0.0107679
R29021 Nand_Gate_4.A.n11 Nand_Gate_4.A 0.00441667
R29022 Nand_Gate_4.A.n16 Nand_Gate_4.A 0.00441667
R29023 Nand_Gate_4.A.n11 Nand_Gate_4.A 0.00406061
R29024 Nand_Gate_4.A.n16 Nand_Gate_4.A 0.00406061
R29025 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 179.256
R29026 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 168.089
R29027 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 150.887
R29028 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 73.6304
R29029 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 60.3943
R29030 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 12.0358
R29031 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 1.05069
R29032 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 0.981478
R29033 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.769522
R29034 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 0.745065
R29035 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.580578
R29036 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 0.533109
R29037 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.428234
R29038 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.063
R29039 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 0.063
R29040 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 0.063
R29041 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.063
R29042 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 0.063
R29043 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 0.063
R29044 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 179.256
R29045 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 168.089
R29046 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 150.887
R29047 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 73.6304
R29048 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 60.3943
R29049 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 12.0358
R29050 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 1.05069
R29051 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.981478
R29052 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.769522
R29053 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 0.745065
R29054 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.580578
R29055 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 0.533109
R29056 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.428234
R29057 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.063
R29058 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 0.063
R29059 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 0.063
R29060 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 0.063
R29061 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 0.063
R29062 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 0.063
R29063 Ring_Counter_0.D_FlipFlop_11.Qbar.n4 Ring_Counter_0.D_FlipFlop_11.Qbar.t0 169.46
R29064 Ring_Counter_0.D_FlipFlop_11.Qbar.n4 Ring_Counter_0.D_FlipFlop_11.Qbar.t3 167.809
R29065 Ring_Counter_0.D_FlipFlop_11.Qbar.n3 Ring_Counter_0.D_FlipFlop_11.Qbar.t1 167.809
R29066 Ring_Counter_0.D_FlipFlop_11.Qbar.n1 Ring_Counter_0.D_FlipFlop_11.Qbar.t5 158.28
R29067 Ring_Counter_0.D_FlipFlop_11.Qbar.t5 Ring_Counter_0.D_FlipFlop_11.Qbar.n0 150.273
R29068 Ring_Counter_0.D_FlipFlop_11.Qbar.n0 Ring_Counter_0.D_FlipFlop_11.Qbar.t4 74.951
R29069 Ring_Counter_0.D_FlipFlop_11.Qbar.n6 Ring_Counter_0.D_FlipFlop_11.Qbar.t2 60.3943
R29070 Ring_Counter_0.D_FlipFlop_11.Qbar.n5 Ring_Counter_0.D_FlipFlop_11.Qbar.n4 11.4489
R29071 Ring_Counter_0.D_FlipFlop_11.Qbar.n3 Ring_Counter_0.D_FlipFlop_11.Qbar 8.5174
R29072 Ring_Counter_0.D_FlipFlop_11.Qbar.n6 Ring_Counter_0.D_FlipFlop_11.Qbar.n5 1.96917
R29073 Ring_Counter_0.D_FlipFlop_11.Qbar.n2 Ring_Counter_0.D_FlipFlop_11.Qbar.n1 0.42585
R29074 Ring_Counter_0.D_FlipFlop_11.Qbar.n1 Ring_Counter_0.D_FlipFlop_11.Qbar 0.390742
R29075 Ring_Counter_0.D_FlipFlop_11.Qbar.n5 Ring_Counter_0.D_FlipFlop_11.Qbar.n3 0.280391
R29076 Ring_Counter_0.D_FlipFlop_11.Qbar.n0 Ring_Counter_0.D_FlipFlop_11.Qbar 0.063
R29077 Ring_Counter_0.D_FlipFlop_11.Qbar Ring_Counter_0.D_FlipFlop_11.Qbar.n6 0.063
R29078 Ring_Counter_0.D_FlipFlop_11.Qbar.n2 Ring_Counter_0.D_FlipFlop_11.Qbar 0.00441667
R29079 Ring_Counter_0.D_FlipFlop_11.Qbar Ring_Counter_0.D_FlipFlop_11.Qbar.n2 0.00406061
R29080 Nand_Gate_7.A.n12 Nand_Gate_7.A.t7 172.387
R29081 Nand_Gate_7.A.n19 Nand_Gate_7.A.t1 169.46
R29082 Nand_Gate_7.A.n18 Nand_Gate_7.A.t3 167.809
R29083 Nand_Gate_7.A.n19 Nand_Gate_7.A.t0 167.809
R29084 Nand_Gate_7.A.n15 Nand_Gate_7.A.t5 158.565
R29085 Nand_Gate_7.A.t5 Nand_Gate_7.A.n14 151.594
R29086 Nand_Gate_7.A.t7 Nand_Gate_7.A.n2 150.293
R29087 Nand_Gate_7.A.n6 Nand_Gate_7.A.t4 150.273
R29088 Nand_Gate_7.A.n3 Nand_Gate_7.A.t11 150.273
R29089 Nand_Gate_7.A Nand_Gate_7.A.t10 99.8701
R29090 Nand_Gate_7.A.n5 Nand_Gate_7.A.t6 74.163
R29091 Nand_Gate_7.A.t10 Nand_Gate_7.A.n10 74.163
R29092 Nand_Gate_7.A.n14 Nand_Gate_7.A.t9 73.6304
R29093 Nand_Gate_7.A.n0 Nand_Gate_7.A.t8 73.6304
R29094 Nand_Gate_7.A.n21 Nand_Gate_7.A.t2 62.1634
R29095 Nand_Gate_7.A.n9 Nand_Gate_7.A.n8 12.6418
R29096 Nand_Gate_7.A.n20 Nand_Gate_7.A.n19 11.4489
R29097 Nand_Gate_7.A.n18 Nand_Gate_7.A.n17 8.21389
R29098 Nand_Gate_7.A.n13 Nand_Gate_7.A 1.2047
R29099 Nand_Gate_7.A.n2 Nand_Gate_7.A.n1 1.19615
R29100 Nand_Gate_7.A.n12 Nand_Gate_7.A.n11 0.922483
R29101 Nand_Gate_7.A.n5 Nand_Gate_7.A 0.851043
R29102 Nand_Gate_7.A.n10 Nand_Gate_7.A 0.851043
R29103 Nand_Gate_7.A.n7 Nand_Gate_7.A.n6 0.61463
R29104 Nand_Gate_7.A.n4 Nand_Gate_7.A.n3 0.61463
R29105 Nand_Gate_7.A.n7 Nand_Gate_7.A 0.486828
R29106 Nand_Gate_7.A.n4 Nand_Gate_7.A 0.486828
R29107 Nand_Gate_7.A.n2 Nand_Gate_7.A 0.447191
R29108 Nand_Gate_7.A.n17 Nand_Gate_7.A.n16 0.425067
R29109 Nand_Gate_7.A.n13 Nand_Gate_7.A.n12 0.399217
R29110 Nand_Gate_7.A.n17 Nand_Gate_7.A 0.39003
R29111 Nand_Gate_7.A.n20 Nand_Gate_7.A.n18 0.280391
R29112 Nand_Gate_7.A.n21 Nand_Gate_7.A.n20 0.200143
R29113 Nand_Gate_7.A.n1 Nand_Gate_7.A 0.1255
R29114 Nand_Gate_7.A.n14 Nand_Gate_7.A 0.063
R29115 Nand_Gate_7.A.n6 Nand_Gate_7.A 0.063
R29116 Nand_Gate_7.A.n8 Nand_Gate_7.A.n5 0.063
R29117 Nand_Gate_7.A.n8 Nand_Gate_7.A.n7 0.063
R29118 Nand_Gate_7.A.n3 Nand_Gate_7.A 0.063
R29119 Nand_Gate_7.A.n10 Nand_Gate_7.A.n9 0.063
R29120 Nand_Gate_7.A.n9 Nand_Gate_7.A.n4 0.063
R29121 Nand_Gate_7.A Nand_Gate_7.A.n21 0.063
R29122 Nand_Gate_7.A.n15 Nand_Gate_7.A.n13 0.024
R29123 Nand_Gate_7.A Nand_Gate_7.A.n15 0.0204394
R29124 Nand_Gate_7.A.n1 Nand_Gate_7.A.n0 0.0107679
R29125 Nand_Gate_7.A.n0 Nand_Gate_7.A 0.0107679
R29126 Nand_Gate_7.A.n11 Nand_Gate_7.A 0.00441667
R29127 Nand_Gate_7.A.n16 Nand_Gate_7.A 0.00441667
R29128 Nand_Gate_7.A.n11 Nand_Gate_7.A 0.00406061
R29129 Nand_Gate_7.A.n16 Nand_Gate_7.A 0.00406061
R29130 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t0 169.46
R29131 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t3 167.809
R29132 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t1 167.809
R29133 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t7 167.226
R29134 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n6 150.273
R29135 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t5 150.273
R29136 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t6 74.951
R29137 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t4 73.6304
R29138 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t2 60.3943
R29139 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n4 12.3891
R29140 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n8 11.4489
R29141 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n10 1.68257
R29142 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n0 1.44615
R29143 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n2 1.2342
R29144 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 1.08448
R29145 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.932141
R29146 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n9 0.3496
R29147 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n7 0.280391
R29148 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.063
R29149 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.063
R29150 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n3 0.063
R29151 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.063
R29152 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n5 0.063
R29153 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n1 0.063
R29154 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t5 316.762
R29155 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t0 169.195
R29156 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t3 150.887
R29157 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n2 150.273
R29158 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t4 74.951
R29159 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t2 73.6304
R29160 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t1 60.3943
R29161 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n6 12.0358
R29162 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n8 0.981478
R29163 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.769522
R29164 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n0 0.745065
R29165 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.580578
R29166 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n4 0.533109
R29167 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.428234
R29168 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.063
R29169 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.063
R29170 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n3 0.063
R29171 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n5 0.063
R29172 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.063
R29173 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n7 0.063
R29174 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n1 0.063
R29175 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 179.256
R29176 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 168.089
R29177 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 150.887
R29178 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 73.6304
R29179 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 60.3943
R29180 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 12.0358
R29181 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 1.05069
R29182 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 0.981478
R29183 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.769522
R29184 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 0.745065
R29185 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.580578
R29186 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 0.533109
R29187 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.428234
R29188 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.063
R29189 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 0.063
R29190 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 0.063
R29191 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.063
R29192 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 0.063
R29193 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 0.063
R29194 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.t2 169.46
R29195 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.t3 167.809
R29196 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.t0 167.809
R29197 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.t7 167.226
R29198 D_FlipFlop_6.3-input-nand_2.C.t7 D_FlipFlop_6.3-input-nand_2.C.n10 150.273
R29199 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C.t4 150.273
R29200 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C.t5 73.6406
R29201 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C.t6 73.6304
R29202 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.C.t1 60.3943
R29203 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C.n5 12.3891
R29204 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C.n12 11.4489
R29205 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C 1.68257
R29206 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C.n0 1.38365
R29207 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C.n8 1.19615
R29208 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C.n3 1.1717
R29209 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C 1.08448
R29210 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C 0.932141
R29211 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.C.n14 0.720633
R29212 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C.n11 0.280391
R29213 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C 0.217464
R29214 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C 0.1255
R29215 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C 0.1255
R29216 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C 0.1255
R29217 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.n7 0.0874565
R29218 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C.n4 0.063
R29219 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C 0.063
R29220 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C.n6 0.063
R29221 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C.n1 0.063
R29222 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.n13 0.0435206
R29223 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C.n9 0.0216397
R29224 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C 0.0216397
R29225 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C.n2 0.0107679
R29226 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C 0.0107679
R29227 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n7 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t2 179.256
R29228 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n7 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t0 168.089
R29229 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n2 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t3 150.273
R29230 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n1 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t4 74.163
R29231 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n0 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t1 61.1389
R29232 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n5 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n4 12.0358
R29233 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n0 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 1.08746
R29234 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n1 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.851043
R29235 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n8 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n6 0.851043
R29236 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n6 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.65675
R29237 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n3 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n2 0.61463
R29238 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n3 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.486828
R29239 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n8 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n7 0.200143
R29240 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n2 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.063
R29241 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n4 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n1 0.063
R29242 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n4 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n3 0.063
R29243 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n5 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n0 0.063
R29244 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n6 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n5 0.063
R29245 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n8 0.063
R29246 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 169.46
R29247 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 167.809
R29248 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 167.809
R29249 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 167.227
R29250 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 151.594
R29251 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 150.273
R29252 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 74.8641
R29253 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 73.6304
R29254 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 61.84
R29255 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 12.3891
R29256 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 11.4489
R29257 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 0.38637
R29258 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 0.280391
R29259 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 0.200143
R29260 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.152844
R29261 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.149957
R29262 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 0.149957
R29263 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.063
R29264 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.063
R29265 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 0.063
R29266 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 0.063
R29267 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.0454219
R29268 Ring_Counter_0.D_FlipFlop_16.Q.n16 Ring_Counter_0.D_FlipFlop_16.Q.t1 169.46
R29269 Ring_Counter_0.D_FlipFlop_16.Q.n15 Ring_Counter_0.D_FlipFlop_16.Q.t2 167.809
R29270 Ring_Counter_0.D_FlipFlop_16.Q.n16 Ring_Counter_0.D_FlipFlop_16.Q.t0 167.809
R29271 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Q.t9 158.585
R29272 Ring_Counter_0.D_FlipFlop_16.Q.t9 Ring_Counter_0.D_FlipFlop_16.Q.n0 151.594
R29273 Ring_Counter_0.D_FlipFlop_16.Q.n8 Ring_Counter_0.D_FlipFlop_16.Q.t5 150.273
R29274 Ring_Counter_0.D_FlipFlop_16.Q.n4 Ring_Counter_0.D_FlipFlop_16.Q.t6 150.273
R29275 Ring_Counter_0.D_FlipFlop_16.Q.n7 Ring_Counter_0.D_FlipFlop_16.Q.t4 74.163
R29276 Ring_Counter_0.D_FlipFlop_16.Q.n3 Ring_Counter_0.D_FlipFlop_16.Q.t7 74.163
R29277 Ring_Counter_0.D_FlipFlop_16.Q.n12 Ring_Counter_0.D_FlipFlop_16.Q.n11 73.9193
R29278 Ring_Counter_0.D_FlipFlop_16.Q.n0 Ring_Counter_0.D_FlipFlop_16.Q.t8 73.6304
R29279 Ring_Counter_0.D_FlipFlop_16.Q.n18 Ring_Counter_0.D_FlipFlop_16.Q.t3 62.1634
R29280 Ring_Counter_0.D_FlipFlop_16.Q.n17 Ring_Counter_0.D_FlipFlop_16.Q.n16 11.4489
R29281 Ring_Counter_0.D_FlipFlop_16.Q.n15 Ring_Counter_0.D_FlipFlop_16.Q.n14 8.21389
R29282 Ring_Counter_0.D_FlipFlop_16.Q.n11 Ring_Counter_0.D_FlipFlop_16.Q.n6 8.12822
R29283 Ring_Counter_0.D_FlipFlop_16.Q.n11 Ring_Counter_0.D_FlipFlop_16.Q.n10 4.5005
R29284 Ring_Counter_0.D_FlipFlop_16.Q.n7 Ring_Counter_0.D_FlipFlop_16.Q 0.851043
R29285 Ring_Counter_0.D_FlipFlop_16.Q.n3 Ring_Counter_0.D_FlipFlop_16.Q 0.851043
R29286 Ring_Counter_0.D_FlipFlop_16.Q.n9 Ring_Counter_0.D_FlipFlop_16.Q.n8 0.61463
R29287 Ring_Counter_0.D_FlipFlop_16.Q.n5 Ring_Counter_0.D_FlipFlop_16.Q.n4 0.61463
R29288 Ring_Counter_0.D_FlipFlop_16.Q.n9 Ring_Counter_0.D_FlipFlop_16.Q 0.486828
R29289 Ring_Counter_0.D_FlipFlop_16.Q.n5 Ring_Counter_0.D_FlipFlop_16.Q 0.486828
R29290 Ring_Counter_0.D_FlipFlop_16.Q.n14 Ring_Counter_0.D_FlipFlop_16.Q 0.39003
R29291 Ring_Counter_0.D_FlipFlop_16.Q.n17 Ring_Counter_0.D_FlipFlop_16.Q.n15 0.280391
R29292 Ring_Counter_0.D_FlipFlop_16.Q.n14 Ring_Counter_0.D_FlipFlop_16.Q.n13 0.224533
R29293 Ring_Counter_0.D_FlipFlop_16.Q.n13 Ring_Counter_0.D_FlipFlop_16.Q 0.20495
R29294 Ring_Counter_0.D_FlipFlop_16.Q.n18 Ring_Counter_0.D_FlipFlop_16.Q.n17 0.200143
R29295 Ring_Counter_0.D_FlipFlop_16.Q.n2 Ring_Counter_0.D_FlipFlop_16.Q.n1 0.149333
R29296 Ring_Counter_0.D_FlipFlop_16.Q.n2 Ring_Counter_0.D_FlipFlop_16.Q 0.139364
R29297 Ring_Counter_0.D_FlipFlop_16.Q.n8 Ring_Counter_0.D_FlipFlop_16.Q 0.063
R29298 Ring_Counter_0.D_FlipFlop_16.Q.n10 Ring_Counter_0.D_FlipFlop_16.Q.n7 0.063
R29299 Ring_Counter_0.D_FlipFlop_16.Q.n10 Ring_Counter_0.D_FlipFlop_16.Q.n9 0.063
R29300 Ring_Counter_0.D_FlipFlop_16.Q.n4 Ring_Counter_0.D_FlipFlop_16.Q 0.063
R29301 Ring_Counter_0.D_FlipFlop_16.Q.n6 Ring_Counter_0.D_FlipFlop_16.Q.n3 0.063
R29302 Ring_Counter_0.D_FlipFlop_16.Q.n6 Ring_Counter_0.D_FlipFlop_16.Q.n5 0.063
R29303 Ring_Counter_0.D_FlipFlop_16.Q.n0 Ring_Counter_0.D_FlipFlop_16.Q 0.063
R29304 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Q.n18 0.063
R29305 Ring_Counter_0.D_FlipFlop_16.Q.n13 Ring_Counter_0.D_FlipFlop_16.Q.n12 0.024
R29306 Ring_Counter_0.D_FlipFlop_16.Q.n12 Ring_Counter_0.D_FlipFlop_16.Q.n2 0.024
R29307 Ring_Counter_0.D_FlipFlop_16.Q.n1 Ring_Counter_0.D_FlipFlop_16.Q 0.00441667
R29308 Ring_Counter_0.D_FlipFlop_16.Q.n1 Ring_Counter_0.D_FlipFlop_16.Q 0.00406061
R29309 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 169.46
R29310 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 167.809
R29311 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 167.809
R29312 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 167.227
R29313 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 151.594
R29314 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 150.273
R29315 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 74.8641
R29316 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 73.6304
R29317 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 61.84
R29318 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 12.3891
R29319 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 11.4489
R29320 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R29321 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 0.280391
R29322 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 0.200143
R29323 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R29324 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R29325 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 0.149957
R29326 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.063
R29327 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 0.063
R29328 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 0.063
R29329 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 0.063
R29330 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R29331 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t0 169.46
R29332 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t2 167.809
R29333 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t3 167.809
R29334 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t5 167.226
R29335 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n6 150.273
R29336 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t4 150.273
R29337 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t7 74.951
R29338 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t6 73.6304
R29339 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t1 60.3943
R29340 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n4 12.3891
R29341 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n8 11.4489
R29342 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n10 1.68257
R29343 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n0 1.44615
R29344 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n2 1.2342
R29345 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 1.08448
R29346 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.932141
R29347 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n9 0.3496
R29348 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n7 0.280391
R29349 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.063
R29350 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.063
R29351 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n3 0.063
R29352 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.063
R29353 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n5 0.063
R29354 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n1 0.063
R29355 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 179.256
R29356 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 168.089
R29357 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 150.887
R29358 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 73.6304
R29359 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 60.3943
R29360 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 12.0358
R29361 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 1.05069
R29362 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 0.981478
R29363 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.769522
R29364 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 0.745065
R29365 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.580578
R29366 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 0.533109
R29367 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.428234
R29368 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.063
R29369 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 0.063
R29370 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 0.063
R29371 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.063
R29372 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 0.063
R29373 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 0.063
R29374 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t1 169.46
R29375 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t2 167.809
R29376 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t0 167.809
R29377 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t4 167.226
R29378 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n6 150.273
R29379 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t5 150.273
R29380 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t6 74.951
R29381 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t7 73.6304
R29382 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t3 60.3943
R29383 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n4 12.3891
R29384 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n8 11.4489
R29385 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n10 1.68257
R29386 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n0 1.44615
R29387 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n2 1.2342
R29388 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 1.08448
R29389 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.932141
R29390 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n9 0.3496
R29391 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n7 0.280391
R29392 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.063
R29393 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.063
R29394 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n3 0.063
R29395 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.063
R29396 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n5 0.063
R29397 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n1 0.063
R29398 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t0 169.46
R29399 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t1 167.809
R29400 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t3 167.809
R29401 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t6 167.226
R29402 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n6 150.273
R29403 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t7 150.273
R29404 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t5 74.951
R29405 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t4 73.6304
R29406 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t2 60.3943
R29407 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n4 12.3891
R29408 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n8 11.4489
R29409 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n10 1.68257
R29410 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n0 1.44615
R29411 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n2 1.2342
R29412 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 1.08448
R29413 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.932141
R29414 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n9 0.3496
R29415 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n7 0.280391
R29416 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.063
R29417 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.063
R29418 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n3 0.063
R29419 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.063
R29420 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n5 0.063
R29421 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n1 0.063
R29422 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.t3 169.46
R29423 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.t2 167.809
R29424 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t0 167.809
R29425 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t4 167.226
R29426 D_FlipFlop_1.3-input-nand_2.C.t4 D_FlipFlop_1.3-input-nand_2.C.n10 150.273
R29427 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C.t5 150.273
R29428 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C.t6 73.6406
R29429 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C.t7 73.6304
R29430 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.C.t1 60.3943
R29431 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C.n5 12.3891
R29432 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.n12 11.4489
R29433 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C 1.68257
R29434 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C.n0 1.38365
R29435 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C.n8 1.19615
R29436 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C.n3 1.1717
R29437 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C 1.08448
R29438 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C 0.932141
R29439 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.C.n14 0.720633
R29440 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.n11 0.280391
R29441 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C 0.217464
R29442 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C 0.1255
R29443 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C 0.1255
R29444 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C 0.1255
R29445 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.n7 0.0874565
R29446 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C.n4 0.063
R29447 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C 0.063
R29448 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C.n6 0.063
R29449 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C.n1 0.063
R29450 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.n13 0.0435206
R29451 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C.n9 0.0216397
R29452 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C 0.0216397
R29453 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C.n2 0.0107679
R29454 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C 0.0107679
R29455 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.t2 169.46
R29456 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.t3 167.809
R29457 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout.t0 167.809
R29458 D_FlipFlop_1.3-input-nand_2.Vout.t4 D_FlipFlop_1.3-input-nand_2.Vout.n11 167.227
R29459 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.t4 150.293
R29460 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.t7 150.273
R29461 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout.t6 73.6406
R29462 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout.t5 73.6304
R29463 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout.t1 60.3809
R29464 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout.n5 12.3891
R29465 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout.n9 11.4489
R29466 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout.n2 1.38365
R29467 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.n1 1.19615
R29468 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.n4 1.1717
R29469 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout 0.848156
R29470 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.Vout.n12 0.447191
R29471 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R29472 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout.n10 0.280391
R29473 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout 0.217464
R29474 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout 0.200143
R29475 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R29476 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R29477 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R29478 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R29479 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout.n7 0.0874565
R29480 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout.n3 0.063
R29481 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout.n6 0.063
R29482 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.Vout.n8 0.063
R29483 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R29484 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout.n0 0.0107679
R29485 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout 0.0107679
R29486 Q2.n8 Q2.t2 169.46
R29487 Q2.n10 Q2.t0 167.809
R29488 Q2.n8 Q2.t3 167.809
R29489 Q2.n16 Q2.t6 158.565
R29490 Q2.n2 Q2.t8 150.543
R29491 Q2.n0 Q2.t7 150.543
R29492 Q2.t6 Q2.n15 150.293
R29493 Q2.n2 Q2.t4 74.4613
R29494 Q2.n0 Q2.t5 74.4613
R29495 Q2.n13 Q2.t9 73.6304
R29496 Q2.n6 Q2.t1 60.3809
R29497 Q2.n5 Q2.n4 12.2652
R29498 Q2.n9 Q2.n8 11.4489
R29499 Q2.n11 Q2.n10 8.21389
R29500 Q2 Q2.n16 5.21615
R29501 Q2.n17 Q2.n5 2.63093
R29502 Q2.n5 Q2 2.39252
R29503 Q2.n7 Q2.n6 1.64452
R29504 Q2.n15 Q2.n14 1.19615
R29505 Q2.n1 Q2 0.984196
R29506 Q2.n6 Q2 0.848156
R29507 Q2.n3 Q2.n2 0.747783
R29508 Q2.n1 Q2.n0 0.747783
R29509 Q2.n3 Q2 0.582531
R29510 Q2.n15 Q2 0.447191
R29511 Q2.n12 Q2.n11 0.425067
R29512 Q2.n11 Q2 0.39003
R29513 Q2.n10 Q2.n9 0.280391
R29514 Q2.n9 Q2 0.200143
R29515 Q2.n14 Q2 0.1255
R29516 Q2.n7 Q2 0.1255
R29517 Q2 Q2.n7 0.063
R29518 Q2.n2 Q2 0.063
R29519 Q2.n4 Q2.n1 0.063
R29520 Q2.n4 Q2.n3 0.063
R29521 Q2.n16 Q2 0.0204394
R29522 Q2.n14 Q2.n13 0.0107679
R29523 Q2.n13 Q2 0.0107679
R29524 Q2.n12 Q2 0.00441667
R29525 Q2 Q2.n12 0.00406061
R29526 Q2.n17 Q2 0.00128333
R29527 Q2.n17 Q2 0.00121212
R29528 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t4 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t2 316.762
R29529 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t0 169.195
R29530 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t4 150.887
R29531 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n2 150.273
R29532 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t5 74.951
R29533 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t3 73.6304
R29534 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t1 60.3943
R29535 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n6 12.0358
R29536 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n8 0.981478
R29537 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.769522
R29538 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n0 0.745065
R29539 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.580578
R29540 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n4 0.533109
R29541 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.428234
R29542 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.063
R29543 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.063
R29544 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n3 0.063
R29545 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n5 0.063
R29546 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.063
R29547 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n7 0.063
R29548 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n1 0.063
R29549 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t0 169.46
R29550 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t1 167.809
R29551 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t2 167.809
R29552 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t6 167.226
R29553 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n6 150.273
R29554 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t5 150.273
R29555 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t7 74.951
R29556 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t4 73.6304
R29557 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t3 60.3943
R29558 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n4 12.3891
R29559 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n8 11.4489
R29560 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n10 1.68257
R29561 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n0 1.44615
R29562 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n2 1.2342
R29563 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 1.08448
R29564 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.932141
R29565 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n9 0.3496
R29566 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n7 0.280391
R29567 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.063
R29568 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.063
R29569 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n3 0.063
R29570 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.063
R29571 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n5 0.063
R29572 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n1 0.063
R29573 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 169.46
R29574 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 168.089
R29575 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 167.809
R29576 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 150.887
R29577 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 73.6304
R29578 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 60.3943
R29579 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 12.0358
R29580 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 11.4489
R29581 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 1.05069
R29582 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 0.981478
R29583 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.769522
R29584 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 0.745065
R29585 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.580578
R29586 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 0.533109
R29587 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.428234
R29588 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.063
R29589 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 0.063
R29590 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 0.063
R29591 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.063
R29592 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 0.063
R29593 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 0.063
R29594 Q3.n2 Q3.t2 169.46
R29595 Q3.n4 Q3.t0 167.809
R29596 Q3.n2 Q3.t3 167.809
R29597 Q3.n10 Q3.t9 158.565
R29598 Q3.n14 Q3.t7 150.543
R29599 Q3.n12 Q3.t8 150.543
R29600 Q3.t9 Q3.n9 150.293
R29601 Q3.n14 Q3.t6 74.4613
R29602 Q3.n12 Q3.t4 74.4613
R29603 Q3.n7 Q3.t5 73.6304
R29604 Q3.n0 Q3.t1 60.3809
R29605 Q3 Q3.n16 12.3648
R29606 Q3.n3 Q3.n2 11.4489
R29607 Q3.n5 Q3.n4 8.21389
R29608 Q3.n11 Q3.n10 5.1166
R29609 Q3.n1 Q3.n0 1.64452
R29610 Q3.n9 Q3.n8 1.19615
R29611 Q3.n17 Q3.n11 1.04077
R29612 Q3.n13 Q3 0.984196
R29613 Q3.n11 Q3 0.946909
R29614 Q3.n0 Q3 0.848156
R29615 Q3.n15 Q3.n14 0.747783
R29616 Q3.n13 Q3.n12 0.747783
R29617 Q3.n15 Q3 0.582531
R29618 Q3.n9 Q3 0.447191
R29619 Q3.n6 Q3.n5 0.425067
R29620 Q3.n5 Q3 0.39003
R29621 Q3.n4 Q3.n3 0.280391
R29622 Q3.n3 Q3 0.200143
R29623 Q3.n8 Q3 0.1255
R29624 Q3.n1 Q3 0.1255
R29625 Q3.n14 Q3 0.063
R29626 Q3.n16 Q3.n13 0.063
R29627 Q3.n16 Q3.n15 0.063
R29628 Q3 Q3.n1 0.063
R29629 Q3.n10 Q3 0.0204394
R29630 Q3.n8 Q3.n7 0.0107679
R29631 Q3.n7 Q3 0.0107679
R29632 Q3.n6 Q3 0.00441667
R29633 Q3 Q3.n6 0.00406061
R29634 Q3.n17 Q3 0.00128333
R29635 Q3.n17 Q3 0.00121212
R29636 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t2 316.762
R29637 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t0 169.195
R29638 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t3 150.887
R29639 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n2 150.273
R29640 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t4 74.951
R29641 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t5 73.6304
R29642 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t1 60.3943
R29643 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n6 12.0358
R29644 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n8 0.981478
R29645 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.769522
R29646 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n0 0.745065
R29647 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.580578
R29648 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n4 0.533109
R29649 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.428234
R29650 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.063
R29651 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.063
R29652 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n3 0.063
R29653 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n5 0.063
R29654 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.063
R29655 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n7 0.063
R29656 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n1 0.063
R29657 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t1 169.46
R29658 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.t2 167.809
R29659 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t0 167.809
R29660 D_FlipFlop_3.3-input-nand_2.Vout.t4 D_FlipFlop_3.3-input-nand_2.Vout.n11 167.227
R29661 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.t4 150.293
R29662 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.t6 150.273
R29663 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout.t7 73.6406
R29664 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout.t5 73.6304
R29665 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout.t3 60.3809
R29666 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n5 12.3891
R29667 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout.n9 11.4489
R29668 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout.n2 1.38365
R29669 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.n1 1.19615
R29670 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.n4 1.1717
R29671 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout 0.848156
R29672 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.Vout.n12 0.447191
R29673 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R29674 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.n10 0.280391
R29675 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout 0.217464
R29676 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout 0.200143
R29677 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R29678 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R29679 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R29680 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R29681 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout.n7 0.0874565
R29682 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n3 0.063
R29683 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout.n6 0.063
R29684 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.Vout.n8 0.063
R29685 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R29686 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout.n0 0.0107679
R29687 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout 0.0107679
R29688 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 169.46
R29689 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 167.809
R29690 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 167.809
R29691 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 167.227
R29692 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 151.594
R29693 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 150.273
R29694 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 74.8641
R29695 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 73.6304
R29696 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 61.84
R29697 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 12.3891
R29698 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 11.4489
R29699 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.38637
R29700 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 0.280391
R29701 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 0.200143
R29702 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.152844
R29703 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.149957
R29704 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 0.149957
R29705 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.063
R29706 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 0.063
R29707 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 0.063
R29708 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 0.063
R29709 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.0454219
R29710 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 169.46
R29711 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 168.089
R29712 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 167.809
R29713 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 150.887
R29714 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 73.6304
R29715 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 60.3943
R29716 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 12.0358
R29717 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 11.4489
R29718 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 1.05069
R29719 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 0.981478
R29720 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.769522
R29721 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 0.745065
R29722 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.580578
R29723 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 0.533109
R29724 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.428234
R29725 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.063
R29726 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 0.063
R29727 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 0.063
R29728 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.063
R29729 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 0.063
R29730 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 0.063
R29731 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t1 169.46
R29732 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.t2 167.809
R29733 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t0 167.809
R29734 D_FlipFlop_3.3-input-nand_2.C.t4 D_FlipFlop_3.3-input-nand_2.C.n13 167.226
R29735 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.t5 150.273
R29736 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.t4 150.273
R29737 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C.t7 73.6406
R29738 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C.t6 73.6304
R29739 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.C.t3 60.3943
R29740 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n7 12.3891
R29741 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n11 11.4489
R29742 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C 1.68257
R29743 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C.n2 1.38365
R29744 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C.n0 1.19615
R29745 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C.n5 1.1717
R29746 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C 1.08448
R29747 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C 0.932141
R29748 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C 0.720633
R29749 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.n12 0.280391
R29750 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C 0.217464
R29751 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29752 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29753 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C 0.1255
R29754 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C.n9 0.0874565
R29755 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.n6 0.063
R29756 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.063
R29757 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C.n8 0.063
R29758 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n3 0.063
R29759 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n10 0.0435206
R29760 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.n1 0.0216397
R29761 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.C.n14 0.0216397
R29762 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C.n4 0.0107679
R29763 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C 0.0107679
R29764 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout.t1 169.46
R29765 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout.t3 167.809
R29766 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout.t2 167.809
R29767 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout.t5 167.227
R29768 D_FlipFlop_5.3-input-nand_2.Vout.t5 D_FlipFlop_5.3-input-nand_2.Vout.n2 150.293
R29769 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.t7 150.273
R29770 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout.t4 73.6406
R29771 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout.t6 73.6304
R29772 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.t0 60.3809
R29773 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n9 12.3891
R29774 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.n4 11.4489
R29775 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.n11 1.38365
R29776 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout.n1 1.19615
R29777 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.n8 1.1717
R29778 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.Vout.n12 0.848156
R29779 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout 0.447191
R29780 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R29781 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.n3 0.280391
R29782 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout 0.217464
R29783 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.Vout.n5 0.200143
R29784 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R29785 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R29786 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R29787 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R29788 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout.n6 0.0874565
R29789 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout 0.063
R29790 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout.n10 0.063
R29791 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n7 0.063
R29792 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R29793 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout.n0 0.0107679
R29794 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout 0.0107679
R29795 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t3 316.762
R29796 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t0 169.195
R29797 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t2 150.887
R29798 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n2 150.273
R29799 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t5 74.951
R29800 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t4 73.6304
R29801 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t1 60.3943
R29802 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n6 12.0358
R29803 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n8 0.981478
R29804 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.769522
R29805 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n0 0.745065
R29806 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.580578
R29807 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n4 0.533109
R29808 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.428234
R29809 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.063
R29810 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.063
R29811 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n3 0.063
R29812 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n5 0.063
R29813 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.063
R29814 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n7 0.063
R29815 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n1 0.063
R29816 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t0 169.46
R29817 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n8 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t1 167.809
R29818 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t2 167.809
R29819 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n7 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t5 167.226
R29820 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n6 150.273
R29821 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t6 150.273
R29822 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t7 74.951
R29823 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t4 73.6304
R29824 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t3 60.3943
R29825 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n4 12.3891
R29826 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n8 11.4489
R29827 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n10 1.68257
R29828 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n0 1.44615
R29829 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n2 1.2342
R29830 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n1 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 1.08448
R29831 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n3 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.932141
R29832 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n9 0.3496
R29833 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n9 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n7 0.280391
R29834 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n6 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.063
R29835 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n2 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.063
R29836 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n4 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n3 0.063
R29837 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n0 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.063
R29838 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n10 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n5 0.063
R29839 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n5 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n1 0.063
R29840 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 179.256
R29841 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 168.089
R29842 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 150.887
R29843 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 73.6304
R29844 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 60.3943
R29845 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 12.0358
R29846 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 1.05069
R29847 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 0.981478
R29848 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.769522
R29849 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 0.745065
R29850 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.580578
R29851 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 0.533109
R29852 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.428234
R29853 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.063
R29854 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 0.063
R29855 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 0.063
R29856 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.063
R29857 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 0.063
R29858 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 0.063
R29859 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 179.256
R29860 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 168.089
R29861 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 150.887
R29862 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 73.6304
R29863 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 60.3943
R29864 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 12.0358
R29865 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 1.05069
R29866 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 0.981478
R29867 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.769522
R29868 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 0.745065
R29869 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.580578
R29870 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 0.533109
R29871 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.428234
R29872 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.063
R29873 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 0.063
R29874 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 0.063
R29875 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.063
R29876 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 0.063
R29877 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 0.063
R29878 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t2 316.762
R29879 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t0 169.195
R29880 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t3 150.887
R29881 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n2 150.273
R29882 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t4 74.951
R29883 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t5 73.6304
R29884 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t1 60.3943
R29885 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n6 12.0358
R29886 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n8 0.981478
R29887 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.769522
R29888 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n0 0.745065
R29889 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.580578
R29890 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n4 0.533109
R29891 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.428234
R29892 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.063
R29893 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.063
R29894 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n3 0.063
R29895 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n5 0.063
R29896 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.063
R29897 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n7 0.063
R29898 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n1 0.063
R29899 Ring_Counter_0.D_FlipFlop_4.Qbar.n4 Ring_Counter_0.D_FlipFlop_4.Qbar.t2 169.46
R29900 Ring_Counter_0.D_FlipFlop_4.Qbar.n4 Ring_Counter_0.D_FlipFlop_4.Qbar.t3 167.809
R29901 Ring_Counter_0.D_FlipFlop_4.Qbar.n6 Ring_Counter_0.D_FlipFlop_4.Qbar.t0 167.809
R29902 Ring_Counter_0.D_FlipFlop_4.Qbar.n1 Ring_Counter_0.D_FlipFlop_4.Qbar.t4 158.28
R29903 Ring_Counter_0.D_FlipFlop_4.Qbar.t4 Ring_Counter_0.D_FlipFlop_4.Qbar.n0 150.273
R29904 Ring_Counter_0.D_FlipFlop_4.Qbar.n0 Ring_Counter_0.D_FlipFlop_4.Qbar.t5 74.951
R29905 Ring_Counter_0.D_FlipFlop_4.Qbar.n3 Ring_Counter_0.D_FlipFlop_4.Qbar.t1 60.3943
R29906 Ring_Counter_0.D_FlipFlop_4.Qbar.n5 Ring_Counter_0.D_FlipFlop_4.Qbar.n4 11.4489
R29907 Ring_Counter_0.D_FlipFlop_4.Qbar Ring_Counter_0.D_FlipFlop_4.Qbar.n6 8.5174
R29908 Ring_Counter_0.D_FlipFlop_4.Qbar.n5 Ring_Counter_0.D_FlipFlop_4.Qbar.n3 1.96917
R29909 Ring_Counter_0.D_FlipFlop_4.Qbar.n2 Ring_Counter_0.D_FlipFlop_4.Qbar.n1 0.42585
R29910 Ring_Counter_0.D_FlipFlop_4.Qbar.n1 Ring_Counter_0.D_FlipFlop_4.Qbar 0.390742
R29911 Ring_Counter_0.D_FlipFlop_4.Qbar.n6 Ring_Counter_0.D_FlipFlop_4.Qbar.n5 0.280391
R29912 Ring_Counter_0.D_FlipFlop_4.Qbar.n3 Ring_Counter_0.D_FlipFlop_4.Qbar 0.063
R29913 Ring_Counter_0.D_FlipFlop_4.Qbar.n0 Ring_Counter_0.D_FlipFlop_4.Qbar 0.063
R29914 Ring_Counter_0.D_FlipFlop_4.Qbar.n2 Ring_Counter_0.D_FlipFlop_4.Qbar 0.00441667
R29915 Ring_Counter_0.D_FlipFlop_4.Qbar Ring_Counter_0.D_FlipFlop_4.Qbar.n2 0.00406061
R29916 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t3 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t5 316.762
R29917 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t0 169.195
R29918 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t3 150.887
R29919 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n2 150.273
R29920 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t4 74.951
R29921 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t2 73.6304
R29922 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t1 60.3943
R29923 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n6 12.0358
R29924 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n8 0.981478
R29925 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.769522
R29926 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n0 0.745065
R29927 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.580578
R29928 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n4 0.533109
R29929 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.428234
R29930 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.063
R29931 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.063
R29932 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n3 0.063
R29933 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n5 0.063
R29934 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.063
R29935 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n7 0.063
R29936 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n1 0.063
R29937 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 179.256
R29938 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 168.089
R29939 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 150.887
R29940 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 73.6304
R29941 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 60.3943
R29942 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 12.0358
R29943 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 1.05069
R29944 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 0.981478
R29945 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.769522
R29946 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 0.745065
R29947 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.580578
R29948 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 0.533109
R29949 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.428234
R29950 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.063
R29951 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 0.063
R29952 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 0.063
R29953 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.063
R29954 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 0.063
R29955 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 0.063
R29956 Nand_Gate_5.A.n12 Nand_Gate_5.A.t7 171.107
R29957 Nand_Gate_5.A.n19 Nand_Gate_5.A.t3 169.46
R29958 Nand_Gate_5.A.n18 Nand_Gate_5.A.t1 167.809
R29959 Nand_Gate_5.A.n19 Nand_Gate_5.A.t0 167.809
R29960 Nand_Gate_5.A.n15 Nand_Gate_5.A.t8 158.565
R29961 Nand_Gate_5.A.t8 Nand_Gate_5.A.n14 151.594
R29962 Nand_Gate_5.A.t7 Nand_Gate_5.A.n2 150.293
R29963 Nand_Gate_5.A.n6 Nand_Gate_5.A.t4 150.273
R29964 Nand_Gate_5.A.n3 Nand_Gate_5.A.t11 150.273
R29965 Nand_Gate_5.A Nand_Gate_5.A.t9 99.8701
R29966 Nand_Gate_5.A.n5 Nand_Gate_5.A.t6 74.163
R29967 Nand_Gate_5.A.t9 Nand_Gate_5.A.n10 74.163
R29968 Nand_Gate_5.A.n14 Nand_Gate_5.A.t5 73.6304
R29969 Nand_Gate_5.A.n0 Nand_Gate_5.A.t10 73.6304
R29970 Nand_Gate_5.A.n21 Nand_Gate_5.A.t2 62.1634
R29971 Nand_Gate_5.A.n9 Nand_Gate_5.A.n8 12.6418
R29972 Nand_Gate_5.A.n20 Nand_Gate_5.A.n19 11.4489
R29973 Nand_Gate_5.A.n18 Nand_Gate_5.A.n17 8.21389
R29974 Nand_Gate_5.A.n13 Nand_Gate_5.A 1.2047
R29975 Nand_Gate_5.A.n2 Nand_Gate_5.A.n1 1.19615
R29976 Nand_Gate_5.A.n12 Nand_Gate_5.A.n11 0.922483
R29977 Nand_Gate_5.A.n5 Nand_Gate_5.A 0.851043
R29978 Nand_Gate_5.A.n10 Nand_Gate_5.A 0.851043
R29979 Nand_Gate_5.A.n7 Nand_Gate_5.A.n6 0.61463
R29980 Nand_Gate_5.A.n4 Nand_Gate_5.A.n3 0.61463
R29981 Nand_Gate_5.A.n7 Nand_Gate_5.A 0.486828
R29982 Nand_Gate_5.A.n4 Nand_Gate_5.A 0.486828
R29983 Nand_Gate_5.A.n2 Nand_Gate_5.A 0.447191
R29984 Nand_Gate_5.A.n17 Nand_Gate_5.A.n16 0.425067
R29985 Nand_Gate_5.A.n13 Nand_Gate_5.A.n12 0.399217
R29986 Nand_Gate_5.A.n17 Nand_Gate_5.A 0.39003
R29987 Nand_Gate_5.A.n20 Nand_Gate_5.A.n18 0.280391
R29988 Nand_Gate_5.A.n21 Nand_Gate_5.A.n20 0.200143
R29989 Nand_Gate_5.A.n1 Nand_Gate_5.A 0.1255
R29990 Nand_Gate_5.A.n14 Nand_Gate_5.A 0.063
R29991 Nand_Gate_5.A.n6 Nand_Gate_5.A 0.063
R29992 Nand_Gate_5.A.n8 Nand_Gate_5.A.n5 0.063
R29993 Nand_Gate_5.A.n8 Nand_Gate_5.A.n7 0.063
R29994 Nand_Gate_5.A.n3 Nand_Gate_5.A 0.063
R29995 Nand_Gate_5.A.n10 Nand_Gate_5.A.n9 0.063
R29996 Nand_Gate_5.A.n9 Nand_Gate_5.A.n4 0.063
R29997 Nand_Gate_5.A Nand_Gate_5.A.n21 0.063
R29998 Nand_Gate_5.A.n15 Nand_Gate_5.A.n13 0.024
R29999 Nand_Gate_5.A Nand_Gate_5.A.n15 0.0204394
R30000 Nand_Gate_5.A.n1 Nand_Gate_5.A.n0 0.0107679
R30001 Nand_Gate_5.A.n0 Nand_Gate_5.A 0.0107679
R30002 Nand_Gate_5.A.n11 Nand_Gate_5.A 0.00441667
R30003 Nand_Gate_5.A.n16 Nand_Gate_5.A 0.00441667
R30004 Nand_Gate_5.A.n11 Nand_Gate_5.A 0.00406061
R30005 Nand_Gate_5.A.n16 Nand_Gate_5.A 0.00406061
R30006 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 169.46
R30007 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 168.089
R30008 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 167.809
R30009 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 150.887
R30010 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 73.6304
R30011 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 60.3943
R30012 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 12.0358
R30013 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 11.4489
R30014 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 1.05069
R30015 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 0.981478
R30016 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.769522
R30017 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 0.745065
R30018 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.580578
R30019 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 0.533109
R30020 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.428234
R30021 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.063
R30022 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 0.063
R30023 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 0.063
R30024 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.063
R30025 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 0.063
R30026 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 0.063
R30027 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 169.46
R30028 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 168.089
R30029 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 167.809
R30030 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 150.887
R30031 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 73.6304
R30032 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 60.3943
R30033 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 12.0358
R30034 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 11.4489
R30035 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 1.05069
R30036 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 0.981478
R30037 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.769522
R30038 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 0.745065
R30039 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.580578
R30040 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 0.533109
R30041 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.428234
R30042 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.063
R30043 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 0.063
R30044 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 0.063
R30045 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.063
R30046 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 0.063
R30047 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 0.063
R30048 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t1 169.46
R30049 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.t2 167.809
R30050 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t0 167.809
R30051 D_FlipFlop_7.3-input-nand_2.Vout.t5 D_FlipFlop_7.3-input-nand_2.Vout.n11 167.227
R30052 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.t5 150.293
R30053 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.t6 150.273
R30054 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout.t4 73.6406
R30055 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout.t7 73.6304
R30056 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout.t3 60.3809
R30057 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n5 12.3891
R30058 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout.n9 11.4489
R30059 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout.n2 1.38365
R30060 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.n1 1.19615
R30061 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.n4 1.1717
R30062 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout 0.848156
R30063 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.Vout.n12 0.447191
R30064 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R30065 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.n10 0.280391
R30066 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout 0.217464
R30067 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout 0.200143
R30068 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R30069 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R30070 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R30071 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R30072 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout.n7 0.0874565
R30073 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n3 0.063
R30074 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout.n6 0.063
R30075 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.Vout.n8 0.063
R30076 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R30077 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout.n0 0.0107679
R30078 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout 0.0107679
R30079 Q4.n2 Q4.t0 169.46
R30080 Q4.n4 Q4.t2 167.809
R30081 Q4.n2 Q4.t1 167.809
R30082 Q4.n10 Q4.t6 158.565
R30083 Q4.n14 Q4.t7 150.543
R30084 Q4.n12 Q4.t8 150.543
R30085 Q4.t6 Q4.n9 150.293
R30086 Q4.n14 Q4.t4 74.4613
R30087 Q4.n12 Q4.t5 74.4613
R30088 Q4.n7 Q4.t9 73.6304
R30089 Q4.n0 Q4.t3 60.3809
R30090 Q4 Q4.n16 12.465
R30091 Q4.n3 Q4.n2 11.4489
R30092 Q4.n5 Q4.n4 8.21389
R30093 Q4.n11 Q4.n10 5.01633
R30094 Q4.n17 Q4.n11 4.81487
R30095 Q4.n11 Q4 4.37791
R30096 Q4.n1 Q4.n0 1.64452
R30097 Q4.n9 Q4.n8 1.19615
R30098 Q4.n13 Q4 0.984196
R30099 Q4.n0 Q4 0.848156
R30100 Q4.n15 Q4.n14 0.747783
R30101 Q4.n13 Q4.n12 0.747783
R30102 Q4.n15 Q4 0.582531
R30103 Q4.n9 Q4 0.447191
R30104 Q4.n6 Q4.n5 0.425067
R30105 Q4.n5 Q4 0.39003
R30106 Q4.n4 Q4.n3 0.280391
R30107 Q4.n3 Q4 0.200143
R30108 Q4.n8 Q4 0.1255
R30109 Q4.n1 Q4 0.1255
R30110 Q4.n14 Q4 0.063
R30111 Q4.n16 Q4.n13 0.063
R30112 Q4.n16 Q4.n15 0.063
R30113 Q4 Q4.n1 0.063
R30114 Q4.n10 Q4 0.0204394
R30115 Q4.n8 Q4.n7 0.0107679
R30116 Q4.n7 Q4 0.0107679
R30117 Q4.n6 Q4 0.00441667
R30118 Q4 Q4.n6 0.00406061
R30119 Q4.n17 Q4 0.00128333
R30120 Q4.n17 Q4 0.00121212
R30121 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 179.256
R30122 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 168.089
R30123 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 150.887
R30124 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 73.6304
R30125 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 60.3943
R30126 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 12.0358
R30127 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 1.05069
R30128 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 0.981478
R30129 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.769522
R30130 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 0.745065
R30131 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.580578
R30132 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 0.533109
R30133 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.428234
R30134 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.063
R30135 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 0.063
R30136 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 0.063
R30137 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.063
R30138 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 0.063
R30139 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 0.063
R30140 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.t3 169.46
R30141 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.t2 167.809
R30142 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t0 167.809
R30143 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t4 167.226
R30144 D_FlipFlop_7.3-input-nand_2.C.t4 D_FlipFlop_7.3-input-nand_2.C.n10 150.273
R30145 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C.t6 150.273
R30146 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C.t5 73.6406
R30147 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C.t7 73.6304
R30148 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.C.t1 60.3943
R30149 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C.n5 12.3891
R30150 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.n12 11.4489
R30151 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C 1.68257
R30152 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C.n0 1.38365
R30153 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C.n8 1.19615
R30154 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C.n3 1.1717
R30155 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C 1.08448
R30156 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C 0.932141
R30157 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.C.n14 0.720633
R30158 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.n11 0.280391
R30159 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C 0.217464
R30160 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30161 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30162 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C 0.1255
R30163 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.n7 0.0874565
R30164 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C.n4 0.063
R30165 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C 0.063
R30166 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C.n6 0.063
R30167 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C.n1 0.063
R30168 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.n13 0.0435206
R30169 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C.n9 0.0216397
R30170 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C 0.0216397
R30171 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C.n2 0.0107679
R30172 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C 0.0107679
R30173 CDAC_v3_0.switch_4.Z.n0 CDAC_v3_0.switch_4.Z.t2 168.075
R30174 CDAC_v3_0.switch_4.Z.n0 CDAC_v3_0.switch_4.Z.t1 168.075
R30175 CDAC_v3_0.switch_4.Z.n20 CDAC_v3_0.switch_4.Z.t0 60.6851
R30176 CDAC_v3_0.switch_4.Z CDAC_v3_0.switch_4.Z.t3 60.6226
R30177 CDAC_v3_0.switch_4.Z.n18 CDAC_v3_0.switch_4.Z.n17 44.8135
R30178 CDAC_v3_0.switch_4.Z.n9 CDAC_v3_0.switch_4.Z.n5 12.0366
R30179 CDAC_v3_0.switch_4.Z.n9 CDAC_v3_0.switch_4.Z.n8 10.5514
R30180 CDAC_v3_0.switch_4.Z.n17 CDAC_v3_0.switch_4.Z.n16 8.6463
R30181 CDAC_v3_0.switch_4.Z.n13 CDAC_v3_0.switch_4.Z.n12 8.08543
R30182 CDAC_v3_0.switch_4.Z.n14 CDAC_v3_0.switch_4.Z.t17 7.92783
R30183 CDAC_v3_0.switch_4.Z.n10 CDAC_v3_0.switch_4.Z.t9 7.92783
R30184 CDAC_v3_0.switch_4.Z.n6 CDAC_v3_0.switch_4.Z.t12 7.92783
R30185 CDAC_v3_0.switch_4.Z.n3 CDAC_v3_0.switch_4.Z.t10 7.92783
R30186 CDAC_v3_0.switch_4.Z.n15 CDAC_v3_0.switch_4.Z.n14 7.62077
R30187 CDAC_v3_0.switch_4.Z.n16 CDAC_v3_0.switch_4.Z.n15 7.62077
R30188 CDAC_v3_0.switch_4.Z.n11 CDAC_v3_0.switch_4.Z.n10 7.62077
R30189 CDAC_v3_0.switch_4.Z.n12 CDAC_v3_0.switch_4.Z.n11 7.62077
R30190 CDAC_v3_0.switch_4.Z.n7 CDAC_v3_0.switch_4.Z.n6 7.62077
R30191 CDAC_v3_0.switch_4.Z.n8 CDAC_v3_0.switch_4.Z.n7 7.62077
R30192 CDAC_v3_0.switch_4.Z.n4 CDAC_v3_0.switch_4.Z.n3 7.62077
R30193 CDAC_v3_0.switch_4.Z.n5 CDAC_v3_0.switch_4.Z.n4 7.62077
R30194 CDAC_v3_0.switch_4.Z.n13 CDAC_v3_0.switch_4.Z.n9 3.80593
R30195 CDAC_v3_0.switch_4.Z.n17 CDAC_v3_0.switch_4.Z.n13 2.04657
R30196 CDAC_v3_0.switch_4.Z.n2 CDAC_v3_0.switch_4.Z.n1 1.34289
R30197 CDAC_v3_0.switch_4.Z.n2 CDAC_v3_0.switch_4.Z 0.42713
R30198 CDAC_v3_0.switch_4.Z.n14 CDAC_v3_0.switch_4.Z.t15 0.307567
R30199 CDAC_v3_0.switch_4.Z.n15 CDAC_v3_0.switch_4.Z.t11 0.307567
R30200 CDAC_v3_0.switch_4.Z.n16 CDAC_v3_0.switch_4.Z.t13 0.307567
R30201 CDAC_v3_0.switch_4.Z.n12 CDAC_v3_0.switch_4.Z.t5 0.307567
R30202 CDAC_v3_0.switch_4.Z.n11 CDAC_v3_0.switch_4.Z.t4 0.307567
R30203 CDAC_v3_0.switch_4.Z.n10 CDAC_v3_0.switch_4.Z.t6 0.307567
R30204 CDAC_v3_0.switch_4.Z.n6 CDAC_v3_0.switch_4.Z.t8 0.307567
R30205 CDAC_v3_0.switch_4.Z.n7 CDAC_v3_0.switch_4.Z.t19 0.307567
R30206 CDAC_v3_0.switch_4.Z.n8 CDAC_v3_0.switch_4.Z.t16 0.307567
R30207 CDAC_v3_0.switch_4.Z.n5 CDAC_v3_0.switch_4.Z.t14 0.307567
R30208 CDAC_v3_0.switch_4.Z.n4 CDAC_v3_0.switch_4.Z.t18 0.307567
R30209 CDAC_v3_0.switch_4.Z.n3 CDAC_v3_0.switch_4.Z.t7 0.307567
R30210 CDAC_v3_0.switch_4.Z.n19 CDAC_v3_0.switch_4.Z 0.182141
R30211 CDAC_v3_0.switch_4.Z.n1 CDAC_v3_0.switch_4.Z 0.178175
R30212 CDAC_v3_0.switch_4.Z.n20 CDAC_v3_0.switch_4.Z.n19 0.128217
R30213 CDAC_v3_0.switch_4.Z.n20 CDAC_v3_0.switch_4.Z 0.1255
R30214 CDAC_v3_0.switch_4.Z.n18 CDAC_v3_0.switch_4.Z.n2 0.063
R30215 CDAC_v3_0.switch_4.Z.n19 CDAC_v3_0.switch_4.Z.n18 0.063
R30216 CDAC_v3_0.switch_4.Z CDAC_v3_0.switch_4.Z.n20 0.063
R30217 CDAC_v3_0.switch_4.Z.n1 CDAC_v3_0.switch_4.Z.n0 0.0130546
R30218 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 169.46
R30219 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 168.089
R30220 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 167.809
R30221 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 150.887
R30222 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 73.6304
R30223 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 60.3943
R30224 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 12.0358
R30225 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 11.4489
R30226 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 1.05069
R30227 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 0.981478
R30228 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.769522
R30229 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 0.745065
R30230 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.580578
R30231 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 0.533109
R30232 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.428234
R30233 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.063
R30234 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 0.063
R30235 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 0.063
R30236 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.063
R30237 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 0.063
R30238 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 0.063
R30239 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 169.46
R30240 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 168.089
R30241 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 167.809
R30242 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 150.887
R30243 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 73.6304
R30244 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 60.3943
R30245 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 12.0358
R30246 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 11.4489
R30247 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 1.05069
R30248 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 0.981478
R30249 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.769522
R30250 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 0.745065
R30251 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.580578
R30252 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 0.533109
R30253 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.428234
R30254 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.063
R30255 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 0.063
R30256 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 0.063
R30257 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.063
R30258 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 0.063
R30259 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 0.063
R30260 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 169.46
R30261 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 168.089
R30262 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 167.809
R30263 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 150.887
R30264 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 73.6304
R30265 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 60.3943
R30266 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 12.0358
R30267 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 11.4489
R30268 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 1.05069
R30269 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 0.981478
R30270 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.769522
R30271 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 0.745065
R30272 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.580578
R30273 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 0.533109
R30274 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.428234
R30275 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.063
R30276 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 0.063
R30277 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 0.063
R30278 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.063
R30279 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 0.063
R30280 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 0.063
R30281 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 169.46
R30282 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 168.089
R30283 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 167.809
R30284 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 150.887
R30285 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 73.6304
R30286 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 60.3943
R30287 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 12.0358
R30288 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 11.4489
R30289 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 1.05069
R30290 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 0.981478
R30291 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.769522
R30292 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 0.745065
R30293 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.580578
R30294 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 0.533109
R30295 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.428234
R30296 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.063
R30297 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 0.063
R30298 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 0.063
R30299 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.063
R30300 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 0.063
R30301 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 0.063
R30302 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 169.46
R30303 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 168.089
R30304 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 167.809
R30305 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 150.887
R30306 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 73.6304
R30307 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 60.3943
R30308 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 12.0358
R30309 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 11.4489
R30310 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 1.05069
R30311 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 0.981478
R30312 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.769522
R30313 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 0.745065
R30314 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.580578
R30315 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 0.533109
R30316 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.428234
R30317 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.063
R30318 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 0.063
R30319 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 0.063
R30320 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.063
R30321 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 0.063
R30322 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 0.063
R30323 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t2 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t5 316.762
R30324 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t0 169.195
R30325 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t2 150.887
R30326 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t5 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n2 150.273
R30327 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t3 74.951
R30328 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t4 73.6304
R30329 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t1 60.3943
R30330 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n6 12.0358
R30331 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n8 0.981478
R30332 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n3 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.769522
R30333 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n0 0.745065
R30334 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n1 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.580578
R30335 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n4 0.533109
R30336 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n5 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.428234
R30337 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n4 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.063
R30338 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n2 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.063
R30339 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n3 0.063
R30340 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n6 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n5 0.063
R30341 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n0 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.063
R30342 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n8 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n7 0.063
R30343 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n7 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n1 0.063
R30344 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.t3 169.46
R30345 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C.t1 167.809
R30346 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.t0 167.809
R30347 D_FlipFlop_5.3-input-nand_2.C.t4 D_FlipFlop_5.3-input-nand_2.C.n13 167.226
R30348 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C.t5 150.273
R30349 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.t4 150.273
R30350 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C.t7 73.6406
R30351 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C.t6 73.6304
R30352 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.C.t2 60.3943
R30353 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C.n7 12.3891
R30354 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n11 11.4489
R30355 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C 1.68257
R30356 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C.n2 1.38365
R30357 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C.n0 1.19615
R30358 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C.n5 1.1717
R30359 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C 1.08448
R30360 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C 0.932141
R30361 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C 0.720633
R30362 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C.n12 0.280391
R30363 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C 0.217464
R30364 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C 0.1255
R30365 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C 0.1255
R30366 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C 0.1255
R30367 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C.n9 0.0874565
R30368 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C.n6 0.063
R30369 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C 0.063
R30370 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C.n8 0.063
R30371 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C.n3 0.063
R30372 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n10 0.0435206
R30373 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.n1 0.0216397
R30374 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.C.n14 0.0216397
R30375 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C.n4 0.0107679
R30376 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C 0.0107679
R30377 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 169.46
R30378 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 168.089
R30379 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 167.809
R30380 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 150.887
R30381 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 73.6304
R30382 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 60.3943
R30383 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 12.0358
R30384 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 11.4489
R30385 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 1.05069
R30386 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 0.981478
R30387 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.769522
R30388 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 0.745065
R30389 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.580578
R30390 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 0.533109
R30391 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.428234
R30392 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.063
R30393 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 0.063
R30394 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 0.063
R30395 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.063
R30396 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 0.063
R30397 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 0.063
R30398 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 169.46
R30399 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 168.089
R30400 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 167.809
R30401 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 150.887
R30402 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 73.6304
R30403 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 60.3943
R30404 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 12.0358
R30405 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 11.4489
R30406 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 1.05069
R30407 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 0.981478
R30408 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.769522
R30409 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 0.745065
R30410 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.580578
R30411 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 0.533109
R30412 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.428234
R30413 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.063
R30414 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 0.063
R30415 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 0.063
R30416 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.063
R30417 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 0.063
R30418 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 0.063
R30419 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 169.46
R30420 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 168.089
R30421 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 167.809
R30422 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 150.887
R30423 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 73.6304
R30424 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 60.3943
R30425 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 12.0358
R30426 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 11.4489
R30427 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 1.05069
R30428 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 0.981478
R30429 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.769522
R30430 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 0.745065
R30431 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.580578
R30432 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 0.533109
R30433 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.428234
R30434 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.063
R30435 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 0.063
R30436 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 0.063
R30437 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.063
R30438 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 0.063
R30439 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 0.063
R30440 a_50454_10637.n0 a_50454_10637.t3 575.905
R30441 a_50454_10637.n1 a_50454_10637.t1 575.905
R30442 a_50454_10637.n0 a_50454_10637.t4 338.675
R30443 a_50454_10637.t0 a_50454_10637.n2 13.268
R30444 a_50454_10637.n2 a_50454_10637.t2 9.51806
R30445 a_50454_10637.n1 a_50454_10637.n0 1.7505
R30446 a_50454_10637.n2 a_50454_10637.n1 0.484196
C0 a_16465_60797# CLK 0.06211f
C1 a_45827_58825# Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.04443f
C2 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout EN 0.61231f
C3 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B a_35135_60797# 0.04443f
C4 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B a_10187_60797# 0.04443f
C5 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.10915f
C6 D_FlipFlop_0.CLK a_50544_48405# 0.04443f
C7 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_2.Vout 0.1215f
C8 a_42263_60797# VDD 0.02865f
C9 a_n9432_51119# a_n8818_51119# 0.05935f
C10 Nand_Gate_6.A a_16465_58825# 0.05925f
C11 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.06935f
C12 a_20029_61411# a_20029_60797# 0.05935f
C13 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.08674f
C14 Nand_Gate_5.A a_41413_54751# 0.06359f
C15 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.01162f
C16 D_FlipFlop_4.nPRE a_16465_55365# 0.01335f
C17 Ring_Counter_0.D_FlipFlop_9.Qbar a_20029_54751# 0.04443f
C18 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_n1355_56723# 0.05964f
C19 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B VDD 1.83506f
C20 a_49391_59439# Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.01335f
C21 D_FlipFlop_5.CLK a_16854_48405# 0.02953f
C22 D_FlipFlop_3.nPRE a_28044_52049# 0.04597f
C23 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.09856f
C24 a_35135_54751# Ring_Counter_0.D_FlipFlop_4.Qbar 0.06113f
C25 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout EN 0.09223f
C26 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C a_10187_56723# 0.04443f
C27 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout EN 0.96763f
C28 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.30156f
C29 a_20029_61411# EN 0.02636f
C30 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout EN 0.78583f
C31 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout VDD 2.29929f
C32 D_FlipFlop_7.nPRE a_n11404_48405# 0.0452f
C33 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 1.09973f
C34 a_41413_60797# CLK 0.06211f
C35 Ring_Counter_0.D_FlipFlop_16.Q a_10187_60797# 0.01768f
C36 a_47214_51119# a_47828_51119# 0.05935f
C37 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.08462f
C38 And_Gate_1.Nand_Gate_0.Vout a_n2995_52049# 0.05964f
C39 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.10034f
C40 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.15413f
C41 a_17468_48405# VDD 0.02521f
C42 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout CLK 0.12427f
C43 Nand_Gate_5.A a_37849_54751# 0.05925f
C44 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout a_44977_59439# 0.04995f
C45 a_17315_55365# a_17315_54751# 0.05935f
C46 D_FlipFlop_4.nPRE a_12901_55365# 0.05925f
C47 a_35135_61411# a_35135_60797# 0.05935f
C48 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout a_34285_60797# 0.05964f
C49 D_FlipFlop_1.Nand_Gate_1.Vout a_45856_48405# 0.05964f
C50 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.06955f
C51 D_FlipFlop_5.3-input-nand_2.Vout a_19570_51119# 0.04443f
C52 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout CLK 0.20785f
C53 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout VDD 2.07898f
C54 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_4.Qbar 0.07122f
C55 Ring_Counter_0.D_FlipFlop_0.Qbar EN 0.1585f
C56 a_n2642_51119# D_FlipFlop_6.3-input-nand_0.Vout 0.01335f
C57 D_FlipFlop_7.nPRE And_Gate_0.A 0.37721f
C58 a_34378_51119# a_34992_51119# 0.05935f
C59 a_19282_52049# VDD 0.02521f
C60 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C EN 0.07565f
C61 D_FlipFlop_5.Nand_Gate_1.Vout a_21542_48405# 0.04444f
C62 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.04109f
C63 a_31486_45397# Q6 0.46416f
C64 And_Gate_7.Nand_Gate_0.Vout VDD 1.39555f
C65 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout EN 0.95226f
C66 a_10808_51119# VDD 0.02521f
C67 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.Nand_Gate_1.Vout 0.1541f
C68 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.Vout 1.01753f
C69 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout EN 0.97707f
C70 a_44977_61411# EN 0.02636f
C71 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout EN 0.087f
C72 a_48541_58825# VDD 0.02521f
C73 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout a_34285_58825# 0.05964f
C74 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.16431f
C75 D_FlipFlop_1.3-input-nand_1.B VDD 1.3477f
C76 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C CLK 0.19664f
C77 CDAC_v3_0.switch_4.Z CDAC_v3_0.switch_7.Z 51.5071f
C78 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_6.Z 36.1389f
C79 CDAC_v3_0.switch_0.Z CDAC_v3_0.OUT 10.2622f
C80 Ring_Counter_0.D_FlipFlop_10.Qbar a_16465_54751# 0.04443f
C81 a_n2028_51119# VDD 0.02521f
C82 Ring_Counter_0.D_FlipFlop_16.Q a_35135_60797# 0.01768f
C83 a_38699_59439# VDD 0.05686f
C84 D_FlipFlop_2.CLK D_FlipFlop_2.3-input-nand_1.B 0.06986f
C85 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.01262f
C86 D_FlipFlop_3.nPRE CLK 0.7173f
C87 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.29165f
C88 D_FlipFlop_3.3-input-nand_2.Vout VDD 2.67043f
C89 a_31571_54751# Ring_Counter_0.D_FlipFlop_5.Qbar 0.06113f
C90 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.07084f
C91 CDAC_v3_0.switch_5.Z VDD 1.07109f
C92 D_FlipFlop_6.3-input-nand_2.C a_n56_48405# 0.05964f
C93 a_28007_58825# VDD 0.02578f
C94 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.04107f
C95 Nand_Gate_4.A EN 0.79742f
C96 a_44977_61411# a_44977_60797# 0.05935f
C97 D_FlipFlop_7.nPRE a_n11404_51119# 0.034f
C98 a_30721_59439# EN 0.045f
C99 a_3059_61411# VDD 0.04448f
C100 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout a_2209_61411# 0.01335f
C101 D_FlipFlop_1.Qbar a_47214_48405# 0.01335f
C102 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout VDD 2.83213f
C103 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.01262f
C104 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.29165f
C105 And_Gate_2.A CLK 1.52489f
C106 CDAC_v3_0.switch_0.Z Q3 0.02962f
C107 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD 1.48403f
C108 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B CLK 0.08407f
C109 a_13751_55365# a_13751_54751# 0.05935f
C110 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.17188f
C111 a_41168_51119# D_FlipFlop_1.3-input-nand_0.Vout 0.01335f
C112 D_FlipFlop_6.nPRE a_9337_55365# 0.01335f
C113 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.01202f
C114 D_FlipFlop_2.Inverter_1.Vout Q7 0.02322f
C115 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout CLK 0.7779f
C116 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout CLK 0.36346f
C117 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.Vout 1.01753f
C118 a_20879_58825# Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.05964f
C119 D_FlipFlop_0.Qbar VDD 1.9032f
C120 D_FlipFlop_7.Qbar Q0 1.1722f
C121 a_17315_59439# CLK 0.03166f
C122 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.21889f
C123 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout VDD 2.29929f
C124 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.06837f
C125 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C VDD 3.50703f
C126 D_FlipFlop_2.3-input-nand_1.B D_FlipFlop_2.3-input-nand_1.Vout 0.08641f
C127 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.01194f
C128 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout CLK 0.01154f
C129 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.01194f
C130 a_6623_58825# CLK 0.03f
C131 D_FlipFlop_5.3-input-nand_1.B a_15496_48405# 0.04443f
C132 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout a_27157_58825# 0.04444f
C133 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_n4069_54751# 0.04444f
C134 D_FlipFlop_1.3-input-nand_2.C VDD 2.67765f
C135 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.01194f
C136 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_8.Qbar 0.11657f
C137 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B VDD 1.78671f
C138 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_n4919_54751# 0.04444f
C139 Nand_Gate_4.A a_30721_58825# 0.05925f
C140 a_28007_61411# VDD 0.04448f
C141 VDD Q4 3.67411f
C142 a_30721_59439# a_30721_58825# 0.05935f
C143 D_FlipFlop_2.CLK D_FlipFlop_2.3-input-nand_2.C 0.19377f
C144 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout CLK 0.12427f
C145 Ring_Counter_0.D_FlipFlop_11.Qbar a_12901_54751# 0.04443f
C146 D_FlipFlop_6.nPRE a_5773_55365# 0.0598f
C147 a_28007_54751# Ring_Counter_0.D_FlipFlop_6.Qbar 0.06113f
C148 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.06837f
C149 D_FlipFlop_7.nPRE a_n1355_58825# 0.05925f
C150 a_30721_56723# VDD 0.02521f
C151 a_37094_48405# VDD 0.02521f
C152 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.Nand_Gate_1.Vout 0.1541f
C153 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout CLK 0.7779f
C154 D_FlipFlop_4.Nand_Gate_1.Vout Q2 0.09808f
C155 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK 0.36346f
C156 a_12901_59439# VDD 0.01186f
C157 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout a_16465_59439# 0.01335f
C158 a_11766_45397# Q1 0.47506f
C159 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_23593_56723# 0.05964f
C160 Ring_Counter_0.D_FlipFlop_16.Q a_n4069_61411# 0.01252f
C161 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout a_16465_56723# 0.04443f
C162 a_2209_58825# VDD 0.02521f
C163 a_10187_59439# a_10187_58825# 0.05935f
C164 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.20923f
C165 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C CLK 0.19397f
C166 a_10187_55365# a_10187_54751# 0.05935f
C167 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.04107f
C168 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.06955f
C169 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout a_27157_61411# 0.01335f
C170 a_n7633_59439# VDD 0.05686f
C171 And_Gate_0.A D_FlipFlop_7.CLK 0.06897f
C172 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout VDD 2.29929f
C173 D_FlipFlop_2.Nand_Gate_1.Vout Q5 0.09982f
C174 a_12166_51119# VDD 0.01186f
C175 a_3059_56723# Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.05964f
C176 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.3-input-nand_2.Vout 0.0846f
C177 a_n505_58825# Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.04443f
C178 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_1.Vout 0.08671f
C179 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.25884f
C180 D_FlipFlop_4.nPRE D_FlipFlop_6.Qbar 0.01961f
C181 a_n670_51119# VDD 0.01186f
C182 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B a_n4069_61411# 0.04995f
C183 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C a_9337_58825# 0.04443f
C184 D_FlipFlop_2.nPRE VDD 7.26608f
C185 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout CLK 0.20785f
C186 Ring_Counter_0.D_FlipFlop_12.Qbar a_9337_54751# 0.04443f
C187 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout VDD 1.46604f
C188 D_FlipFlop_7.nPRE a_2209_55365# 0.01335f
C189 Ring_Counter_0.D_FlipFlop_16.Q a_20879_61411# 0.01252f
C190 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.07084f
C191 a_3059_59439# Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.01335f
C192 D_FlipFlop_7.nPRE D_FlipFlop_7.3-input-nand_1.B 0.27142f
C193 a_24443_54751# Ring_Counter_0.D_FlipFlop_7.Qbar 0.06113f
C194 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Qbar 0.06863f
C195 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.01194f
C196 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout a_10187_59439# 0.04543f
C197 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.04109f
C198 D_FlipFlop_6.3-input-nand_1.B D_FlipFlop_6.3-input-nand_1.Vout 0.08641f
C199 And_Gate_0.Nand_Gate_0.Vout a_n11757_52049# 0.05964f
C200 And_Gate_4.A And_Gate_4.Nand_Gate_0.Vout 0.24482f
C201 a_49930_51119# EN 0.04501f
C202 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.06837f
C203 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 1.01604f
C204 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B VDD 1.71455f
C205 a_2046_48405# VDD 0.02521f
C206 Vbias Vin 0.78432f
C207 a_6623_56723# VDD 0.02578f
C208 D_FlipFlop_6.Qbar Q1 1.17251f
C209 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.3-input-nand_2.C 0.06863f
C210 D_FlipFlop_5.nPRE D_FlipFlop_5.Inverter_1.Vout 0.07033f
C211 a_6623_55365# a_6623_54751# 0.05935f
C212 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B CLK 0.08407f
C213 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.3-input-nand_2.Vout 0.0846f
C214 D_FlipFlop_3.3-input-nand_1.Vout a_24258_48405# 0.05964f
C215 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.25966f
C216 D_FlipFlop_7.nPRE a_n1355_55365# 0.05925f
C217 D_FlipFlop_0.Nand_Gate_0.Vout VDD 1.48317f
C218 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout EN 0.61231f
C219 Nand_Gate_4.A a_30721_61411# 0.04995f
C220 D_FlipFlop_7.Nand_Gate_0.Vout Q0 0.11094f
C221 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_3059_55365# 0.04995f
C222 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_28007_54751# 0.04444f
C223 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_2209_55365# 0.04995f
C224 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_27157_54751# 0.04444f
C225 a_n7633_60797# CLK 0.04443f
C226 CDAC_v3_0.switch_5.Z m3_3428_4751# 1.89962f
C227 Ring_Counter_0.D_FlipFlop_16.Q a_45827_61411# 0.01252f
C228 D_FlipFlop_6.3-input-nand_1.Vout a_n56_48405# 0.04444f
C229 D_FlipFlop_1.3-input-nand_0.Vout VDD 1.74442f
C230 D_FlipFlop_4.CLK D_FlipFlop_4.3-input-nand_2.Vout 0.1192f
C231 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.21575f
C232 And_Gate_1.A VDD 1.33887f
C233 D_FlipFlop_5.nPRE a_20029_61411# 0.04995f
C234 D_FlipFlop_2.CLK D_FlipFlop_2.3-input-nand_0.Vout 0.25957f
C235 D_FlipFlop_1.nPRE a_41413_60797# 0.10368f
C236 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout a_6623_56723# 0.04995f
C237 a_15710_45397# CDAC_v3_0.switch_2.Z 0.27028f
C238 CDAC_v3_0.switch_0.Z a_19654_45397# 0.022f
C239 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout a_52105_61411# 0.01335f
C240 a_10187_60797# Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.05964f
C241 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.25966f
C242 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Qbar 0.07122f
C243 a_12901_60797# VDD 0.02521f
C244 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.01162f
C245 Ring_Counter_0.D_FlipFlop_13.Qbar a_5773_54751# 0.04443f
C246 a_55976_48405# VDD 0.01186f
C247 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.06935f
C248 D_FlipFlop_7.nPRE D_FlipFlop_7.3-input-nand_2.C 0.05823f
C249 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B CLK 0.08407f
C250 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.08582f
C251 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_1.Vout 0.08671f
C252 a_20879_54751# Ring_Counter_0.D_FlipFlop_8.Qbar 0.06113f
C253 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C a_38699_56723# 0.04443f
C254 a_n4069_61411# EN 0.07048f
C255 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.3-input-nand_2.C 0.06863f
C256 D_FlipFlop_4.3-input-nand_2.C a_8706_48405# 0.05964f
C257 a_17315_60797# CLK 0.06211f
C258 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.25966f
C259 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout 0.25855f
C260 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.06837f
C261 D_FlipFlop_3.nPRE a_30721_55365# 0.01335f
C262 D_FlipFlop_0.Qbar a_55976_48405# 0.01335f
C263 D_FlipFlop_0.CLK a_52516_48405# 0.02953f
C264 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.09851f
C265 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.10034f
C266 a_3059_55365# a_3059_54751# 0.05935f
C267 D_FlipFlop_3.nPRE a_23644_48405# 0.0452f
C268 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout a_n7633_58825# 0.04444f
C269 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.15413f
C270 a_n8818_51119# D_FlipFlop_7.3-input-nand_2.Vout 0.05964f
C271 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B CLK 0.08407f
C272 a_37849_60797# VDD 0.02521f
C273 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.01202f
C274 D_FlipFlop_3.nPRE D_FlipFlop_3.Nand_Gate_0.Vout 0.5831f
C275 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 1.09983f
C276 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.01262f
C277 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.29165f
C278 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_48541_56723# 0.05964f
C279 Nand_Gate_3.A D_FlipFlop_3.nPRE 2.13698f
C280 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C281 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.01323f
C282 D_FlipFlop_3.nPRE a_27157_55365# 0.05925f
C283 a_20879_61411# EN 0.07048f
C284 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout VDD 2.29929f
C285 D_FlipFlop_5.nPRE a_20029_58825# 0.05925f
C286 a_42263_60797# CLK 0.06211f
C287 D_FlipFlop_3.3-input-nand_1.B a_24258_48405# 0.04443f
C288 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.01202f
C289 D_FlipFlop_4.Qbar a_12780_51119# 0.04443f
C290 Ring_Counter_0.D_FlipFlop_14.Qbar a_2209_54751# 0.04443f
C291 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.16431f
C292 D_FlipFlop_7.CLK D_FlipFlop_7.3-input-nand_1.B 0.06986f
C293 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B 0.29684f
C294 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout a_45827_59439# 0.04543f
C295 Ring_Counter_0.D_FlipFlop_16.Q a_5773_60797# 0.01768f
C296 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B CLK 0.06986f
C297 a_28007_56723# Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.05964f
C298 a_20928_48405# VDD 0.01186f
C299 Nand_Gate_5.A a_38699_54751# 0.05987f
C300 a_17315_54751# Ring_Counter_0.D_FlipFlop_9.Qbar 0.06113f
C301 D_FlipFlop_0.3-input-nand_1.B EN 0.33109f
C302 a_6120_51119# a_6734_51119# 0.05935f
C303 a_35135_60797# Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.05964f
C304 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.08674f
C305 D_FlipFlop_4.Qbar Q2 1.17288f
C306 D_FlipFlop_6.nPRE D_FlipFlop_6.Nand_Gate_0.Vout 0.5831f
C307 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.10915f
C308 D_FlipFlop_1.Nand_Gate_1.Vout a_47828_48405# 0.04444f
C309 D_FlipFlop_6.3-input-nand_2.C a_n56_51119# 0.04443f
C310 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout CLK 0.20785f
C311 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD 1.48403f
C312 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout a_44977_58825# 0.05964f
C313 Nand_Gate_7.A a_44977_59439# 0.05925f
C314 D_FlipFlop_6.Nand_Gate_0.Vout Q1 0.11094f
C315 a_34992_51119# D_FlipFlop_2.3-input-nand_2.Vout 0.05964f
C316 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_35135_55365# 0.04995f
C317 a_28044_52049# VDD 0.02521f
C318 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_34285_55365# 0.04995f
C319 a_56590_51119# VDD 0.02521f
C320 a_n4744_51119# Q0 0.05964f
C321 a_14882_51119# VDD 0.01186f
C322 a_n505_55365# a_n505_54751# 0.05935f
C323 a_45827_61411# EN 0.07048f
C324 a_43754_51119# VDD 0.02521f
C325 a_49391_58825# VDD 0.02521f
C326 Nand_Gate_0.A a_2209_60797# 0.10368f
C327 CDAC_v3_0.switch_5.Z CDAC_v3_0.switch_7.Z 56.6053f
C328 CDAC_v3_0.switch_2.Z CDAC_v3_0.OUT 19.1158f
C329 CDAC_v3_0.switch_4.Z CDAC_v3_0.switch_6.Z 39.3126f
C330 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.08462f
C331 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout VDD 2.8343f
C332 Ring_Counter_0.D_FlipFlop_16.Q a_30721_60797# 0.01768f
C333 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout a_20029_59439# 0.04995f
C334 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B a_13751_60797# 0.04443f
C335 D_FlipFlop_0.Qbar a_56590_51119# 0.04443f
C336 CDAC_v3_0.switch_7.Z VDD 1.07386f
C337 And_Gate_7.Nand_Gate_0.Vout CLK 0.62717f
C338 And_Gate_7.Nand_Gate_0.Vout D_FlipFlop_0.CLK 0.25559f
C339 Nand_Gate_7.A a_48541_54751# 0.06359f
C340 D_FlipFlop_7.nPRE D_FlipFlop_7.3-input-nand_0.Vout 0.94513f
C341 a_3059_61411# Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.01335f
C342 D_FlipFlop_7.CLK D_FlipFlop_7.3-input-nand_2.C 0.19377f
C343 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout VDD 2.72531f
C344 a_49930_51119# a_50544_51119# 0.05935f
C345 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD 1.89599f
C346 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout EN 0.61231f
C347 Ring_Counter_0.D_FlipFlop_15.Qbar a_n1355_54751# 0.04443f
C348 a_n1355_61411# VDD 0.08862f
C349 D_FlipFlop_0.3-input-nand_2.C EN 0.81235f
C350 a_31571_58825# Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.05964f
C351 a_38699_59439# CLK 0.03166f
C352 D_FlipFlop_1.3-input-nand_2.C a_43754_51119# 0.04443f
C353 a_12901_56723# VDD 0.02521f
C354 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.26069f
C355 a_13751_54751# Ring_Counter_0.D_FlipFlop_10.Qbar 0.06113f
C356 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.20923f
C357 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout EN 0.78583f
C358 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C VDD 3.50703f
C359 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.01194f
C360 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.01194f
C361 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.01323f
C362 a_28007_58825# CLK 0.03f
C363 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.01202f
C364 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C365 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.1143f
C366 a_41413_59439# a_41413_58825# 0.05935f
C367 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout CLK 0.53027f
C368 VDD CLK 53.0347f
C369 D_FlipFlop_0.CLK VDD 2.17541f
C370 Nand_Gate_7.A a_44977_54751# 0.05925f
C371 D_FlipFlop_3.Nand_Gate_1.Vout Q5 0.01969f
C372 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout a_28007_58825# 0.04444f
C373 D_FlipFlop_6.Nand_Gate_1.Vout a_3404_48405# 0.04995f
C374 a_n4069_55365# a_n4069_54751# 0.05935f
C375 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout a_44977_56723# 0.04443f
C376 D_FlipFlop_3.CLK a_24258_48405# 0.04443f
C377 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout VDD 2.72531f
C378 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD 1.89599f
C379 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.06837f
C380 a_52105_55365# VDD 0.0563f
C381 a_23593_61411# VDD 0.08862f
C382 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C EN 0.07565f
C383 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B EN 0.37578f
C384 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout a_27157_59439# 0.01335f
C385 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.09856f
C386 a_34285_59439# VDD 0.01186f
C387 Nand_Gate_0.A a_2209_59439# 0.05925f
C388 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout CLK 0.20785f
C389 D_FlipFlop_7.CLK a_n9432_48405# 0.02953f
C390 a_20879_59439# a_20879_58825# 0.05935f
C391 a_23593_58825# VDD 0.02521f
C392 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Qbar 1.14393f
C393 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.26069f
C394 D_FlipFlop_4.Nand_Gate_0.Vout a_12780_51119# 0.04444f
C395 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C CLK 0.19664f
C396 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout VDD 2.07898f
C397 a_39066_48405# VDD 0.02521f
C398 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C a_n505_56723# 0.04443f
C399 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B CLK 0.08407f
C400 D_FlipFlop_7.nPRE a_n11757_52049# 0.02193f
C401 D_FlipFlop_5.Qbar Q3 1.17143f
C402 a_13751_59439# VDD 0.05686f
C403 D_FlipFlop_0.3-input-nand_2.Vout Q7 0.01585f
C404 Ring_Counter_0.D_FlipFlop_16.Qbar a_n4919_54751# 0.04443f
C405 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.06935f
C406 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.01202f
C407 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_9.Qbar 0.07122f
C408 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.0646f
C409 D_FlipFlop_4.Nand_Gate_0.Vout Q2 0.11094f
C410 a_10187_58825# Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.04443f
C411 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.13492f
C412 a_3059_58825# VDD 0.02578f
C413 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout a_2209_58825# 0.04444f
C414 a_48541_55365# VDD 0.01186f
C415 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.01262f
C416 a_10187_54751# Ring_Counter_0.D_FlipFlop_11.Qbar 0.06113f
C417 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.29165f
C418 a_5773_59439# EN 0.045f
C419 a_4018_51119# Q1 0.05964f
C420 D_FlipFlop_6.3-input-nand_0.Vout a_n56_51119# 0.04444f
C421 a_28007_61411# Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.01335f
C422 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout VDD 2.74716f
C423 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout VDD 2.75736f
C424 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout VDD 2.29929f
C425 a_48541_61411# VDD 0.07045f
C426 D_FlipFlop_5.3-input-nand_1.B VDD 1.34773f
C427 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C a_20029_58825# 0.04443f
C428 D_FlipFlop_5.3-input-nand_2.C a_17468_48405# 0.05964f
C429 a_13751_59439# Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.01335f
C430 D_FlipFlop_6.3-input-nand_2.Vout VDD 2.67043f
C431 a_n7633_55365# a_n7633_54751# 0.05935f
C432 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.08582f
C433 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout a_5773_56723# 0.04443f
C434 a_n7633_59439# CLK 0.02953f
C435 a_44977_55365# VDD 0.01186f
C436 And_Gate_7.A a_49577_52049# 0.04995f
C437 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout CLK 0.20785f
C438 D_FlipFlop_0.Nand_Gate_0.Vout a_56590_51119# 0.04444f
C439 D_FlipFlop_1.nPRE a_41168_51119# 0.034f
C440 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.48403f
C441 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.0646f
C442 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 1.09973f
C443 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.06462f
C444 Ring_Counter_0.D_FlipFlop_16.Q a_16465_61411# 0.01252f
C445 D_FlipFlop_7.CLK D_FlipFlop_7.3-input-nand_0.Vout 0.25957f
C446 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.06955f
C447 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.01323f
C448 D_FlipFlop_0.3-input-nand_0.Vout EN 0.18661f
C449 D_FlipFlop_5.nPRE Q3 0.03683f
C450 a_n4069_61411# a_n4069_60797# 0.05935f
C451 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout a_n4919_60797# 0.05964f
C452 a_4018_48405# VDD 0.02521f
C453 D_FlipFlop_1.3-input-nand_0.Vout a_43754_51119# 0.04444f
C454 D_FlipFlop_0.3-input-nand_1.Vout a_50544_48405# 0.05964f
C455 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.06955f
C456 D_FlipFlop_2.nPRE CLK 0.70981f
C457 D_FlipFlop_3.Qbar VDD 1.96371f
C458 D_FlipFlop_2.3-input-nand_1.B a_33020_48405# 0.04443f
C459 a_41413_55365# VDD 0.01186f
C460 a_6623_54751# Ring_Counter_0.D_FlipFlop_12.Qbar 0.06113f
C461 Nand_Gate_5.A EN 0.79742f
C462 D_FlipFlop_3.3-input-nand_1.Vout a_26230_48405# 0.04444f
C463 D_FlipFlop_5.3-input-nand_2.C VDD 2.67794f
C464 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.Qbar 1.27496f
C465 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_13.Qbar 0.11657f
C466 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout 0.30046f
C467 And_Gate_6.Nand_Gate_0.Vout VDD 1.39327f
C468 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.Inverter_1.Vout 0.06895f
C469 CDAC_v3_0.switch_6.Z m3_3428_33935# 16.1764f
C470 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.07084f
C471 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.0646f
C472 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout a_n1355_58825# 0.05964f
C473 D_FlipFlop_2.nPRE a_34285_59439# 0.05925f
C474 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.06462f
C475 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B CLK 0.08407f
C476 Ring_Counter_0.D_FlipFlop_16.Q a_41413_61411# 0.01252f
C477 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.09397f
C478 CDAC_v3_0.switch_0.Z a_23598_45397# 0.02212f
C479 VDD Q0 3.77344f
C480 a_13751_60797# VDD 0.02865f
C481 a_37849_55365# VDD 0.01186f
C482 a_5773_61411# a_5773_60797# 0.05935f
C483 a_7822_45397# VDD 1.17814f
C484 D_FlipFlop_3.Qbar Q4 1.17143f
C485 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.Qbar 0.13504f
C486 D_FlipFlop_3.Inverter_1.Vout a_28332_51119# 0.04443f
C487 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_0.Qbar 0.07122f
C488 D_FlipFlop_5.Nand_Gate_0.Vout Q3 0.11094f
C489 And_Gate_1.A CLK 1.52489f
C490 And_Gate_4.A D_FlipFlop_3.CLK 0.06897f
C491 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B a_n505_61411# 0.04995f
C492 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.06837f
C493 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout EN 0.09223f
C494 a_12780_51119# Q2 0.05964f
C495 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout EN 0.96763f
C496 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.09856f
C497 a_n670_51119# D_FlipFlop_6.3-input-nand_2.Vout 0.01335f
C498 a_12901_60797# CLK 0.06211f
C499 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.Inverter_1.Vout 0.26069f
C500 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout a_37849_58825# 0.04444f
C501 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.Inverter_1.Vout 0.06895f
C502 a_34285_55365# VDD 0.01186f
C503 a_3059_54751# Ring_Counter_0.D_FlipFlop_13.Qbar 0.06113f
C504 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout a_5773_56723# 0.04443f
C505 a_20879_61411# a_20879_60797# 0.05935f
C506 D_FlipFlop_4.3-input-nand_1.Vout a_6120_48405# 0.01335f
C507 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_10.Qbar 0.01625f
C508 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout a_20029_60797# 0.05964f
C509 a_38699_60797# VDD 0.02865f
C510 And_Gate_7.A EN 0.06541f
C511 D_FlipFlop_1.Inverter_1.Vout VDD 1.70303f
C512 VDD Vbias 0.3571p
C513 a_n4919_59439# a_n4919_58825# 0.05935f
C514 D_FlipFlop_2.CLK D_FlipFlop_2.Inverter_1.Vout 0.20785f
C515 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout 0.01202f
C516 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.06734f
C517 a_19570_51119# D_FlipFlop_5.Nand_Gate_0.Vout 0.05964f
C518 D_FlipFlop_1.nPRE D_FlipFlop_1.3-input-nand_1.B 0.27142f
C519 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout EN 0.09223f
C520 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout EN 0.96763f
C521 a_47214_48405# a_47828_48405# 0.05935f
C522 a_16465_61411# EN 0.02636f
C523 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout VDD 2.29929f
C524 a_30721_55365# VDD 0.01186f
C525 a_38699_56723# VDD 0.02578f
C526 a_37849_60797# CLK 0.06211f
C527 D_FlipFlop_4.CLK D_FlipFlop_4.3-input-nand_1.Vout 0.67419f
C528 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout 0.30046f
C529 D_FlipFlop_5.CLK a_15496_51119# 0.04443f
C530 D_FlipFlop_2.nPRE D_FlipFlop_3.Qbar 0.01961f
C531 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.Nand_Gate_0.Vout 0.16429f
C532 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.06955f
C533 Ring_Counter_0.D_FlipFlop_16.Q a_6623_60797# 0.01768f
C534 a_23644_48405# VDD 0.01212f
C535 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.Qbar 1.27496f
C536 a_6734_51119# D_FlipFlop_4.3-input-nand_0.Vout 0.05964f
C537 a_43140_51119# D_FlipFlop_1.3-input-nand_2.Vout 0.01335f
C538 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.Inverter_1.Vout 0.26069f
C539 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.26069f
C540 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout EN 0.61231f
C541 D_FlipFlop_1.nPRE VDD 7.2893f
C542 a_30721_61411# a_30721_60797# 0.05935f
C543 D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.43587f
C544 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_10187_54751# 0.04444f
C545 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout CLK 0.20785f
C546 a_n4919_56723# VDD 0.02521f
C547 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_4.Qbar 0.11657f
C548 a_36806_52049# VDD 0.02521f
C549 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_9337_54751# 0.04444f
C550 Nand_Gate_3.A VDD 4.36236f
C551 D_FlipFlop_5.3-input-nand_0.Vout VDD 1.74442f
C552 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_5773_56723# 0.05964f
C553 a_27157_55365# VDD 0.01186f
C554 a_n505_54751# Ring_Counter_0.D_FlipFlop_14.Qbar 0.06113f
C555 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout a_24443_56723# 0.04995f
C556 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout EN 0.09223f
C557 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout EN 0.96763f
C558 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.10915f
C559 a_41413_61411# EN 0.02636f
C560 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.07084f
C561 CDAC_v3_0.switch_5.Z CDAC_v3_0.switch_6.Z 36.1069f
C562 CDAC_v3_0.switch_3.Z CDAC_v3_0.OUT 37.6729f
C563 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.Qbar 0.14329f
C564 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout EN 0.08727f
C565 D_FlipFlop_2.nPRE a_37849_55365# 0.01335f
C566 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout a_20879_59439# 0.04543f
C567 Ring_Counter_0.D_FlipFlop_16.Q a_31571_60797# 0.01768f
C568 D_FlipFlop_2.Qbar Q5 1.17195f
C569 D_FlipFlop_5.nPRE a_20928_51119# 0.04443f
C570 D_FlipFlop_1.nPRE D_FlipFlop_1.3-input-nand_2.C 0.05823f
C571 CDAC_v3_0.switch_6.Z VDD 1.0692f
C572 And_Gate_6.A a_40815_52049# 0.04995f
C573 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.08674f
C574 a_42263_58825# Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.05964f
C575 D_FlipFlop_3.3-input-nand_2.C a_26230_48405# 0.05964f
C576 a_45827_61411# a_45827_60797# 0.05935f
C577 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout a_44977_60797# 0.05964f
C578 D_FlipFlop_3.Nand_Gate_0.Vout Q4 0.11094f
C579 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout EN 0.78583f
C580 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout a_30721_56723# 0.04443f
C581 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.01194f
C582 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.01194f
C583 a_50544_51119# D_FlipFlop_0.3-input-nand_0.Vout 0.05964f
C584 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.01194f
C585 a_23593_55365# VDD 0.01186f
C586 a_49391_58825# CLK 0.03f
C587 a_n505_61411# VDD 0.04448f
C588 a_21542_51119# Q3 0.05964f
C589 CDAC_v3_0.switch_3.Z Q3 0.17576f
C590 a_29690_48405# a_30304_48405# 0.05935f
C591 a_52105_59439# a_52105_58825# 0.05935f
C592 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout CLK 0.12427f
C593 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_12.Qbar 0.02118f
C594 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout VDD 2.07898f
C595 D_FlipFlop_2.nPRE a_34285_55365# 0.05925f
C596 a_n11404_48405# VDD 0.01186f
C597 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.04109f
C598 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.01202f
C599 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.08462f
C600 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout a_38699_56723# 0.04995f
C601 D_FlipFlop_3.Nand_Gate_1.Vout a_29690_48405# 0.04995f
C602 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C a_28007_56723# 0.04443f
C603 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout CLK 0.7779f
C604 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout a_n4919_59439# 0.04995f
C605 D_FlipFlop_3.nPRE a_27157_56723# 0.05925f
C606 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout CLK 0.36346f
C607 Nand_Gate_7.A a_45827_54751# 0.05987f
C608 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C EN 0.07565f
C609 D_FlipFlop_6.nPRE a_n2995_52049# 0.02193f
C610 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.17193f
C611 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout a_37849_59439# 0.01335f
C612 D_FlipFlop_4.nPRE a_8092_51119# 0.045f
C613 a_20029_55365# VDD 0.01186f
C614 a_n4069_54751# Ring_Counter_0.D_FlipFlop_15.Qbar 0.06113f
C615 D_FlipFlop_3.CLK a_26230_48405# 0.02953f
C616 D_FlipFlop_1.3-input-nand_1.B a_41782_48405# 0.04443f
C617 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.09856f
C618 a_44977_58825# VDD 0.02521f
C619 a_31571_59439# a_31571_58825# 0.05935f
C620 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.04107f
C621 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C CLK 0.19664f
C622 And_Gate_0.A VDD 1.37593f
C623 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.15413f
C624 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B a_17315_61411# 0.04995f
C625 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.01323f
C626 a_24443_61411# VDD 0.04448f
C627 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout a_12901_61411# 0.01335f
C628 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B a_38699_60797# 0.04443f
C629 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.Qbar 1.27567f
C630 D_FlipFlop_5.Nand_Gate_0.Vout a_20928_51119# 0.04543f
C631 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout a_44977_56723# 0.04443f
C632 a_35135_59439# VDD 0.05686f
C633 D_FlipFlop_0.CLK CLK 0.01125f
C634 D_FlipFlop_2.3-input-nand_1.B Q6 0.01803f
C635 D_FlipFlop_7.nPRE D_FlipFlop_7.Inverter_1.Vout 0.07033f
C636 a_24443_58825# VDD 0.02578f
C637 a_20879_58825# Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.04443f
C638 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B a_28007_60797# 0.04443f
C639 a_41782_48405# VDD 0.02521f
C640 a_27157_59439# EN 0.045f
C641 D_FlipFlop_6.nPRE a_5773_60797# 0.10368f
C642 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.48403f
C643 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.01202f
C644 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout VDD 2.8343f
C645 a_16465_55365# VDD 0.01186f
C646 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B a_45827_60797# 0.04443f
C647 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout CLK 0.7779f
C648 D_FlipFlop_4.3-input-nand_0.Vout a_8092_51119# 0.04543f
C649 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK 0.36346f
C650 D_FlipFlop_2.nPRE a_36806_52049# 0.04443f
C651 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout a_3059_58825# 0.04444f
C652 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C a_30721_58825# 0.04443f
C653 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_17315_55365# 0.04995f
C654 D_FlipFlop_3.nPRE Nand_Gate_4.A 0.04143f
C655 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_42263_54751# 0.04444f
C656 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.16431f
C657 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_16465_55365# 0.04995f
C658 a_49391_55365# VDD 0.01186f
C659 a_30304_51119# VDD 0.02521f
C660 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_41413_54751# 0.04444f
C661 D_FlipFlop_6.nPRE a_5773_59439# 0.05925f
C662 a_12166_48405# a_12780_48405# 0.05935f
C663 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.Qbar 0.14772f
C664 a_n11404_51119# VDD 0.01186f
C665 a_24443_59439# Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.01335f
C666 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.01194f
C667 a_17468_51119# VDD 0.02521f
C668 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B 0.29684f
C669 a_49391_61411# VDD 0.07122f
C670 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout VDD 2.29929f
C671 a_13751_59439# CLK 0.03166f
C672 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B 0.02535f
C673 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.30156f
C674 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C VDD 3.50703f
C675 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 1.09973f
C676 a_12901_55365# VDD 0.01186f
C677 a_n7633_54751# Ring_Counter_0.D_FlipFlop_16.Qbar 0.06113f
C678 a_3059_58825# CLK 0.03f
C679 D_FlipFlop_1.Qbar Q6 1.17198f
C680 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout CLK 0.12198f
C681 a_45827_55365# VDD 0.0563f
C682 D_FlipFlop_2.Nand_Gate_0.Vout Q5 0.11094f
C683 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_14.Qbar 0.03196f
C684 D_FlipFlop_1.nPRE D_FlipFlop_1.3-input-nand_0.Vout 0.94459f
C685 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout CLK 0.25966f
C686 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout CLK 0.20785f
C687 a_30304_51119# Q4 0.05964f
C688 a_44977_56723# VDD 0.02521f
C689 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.08674f
C690 Ring_Counter_0.D_FlipFlop_16.Q a_17315_61411# 0.01252f
C691 D_FlipFlop_0.3-input-nand_0.Vout a_51902_51119# 0.04995f
C692 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B a_49391_61411# 0.04995f
C693 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.04107f
C694 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_30721_56723# 0.05964f
C695 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout a_37849_61411# 0.01335f
C696 a_n4069_60797# Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.05964f
C697 a_9337_59439# VDD 0.01186f
C698 a_9337_55365# VDD 0.01186f
C699 a_6734_48405# VDD 0.02521f
C700 D_FlipFlop_0.3-input-nand_1.Vout a_52516_48405# 0.04444f
C701 D_FlipFlop_0.Nand_Gate_1.Vout VDD 1.46558f
C702 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout a_9337_58825# 0.05964f
C703 a_n1355_58825# VDD 0.02521f
C704 a_42263_55365# VDD 0.0563f
C705 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_15.Qbar 0.01691f
C706 a_10187_56723# Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.05964f
C707 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.Qbar 1.27148f
C708 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.30156f
C709 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.08462f
C710 a_n5358_48405# a_n4744_48405# 0.05935f
C711 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.01262f
C712 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.29165f
C713 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout a_30721_59439# 0.04995f
C714 CDAC_v3_0.switch_0.Z Q6 0.02956f
C715 CDAC_v3_0.switch_6.Z m3_3428_4751# 16.1792f
C716 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout EN 0.08727f
C717 Ring_Counter_0.D_FlipFlop_16.Q a_42263_61411# 0.01252f
C718 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.01262f
C719 D_FlipFlop_0.Qbar D_FlipFlop_0.Nand_Gate_1.Vout 0.11654f
C720 a_5773_55365# VDD 0.01186f
C721 CDAC_v3_0.switch_0.Z a_27542_45397# 0.02212f
C722 a_20928_51119# a_21542_51119# 0.05935f
C723 a_19654_45397# CDAC_v3_0.switch_3.Z 0.27076f
C724 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.29165f
C725 D_FlipFlop_1.3-input-nand_1.B Q7 0.02377f
C726 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.30156f
C727 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout a_34285_56723# 0.04443f
C728 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.12285f
C729 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C730 a_38699_55365# VDD 0.0563f
C731 D_FlipFlop_6.CLK a_n2028_48405# 0.04443f
C732 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.04109f
C733 a_11766_45397# VDD 1.17814f
C734 And_Gate_5.A a_32053_52049# 0.04995f
C735 And_Gate_6.Nand_Gate_0.Vout CLK 0.79128f
C736 a_9337_60797# VDD 0.02521f
C737 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.Qbar 0.12528f
C738 D_FlipFlop_7.CLK D_FlipFlop_7.Inverter_1.Vout 0.20785f
C739 D_FlipFlop_7.3-input-nand_2.Vout a_n6716_51119# 0.04443f
C740 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_14.Qbar 0.07122f
C741 D_FlipFlop_0.Inverter_1.Vout EN 0.56808f
C742 a_8092_51119# a_8706_51119# 0.05935f
C743 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout a_49391_55365# 0.04995f
C744 a_n4069_58825# Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.05964f
C745 D_FlipFlop_1.CLK D_FlipFlop_1.3-input-nand_1.B 0.06986f
C746 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.08582f
C747 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_48541_55365# 0.04995f
C748 a_20879_56723# VDD 0.02578f
C749 VDD Q7 3.93306f
C750 a_n7633_61411# EN 0.0452f
C751 D_FlipFlop_2.3-input-nand_2.C a_34992_48405# 0.05964f
C752 a_2209_55365# VDD 0.01186f
C753 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout a_38699_58825# 0.04444f
C754 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.30156f
C755 a_13751_60797# CLK 0.06211f
C756 D_FlipFlop_7.3-input-nand_1.B VDD 1.38856f
C757 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout EN 0.61231f
C758 D_FlipFlop_2.3-input-nand_1.Vout a_32406_48405# 0.01335f
C759 a_5773_59439# a_5773_58825# 0.05935f
C760 CDAC_v3_0.OUT Vin 0.01779f
C761 a_35135_55365# VDD 0.0563f
C762 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_16.Qbar 0.01148f
C763 D_FlipFlop_1.CLK VDD 2.17721f
C764 a_20879_60797# Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.05964f
C765 D_FlipFlop_4.3-input-nand_1.Vout a_8092_48405# 0.04543f
C766 D_FlipFlop_0.Qbar Q7 1.22378f
C767 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout VDD 2.29929f
C768 a_34285_60797# VDD 0.02521f
C769 D_FlipFlop_1.Nand_Gate_0.Vout Q6 0.11094f
C770 D_FlipFlop_1.3-input-nand_2.C Q7 0.02769f
C771 Nand_Gate_3.A a_28044_52049# 0.04443f
C772 a_39066_51119# Q5 0.05964f
C773 a_n1355_55365# VDD 0.01186f
C774 Q5 Q6 3.81026f
C775 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.Qbar 1.28455f
C776 D_FlipFlop_2.3-input-nand_2.Vout a_37094_51119# 0.04443f
C777 a_14882_51119# D_FlipFlop_5.3-input-nand_0.Vout 0.01335f
C778 a_17315_61411# EN 0.07048f
C779 a_51902_51119# a_52516_51119# 0.05935f
C780 a_31571_55365# VDD 0.0563f
C781 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout a_12901_58825# 0.04444f
C782 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.10915f
C783 D_FlipFlop_0.3-input-nand_1.B a_50544_48405# 0.04443f
C784 a_38699_60797# CLK 0.06211f
C785 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout VDD 2.29929f
C786 a_27542_45397# Q5 0.46416f
C787 a_51902_48405# EN 0.045f
C788 a_45856_51119# VDD 0.02521f
C789 D_FlipFlop_5.nPRE a_14882_48405# 0.0452f
C790 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_2.Vout 1.01753f
C791 D_FlipFlop_1.CLK D_FlipFlop_1.3-input-nand_2.C 0.19377f
C792 a_25616_48405# VDD 0.01186f
C793 D_FlipFlop_6.Qbar VDD 1.96371f
C794 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.06837f
C795 Ring_Counter_0.D_FlipFlop_16.Q a_2209_60797# 0.01768f
C796 D_FlipFlop_5.Qbar D_FlipFlop_5.Nand_Gate_1.Vout 0.11654f
C797 And_Gate_2.Nand_Gate_0.Vout D_FlipFlop_4.CLK 0.25559f
C798 a_33020_51119# VDD 0.02521f
C799 D_FlipFlop_0.3-input-nand_1.Vout VDD 1.78027f
C800 D_FlipFlop_7.3-input-nand_2.C VDD 2.67765f
C801 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.01162f
C802 a_n4919_55365# VDD 0.01186f
C803 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout VDD 2.07898f
C804 a_45568_52049# VDD 0.02521f
C805 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.Qbar 0.12814f
C806 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout CLK 0.20785f
C807 a_28007_55365# VDD 0.0563f
C808 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.01202f
C809 a_42263_61411# EN 0.07048f
C810 CDAC_v3_0.switch_4.Z CDAC_v3_0.OUT 75.3701f
C811 CDAC_v3_0.switch_7.Z CDAC_v3_0.switch_6.Z 42.291f
C812 D_FlipFlop_1.nPRE CLK 0.7153f
C813 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.01194f
C814 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.01194f
C815 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.04109f
C816 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.06955f
C817 Nand_Gate_7.A EN 0.8565f
C818 Ring_Counter_0.D_FlipFlop_16.Q a_27157_60797# 0.01768f
C819 Nand_Gate_3.A CLK 0.51831f
C820 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.10034f
C821 a_45827_60797# Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.05964f
C822 D_FlipFlop_4.nPRE a_5767_52049# 0.02193f
C823 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_5.Qbar 0.07122f
C824 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_2.Vout 1.09975f
C825 a_35135_56723# Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.05964f
C826 a_24443_55365# VDD 0.0563f
C827 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout VDD 2.72531f
C828 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD 1.89599f
C829 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.15413f
C830 a_n4919_61411# VDD 0.08862f
C831 Nand_Gate_3.A a_23593_61411# 0.04995f
C832 Nand_Gate_7.A a_44977_60797# 0.10368f
C833 D_FlipFlop_0.Nand_Gate_1.Vout a_55976_48405# 0.04995f
C834 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C EN 0.76213f
C835 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD 1.48403f
C836 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout a_48541_59439# 0.01335f
C837 a_n9432_48405# VDD 0.01186f
C838 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.07084f
C839 Nand_Gate_3.A a_23593_58825# 0.05925f
C840 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.01202f
C841 a_42263_59439# a_42263_58825# 0.05935f
C842 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout a_n4069_59439# 0.04543f
C843 D_FlipFlop_2.nPRE a_34285_60797# 0.10368f
C844 D_FlipFlop_5.Inverter_1.Vout VDD 1.70539f
C845 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.16973f
C846 Ring_Counter_0.D_FlipFlop_16.Q a_52105_60797# 0.04443f
C847 D_FlipFlop_4.nPRE D_FlipFlop_4.3-input-nand_2.Vout 0.76528f
C848 And_Gate_5.Nand_Gate_0.Vout VDD 1.39377f
C849 a_20879_55365# VDD 0.0563f
C850 D_FlipFlop_0.Nand_Gate_0.Vout Q7 0.11443f
C851 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.16431f
C852 a_7822_45397# Q0 0.47798f
C853 a_45827_58825# VDD 0.02578f
C854 a_47828_51119# Q6 0.05964f
C855 a_31571_58825# Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.04443f
C856 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout a_n4919_56723# 0.04443f
C857 a_13751_61411# Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.01335f
C858 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.08582f
C859 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout VDD 2.72531f
C860 a_48541_59439# EN 0.045f
C861 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.06935f
C862 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD 1.89599f
C863 a_20029_61411# VDD 0.08862f
C864 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout VDD 2.8343f
C865 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.01162f
C866 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C a_41413_58825# 0.04443f
C867 And_Gate_4.A a_23291_52049# 0.04995f
C868 D_FlipFlop_5.CLK D_FlipFlop_5.3-input-nand_2.Vout 0.1192f
C869 a_43754_48405# VDD 0.02521f
C870 D_FlipFlop_1.nPRE a_44977_55365# 0.01335f
C871 a_47214_51119# VDD 0.01186f
C872 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout a_48541_58825# 0.04444f
C873 a_35135_59439# Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.01335f
C874 a_27157_56723# VDD 0.02521f
C875 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.3-input-nand_2.Vout 0.0846f
C876 a_17315_55365# VDD 0.0563f
C877 D_FlipFlop_1.CLK D_FlipFlop_1.3-input-nand_0.Vout 0.25957f
C878 D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.43587f
C879 And_Gate_0.A CLK 1.35158f
C880 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_n7633_54751# 0.04444f
C881 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_9.Qbar 0.11657f
C882 a_34378_51119# VDD 0.01186f
C883 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.07152f
C884 a_35135_59439# CLK 0.03166f
C885 Ring_Counter_0.D_FlipFlop_0.Qbar VDD 1.95435f
C886 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout EN 0.78583f
C887 D_FlipFlop_7.3-input-nand_0.Vout VDD 1.74441f
C888 D_FlipFlop_1.Nand_Gate_1.Vout VDD 1.44304f
C889 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 1.09973f
C890 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C VDD 3.50703f
C891 a_24443_58825# CLK 0.03f
C892 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.10034f
C893 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout VDD 1.86486f
C894 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD 1.88044f
C895 a_44977_61411# VDD 0.08862f
C896 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout VDD 2.29893f
C897 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.06935f
C898 D_FlipFlop_4.Nand_Gate_1.Vout a_10808_48405# 0.05964f
C899 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout CLK 0.12427f
C900 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Qbar 0.06863f
C901 D_FlipFlop_1.nPRE a_41413_55365# 0.05925f
C902 D_FlipFlop_1.3-input-nand_2.C a_43754_48405# 0.05964f
C903 a_13751_55365# VDD 0.0563f
C904 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout a_10187_56723# 0.04995f
C905 D_FlipFlop_1.nPRE And_Gate_6.Nand_Gate_0.Vout 0.12437f
C906 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.25966f
C907 Ring_Counter_0.D_FlipFlop_1.Qbar VDD 1.99811f
C908 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C EN 0.07565f
C909 Nand_Gate_4.A VDD 4.53917f
C910 a_30721_59439# VDD 0.01186f
C911 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.1143f
C912 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.3-input-nand_2.C 0.06863f
C913 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.Nand_Gate_1.Vout 0.1541f
C914 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout CLK 0.20785f
C915 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout VDD 2.07898f
C916 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.0646f
C917 Nand_Gate_2.A a_9337_61411# 0.04995f
C918 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_2.Vout 0.0846f
C919 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout 0.25855f
C920 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.06462f
C921 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.01202f
C922 Ring_Counter_0.D_FlipFlop_16.Q a_12901_61411# 0.01252f
C923 a_20029_58825# VDD 0.02521f
C924 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout a_20029_58825# 0.05964f
C925 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.09856f
C926 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C927 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout 0.08377f
C928 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.01202f
C929 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C CLK 0.19664f
C930 a_38699_61411# Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.01335f
C931 a_10187_59439# VDD 0.05686f
C932 a_8706_48405# VDD 0.02521f
C933 a_10187_55365# VDD 0.0563f
C934 a_n505_58825# VDD 0.02578f
C935 a_3059_56723# VDD 0.02578f
C936 D_FlipFlop_5.nPRE D_FlipFlop_5.3-input-nand_1.Vout 0.06632f
C937 Ring_Counter_0.D_FlipFlop_2.Qbar VDD 1.99882f
C938 D_FlipFlop_2.nPRE And_Gate_5.Nand_Gate_0.Vout 0.12031f
C939 D_FlipFlop_6.CLK D_FlipFlop_6.3-input-nand_1.B 0.06986f
C940 a_2209_59439# EN 0.045f
C941 a_n11757_52049# VDD 0.02693f
C942 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout a_31571_59439# 0.04543f
C943 a_56590_51119# Q7 0.06113f
C944 D_FlipFlop_2.CLK a_34378_48405# 0.02953f
C945 CDAC_v3_0.OUT m3_3428_33935# 1.25228f
C946 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.08674f
C947 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.01162f
C948 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.0646f
C949 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.06462f
C950 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C a_17315_56723# 0.04443f
C951 Ring_Counter_0.D_FlipFlop_16.Q a_37849_61411# 0.01252f
C952 a_6623_55365# VDD 0.0563f
C953 CDAC_v3_0.switch_0.Z a_31486_45397# 0.022f
C954 D_FlipFlop_1.nPRE D_FlipFlop_1.Inverter_1.Vout 0.07033f
C955 a_6623_58825# Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.05964f
C956 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout 0.25855f
C957 D_FlipFlop_6.CLK a_n56_48405# 0.02953f
C958 Nand_Gate_4.A a_30721_56723# 0.05925f
C959 Ring_Counter_0.D_FlipFlop_3.Qbar VDD 2.00188f
C960 a_6623_61411# a_6623_60797# 0.05935f
C961 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout a_5773_60797# 0.05964f
C962 a_10187_60797# VDD 0.02865f
C963 a_15710_45397# VDD 1.17814f
C964 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout a_n7633_56723# 0.04995f
C965 D_FlipFlop_1.3-input-nand_1.B D_FlipFlop_1.3-input-nand_1.Vout 0.08641f
C966 D_FlipFlop_3.nPRE And_Gate_4.Nand_Gate_0.Vout 0.12031f
C967 D_FlipFlop_3.Inverter_1.Vout Q5 0.01387f
C968 D_FlipFlop_7.Qbar a_n4744_48405# 0.06113f
C969 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.01194f
C970 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.01194f
C971 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.15413f
C972 D_FlipFlop_2.nPRE a_34378_51119# 0.045f
C973 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_n505_55365# 0.04995f
C974 a_8706_51119# D_FlipFlop_4.3-input-nand_2.Vout 0.05964f
C975 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_24443_54751# 0.04444f
C976 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_n1355_55365# 0.04995f
C977 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.08462f
C978 a_16465_59439# a_16465_58825# 0.05935f
C979 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_0.Qbar 0.11657f
C980 a_4018_51119# VDD 0.02521f
C981 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_23593_54751# 0.04444f
C982 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.10034f
C983 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout a_5773_59439# 0.04995f
C984 And_Gate_3.A And_Gate_3.Nand_Gate_0.Vout 0.24482f
C985 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout EN 0.06639f
C986 a_3059_55365# VDD 0.0563f
C987 a_n8818_51119# VDD 0.02521f
C988 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.1143f
C989 D_FlipFlop_6.CLK D_FlipFlop_6.3-input-nand_2.C 0.19377f
C990 D_FlipFlop_1.3-input-nand_1.Vout VDD 1.76485f
C991 a_9337_60797# CLK 0.06211f
C992 D_FlipFlop_2.3-input-nand_1.Vout a_34378_48405# 0.04543f
C993 D_FlipFlop_7.nPRE a_n5358_51119# 0.04443f
C994 Ring_Counter_0.D_FlipFlop_4.Qbar VDD 2.00088f
C995 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.Nand_Gate_1.Vout 0.1541f
C996 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.16431f
C997 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.01323f
C998 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout a_2209_59439# 0.01335f
C999 D_FlipFlop_3.Qbar a_30304_51119# 0.04443f
C1000 D_FlipFlop_5.nPRE And_Gate_3.Nand_Gate_0.Vout 0.12031f
C1001 D_FlipFlop_0.CLK Q7 0.05341f
C1002 a_35135_60797# VDD 0.02865f
C1003 a_16465_61411# a_16465_60797# 0.05935f
C1004 Nand_Gate_4.A D_FlipFlop_2.nPRE 2.51364f
C1005 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.04109f
C1006 a_n4069_59439# a_n4069_58825# 0.05935f
C1007 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B a_42263_61411# 0.04995f
C1008 a_23644_51119# a_24258_51119# 0.05935f
C1009 a_n505_55365# VDD 0.0563f
C1010 D_FlipFlop_5.3-input-nand_2.C a_17468_51119# 0.04443f
C1011 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B 0.29684f
C1012 Nand_Gate_3.A a_27157_55365# 0.0139f
C1013 a_49930_48405# a_50544_48405# 0.05935f
C1014 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_1.Vout 0.08671f
C1015 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout EN 0.09223f
C1016 D_FlipFlop_1.CLK CLK 0.07954f
C1017 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout a_13751_58825# 0.04444f
C1018 Ring_Counter_0.D_FlipFlop_5.Qbar VDD 2.00117f
C1019 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout EN 0.96763f
C1020 a_52516_51119# D_FlipFlop_0.3-input-nand_2.Vout 0.05964f
C1021 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout CLK 0.20785f
C1022 a_12901_61411# EN 0.02636f
C1023 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B EN 0.3979f
C1024 And_Gate_3.A a_14529_52049# 0.04995f
C1025 Nand_Gate_5.A a_37849_59439# 0.05925f
C1026 a_49930_51119# VDD 0.01186f
C1027 a_34285_60797# CLK 0.06211f
C1028 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B a_3059_60797# 0.04443f
C1029 Nand_Gate_6.A a_20029_54751# 0.06113f
C1030 a_28332_48405# VDD 0.02521f
C1031 Ring_Counter_0.D_FlipFlop_16.Q a_3059_60797# 0.01768f
C1032 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C a_n4919_58825# 0.04443f
C1033 a_31571_61411# a_31571_60797# 0.05935f
C1034 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout a_30721_60797# 0.05964f
C1035 a_n4069_55365# VDD 0.0563f
C1036 D_FlipFlop_5.nPRE a_14529_52049# 0.02193f
C1037 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD 1.45175f
C1038 a_54330_52049# VDD 0.02521f
C1039 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout CLK 0.21133f
C1040 Nand_Gate_3.A a_23593_55365# 0.05925f
C1041 D_FlipFlop_4.3-input-nand_1.B D_FlipFlop_4.3-input-nand_1.Vout 0.08641f
C1042 Ring_Counter_0.D_FlipFlop_6.Qbar VDD 1.99776f
C1043 Nand_Gate_6.A a_16465_54751# 0.05925f
C1044 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout EN 0.09223f
C1045 CDAC_v3_0.switch_0.Z Q2 0.02962f
C1046 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout EN 0.96763f
C1047 CDAC_v3_0.switch_5.Z CDAC_v3_0.OUT 0.14574p
C1048 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.08674f
C1049 a_37849_61411# EN 0.02636f
C1050 D_FlipFlop_7.3-input-nand_1.Vout a_n10790_48405# 0.05964f
C1051 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.06935f
C1052 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_1.Vout 0.67481f
C1053 CDAC_v3_0.OUT VDD 0.1543f
C1054 Ring_Counter_0.D_FlipFlop_16.Q a_28007_60797# 0.01768f
C1055 a_n7633_55365# VDD 0.0563f
C1056 D_FlipFlop_0.3-input-nand_2.C a_52516_48405# 0.05964f
C1057 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_31571_55365# 0.04995f
C1058 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_30721_55365# 0.04995f
C1059 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.25966f
C1060 Ring_Counter_0.D_FlipFlop_7.Qbar VDD 1.99815f
C1061 a_41413_61411# a_41413_60797# 0.05935f
C1062 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.04107f
C1063 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout a_23593_56723# 0.04443f
C1064 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout EN 0.61231f
C1065 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout a_n1355_61411# 0.01335f
C1066 a_n4069_61411# VDD 0.04448f
C1067 a_32406_48405# a_33020_48405# 0.05935f
C1068 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.08462f
C1069 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.Qbar 1.27275f
C1070 VDD Q3 3.54595f
C1071 D_FlipFlop_3.nPRE a_23644_51119# 0.034f
C1072 a_9337_56723# VDD 0.02521f
C1073 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout a_41413_59439# 0.04995f
C1074 a_n6716_48405# VDD 0.02521f
C1075 D_FlipFlop_6.CLK D_FlipFlop_6.3-input-nand_0.Vout 0.25957f
C1076 D_FlipFlop_2.Nand_Gate_1.Vout VDD 1.44304f
C1077 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.06955f
C1078 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_12901_56723# 0.05964f
C1079 a_42263_58825# Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.04443f
C1080 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.01202f
C1081 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_1.Vout 0.08671f
C1082 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.20928f
C1083 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout CLK 0.7779f
C1084 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout CLK 0.36346f
C1085 D_FlipFlop_3.Nand_Gate_0.Vout a_30304_51119# 0.04444f
C1086 Ring_Counter_0.D_FlipFlop_8.Qbar VDD 2.00026f
C1087 a_47828_48405# Q6 0.05747f
C1088 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C a_52105_58825# 0.04443f
C1089 Nand_Gate_2.A a_12901_54751# 0.06113f
C1090 a_49391_59439# EN 0.045f
C1091 D_FlipFlop_3.nPRE D_FlipFlop_3.3-input-nand_1.Vout 0.06632f
C1092 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.01194f
C1093 a_n7633_56723# Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.05964f
C1094 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.Qbar 0.12029f
C1095 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout a_9337_56723# 0.04443f
C1096 D_FlipFlop_6.nPRE a_n2642_51119# 0.034f
C1097 a_20879_61411# VDD 0.04448f
C1098 a_45827_59439# Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.01335f
C1099 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.25966f
C1100 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.06837f
C1101 D_FlipFlop_5.3-input-nand_0.Vout a_17468_51119# 0.04444f
C1102 a_19570_51119# VDD 0.02521f
C1103 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.06863f
C1104 And_Gate_5.Nand_Gate_0.Vout CLK 0.79128f
C1105 And_Gate_6.Nand_Gate_0.Vout D_FlipFlop_1.CLK 0.25559f
C1106 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout EN 0.78583f
C1107 a_47214_48405# VDD 0.01186f
C1108 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout a_49391_58825# 0.04444f
C1109 D_FlipFlop_0.3-input-nand_1.B VDD 1.2956f
C1110 D_FlipFlop_6.CLK D_FlipFlop_6.3-input-nand_1.Vout 0.67419f
C1111 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout VDD 2.07898f
C1112 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 1.09973f
C1113 Ring_Counter_0.D_FlipFlop_9.Qbar VDD 1.9996f
C1114 a_45827_58825# CLK 0.03f
C1115 a_6734_51119# VDD 0.02521f
C1116 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout CLK 0.7779f
C1117 Nand_Gate_2.A a_9337_58825# 0.05925f
C1118 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout CLK 0.36346f
C1119 Nand_Gate_2.A a_9337_54751# 0.05925f
C1120 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout CLK 0.12427f
C1121 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.04109f
C1122 D_FlipFlop_2.3-input-nand_2.Vout VDD 2.67108f
C1123 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.01162f
C1124 a_14882_48405# a_15496_48405# 0.05935f
C1125 D_FlipFlop_6.Qbar a_4018_48405# 0.06113f
C1126 D_FlipFlop_2.Nand_Gate_1.Vout a_37094_48405# 0.05964f
C1127 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B 0.02535f
C1128 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.04107f
C1129 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout a_23593_61411# 0.01335f
C1130 a_45827_61411# VDD 0.04448f
C1131 D_FlipFlop_4.Nand_Gate_1.Vout a_12780_48405# 0.04444f
C1132 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C EN 0.07565f
C1133 D_FlipFlop_2.CLK VDD 2.17782f
C1134 a_52105_59439# VDD 0.05686f
C1135 Ring_Counter_0.D_FlipFlop_10.Qbar VDD 2.00254f
C1136 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout a_23593_58825# 0.04444f
C1137 D_FlipFlop_1.Inverter_1.Vout Q7 0.02777f
C1138 a_41413_58825# VDD 0.02521f
C1139 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.01323f
C1140 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout a_30721_58825# 0.05964f
C1141 D_FlipFlop_6.Inverter_1.Vout a_2046_51119# 0.04443f
C1142 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C CLK 0.19664f
C1143 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_10.Qbar 0.07122f
C1144 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.10034f
C1145 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout CLK 0.7779f
C1146 a_31571_59439# VDD 0.05686f
C1147 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK 0.36346f
C1148 Nand_Gate_0.A a_2209_56723# 0.05925f
C1149 D_FlipFlop_4.nPRE D_FlipFlop_4.3-input-nand_1.Vout 0.06632f
C1150 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout CLK 0.2743f
C1151 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.48403f
C1152 Ring_Counter_0.D_FlipFlop_16.Q a_13751_61411# 0.01252f
C1153 a_20879_58825# VDD 0.02578f
C1154 D_FlipFlop_0.3-input-nand_2.C VDD 2.73475f
C1155 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C a_45827_56723# 0.04443f
C1156 And_Gate_2.A a_5767_52049# 0.04995f
C1157 D_FlipFlop_1.CLK D_FlipFlop_1.Inverter_1.Vout 0.20785f
C1158 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.Inverter_1.Vout 0.06895f
C1159 a_23593_59439# EN 0.045f
C1160 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.01194f
C1161 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout VDD 2.8343f
C1162 Ring_Counter_0.D_FlipFlop_11.Qbar VDD 2.00063f
C1163 a_12166_48405# VDD 0.01186f
C1164 D_FlipFlop_3.nPRE D_FlipFlop_3.3-input-nand_1.B 0.27142f
C1165 D_FlipFlop_7.Inverter_1.Vout VDD 1.70303f
C1166 Nand_Gate_4.A CLK 0.52614f
C1167 D_FlipFlop_3.nPRE a_27157_59439# 0.05925f
C1168 Nand_Gate_0.A a_5773_54751# 0.06113f
C1169 D_FlipFlop_2.3-input-nand_1.Vout VDD 1.76485f
C1170 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.15413f
C1171 D_FlipFlop_1.nPRE Q7 0.01779f
C1172 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.26069f
C1173 D_FlipFlop_3.CLK a_24258_51119# 0.04443f
C1174 a_n2642_48405# a_n2028_48405# 0.05935f
C1175 a_n2995_52049# VDD 0.02521f
C1176 D_FlipFlop_5.nPRE D_FlipFlop_4.Qbar 0.01961f
C1177 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.06955f
C1178 a_n6716_51119# D_FlipFlop_7.Nand_Gate_0.Vout 0.05964f
C1179 a_17315_58825# Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.05964f
C1180 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B 0.02535f
C1181 CDAC_v3_0.OUT m3_3428_4751# 1.25228f
C1182 a_10187_59439# CLK 0.03166f
C1183 D_FlipFlop_1.Inverter_1.Vout a_45856_51119# 0.04443f
C1184 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C1185 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C VDD 3.50703f
C1186 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.01194f
C1187 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B VDD 1.74109f
C1188 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.01194f
C1189 Ring_Counter_0.D_FlipFlop_16.Q a_38699_61411# 0.01252f
C1190 Ring_Counter_0.D_FlipFlop_12.Qbar VDD 1.99817f
C1191 a_n505_58825# CLK 0.03f
C1192 D_FlipFlop_1.nPRE D_FlipFlop_1.CLK 0.16746f
C1193 a_23598_45397# CDAC_v3_0.switch_4.Z 0.27028f
C1194 CDAC_v3_0.switch_0.Z a_35430_45397# 0.02212f
C1195 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.Nand_Gate_0.Vout 0.16429f
C1196 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.26069f
C1197 a_27157_59439# a_27157_58825# 0.05935f
C1198 D_FlipFlop_6.nPRE D_FlipFlop_6.3-input-nand_1.B 0.27142f
C1199 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.04107f
C1200 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B 0.02535f
C1201 Nand_Gate_0.A a_2209_54751# 0.05957f
C1202 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.Inverter_1.Vout 0.26069f
C1203 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.16431f
C1204 a_16854_51119# D_FlipFlop_5.3-input-nand_2.Vout 0.01335f
C1205 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.17188f
C1206 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout a_48541_61411# 0.01335f
C1207 a_6623_60797# Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.05964f
C1208 a_n11757_52049# CLK 0.04443f
C1209 a_20928_51119# VDD 0.01186f
C1210 a_19654_45397# VDD 1.17814f
C1211 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.Inverter_1.Vout 0.06935f
C1212 CDAC_v3_0.switch_6.Z Q7 0.17554f
C1213 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_37849_56723# 0.05964f
C1214 a_5773_60797# VDD 0.02521f
C1215 D_FlipFlop_2.nPRE D_FlipFlop_2.3-input-nand_2.Vout 0.76528f
C1216 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.07084f
C1217 a_8092_51119# VDD 0.01186f
C1218 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_14.Qbar 0.11657f
C1219 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout a_6623_59439# 0.04543f
C1220 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.26069f
C1221 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C1222 a_5773_59439# VDD 0.01186f
C1223 D_FlipFlop_3.nPRE D_FlipFlop_3.3-input-nand_2.C 0.05823f
C1224 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout a_12901_59439# 0.01335f
C1225 Ring_Counter_0.D_FlipFlop_13.Qbar VDD 1.99978f
C1226 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.06837f
C1227 a_17315_56723# Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.05964f
C1228 D_FlipFlop_2.nPRE D_FlipFlop_2.CLK 0.1668f
C1229 D_FlipFlop_6.nPRE a_5773_56723# 0.05925f
C1230 a_37094_51119# D_FlipFlop_2.Nand_Gate_0.Vout 0.05964f
C1231 a_10187_60797# CLK 0.06211f
C1232 a_6623_59439# a_6623_58825# 0.05935f
C1233 a_n4919_58825# VDD 0.02521f
C1234 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.09856f
C1235 D_FlipFlop_4.nPRE a_12901_61411# 0.04995f
C1236 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B a_31571_60797# 0.04443f
C1237 D_FlipFlop_7.3-input-nand_1.B a_n11404_48405# 0.04995f
C1238 And_Gate_4.Nand_Gate_0.Vout VDD 1.39123f
C1239 D_FlipFlop_1.nPRE a_45568_52049# 0.04443f
C1240 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.Nand_Gate_0.Vout 0.16429f
C1241 a_n4069_58825# Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.04443f
C1242 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B a_20879_60797# 0.04443f
C1243 a_30721_60797# VDD 0.02521f
C1244 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.08582f
C1245 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_1.Qbar 0.07122f
C1246 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B 0.02535f
C1247 a_24258_51119# D_FlipFlop_3.3-input-nand_0.Vout 0.05964f
C1248 D_FlipFlop_6.nPRE D_FlipFlop_6.3-input-nand_2.C 0.05823f
C1249 Ring_Counter_0.D_FlipFlop_14.Qbar VDD 2.00097f
C1250 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C1251 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.04109f
C1252 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C a_5773_58825# 0.04443f
C1253 D_FlipFlop_3.nPRE D_FlipFlop_3.CLK 0.1668f
C1254 Nand_Gate_1.A a_n1355_54751# 0.06113f
C1255 a_13751_61411# EN 0.07048f
C1256 D_FlipFlop_0.3-input-nand_0.Vout VDD 1.77947f
C1257 a_35135_56723# VDD 0.02578f
C1258 a_35135_60797# CLK 0.06211f
C1259 a_n505_59439# Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.01335f
C1260 a_30304_48405# VDD 0.02521f
C1261 D_FlipFlop_2.nPRE D_FlipFlop_2.3-input-nand_1.Vout 0.06632f
C1262 Ring_Counter_0.D_FlipFlop_16.Q a_n1355_60797# 0.01768f
C1263 And_Gate_3.A D_FlipFlop_5.CLK 0.06897f
C1264 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout EN 0.61231f
C1265 a_31571_60797# Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.05964f
C1266 Nand_Gate_5.A VDD 4.5982f
C1267 Ring_Counter_0.D_FlipFlop_15.Qbar VDD 2.00272f
C1268 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.Q 0.26977f
C1269 D_FlipFlop_3.Nand_Gate_1.Vout VDD 1.44304f
C1270 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout a_52105_56723# 0.04443f
C1271 D_FlipFlop_7.Nand_Gate_0.Vout a_n5358_51119# 0.04543f
C1272 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1273 D_FlipFlop_1.CLK a_41782_48405# 0.04443f
C1274 D_FlipFlop_5.3-input-nand_1.Vout a_15496_48405# 0.05964f
C1275 Nand_Gate_1.A a_n4919_54751# 0.06171f
C1276 D_FlipFlop_5.nPRE D_FlipFlop_5.CLK 0.1668f
C1277 Nand_Gate_6.A a_17315_54751# 0.05987f
C1278 Nand_Gate_6.A EN 0.79742f
C1279 CDAC_v3_0.switch_2.Z Q2 0.17946f
C1280 CDAC_v3_0.switch_7.Z CDAC_v3_0.OUT 0.28889p
C1281 D_FlipFlop_6.Nand_Gate_1.Vout Q1 0.09808f
C1282 D_FlipFlop_4.Qbar a_12780_48405# 0.06113f
C1283 D_FlipFlop_7.3-input-nand_1.Vout a_n8818_48405# 0.04444f
C1284 a_38699_61411# EN 0.07048f
C1285 a_30304_48405# Q4 0.05747f
C1286 D_FlipFlop_4.CLK a_8092_48405# 0.02953f
C1287 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B 0.02535f
C1288 Ring_Counter_0.D_FlipFlop_16.Qbar VDD 1.96531f
C1289 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout 0.30046f
C1290 Ring_Counter_0.D_FlipFlop_16.Q a_23593_60797# 0.01768f
C1291 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C a_6623_56723# 0.04443f
C1292 And_Gate_7.A And_Gate_7.Nand_Gate_0.Vout 0.26587f
C1293 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_6623_54751# 0.04444f
C1294 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_5.Qbar 0.11657f
C1295 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_5773_54751# 0.04444f
C1296 D_FlipFlop_4.nPRE D_FlipFlop_4.Nand_Gate_0.Vout 0.5831f
C1297 D_FlipFlop_3.Nand_Gate_1.Vout Q4 0.09956f
C1298 a_n505_61411# Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.01335f
C1299 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout VDD 2.72531f
C1300 And_Gate_1.A a_n2995_52049# 0.04995f
C1301 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD 1.87537f
C1302 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.01262f
C1303 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.29165f
C1304 Nand_Gate_2.A EN 0.79742f
C1305 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout a_42263_59439# 0.04543f
C1306 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.15413f
C1307 D_FlipFlop_3.nPRE D_FlipFlop_3.3-input-nand_0.Vout 0.94459f
C1308 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout VDD 2.07898f
C1309 a_n4744_48405# VDD 0.02521f
C1310 Nand_Gate_4.A a_34285_55365# 0.0139f
C1311 Nand_Gate_1.A a_n4919_60797# 0.10368f
C1312 D_FlipFlop_1.nPRE a_47214_51119# 0.04443f
C1313 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.08674f
C1314 D_FlipFlop_2.Nand_Gate_0.Vout a_38452_51119# 0.04543f
C1315 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.01202f
C1316 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.10915f
C1317 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.01202f
C1318 D_FlipFlop_0.Nand_Gate_1.Vout Q7 0.13061f
C1319 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B a_6623_60797# 0.04443f
C1320 And_Gate_7.A VDD 1.45624f
C1321 Ring_Counter_0.D_FlipFlop_16.Q a_48541_60797# 0.01768f
C1322 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout EN 0.08727f
C1323 D_FlipFlop_3.3-input-nand_0.Vout a_25616_51119# 0.04543f
C1324 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.06837f
C1325 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.16431f
C1326 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout EN 0.0649f
C1327 Nand_Gate_0.A EN 0.79742f
C1328 D_FlipFlop_6.nPRE D_FlipFlop_6.3-input-nand_0.Vout 0.94459f
C1329 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 1.09973f
C1330 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.09856f
C1331 Nand_Gate_4.A a_30721_55365# 0.05925f
C1332 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout VDD 2.72531f
C1333 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_0.Z 7.19346f
C1334 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD 1.89599f
C1335 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.08462f
C1336 a_16465_61411# VDD 0.08862f
C1337 a_42263_56723# Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.05964f
C1338 a_23644_51119# VDD 0.01186f
C1339 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout a_16465_59439# 0.04995f
C1340 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout 0.26069f
C1341 a_49930_48405# VDD 0.01205f
C1342 a_52516_51119# VDD 0.02521f
C1343 D_FlipFlop_2.nPRE Nand_Gate_5.A 0.04143f
C1344 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.48403f
C1345 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.06734f
C1346 Nand_Gate_2.A a_10187_54751# 0.05987f
C1347 Nand_Gate_4.A a_36806_52049# 0.0451f
C1348 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C EN 0.07565f
C1349 D_FlipFlop_6.CLK D_FlipFlop_6.Inverter_1.Vout 0.20785f
C1350 Nand_Gate_1.A EN 0.79742f
C1351 D_FlipFlop_2.Nand_Gate_1.Vout a_39066_48405# 0.04444f
C1352 D_FlipFlop_3.3-input-nand_1.Vout VDD 1.76485f
C1353 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout 0.30046f
C1354 a_n5358_51119# a_n4744_51119# 0.05935f
C1355 a_24443_61411# Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.01335f
C1356 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B EN 0.3979f
C1357 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout a_41413_58825# 0.05964f
C1358 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout VDD 2.72531f
C1359 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_1.B 0.06986f
C1360 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B 0.02535f
C1361 D_FlipFlop_6.nPRE D_FlipFlop_6.3-input-nand_1.Vout 0.06632f
C1362 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD 1.89599f
C1363 Ring_Counter_0.D_FlipFlop_9.Qbar CLK 0.07015f
C1364 a_41413_61411# VDD 0.08862f
C1365 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.Qbar 1.27332f
C1366 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout VDD 2.26641f
C1367 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.11774f
C1368 D_FlipFlop_4.nPRE a_12901_58825# 0.05925f
C1369 D_FlipFlop_1.CLK Q7 0.05341f
C1370 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout a_24443_58825# 0.04444f
C1371 D_FlipFlop_5.nPRE Q2 0.01495f
C1372 a_42263_58825# VDD 0.02578f
C1373 a_44977_59439# EN 0.045f
C1374 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.30156f
C1375 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_13751_55365# 0.04995f
C1376 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_38699_54751# 0.04444f
C1377 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_12901_55365# 0.04995f
C1378 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout VDD 2.8343f
C1379 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_37849_54751# 0.04444f
C1380 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.10915f
C1381 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.16917f
C1382 D_FlipFlop_6.3-input-nand_1.B a_n2642_48405# 0.04995f
C1383 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.01262f
C1384 a_41413_56723# VDD 0.02521f
C1385 D_FlipFlop_2.CLK CLK 0.07954f
C1386 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.29165f
C1387 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.0646f
C1388 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.06462f
C1389 D_FlipFlop_3.3-input-nand_1.Vout Q4 0.01372f
C1390 Ring_Counter_0.D_FlipFlop_16.Q a_9337_61411# 0.01252f
C1391 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.Qbar 0.11848f
C1392 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout a_20879_56723# 0.04995f
C1393 a_14882_48405# VDD 0.01186f
C1394 D_FlipFlop_4.nPRE And_Gate_2.Nand_Gate_0.Vout 0.12031f
C1395 D_FlipFlop_4.nPRE Q2 0.03683f
C1396 a_n7633_61411# a_n7633_60797# 0.05935f
C1397 a_28007_58825# Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.05964f
C1398 a_31571_59439# CLK 0.03166f
C1399 a_38452_51119# a_39066_51119# 0.05935f
C1400 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout a_12901_56723# 0.04443f
C1401 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout a_n1355_58825# 0.04444f
C1402 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout EN 0.78583f
C1403 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.01194f
C1404 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C VDD 3.50703f
C1405 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.01194f
C1406 D_FlipFlop_0.3-input-nand_1.Vout Q7 0.02726f
C1407 a_20879_58825# CLK 0.03057f
C1408 a_5767_52049# VDD 0.02521f
C1409 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_2.C 0.19377f
C1410 a_49391_55365# Ring_Counter_0.D_FlipFlop_0.Qbar 0.01335f
C1411 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout a_27157_56723# 0.04443f
C1412 a_37849_59439# a_37849_58825# 0.05935f
C1413 D_FlipFlop_1.nPRE D_FlipFlop_1.3-input-nand_1.Vout 0.06632f
C1414 D_FlipFlop_4.3-input-nand_2.Vout a_10808_51119# 0.04443f
C1415 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout CLK 0.12427f
C1416 a_n11404_51119# D_FlipFlop_7.3-input-nand_0.Vout 0.01335f
C1417 Nand_Gate_1.A a_n7004_52049# 0.04443f
C1418 a_25616_51119# a_26230_51119# 0.05935f
C1419 D_FlipFlop_7.Nand_Gate_1.Vout a_n5358_48405# 0.04995f
C1420 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.06734f
C1421 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.0646f
C1422 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.06462f
C1423 D_FlipFlop_6.nPRE And_Gate_2.Nand_Gate_0.Vout 0.01462f
C1424 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.06837f
C1425 Ring_Counter_0.D_FlipFlop_16.Q a_34285_61411# 0.01252f
C1426 a_n6716_51119# VDD 0.02521f
C1427 a_49391_61411# Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout 0.01335f
C1428 Nand_Gate_5.A a_37849_60797# 0.10368f
C1429 Nand_Gate_0.A a_3059_54751# 0.05987f
C1430 a_n2995_52049# CLK 0.04479f
C1431 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.20923f
C1432 D_FlipFlop_3.3-input-nand_1.B VDD 1.34831f
C1433 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C EN 0.07565f
C1434 a_23598_45397# VDD 1.17814f
C1435 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout a_35135_56723# 0.04995f
C1436 a_27157_59439# VDD 0.01186f
C1437 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout a_23593_59439# 0.01335f
C1438 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.01202f
C1439 a_6623_60797# VDD 0.02865f
C1440 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout a_52105_59439# 0.04995f
C1441 D_FlipFlop_5.Qbar a_21542_48405# 0.06113f
C1442 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.01323f
C1443 a_2209_61411# a_2209_60797# 0.05935f
C1444 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.1143f
C1445 D_FlipFlop_4.3-input-nand_2.Vout VDD 2.67107f
C1446 a_17315_59439# a_17315_58825# 0.05935f
C1447 a_16465_58825# VDD 0.02521f
C1448 D_FlipFlop_3.nPRE a_27157_60797# 0.10368f
C1449 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.06837f
C1450 Nand_Gate_6.A And_Gate_3.A 0.0808f
C1451 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.06955f
C1452 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C CLK 0.19664f
C1453 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B CLK 0.08407f
C1454 And_Gate_0.A a_n11757_52049# 0.04995f
C1455 a_17315_56723# VDD 0.02578f
C1456 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout 0.09856f
C1457 a_6623_59439# VDD 0.05686f
C1458 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.17551f
C1459 a_6623_58825# Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.04443f
C1460 a_n4069_58825# VDD 0.02578f
C1461 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout a_41413_56723# 0.04443f
C1462 D_FlipFlop_5.Nand_Gate_1.Vout VDD 1.44333f
C1463 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout EN 0.61231f
C1464 a_5773_60797# CLK 0.06211f
C1465 D_FlipFlop_0.3-input-nand_2.Vout a_54618_51119# 0.04443f
C1466 a_n1355_59439# EN 0.045f
C1467 CDAC_v3_0.OUT Vbias 1.07744f
C1468 Nand_Gate_6.A D_FlipFlop_5.nPRE 1.14848f
C1469 a_32406_51119# D_FlipFlop_2.3-input-nand_0.Vout 0.01335f
C1470 Nand_Gate_1.A a_n4919_59439# 0.05925f
C1471 a_23598_45397# Q4 0.46608f
C1472 a_45827_55365# Ring_Counter_0.D_FlipFlop_1.Qbar 0.01335f
C1473 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C a_16465_58825# 0.04443f
C1474 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_15.Qbar 0.07122f
C1475 a_17315_61411# a_17315_60797# 0.05935f
C1476 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.Vout 1.01753f
C1477 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.10915f
C1478 a_31571_60797# VDD 0.02865f
C1479 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout a_16465_60797# 0.05964f
C1480 D_FlipFlop_2.Qbar VDD 1.96371f
C1481 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.07084f
C1482 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_45827_55365# 0.04995f
C1483 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_n4919_56723# 0.05964f
C1484 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_44977_55365# 0.04995f
C1485 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout a_49391_56723# 0.04995f
C1486 a_10187_59439# Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.01335f
C1487 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B a_n7633_61411# 0.04975f
C1488 D_FlipFlop_3.3-input-nand_2.C VDD 2.6783f
C1489 a_12780_48405# Q2 0.05747f
C1490 a_51902_48405# a_52516_48405# 0.05935f
C1491 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.09856f
C1492 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout EN 0.09223f
C1493 D_FlipFlop_4.nPRE Nand_Gate_6.A 0.04143f
C1494 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout EN 0.96763f
C1495 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.01162f
C1496 And_Gate_4.Nand_Gate_0.Vout CLK 0.79128f
C1497 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 1.09973f
C1498 a_9337_61411# EN 0.02636f
C1499 a_33020_48405# VDD 0.02521f
C1500 a_30721_60797# CLK 0.06211f
C1501 Ring_Counter_0.D_FlipFlop_16.Q a_n505_60797# 0.01768f
C1502 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C a_35135_56723# 0.04443f
C1503 D_FlipFlop_1.3-input-nand_1.Vout a_41782_48405# 0.05964f
C1504 D_FlipFlop_3.CLK D_FlipFlop_3.3-input-nand_2.Vout 0.1192f
C1505 a_27157_61411# a_27157_60797# 0.05935f
C1506 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout VDD 2.04725f
C1507 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.Qbar 1.29337f
C1508 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout a_34285_58825# 0.04444f
C1509 D_FlipFlop_1.Nand_Gate_1.Vout Q7 0.02995f
C1510 D_FlipFlop_0.CLK D_FlipFlop_0.3-input-nand_0.Vout 0.25974f
C1511 D_FlipFlop_5.3-input-nand_1.Vout a_17468_48405# 0.04444f
C1512 D_FlipFlop_1.CLK a_43754_48405# 0.02953f
C1513 Nand_Gate_1.A a_n4069_54751# 0.06233f
C1514 D_FlipFlop_3.3-input-nand_2.C Q4 0.01368f
C1515 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout VDD 2.29929f
C1516 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.04109f
C1517 D_FlipFlop_7.3-input-nand_2.C a_n9432_48405# 0.01335f
C1518 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.10034f
C1519 Nand_Gate_2.A D_FlipFlop_4.nPRE 0.28905f
C1520 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.15413f
C1521 D_FlipFlop_3.CLK VDD 2.17842f
C1522 CDAC_v3_0.switch_6.Z CDAC_v3_0.OUT 0.57904p
C1523 a_42263_55365# Ring_Counter_0.D_FlipFlop_2.Qbar 0.01335f
C1524 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout EN 0.09223f
C1525 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout EN 0.96763f
C1526 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout a_n4919_58825# 0.05964f
C1527 Nand_Gate_5.A CLK 0.52845f
C1528 a_n5358_51119# VDD 0.01186f
C1529 a_34285_61411# EN 0.02636f
C1530 Ring_Counter_0.D_FlipFlop_16.Q a_24443_60797# 0.01768f
C1531 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.Qbar 0.11806f
C1532 D_FlipFlop_0.Inverter_1.Vout VDD 1.73165f
C1533 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.30156f
C1534 a_42263_61411# a_42263_60797# 0.05935f
C1535 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.01202f
C1536 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout a_41413_60797# 0.05964f
C1537 a_34378_48405# a_34992_48405# 0.05935f
C1538 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.16431f
C1539 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.01194f
C1540 D_FlipFlop_6.nPRE Nand_Gate_2.A 0.04125f
C1541 a_n7633_61411# VDD 0.09865f
C1542 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.06955f
C1543 a_n2028_48405# VDD 0.02521f
C1544 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Qbar 0.06863f
C1545 D_FlipFlop_3.CLK Q4 0.03348f
C1546 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD 1.48403f
C1547 D_FlipFlop_4.3-input-nand_1.B a_6120_48405# 0.04995f
C1548 And_Gate_1.Nand_Gate_0.Vout D_FlipFlop_6.CLK 0.25559f
C1549 D_FlipFlop_5.3-input-nand_1.Vout VDD 1.76541f
C1550 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.01202f
C1551 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_6.Qbar 0.07122f
C1552 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout CLK 0.7779f
C1553 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout CLK 0.36238f
C1554 Ring_Counter_0.D_FlipFlop_16.Q a_49391_60797# 0.01768f
C1555 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.3-input-nand_2.C 0.06863f
C1556 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.09856f
C1557 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.09856f
C1558 CDAC_v3_0.switch_5.Z m3_3428_38799# 1.89962f
C1559 D_FlipFlop_6.3-input-nand_1.Vout a_n2642_48405# 0.01335f
C1560 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.3-input-nand_2.Vout 0.0846f
C1561 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout a_13751_56723# 0.04995f
C1562 D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.43587f
C1563 a_38699_55365# Ring_Counter_0.D_FlipFlop_3.Qbar 0.01335f
C1564 Nand_Gate_0.A D_FlipFlop_6.nPRE 1.10458f
C1565 D_FlipFlop_4.CLK D_FlipFlop_4.3-input-nand_1.B 0.06986f
C1566 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.25966f
C1567 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.07084f
C1568 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.04107f
C1569 a_52105_61411# a_52105_60797# 0.05935f
C1570 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_2.Z 23.4364f
C1571 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.30156f
C1572 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout a_17315_59439# 0.04543f
C1573 a_17315_61411# VDD 0.04448f
C1574 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout a_9337_61411# 0.01335f
C1575 D_FlipFlop_3.3-input-nand_0.Vout VDD 1.74442f
C1576 And_Gate_7.A CLK 0.34279f
C1577 And_Gate_7.A D_FlipFlop_0.CLK 0.07237f
C1578 D_FlipFlop_1.nPRE a_41413_58825# 0.05925f
C1579 a_51902_48405# VDD 0.01186f
C1580 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.08674f
C1581 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.01323f
C1582 D_FlipFlop_7.nPRE D_FlipFlop_7.3-input-nand_1.Vout 0.06632f
C1583 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Qbar 0.06863f
C1584 a_23593_56723# VDD 0.02521f
C1585 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout a_52105_58825# 0.05964f
C1586 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.11436f
C1587 D_FlipFlop_3.nPRE D_FlipFlop_3.Inverter_1.Vout 0.07033f
C1588 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout CLK 0.78138f
C1589 a_16854_48405# a_17468_48405# 0.05935f
C1590 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout CLK 0.46165f
C1591 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_20029_56723# 0.05964f
C1592 D_FlipFlop_7.nPRE Nand_Gate_0.A 0.04305f
C1593 Nand_Gate_1.A D_FlipFlop_6.nPRE 0.03898f
C1594 D_FlipFlop_3.Qbar a_30304_48405# 0.06113f
C1595 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B a_35135_61411# 0.04995f
C1596 D_FlipFlop_5.nPRE a_16854_51119# 0.045f
C1597 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B a_10187_61411# 0.04995f
C1598 D_FlipFlop_1.3-input-nand_1.Vout Q7 0.02726f
C1599 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.3-input-nand_2.C 0.06863f
C1600 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.01194f
C1601 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.08462f
C1602 Nand_Gate_6.A a_16465_59439# 0.05925f
C1603 a_42263_61411# VDD 0.04448f
C1604 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_0.Vout 0.25855f
C1605 D_FlipFlop_3.Qbar D_FlipFlop_3.Nand_Gate_1.Vout 0.11654f
C1606 a_n505_56723# Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.05964f
C1607 Nand_Gate_5.A a_41413_55365# 0.0139f
C1608 And_Gate_3.Nand_Gate_0.Vout VDD 1.39634f
C1609 Nand_Gate_6.A a_16465_56723# 0.05925f
C1610 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout a_41413_56723# 0.04443f
C1611 D_FlipFlop_4.CLK D_FlipFlop_4.3-input-nand_2.C 0.19377f
C1612 D_FlipFlop_7.nPRE a_n1355_60797# 0.10368f
C1613 Nand_Gate_7.A VDD 4.59623f
C1614 D_FlipFlop_6.nPRE D_FlipFlop_6.Inverter_1.Vout 0.07033f
C1615 D_FlipFlop_5.CLK a_15496_48405# 0.04443f
C1616 D_FlipFlop_3.nPRE a_23291_52049# 0.02193f
C1617 Nand_Gate_5.A And_Gate_6.Nand_Gate_0.Vout 0.01068f
C1618 a_35135_55365# Ring_Counter_0.D_FlipFlop_4.Qbar 0.01335f
C1619 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_10.Qbar 0.11657f
C1620 D_FlipFlop_1.CLK D_FlipFlop_1.3-input-nand_1.Vout 0.67419f
C1621 Nand_Gate_1.A D_FlipFlop_7.nPRE 1.92259f
C1622 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout a_n4069_56723# 0.04995f
C1623 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout CLK 0.7779f
C1624 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1625 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.21032f
C1626 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK 0.36346f
C1627 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout VDD 2.07898f
C1628 a_38699_58825# Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.05964f
C1629 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout CLK 0.20785f
C1630 Nand_Gate_0.A a_1758_52049# 0.04443f
C1631 CDAC_v3_0.switch_0.Z Q5 0.02961f
C1632 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout EN 0.78583f
C1633 Ring_Counter_0.D_FlipFlop_16.Q a_10187_61411# 0.01252f
C1634 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1635 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.04109f
C1636 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C VDD 2.82117f
C1637 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.01194f
C1638 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.01194f
C1639 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C a_n4069_56723# 0.04443f
C1640 a_16854_48405# VDD 0.01186f
C1641 a_42263_58825# CLK 0.03f
C1642 Nand_Gate_5.A a_37849_55365# 0.05925f
C1643 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.04107f
C1644 D_FlipFlop_6.Qbar a_4018_51119# 0.04443f
C1645 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout a_34285_61411# 0.01335f
C1646 a_n7633_60797# Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.05964f
C1647 a_48541_59439# a_48541_58825# 0.05935f
C1648 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.01162f
C1649 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout CLK 0.12427f
C1650 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout a_n505_58825# 0.04444f
C1651 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.10915f
C1652 a_n505_56723# VDD 0.02578f
C1653 a_n2642_51119# a_n2028_51119# 0.05935f
C1654 D_FlipFlop_4.Nand_Gate_1.Vout VDD 1.44366f
C1655 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_0.Vout 0.25963f
C1656 a_14529_52049# VDD 0.02521f
C1657 a_n670_48405# a_n56_48405# 0.05935f
C1658 D_FlipFlop_5.Nand_Gate_1.Vout a_20928_48405# 0.04995f
C1659 D_FlipFlop_2.nPRE D_FlipFlop_2.Nand_Gate_0.Vout 0.5831f
C1660 D_FlipFlop_7.3-input-nand_2.C a_n8818_51119# 0.04443f
C1661 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C EN 0.07565f
C1662 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1663 a_26230_51119# D_FlipFlop_3.3-input-nand_2.Vout 0.05964f
C1664 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout a_34285_59439# 0.01335f
C1665 a_48541_59439# VDD 0.01186f
C1666 a_39066_51119# VDD 0.02521f
C1667 VDD Q6 3.6128f
C1668 D_FlipFlop_4.nPRE a_6120_48405# 0.0452f
C1669 a_27542_45397# CDAC_v3_0.switch_5.Z 0.27062f
C1670 a_n2642_51119# VDD 0.01186f
C1671 Ring_Counter_0.D_FlipFlop_16.Q a_35135_61411# 0.01252f
C1672 a_37849_58825# VDD 0.02521f
C1673 a_28007_59439# a_28007_58825# 0.05935f
C1674 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.10034f
C1675 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C CLK 0.19664f
C1676 a_26230_51119# VDD 0.02521f
C1677 a_5767_52049# CLK 0.04479f
C1678 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout 0.01194f
C1679 a_31571_55365# Ring_Counter_0.D_FlipFlop_5.Qbar 0.01335f
C1680 a_27542_45397# VDD 1.17814f
C1681 D_FlipFlop_6.3-input-nand_2.C a_n670_48405# 0.01335f
C1682 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout 0.06895f
C1683 a_28007_59439# VDD 0.05686f
C1684 a_n4744_48405# Q0 0.05747f
C1685 a_2209_60797# VDD 0.02521f
C1686 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.08674f
C1687 a_17315_58825# Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.04443f
C1688 a_17315_58825# VDD 0.02578f
C1689 D_FlipFlop_1.Qbar a_47828_51119# 0.04443f
C1690 D_FlipFlop_5.nPRE a_20029_56723# 0.05925f
C1691 D_FlipFlop_7.CLK D_FlipFlop_7.3-input-nand_1.Vout 0.67419f
C1692 D_FlipFlop_7.Qbar D_FlipFlop_7.Nand_Gate_1.Vout 0.11654f
C1693 a_20029_59439# EN 0.045f
C1694 D_FlipFlop_4.nPRE D_FlipFlop_4.CLK 0.1668f
C1695 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.01323f
C1696 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1697 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout VDD 2.8343f
C1698 a_41168_51119# a_41782_51119# 0.05935f
C1699 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout 0.06935f
C1700 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C a_27157_58825# 0.04443f
C1701 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.21777f
C1702 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.01262f
C1703 a_6623_60797# CLK 0.06211f
C1704 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.29165f
C1705 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.01323f
C1706 D_FlipFlop_2.3-input-nand_2.C a_34992_51119# 0.04443f
C1707 D_FlipFlop_2.Nand_Gate_1.Vout Q7 0.02995f
C1708 Ring_Counter_0.D_FlipFlop_16.Q a_n4919_54751# 0.06113f
C1709 a_20879_59439# Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.01335f
C1710 Nand_Gate_5.A D_FlipFlop_1.nPRE 2.52951f
C1711 And_Gate_6.A VDD 1.33624f
C1712 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.08462f
C1713 D_FlipFlop_5.3-input-nand_1.B a_14882_48405# 0.04995f
C1714 a_17315_60797# Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.05964f
C1715 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout a_27157_59439# 0.04995f
C1716 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_n4069_55365# 0.04995f
C1717 a_6623_59439# CLK 0.03166f
C1718 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_20879_54751# 0.04444f
C1719 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_n4919_55365# 0.04995f
C1720 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_1.Qbar 0.11657f
C1721 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.06935f
C1722 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.01202f
C1723 D_FlipFlop_4.CLK D_FlipFlop_4.3-input-nand_0.Vout 0.25957f
C1724 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_20029_54751# 0.04444f
C1725 a_27157_60797# VDD 0.02521f
C1726 Nand_Gate_4.A a_30721_59439# 0.05925f
C1727 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C VDD 3.50703f
C1728 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 1.09973f
C1729 a_n4069_58825# CLK 0.03f
C1730 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1731 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.08643f
C1732 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_44977_56723# 0.05964f
C1733 D_FlipFlop_4.CLK Q1 0.01843f
C1734 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B EN 0.3979f
C1735 a_28007_55365# Ring_Counter_0.D_FlipFlop_6.Qbar 0.01335f
C1736 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout 0.15413f
C1737 D_FlipFlop_7.nPRE a_n1355_59439# 0.05925f
C1738 a_10187_61411# EN 0.07048f
C1739 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B EN 0.3979f
C1740 a_34992_48405# VDD 0.02521f
C1741 a_31571_60797# CLK 0.06211f
C1742 D_FlipFlop_0.3-input-nand_1.B Q7 0.02377f
C1743 a_24443_56723# Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.05964f
C1744 D_FlipFlop_6.Nand_Gate_0.Vout a_4018_51119# 0.04444f
C1745 Ring_Counter_0.D_FlipFlop_16.Q a_n4919_60797# 0.01768f
C1746 a_2209_59439# VDD 0.01186f
C1747 And_Gate_2.A And_Gate_2.Nand_Gate_0.Vout 0.24482f
C1748 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.Nand_Gate_1.Vout 0.1541f
C1749 D_FlipFlop_1.3-input-nand_1.Vout a_43754_48405# 0.04444f
C1750 Nand_Gate_6.A a_16465_60797# 0.10368f
C1751 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout a_35135_58825# 0.04444f
C1752 D_FlipFlop_4.3-input-nand_1.Vout VDD 1.76545f
C1753 a_52105_60797# VDD 0.0304f
C1754 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout a_5773_58825# 0.05964f
C1755 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.16431f
C1756 D_FlipFlop_7.3-input-nand_2.C a_n6716_48405# 0.04443f
C1757 D_FlipFlop_7.3-input-nand_0.Vout a_n8818_51119# 0.04444f
C1758 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout a_2209_56723# 0.04443f
C1759 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B EN 0.3979f
C1760 D_FlipFlop_2.Qbar a_39066_48405# 0.06113f
C1761 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout a_12901_56723# 0.04443f
C1762 a_35135_61411# EN 0.07048f
C1763 D_FlipFlop_6.3-input-nand_1.B VDD 1.3477f
C1764 a_49391_56723# VDD 0.02521f
C1765 Ring_Counter_0.D_FlipFlop_16.Q a_20029_60797# 0.01768f
C1766 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout CLK 0.20785f
C1767 D_FlipFlop_5.nPRE a_23593_54751# 0.06113f
C1768 a_42263_60797# Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.05964f
C1769 a_24443_55365# Ring_Counter_0.D_FlipFlop_7.Qbar 0.01335f
C1770 D_FlipFlop_3.CLK CLK 0.07954f
C1771 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout a_9337_58825# 0.04444f
C1772 D_FlipFlop_1.Nand_Gate_0.Vout a_47828_51119# 0.04444f
C1773 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout EN 0.61231f
C1774 D_FlipFlop_0.3-input-nand_2.C Q7 0.02769f
C1775 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout VDD 2.71849f
C1776 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B EN 0.3979f
C1777 a_n7633_58825# Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.05964f
C1778 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_4.Qbar 0.02097f
C1779 a_n56_48405# VDD 0.02521f
C1780 Ring_Counter_0.D_FlipFlop_16.Q EN 1.92162f
C1781 a_5773_56723# VDD 0.02521f
C1782 D_FlipFlop_0.3-input-nand_1.B D_FlipFlop_0.3-input-nand_1.Vout 0.08641f
C1783 D_FlipFlop_0.CLK D_FlipFlop_0.Inverter_1.Vout 0.20785f
C1784 D_FlipFlop_3.3-input-nand_1.Vout a_23644_48405# 0.01335f
C1785 D_FlipFlop_2.3-input-nand_0.Vout a_34992_51119# 0.04444f
C1786 a_54618_51119# VDD 0.02521f
C1787 a_2209_59439# a_2209_58825# 0.05935f
C1788 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.12285f
C1789 D_FlipFlop_5.nPRE a_20029_54751# 0.06135f
C1790 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_28007_55365# 0.04995f
C1791 D_FlipFlop_4.Qbar VDD 1.96371f
C1792 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_27157_55365# 0.04995f
C1793 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout a_52105_54751# 0.04444f
C1794 Ring_Counter_0.D_FlipFlop_16.Q a_44977_60797# 0.01768f
C1795 D_FlipFlop_6.3-input-nand_1.Vout a_n670_48405# 0.04543f
C1796 CDAC_v3_0.switch_5.Z m3_3428_9615# 1.89962f
C1797 a_41782_51119# VDD 0.02521f
C1798 D_FlipFlop_6.3-input-nand_2.C VDD 2.67765f
C1799 D_FlipFlop_2.CLK a_33020_51119# 0.04443f
C1800 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B EN 0.3979f
C1801 D_FlipFlop_1.nPRE a_41413_61411# 0.04995f
C1802 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.Qbar 1.29337f
C1803 D_FlipFlop_6.nPRE And_Gate_1.Nand_Gate_0.Vout 0.10314f
C1804 a_10187_61411# Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.01335f
C1805 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_2.Z 6.50533f
C1806 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.Nand_Gate_1.Vout 0.1541f
C1807 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout VDD 2.72531f
C1808 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.06955f
C1809 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD 1.89599f
C1810 a_12901_61411# VDD 0.08862f
C1811 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B VDD 1.71455f
C1812 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout a_n4919_56723# 0.04443f
C1813 a_54618_48405# VDD 0.02521f
C1814 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B a_24443_60797# 0.04443f
C1815 a_20879_55365# Ring_Counter_0.D_FlipFlop_8.Qbar 0.01335f
C1816 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout VDD 2.07898f
C1817 D_FlipFlop_1.nPRE a_41413_56723# 0.05925f
C1818 D_FlipFlop_4.3-input-nand_2.C a_8092_48405# 0.01335f
C1819 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.01202f
C1820 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_1.Vout 0.08671f
C1821 D_FlipFlop_5.Inverter_1.Vout a_19570_51119# 0.04443f
C1822 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.Qbar 0.11806f
C1823 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.26069f
C1824 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.08582f
C1825 D_FlipFlop_7.nPRE And_Gate_1.Nand_Gate_0.Vout 0.02463f
C1826 D_FlipFlop_5.nPRE D_FlipFlop_5.3-input-nand_2.Vout 0.76528f
C1827 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.08582f
C1828 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.01323f
C1829 D_FlipFlop_0.CLK a_51902_48405# 0.02953f
C1830 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.07084f
C1831 D_FlipFlop_6.Nand_Gate_1.Vout VDD 1.44304f
C1832 Nand_Gate_2.A a_10520_52049# 0.04443f
C1833 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout 0.06935f
C1834 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout a_n7633_59439# 0.04543f
C1835 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C a_24443_56723# 0.04443f
C1836 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout VDD 2.72531f
C1837 a_n9432_51119# D_FlipFlop_7.3-input-nand_2.Vout 0.01335f
C1838 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.Inverter_1.Vout 0.26069f
C1839 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD 1.89599f
C1840 a_37849_61411# VDD 0.08862f
C1841 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.Inverter_1.Vout 0.06895f
C1842 D_FlipFlop_4.nPRE a_16465_54751# 0.06113f
C1843 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.17188f
C1844 a_49391_58825# Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.05964f
C1845 Nand_Gate_2.A And_Gate_2.A 0.07775f
C1846 D_FlipFlop_5.CLK a_17468_48405# 0.02953f
C1847 a_49391_56723# Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout 0.05964f
C1848 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout EN 0.78583f
C1849 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.01194f
C1850 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.01194f
C1851 D_FlipFlop_3.Inverter_1.Vout VDD 1.70372f
C1852 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.15413f
C1853 D_FlipFlop_5.3-input-nand_1.B D_FlipFlop_5.3-input-nand_1.Vout 0.08641f
C1854 D_FlipFlop_5.nPRE a_20029_59439# 0.05925f
C1855 D_FlipFlop_3.3-input-nand_1.B a_23644_48405# 0.04995f
C1856 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.48403f
C1857 a_10808_51119# D_FlipFlop_4.Nand_Gate_0.Vout 0.05964f
C1858 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.0646f
C1859 And_Gate_5.Nand_Gate_0.Vout D_FlipFlop_2.CLK 0.25559f
C1860 And_Gate_3.Nand_Gate_0.Vout CLK 0.79128f
C1861 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.06462f
C1862 Ring_Counter_0.D_FlipFlop_16.Q a_5773_61411# 0.01252f
C1863 a_19570_48405# VDD 0.02521f
C1864 Nand_Gate_7.A CLK 0.45134f
C1865 D_FlipFlop_4.nPRE a_12901_54751# 0.06135f
C1866 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout a_44977_58825# 0.04444f
C1867 a_17315_55365# Ring_Counter_0.D_FlipFlop_9.Qbar 0.01335f
C1868 a_35135_61411# Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.01335f
C1869 D_FlipFlop_1.Nand_Gate_1.Vout a_47214_48405# 0.04995f
C1870 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C EN 0.07565f
C1871 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.Nand_Gate_0.Vout 0.16429f
C1872 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.16431f
C1873 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_11.Qbar 0.07122f
C1874 a_n2028_51119# D_FlipFlop_6.3-input-nand_0.Vout 0.05964f
C1875 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout a_44977_59439# 0.01335f
C1876 a_34378_51119# D_FlipFlop_2.3-input-nand_2.Vout 0.01335f
C1877 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.Inverter_1.Vout 0.26069f
C1878 a_23291_52049# VDD 0.02521f
C1879 a_55976_51119# VDD 0.01186f
C1880 a_n5358_51119# Q0 0.01335f
C1881 CDAC_v3_0.switch_7.Z Q6 0.17526f
C1882 a_38699_59439# a_38699_58825# 0.05935f
C1883 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.25966f
C1884 D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.43587f
C1885 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C CLK 0.19645f
C1886 D_FlipFlop_5.CLK VDD 2.17957f
C1887 a_43140_51119# VDD 0.01186f
C1888 Nand_Gate_0.A a_2209_61411# 0.04995f
C1889 a_49391_59439# VDD 0.01186f
C1890 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B 0.02535f
C1891 D_FlipFlop_6.3-input-nand_0.Vout VDD 1.74442f
C1892 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.0646f
C1893 a_38699_58825# VDD 0.02578f
C1894 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.06462f
C1895 a_28007_58825# Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.04443f
C1896 Ring_Counter_0.D_FlipFlop_16.Q a_30721_61411# 0.01252f
C1897 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_1.Vout 0.08671f
C1898 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B a_13751_61411# 0.04995f
C1899 a_41413_59439# EN 0.045f
C1900 a_14529_52049# CLK 0.04479f
C1901 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B 0.29684f
C1902 a_31486_45397# VDD 1.17814f
C1903 D_FlipFlop_6.3-input-nand_2.C a_2046_48405# 0.04443f
C1904 a_54618_51119# D_FlipFlop_0.Nand_Gate_0.Vout 0.05964f
C1905 D_FlipFlop_1.nPRE D_FlipFlop_2.Qbar 0.01961f
C1906 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout VDD 2.8343f
C1907 Nand_Gate_7.A a_48541_55365# 0.0139f
C1908 a_3059_61411# a_3059_60797# 0.05935f
C1909 a_3059_60797# VDD 0.02865f
C1910 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout a_2209_60797# 0.05964f
C1911 D_FlipFlop_1.Qbar a_47828_48405# 0.06113f
C1912 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C a_37849_58825# 0.04443f
C1913 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.17364f
C1914 a_31571_59439# Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.01335f
C1915 a_41782_51119# D_FlipFlop_1.3-input-nand_0.Vout 0.05964f
C1916 a_13751_55365# Ring_Counter_0.D_FlipFlop_10.Qbar 0.01335f
C1917 D_FlipFlop_6.nPRE a_9337_54751# 0.06113f
C1918 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.04107f
C1919 a_28007_59439# CLK 0.03166f
C1920 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.25966f
C1921 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout EN 0.78583f
C1922 D_FlipFlop_6.3-input-nand_1.Vout VDD 1.76485f
C1923 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C VDD 3.50703f
C1924 a_2209_60797# CLK 0.06211f
C1925 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B 0.29684f
C1926 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 1.09973f
C1927 a_17315_58825# CLK 0.03f
C1928 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.07084f
C1929 Nand_Gate_7.A a_44977_55365# 0.05925f
C1930 D_FlipFlop_7.3-input-nand_2.Vout a_n8818_48405# 0.04443f
C1931 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.01162f
C1932 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout a_28007_59439# 0.04543f
C1933 D_FlipFlop_6.Nand_Gate_1.Vout a_2046_48405# 0.05964f
C1934 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.12285f
C1935 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout CLK 0.12427f
C1936 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_15.Qbar 0.11657f
C1937 Nand_Gate_5.A a_45568_52049# 0.0451f
C1938 D_FlipFlop_3.nPRE a_29690_51119# 0.04443f
C1939 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout EN 0.08727f
C1940 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.08674f
C1941 a_28007_60797# VDD 0.02865f
C1942 a_12901_61411# a_12901_60797# 0.05935f
C1943 D_FlipFlop_6.nPRE a_5773_54751# 0.06171f
C1944 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.01202f
C1945 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C EN 0.07565f
C1946 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout a_30721_56723# 0.04443f
C1947 And_Gate_6.A CLK 1.52489f
C1948 D_FlipFlop_7.CLK a_n10790_48405# 0.04443f
C1949 a_23593_59439# VDD 0.01186f
C1950 Ring_Counter_0.D_FlipFlop_16.Q a_n7633_54751# 0.04443f
C1951 D_FlipFlop_4.Nand_Gate_0.Vout a_12166_51119# 0.04543f
C1952 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout EN 0.09223f
C1953 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B 0.29684f
C1954 a_38452_48405# VDD 0.01186f
C1955 a_31571_56723# VDD 0.02578f
C1956 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.10034f
C1957 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout EN 0.96763f
C1958 a_5773_61411# EN 0.02636f
C1959 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C1960 a_12901_58825# VDD 0.02521f
C1961 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout a_16465_58825# 0.05964f
C1962 CDAC_v3_0.switch_0.Z Q1 0.21005f
C1963 a_27157_60797# CLK 0.06211f
C1964 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C CLK 0.19664f
C1965 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.08462f
C1966 D_FlipFlop_6.nPRE a_3404_51119# 0.04443f
C1967 Ring_Counter_0.D_FlipFlop_16.Q a_n4069_60797# 0.01768f
C1968 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_2.Qbar 0.07122f
C1969 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout EN 0.61231f
C1970 a_3059_59439# VDD 0.05686f
C1971 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout a_2209_59439# 0.04995f
C1972 a_10187_55365# Ring_Counter_0.D_FlipFlop_11.Qbar 0.01335f
C1973 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1974 D_FlipFlop_6.3-input-nand_0.Vout a_n670_51119# 0.04543f
C1975 a_3404_51119# Q1 0.01335f
C1976 a_28007_61411# a_28007_60797# 0.05935f
C1977 a_n7633_58825# VDD 0.02578f
C1978 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout a_27157_60797# 0.05964f
C1979 a_n4919_59439# EN 0.045f
C1980 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C1981 a_12780_51119# VDD 0.02521f
C1982 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.26069f
C1983 D_FlipFlop_5.3-input-nand_2.C a_16854_48405# 0.01335f
C1984 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B 0.29684f
C1985 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_2209_56723# 0.05964f
C1986 And_Gate_2.Nand_Gate_0.Vout VDD 1.38895f
C1987 D_FlipFlop_4.CLK D_FlipFlop_4.Inverter_1.Vout 0.20785f
C1988 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C1989 a_n56_51119# VDD 0.02521f
C1990 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout EN 0.09223f
C1991 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B a_n4069_60797# 0.04443f
C1992 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout EN 0.96763f
C1993 VDD Q2 3.61866f
C1994 a_30721_61411# EN 0.02636f
C1995 a_52105_60797# CLK 0.04443f
C1996 D_FlipFlop_0.Nand_Gate_0.Vout a_55976_51119# 0.04995f
C1997 D_FlipFlop_7.nPRE a_2209_54751# 0.06113f
C1998 Ring_Counter_0.D_FlipFlop_16.Q a_20879_60797# 0.01768f
C1999 a_3059_58825# Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C 0.05964f
C2000 D_FlipFlop_7.nPRE a_n9432_51119# 0.045f
C2001 D_FlipFlop_7.CLK a_n10790_51119# 0.04443f
C2002 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout a_10187_58825# 0.04444f
C2003 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.10915f
C2004 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.01194f
C2005 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.01194f
C2006 a_37849_61411# a_37849_60797# 0.05935f
C2007 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.04107f
C2008 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B 0.29684f
C2009 a_12901_59439# a_12901_58825# 0.05935f
C2010 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout a_n4919_61411# 0.01335f
C2011 D_FlipFlop_1.3-input-nand_0.Vout a_43140_51119# 0.04543f
C2012 a_3404_48405# VDD 0.01186f
C2013 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C2014 D_FlipFlop_0.3-input-nand_1.Vout a_49930_48405# 0.01335f
C2015 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout VDD 2.07898f
C2016 And_Gate_2.A D_FlipFlop_4.CLK 0.06897f
C2017 D_FlipFlop_2.3-input-nand_1.B a_32406_48405# 0.04995f
C2018 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.26069f
C2019 a_6623_55365# Ring_Counter_0.D_FlipFlop_12.Qbar 0.01335f
C2020 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.04109f
C2021 D_FlipFlop_3.3-input-nand_1.Vout a_25616_48405# 0.04543f
C2022 D_FlipFlop_7.nPRE a_n1355_54751# 0.05925f
C2023 D_FlipFlop_7.Nand_Gate_1.Vout VDD 1.44304f
C2024 Nand_Gate_4.A a_30721_60797# 0.10368f
C2025 D_FlipFlop_5.nPRE a_20879_54751# 0.06196f
C2026 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_3059_54751# 0.04444f
C2027 Nand_Gate_3.A a_23593_56723# 0.05925f
C2028 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_6.Qbar 0.11657f
C2029 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_2209_54751# 0.04444f
C2030 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout CLK 0.67422f
C2031 Ring_Counter_0.D_FlipFlop_16.Q a_45827_60797# 0.01768f
C2032 CDAC_v3_0.switch_6.Z m3_3428_38799# 16.1764f
C2033 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout a_n1355_59439# 0.01335f
C2034 D_FlipFlop_5.nPRE a_20029_60797# 0.10368f
C2035 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B 0.29684f
C2036 a_n7633_59439# a_n7633_58825# 0.05935f
C2037 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.30156f
C2038 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.08674f
C2039 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_4.Z 0.28068f
C2040 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_3.Z 19.6021f
C2041 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout a_52105_60797# 0.05964f
C2042 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.21542f
C2043 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.01194f
C2044 a_13751_61411# VDD 0.04448f
C2045 Nand_Gate_6.A a_19282_52049# 0.04443f
C2046 D_FlipFlop_1.nPRE Nand_Gate_7.A 0.05024f
C2047 a_56590_48405# VDD 0.02521f
C2048 a_12166_51119# a_12780_51119# 0.05935f
C2049 And_Gate_6.A And_Gate_6.Nand_Gate_0.Vout 0.24482f
C2050 D_FlipFlop_5.nPRE EN 0.79742f
C2051 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.26069f
C2052 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD 1.48403f
C2053 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.16917f
C2054 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.15413f
C2055 D_FlipFlop_4.3-input-nand_2.C a_10808_48405# 0.04443f
C2056 a_12166_51119# Q2 0.01335f
C2057 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout CLK 0.78664f
C2058 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.08462f
C2059 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout CLK 0.36346f
C2060 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B EN 0.3979f
C2061 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B 0.29684f
C2062 D_FlipFlop_3.nPRE a_30721_54751# 0.06113f
C2063 a_n670_51119# a_n56_51119# 0.05935f
C2064 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout a_37849_59439# 0.04995f
C2065 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B CLK 0.08407f
C2066 D_FlipFlop_0.Qbar a_56590_48405# 0.06113f
C2067 a_3059_55365# Ring_Counter_0.D_FlipFlop_13.Qbar 0.01335f
C2068 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B EN 0.3979f
C2069 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.06734f
C2070 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.01162f
C2071 Nand_Gate_6.A VDD 4.32137f
C2072 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.04107f
C2073 And_Gate_5.A VDD 1.34097f
C2074 a_38699_61411# VDD 0.04448f
C2075 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout a_20029_61411# 0.01335f
C2076 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_2.Qbar 0.02966f
C2077 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout EN 0.08727f
C2078 D_FlipFlop_4.nPRE a_6120_51119# 0.034f
C2079 D_FlipFlop_4.nPRE EN 0.79742f
C2080 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.20923f
C2081 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.16431f
C2082 D_FlipFlop_6.nPRE D_FlipFlop_6.CLK 0.16209f
C2083 a_55976_51119# a_56590_51119# 0.05935f
C2084 D_FlipFlop_6.3-input-nand_2.Vout a_n56_48405# 0.04443f
C2085 D_FlipFlop_3.nPRE a_27157_54751# 0.05925f
C2086 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B 0.29684f
C2087 D_FlipFlop_1.nPRE Q6 0.03712f
C2088 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout CLK 0.7779f
C2089 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK 0.36346f
C2090 a_37849_56723# VDD 0.02521f
C2091 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.10034f
C2092 Nand_Gate_2.A VDD 4.25845f
C2093 Ring_Counter_0.D_FlipFlop_16.Q a_6623_61411# 0.01252f
C2094 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout a_45827_58825# 0.04444f
C2095 D_FlipFlop_3.3-input-nand_2.Vout a_28332_51119# 0.04443f
C2096 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.Qbar 1.29337f
C2097 a_51902_51119# EN 0.01768f
C2098 a_21542_48405# VDD 0.02521f
C2099 D_FlipFlop_4.nPRE a_13751_54751# 0.06196f
C2100 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_27157_56723# 0.05964f
C2101 a_6120_51119# D_FlipFlop_4.3-input-nand_0.Vout 0.01335f
C2102 a_43140_51119# a_43754_51119# 0.05935f
C2103 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.01194f
C2104 a_49391_59439# a_49391_58825# 0.05935f
C2105 D_FlipFlop_6.nPRE EN 0.79742f
C2106 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.30154f
C2107 a_28332_51119# VDD 0.02521f
C2108 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.Vout 1.01753f
C2109 Nand_Gate_7.A a_44977_58825# 0.05925f
C2110 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_10187_55365# 0.04995f
C2111 a_32053_52049# VDD 0.02521f
C2112 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_35135_54751# 0.04444f
C2113 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_9337_55365# 0.04995f
C2114 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_34285_54751# 0.04444f
C2115 D_FlipFlop_7.3-input-nand_1.Vout VDD 1.76484f
C2116 D_FlipFlop_6.3-input-nand_1.B Q0 0.01488f
C2117 a_38699_58825# Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.04443f
C2118 a_15496_51119# VDD 0.02521f
C2119 D_FlipFlop_7.Inverter_1.Vout a_n6716_48405# 0.04995f
C2120 a_6623_56723# Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.05964f
C2121 a_n505_55365# Ring_Counter_0.D_FlipFlop_14.Qbar 0.01335f
C2122 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout VDD 2.29929f
C2123 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.09856f
C2124 D_FlipFlop_1.3-input-nand_2.Vout VDD 2.67043f
C2125 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout VDD 3.55971f
C2126 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_4.Qbar 0.11806f
C2127 Nand_Gate_0.A VDD 4.27383f
C2128 a_31486_45397# CDAC_v3_0.switch_7.Z 0.27022f
C2129 D_FlipFlop_2.CLK D_FlipFlop_2.3-input-nand_2.Vout 0.1192f
C2130 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C a_48541_58825# 0.04443f
C2131 D_FlipFlop_1.nPRE And_Gate_6.A 0.38333f
C2132 D_FlipFlop_7.nPRE EN 0.79742f
C2133 Ring_Counter_0.D_FlipFlop_16.Q a_31571_61411# 0.01252f
C2134 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout a_20029_58825# 0.04444f
C2135 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.08582f
C2136 a_23291_52049# CLK 0.04479f
C2137 a_35430_45397# VDD 1.17814f
C2138 a_42263_59439# Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.01335f
C2139 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.04107f
C2140 D_FlipFlop_3.3-input-nand_2.C a_25616_48405# 0.01335f
C2141 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout a_44977_61411# 0.01335f
C2142 a_3059_60797# Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.05964f
C2143 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.04109f
C2144 a_49930_51119# D_FlipFlop_0.3-input-nand_0.Vout 0.01335f
C2145 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.01202f
C2146 D_FlipFlop_5.CLK CLK 0.07954f
C2147 a_49391_59439# CLK 0.03166f
C2148 a_n1355_60797# VDD 0.02521f
C2149 a_20928_51119# Q3 0.01335f
C2150 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.21297f
C2151 a_19654_45397# Q3 0.46777f
C2152 D_FlipFlop_0.Inverter_1.Vout Q7 0.02777f
C2153 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout EN 0.78583f
C2154 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 1.09973f
C2155 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C VDD 3.50703f
C2156 a_38699_58825# CLK 0.03f
C2157 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.Vout 1.01753f
C2158 a_13751_56723# VDD 0.02578f
C2159 Nand_Gate_1.A VDD 4.36672f
C2160 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.10915f
C2161 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout CLK 0.12427f
C2162 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B VDD 1.71455f
C2163 D_FlipFlop_2.nPRE And_Gate_5.A 0.3733f
C2164 D_FlipFlop_3.Nand_Gate_1.Vout a_28332_48405# 0.05964f
C2165 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout EN 0.61231f
C2166 a_3059_60797# CLK 0.06211f
C2167 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.06734f
C2168 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.06955f
C2169 D_FlipFlop_6.Nand_Gate_1.Vout a_4018_48405# 0.04444f
C2170 D_FlipFlop_4.nPRE D_FlipFlop_4.3-input-nand_1.B 0.27142f
C2171 Nand_Gate_7.A a_44977_56723# 0.05925f
C2172 a_n4069_55365# Ring_Counter_0.D_FlipFlop_15.Qbar 0.01335f
C2173 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C EN 0.07537f
C2174 D_FlipFlop_3.CLK a_25616_48405# 0.02953f
C2175 D_FlipFlop_1.3-input-nand_1.B a_41168_48405# 0.04995f
C2176 D_FlipFlop_6.Inverter_1.Vout VDD 1.70303f
C2177 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.01162f
C2178 a_44977_59439# VDD 0.01186f
C2179 a_52105_54751# VDD 0.02521f
C2180 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C a_13751_56723# 0.04443f
C2181 a_23593_60797# VDD 0.02521f
C2182 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout 0.30046f
C2183 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B a_38699_61411# 0.04995f
C2184 D_FlipFlop_6.nPRE a_6623_54751# 0.06233f
C2185 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout a_27157_58825# 0.05964f
C2186 a_34285_58825# VDD 0.02521f
C2187 a_55976_48405# a_56590_48405# 0.05935f
C2188 D_FlipFlop_2.CLK D_FlipFlop_2.3-input-nand_1.Vout 0.67419f
C2189 Nand_Gate_0.A a_2209_58825# 0.05925f
C2190 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C CLK 0.19664f
C2191 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.01162f
C2192 D_FlipFlop_3.nPRE And_Gate_4.A 0.37768f
C2193 D_FlipFlop_7.CLK a_n8818_48405# 0.02953f
C2194 a_24443_59439# VDD 0.05686f
C2195 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B a_28007_61411# 0.04995f
C2196 a_41168_48405# VDD 0.01186f
C2197 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.15413f
C2198 D_FlipFlop_6.nPRE a_5773_61411# 0.04995f
C2199 D_FlipFlop_5.CLK D_FlipFlop_5.3-input-nand_1.B 0.06986f
C2200 a_6623_61411# EN 0.07048f
C2201 D_FlipFlop_7.nPRE a_n7004_52049# 0.04597f
C2202 a_13751_58825# VDD 0.02578f
C2203 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B a_45827_61411# 0.04995f
C2204 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.07084f
C2205 a_28007_60797# CLK 0.06211f
C2206 D_FlipFlop_2.nPRE a_32053_52049# 0.02193f
C2207 a_16465_59439# EN 0.045f
C2208 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_16.Qbar 0.06863f
C2209 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout a_3059_59439# 0.04543f
C2210 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.10034f
C2211 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.09856f
C2212 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout VDD 2.8343f
C2213 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_42263_55365# 0.04995f
C2214 a_29690_51119# VDD 0.01186f
C2215 a_48541_54751# VDD 0.02521f
C2216 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_41413_55365# 0.04995f
C2217 D_FlipFlop_4.3-input-nand_1.B Q1 0.01615f
C2218 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.3-input-nand_2.Vout 0.0846f
C2219 a_28007_60797# Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.05964f
C2220 D_FlipFlop_7.nPRE And_Gate_0.Nand_Gate_0.Vout 0.12621f
C2221 a_16854_51119# VDD 0.01186f
C2222 a_48541_60797# VDD 0.02521f
C2223 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.10034f
C2224 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.01202f
C2225 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.16431f
C2226 D_FlipFlop_5.nPRE And_Gate_3.A 0.3744f
C2227 D_FlipFlop_5.3-input-nand_2.C a_19570_48405# 0.04443f
C2228 D_FlipFlop_4.nPRE D_FlipFlop_4.3-input-nand_2.C 0.05823f
C2229 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout a_17315_56723# 0.04995f
C2230 a_13751_58825# Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.05964f
C2231 a_n7633_55365# Ring_Counter_0.D_FlipFlop_16.Qbar 0.01335f
C2232 a_3059_59439# CLK 0.03166f
C2233 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.25966f
C2234 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout a_52105_56723# 0.05964f
C2235 a_31571_61411# EN 0.07048f
C2236 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C VDD 3.50703f
C2237 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.01194f
C2238 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Qbar 0.06863f
C2239 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.01194f
C2240 a_44977_54751# VDD 0.02521f
C2241 And_Gate_7.A a_54330_52049# 0.06113f
C2242 a_n7633_58825# CLK 0.02953f
C2243 a_23593_59439# a_23593_58825# 0.05935f
C2244 D_FlipFlop_7.nPRE D_FlipFlop_7.3-input-nand_2.Vout 0.76528f
C2245 a_29690_51119# Q4 0.01335f
C2246 Ring_Counter_0.D_FlipFlop_16.Q a_16465_60797# 0.01768f
C2247 a_38452_48405# a_39066_48405# 0.05935f
C2248 a_31571_56723# Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.05964f
C2249 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.06734f
C2250 D_FlipFlop_5.CLK D_FlipFlop_5.3-input-nand_2.C 0.19377f
C2251 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout a_23593_56723# 0.04443f
C2252 And_Gate_2.Nand_Gate_0.Vout CLK 0.79128f
C2253 D_FlipFlop_4.nPRE And_Gate_3.A 0.01999f
C2254 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.3-input-nand_2.C 0.06863f
C2255 a_n4069_61411# Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.01335f
C2256 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.3-input-nand_2.Vout 0.0846f
C2257 D_FlipFlop_4.3-input-nand_2.Vout a_8706_48405# 0.04443f
C2258 a_6120_48405# VDD 0.01186f
C2259 D_FlipFlop_0.3-input-nand_1.Vout a_51902_48405# 0.04543f
C2260 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD 1.48403f
C2261 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B 0.29684f
C2262 Nand_Gate_0.A And_Gate_1.A 0.07817f
C2263 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout a_9337_59439# 0.01335f
C2264 a_n1355_59439# VDD 0.01186f
C2265 a_41413_54751# VDD 0.02521f
C2266 D_FlipFlop_7.nPRE a_n505_54751# 0.05987f
C2267 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout a_31571_56723# 0.04995f
C2268 a_3059_59439# a_3059_58825# 0.05935f
C2269 D_FlipFlop_4.nPRE D_FlipFlop_5.nPRE 0.04585f
C2270 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.17188f
C2271 CDAC_v3_0.switch_6.Z m3_3428_9615# 16.1792f
C2272 D_FlipFlop_2.nPRE a_34285_58825# 0.05925f
C2273 D_FlipFlop_4.CLK VDD 2.17721f
C2274 Ring_Counter_0.D_FlipFlop_16.Q a_41413_60797# 0.01768f
C2275 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.01262f
C2276 a_n7633_58825# Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.04443f
C2277 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_4.Z 2.32723f
C2278 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.29165f
C2279 Q6 Q7 6.30379f
C2280 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout a_n505_56723# 0.04995f
C2281 D_FlipFlop_6.Inverter_1.Vout a_2046_48405# 0.04995f
C2282 D_FlipFlop_5.nPRE D_FlipFlop_5.Nand_Gate_0.Vout 0.5831f
C2283 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout VDD 2.72531f
C2284 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout a_37849_56723# 0.04443f
C2285 a_37849_54751# VDD 0.02521f
C2286 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.25858f
C2287 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD 1.89599f
C2288 CDAC_v3_0.switch_8.Z VDD 1.08716f
C2289 a_9337_61411# VDD 0.08862f
C2290 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout EN 0.19184f
C2291 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_2.C 0.07084f
C2292 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C a_2209_58825# 0.04443f
C2293 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.06837f
C2294 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_7.Qbar 0.07122f
C2295 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout 0.25855f
C2296 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B a_n505_60797# 0.04443f
C2297 a_n4069_59439# Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.01335f
C2298 a_20029_56723# VDD 0.02521f
C2299 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout a_20029_56723# 0.04443f
C2300 D_FlipFlop_5.3-input-nand_1.B Q2 0.0191f
C2301 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.20931f
C2302 a_20928_48405# a_21542_48405# 0.05935f
C2303 D_FlipFlop_2.3-input-nand_2.C a_34378_48405# 0.01335f
C2304 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout a_38699_59439# 0.04543f
C2305 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout a_45827_56723# 0.04995f
C2306 a_n56_51119# D_FlipFlop_6.3-input-nand_2.Vout 0.05964f
C2307 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.08674f
C2308 And_Gate_0.Nand_Gate_0.Vout D_FlipFlop_7.CLK 0.25559f
C2309 a_34285_54751# VDD 0.02521f
C2310 a_20879_61411# Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.01335f
C2311 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C2312 D_FlipFlop_4.3-input-nand_1.Vout a_6734_48405# 0.05964f
C2313 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout VDD 2.72531f
C2314 D_FlipFlop_4.nPRE D_FlipFlop_4.3-input-nand_0.Vout 0.94459f
C2315 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD 1.89599f
C2316 D_FlipFlop_6.nPRE D_FlipFlop_4.nPRE 0.68069f
C2317 a_34285_61411# VDD 0.08862f
C2318 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout a_52105_56723# 0.04443f
C2319 D_FlipFlop_4.nPRE Q1 0.01391f
C2320 D_FlipFlop_5.Qbar a_21542_51119# 0.04443f
C2321 a_38452_51119# Q5 0.01335f
C2322 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout 0.06935f
C2323 D_FlipFlop_1.nPRE a_43140_51119# 0.045f
C2324 D_FlipFlop_3.nPRE a_28007_54751# 0.05987f
C2325 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.08462f
C2326 Nand_Gate_6.A CLK 0.95447f
C2327 a_14882_51119# a_15496_51119# 0.05935f
C2328 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C2329 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.01162f
C2330 D_FlipFlop_7.CLK D_FlipFlop_7.3-input-nand_2.Vout 0.1192f
C2331 a_30721_54751# VDD 0.02521f
C2332 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout VDD 2.07898f
C2333 D_FlipFlop_0.3-input-nand_1.B a_49930_48405# 0.04995f
C2334 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout a_12901_59439# 0.04995f
C2335 And_Gate_5.A CLK 1.52489f
C2336 And_Gate_6.A D_FlipFlop_1.CLK 0.06897f
C2337 D_FlipFlop_5.CLK D_FlipFlop_5.3-input-nand_0.Vout 0.25957f
C2338 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.0646f
C2339 D_FlipFlop_0.3-input-nand_2.Vout EN 0.09383f
C2340 a_24258_48405# VDD 0.02521f
C2341 D_FlipFlop_4.3-input-nand_2.C a_8706_51119# 0.04443f
C2342 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.01202f
C2343 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.06462f
C2344 Ring_Counter_0.D_FlipFlop_16.Q a_2209_61411# 0.01252f
C2345 a_43754_51119# D_FlipFlop_1.3-input-nand_2.Vout 0.05964f
C2346 a_49391_58825# Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.04443f
C2347 a_32406_51119# VDD 0.01186f
C2348 D_FlipFlop_6.nPRE Q1 0.03683f
C2349 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_11.Qbar 0.11657f
C2350 a_n4069_56723# VDD 0.02578f
C2351 a_40815_52049# VDD 0.02521f
C2352 a_3404_48405# a_4018_48405# 0.05935f
C2353 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.10029f
C2354 a_27157_54751# VDD 0.02521f
C2355 Nand_Gate_2.A CLK 0.5121f
C2356 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.1143f
C2357 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.30156f
C2358 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.01262f
C2359 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.29165f
C2360 D_FlipFlop_2.nPRE a_37849_54751# 0.06113f
C2361 And_Gate_1.Nand_Gate_0.Vout VDD 1.39709f
C2362 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout a_20879_58825# 0.04444f
C2363 D_FlipFlop_7.nPRE D_FlipFlop_6.nPRE 1.66474f
C2364 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.0646f
C2365 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.06462f
C2366 a_32053_52049# CLK 0.04479f
C2367 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout EN 0.78583f
C2368 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.01323f
C2369 Ring_Counter_0.D_FlipFlop_16.Q a_27157_61411# 0.01252f
C2370 And_Gate_6.A a_45568_52049# 0.05964f
C2371 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 1.09973f
C2372 D_FlipFlop_3.3-input-nand_2.C a_28332_48405# 0.04443f
C2373 a_45827_61411# Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.01335f
C2374 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_0.Qbar 0.03069f
C2375 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout CLK 0.20785f
C2376 D_FlipFlop_0.3-input-nand_2.C a_52516_51119# 0.04443f
C2377 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.22118f
C2378 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout EN 0.63795f
C2379 a_23593_54751# VDD 0.02521f
C2380 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout CLK 0.1215f
C2381 a_n505_60797# VDD 0.02865f
C2382 Nand_Gate_0.A CLK 0.52304f
C2383 a_n1355_61411# a_n1355_60797# 0.05935f
C2384 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C a_42263_56723# 0.04443f
C2385 D_FlipFlop_7.Nand_Gate_1.Vout Q0 0.09808f
C2386 Nand_Gate_7.A a_44977_61411# 0.04995f
C2387 D_FlipFlop_2.nPRE a_34285_54751# 0.05925f
C2388 D_FlipFlop_0.Nand_Gate_1.Vout a_54618_48405# 0.05964f
C2389 a_n10790_48405# VDD 0.02521f
C2390 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C EN 0.07565f
C2391 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.30156f
C2392 Nand_Gate_3.A a_23593_59439# 0.05925f
C2393 D_FlipFlop_3.Nand_Gate_1.Vout a_30304_48405# 0.04444f
C2394 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.15413f
C2395 D_FlipFlop_2.nPRE a_34285_61411# 0.04995f
C2396 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout a_n4919_58825# 0.04444f
C2397 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.Qbar 1.29337f
C2398 a_n1355_60797# CLK 0.06211f
C2399 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C 0.08674f
C2400 D_FlipFlop_3.nPRE EN 0.79742f
C2401 D_FlipFlop_6.nPRE a_1758_52049# 0.0451f
C2402 D_FlipFlop_5.Nand_Gate_1.Vout Q3 0.10859f
C2403 Ring_Counter_0.D_FlipFlop_16.Q a_52105_61411# 0.04794f
C2404 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout a_37849_58825# 0.05964f
C2405 D_FlipFlop_5.3-input-nand_2.Vout a_17468_48405# 0.04443f
C2406 a_20029_54751# VDD 0.02521f
C2407 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C CLK 0.19664f
C2408 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.17188f
C2409 Nand_Gate_1.A CLK 0.51983f
C2410 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout a_16465_56723# 0.04443f
C2411 a_45827_59439# VDD 0.05686f
C2412 a_47214_51119# Q6 0.01335f
C2413 a_13751_61411# a_13751_60797# 0.05935f
C2414 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B a_17315_60797# 0.04443f
C2415 a_24443_60797# VDD 0.02865f
C2416 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout a_12901_60797# 0.05964f
C2417 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.08582f
C2418 D_FlipFlop_5.Nand_Gate_0.Vout a_21542_51119# 0.04444f
C2419 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B CLK 0.08407f
C2420 a_35135_58825# VDD 0.02578f
C2421 a_37849_59439# EN 0.045f
C2422 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B EN 0.3979f
C2423 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.16431f
C2424 D_FlipFlop_1.Nand_Gate_1.Vout Q6 0.10016f
C2425 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.1143f
C2426 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout VDD 2.8343f
C2427 D_FlipFlop_2.Qbar D_FlipFlop_2.Nand_Gate_1.Vout 0.11654f
C2428 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.08582f
C2429 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.08462f
C2430 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.Qbar 0.11806f
C2431 a_43140_48405# VDD 0.01186f
C2432 D_FlipFlop_2.nPRE a_32406_51119# 0.034f
C2433 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout a_48541_59439# 0.04995f
C2434 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout EN 0.09223f
C2435 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout EN 0.96763f
C2436 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C2437 a_16465_54751# VDD 0.02521f
C2438 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.08582f
C2439 D_FlipFlop_1.CLK a_41782_51119# 0.04443f
C2440 D_FlipFlop_4.3-input-nand_0.Vout a_8706_51119# 0.04444f
C2441 a_2209_61411# EN 0.02636f
C2442 a_2046_51119# VDD 0.02521f
C2443 D_FlipFlop_4.Inverter_1.Vout a_10808_48405# 0.04995f
C2444 a_23593_60797# CLK 0.06211f
C2445 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.06955f
C2446 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_n7633_55365# 0.04995f
C2447 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_17315_54751# 0.04444f
C2448 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_2.Qbar 0.11657f
C2449 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_16465_54751# 0.04444f
C2450 D_FlipFlop_2.3-input-nand_1.B VDD 1.34831f
C2451 a_49391_54751# VDD 0.02521f
C2452 D_FlipFlop_6.nPRE a_5773_58825# 0.05925f
C2453 a_n10790_51119# VDD 0.02521f
C2454 a_24443_58825# Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.05964f
C2455 a_24443_59439# CLK 0.03166f
C2456 a_52105_55365# a_52105_54751# 0.05935f
C2457 a_49391_60797# VDD 0.02521f
C2458 D_FlipFlop_5.3-input-nand_2.Vout VDD 2.67043f
C2459 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout EN 0.78583f
C2460 a_23593_61411# a_23593_60797# 0.05935f
C2461 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.01194f
C2462 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C VDD 3.50703f
C2463 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.01194f
C2464 a_13751_58825# CLK 0.03f
C2465 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.10915f
C2466 D_FlipFlop_1.3-input-nand_2.C a_43140_48405# 0.01335f
C2467 And_Gate_4.A VDD 1.33669f
C2468 a_34285_59439# a_34285_58825# 0.05935f
C2469 a_12901_54751# VDD 0.02521f
C2470 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout CLK 0.12427f
C2471 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C2472 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout EN 0.09223f
C2473 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.07084f
C2474 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout EN 0.96763f
C2475 a_45827_54751# VDD 0.02521f
C2476 a_27157_61411# EN 0.02636f
C2477 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout a_n1355_56723# 0.04443f
C2478 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.26069f
C2479 a_48541_60797# CLK 0.06211f
C2480 a_45827_56723# VDD 0.02578f
C2481 Ring_Counter_0.D_FlipFlop_16.Q a_17315_60797# 0.01768f
C2482 D_FlipFlop_0.3-input-nand_0.Vout a_52516_51119# 0.04444f
C2483 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C EN 0.07517f
C2484 D_FlipFlop_7.Inverter_1.Vout a_n6716_51119# 0.04443f
C2485 a_20029_59439# VDD 0.01186f
C2486 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout a_20029_59439# 0.01335f
C2487 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.06935f
C2488 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B a_49391_60797# 0.04443f
C2489 D_FlipFlop_1.Qbar VDD 1.96179f
C2490 a_38699_61411# a_38699_60797# 0.05935f
C2491 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout a_37849_60797# 0.05964f
C2492 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout EN 0.61231f
C2493 a_9337_58825# VDD 0.02521f
C2494 a_13751_59439# a_13751_58825# 0.05935f
C2495 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.01194f
C2496 a_9337_54751# VDD 0.02521f
C2497 a_8092_48405# VDD 0.0123f
C2498 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C CLK 0.19664f
C2499 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C2500 D_FlipFlop_2.3-input-nand_2.C VDD 2.67826f
C2501 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.Inverter_1.Vout 0.06895f
C2502 a_n505_59439# VDD 0.05686f
C2503 a_2209_56723# VDD 0.02521f
C2504 And_Gate_1.A And_Gate_1.Nand_Gate_0.Vout 0.24482f
C2505 a_42263_54751# VDD 0.02521f
C2506 D_FlipFlop_7.nPRE D_FlipFlop_7.CLK 0.1668f
C2507 a_3059_58825# Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.04443f
C2508 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_9337_56723# 0.05964f
C2509 D_FlipFlop_6.Qbar D_FlipFlop_6.Nand_Gate_1.Vout 0.11654f
C2510 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout a_30721_58825# 0.04444f
C2511 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout EN 0.08731f
C2512 a_52105_61411# EN 0.04454f
C2513 a_48541_55365# a_48541_54751# 0.05935f
C2514 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.20923f
C2515 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout a_48541_56723# 0.04443f
C2516 a_55976_51119# Q7 0.01335f
C2517 CDAC_v3_0.OUT m3_3428_38799# 1.25228f
C2518 D_FlipFlop_2.CLK a_33020_48405# 0.04443f
C2519 Ring_Counter_0.D_FlipFlop_16.Q a_42263_60797# 0.01768f
C2520 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C a_12901_58825# 0.04443f
C2521 a_5773_54751# VDD 0.02521f
C2522 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_7.Z 0.05555f
C2523 CDAC_v3_0.switch_2.Z CDAC_v3_0.switch_4.Z 21.4938f
C2524 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_5.Z 0.10871f
C2525 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B VDD 1.71455f
C2526 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.01764f
C2527 a_6623_59439# Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.01335f
C2528 D_FlipFlop_2.Inverter_1.Vout a_37094_51119# 0.04443f
C2529 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.04107f
C2530 a_48541_61411# a_48541_60797# 0.05935f
C2531 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout 0.06935f
C2532 a_38699_54751# VDD 0.02521f
C2533 D_FlipFlop_6.CLK a_n670_48405# 0.02953f
C2534 And_Gate_5.A a_36806_52049# 0.05964f
C2535 CDAC_v3_0.switch_0.Z VDD 1.31192f
C2536 a_10187_61411# VDD 0.04448f
C2537 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B VDD 1.71455f
C2538 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout a_5773_61411# 0.01335f
C2539 D_FlipFlop_7.Qbar a_n5358_48405# 0.01335f
C2540 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C a_3059_56723# 0.04443f
C2541 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.Nand_Gate_0.Vout 0.16429f
C2542 Nand_Gate_7.A a_54330_52049# 0.0451f
C2543 D_FlipFlop_2.nPRE D_FlipFlop_2.3-input-nand_1.B 0.27142f
C2544 D_FlipFlop_4.CLK CLK 0.07954f
C2545 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B EN 0.3979f
C2546 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.Inverter_1.Vout 0.26069f
C2547 a_8092_51119# D_FlipFlop_4.3-input-nand_2.Vout 0.01335f
C2548 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_24443_55365# 0.04995f
C2549 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout a_49391_54751# 0.04444f
C2550 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_23593_55365# 0.04995f
C2551 a_3404_51119# VDD 0.01186f
C2552 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 1.09973f
C2553 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout VDD 2.07898f
C2554 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_48541_54751# 0.04444f
C2555 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.Inverter_1.Vout 0.06895f
C2556 D_FlipFlop_2.3-input-nand_2.C a_37094_48405# 0.04443f
C2557 a_2209_54751# VDD 0.02521f
C2558 D_FlipFlop_3.nPRE D_FlipFlop_5.Qbar 0.01961f
C2559 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.04109f
C2560 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.06955f
C2561 a_n9432_51119# VDD 0.01186f
C2562 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout CLK 0.7779f
C2563 D_FlipFlop_6.nPRE a_n2642_48405# 0.0452f
C2564 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout CLK 0.36346f
C2565 D_FlipFlop_2.3-input-nand_1.Vout a_33020_48405# 0.05964f
C2566 a_35135_54751# VDD 0.02521f
C2567 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B VDD 1.71455f
C2568 D_FlipFlop_4.3-input-nand_1.Vout a_8706_48405# 0.04444f
C2569 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.01194f
C2570 a_28332_51119# D_FlipFlop_3.Nand_Gate_0.Vout 0.05964f
C2571 CDAC_v3_0.switch_0.Z Q4 0.02962f
C2572 a_44977_55365# a_44977_54751# 0.05935f
C2573 a_35135_61411# VDD 0.04448f
C2574 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout 0.06935f
C2575 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B EN 0.3979f
C2576 a_n1355_54751# VDD 0.02521f
C2577 And_Gate_7.Nand_Gate_0.Vout a_49577_52049# 0.05964f
C2578 D_FlipFlop_1.nPRE D_FlipFlop_1.3-input-nand_2.Vout 0.76528f
C2579 D_FlipFlop_6.nPRE D_FlipFlop_7.Qbar 0.01961f
C2580 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.07084f
C2581 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.Nand_Gate_0.Vout 0.16429f
C2582 D_FlipFlop_3.3-input-nand_2.Vout a_26230_48405# 0.04443f
C2583 a_15496_51119# D_FlipFlop_5.3-input-nand_0.Vout 0.05964f
C2584 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout a_13751_59439# 0.04543f
C2585 a_51902_51119# D_FlipFlop_0.3-input-nand_2.Vout 0.01335f
C2586 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.Inverter_1.Vout 0.26069f
C2587 a_31571_54751# VDD 0.02521f
C2588 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout CLK 0.7779f
C2589 CDAC_v3_0.switch_5.Z Q5 0.17562f
C2590 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.48403f
C2591 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK 0.36346f
C2592 D_FlipFlop_2.nPRE D_FlipFlop_2.3-input-nand_2.C 0.05823f
C2593 Nand_Gate_6.A a_20029_55365# 0.01335f
C2594 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B a_3059_61411# 0.04995f
C2595 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B VDD 1.71455f
C2596 D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.43587f
C2597 a_26230_48405# VDD 0.02521f
C2598 Ring_Counter_0.D_FlipFlop_16.Q a_3059_61411# 0.01252f
C2599 Ring_Counter_0.D_FlipFlop_16.Q VDD 24.0851f
C2600 VDD Q5 3.73573f
C2601 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B EN 0.3979f
C2602 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.04107f
C2603 D_FlipFlop_2.3-input-nand_0.Vout VDD 1.74442f
C2604 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout a_30721_61411# 0.01335f
C2605 a_n4919_54751# VDD 0.02521f
C2606 a_49577_52049# VDD 0.02521f
C2607 a_28007_54751# VDD 0.02521f
C2608 D_FlipFlop_5.Inverter_1.Vout a_19570_48405# 0.04995f
C2609 D_FlipFlop_4.nPRE D_FlipFlop_4.Inverter_1.Vout 0.07033f
C2610 Nand_Gate_1.A a_n4919_56723# 0.05925f
C2611 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B 0.02535f
C2612 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.10915f
C2613 Nand_Gate_6.A a_16465_55365# 0.05925f
C2614 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B VDD 1.71455f
C2615 a_35430_45397# CDAC_v3_0.switch_6.Z 0.27006f
C2616 a_41413_55365# a_41413_54751# 0.05935f
C2617 D_FlipFlop_7.3-input-nand_1.Vout a_n11404_48405# 0.01335f
C2618 D_FlipFlop_3.nPRE Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B 0.29684f
C2619 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B 0.45531f
C2620 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B EN 0.27162f
C2621 a_40815_52049# CLK 0.04479f
C2622 Ring_Counter_0.D_FlipFlop_16.Q a_28007_61411# 0.01252f
C2623 Q4 Q5 1.34643f
C2624 a_52105_56723# VDD 0.02865f
C2625 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_12.Qbar 0.07122f
C2626 D_FlipFlop_4.nPRE a_10520_52049# 0.04597f
C2627 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.01194f
C2628 D_FlipFlop_0.3-input-nand_2.C a_51902_48405# 0.01335f
C2629 D_FlipFlop_5.CLK D_FlipFlop_5.Inverter_1.Vout 0.20785f
C2630 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_34285_56723# 0.05964f
C2631 a_24443_54751# VDD 0.02521f
C2632 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout EN 0.08727f
C2633 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.26069f
C2634 a_n4919_60797# VDD 0.02521f
C2635 And_Gate_1.Nand_Gate_0.Vout CLK 0.79128f
C2636 And_Gate_4.Nand_Gate_0.Vout D_FlipFlop_3.CLK 0.25559f
C2637 Nand_Gate_3.A a_23593_60797# 0.10368f
C2638 D_FlipFlop_4.nPRE And_Gate_2.A 0.37487f
C2639 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.Nand_Gate_1.Vout 0.1541f
C2640 D_FlipFlop_0.Nand_Gate_1.Vout a_56590_48405# 0.04444f
C2641 D_FlipFlop_2.nPRE a_35135_54751# 0.05987f
C2642 D_FlipFlop_1.nPRE a_41168_48405# 0.0452f
C2643 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout a_48541_58825# 0.05964f
C2644 a_n8818_48405# VDD 0.02521f
C2645 D_FlipFlop_6.CLK a_n2028_51119# 0.04443f
C2646 a_13751_56723# Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.05964f
C2647 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout a_n4069_58825# 0.04444f
C2648 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout a_9337_56723# 0.04443f
C2649 a_n505_60797# CLK 0.06211f
C2650 D_FlipFlop_3.Nand_Gate_0.Vout a_29690_51119# 0.04543f
C2651 a_20879_54751# VDD 0.02521f
C2652 And_Gate_7.Nand_Gate_0.Vout EN 0.01133f
C2653 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.20923f
C2654 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.01323f
C2655 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout VDD 2.8343f
C2656 CDAC_v3_0.switch_8.Z Q0 0.18158f
C2657 Nand_Gate_2.A a_12901_55365# 0.01335f
C2658 a_13751_60797# Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.05964f
C2659 D_FlipFlop_6.CLK VDD 2.17721f
C2660 a_37849_55365# a_37849_54751# 0.05935f
C2661 D_FlipFlop_6.nPRE And_Gate_2.A 0.01015f
C2662 a_20029_60797# VDD 0.02521f
C2663 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.1143f
C2664 a_7822_45397# CDAC_v3_0.switch_8.Z 0.28688f
C2665 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.04109f
C2666 D_FlipFlop_2.3-input-nand_2.Vout Q6 0.01377f
C2667 D_FlipFlop_5.3-input-nand_0.Vout a_16854_51119# 0.04543f
C2668 Nand_Gate_1.A And_Gate_0.A 0.07559f
C2669 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C2670 And_Gate_4.A a_28044_52049# 0.05964f
C2671 D_FlipFlop_2.nPRE Q5 0.0494f
C2672 D_FlipFlop_7.nPRE a_n1355_56723# 0.05925f
C2673 a_45856_48405# VDD 0.02521f
C2674 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.01262f
C2675 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout a_49391_59439# 0.04543f
C2676 D_FlipFlop_1.nPRE a_44977_54751# 0.06113f
C2677 D_FlipFlop_2.nPRE D_FlipFlop_2.3-input-nand_0.Vout 0.94459f
C2678 a_56590_48405# Q7 0.06303f
C2679 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.29165f
C2680 a_47828_51119# VDD 0.02521f
C2681 a_28007_56723# VDD 0.02578f
C2682 a_35135_58825# Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.05964f
C2683 a_17315_54751# VDD 0.02521f
C2684 a_45827_59439# CLK 0.03166f
C2685 a_6120_51119# VDD 0.01186f
C2686 a_3059_61411# EN 0.07048f
C2687 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C 0.08674f
C2688 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout EN 0.78543f
C2689 VDD EN 80.3866f
C2690 a_24443_60797# CLK 0.06211f
C2691 D_FlipFlop_2.CLK Q6 0.04416f
C2692 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_16.Qbar 0.11657f
C2693 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C VDD 3.50703f
C2694 Nand_Gate_2.A a_9337_59439# 0.05925f
C2695 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.01194f
C2696 D_FlipFlop_3.3-input-nand_1.B D_FlipFlop_3.3-input-nand_1.Vout 0.08641f
C2697 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C 0.01194f
C2698 a_34992_51119# VDD 0.02521f
C2699 Nand_Gate_2.A a_9337_55365# 0.05925f
C2700 a_35135_58825# CLK 0.03f
C2701 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout EN 0.61231f
C2702 D_FlipFlop_6.Qbar a_3404_48405# 0.01335f
C2703 a_44977_59439# a_44977_58825# 0.05935f
C2704 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_16.Q 0.15834f
C2705 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B 0.02535f
C2706 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout CLK 0.12427f
C2707 D_FlipFlop_7.nPRE D_FlipFlop_7.Nand_Gate_0.Vout 0.5831f
C2708 a_44977_60797# VDD 0.02521f
C2709 D_FlipFlop_4.Nand_Gate_1.Vout a_12166_48405# 0.04995f
C2710 D_FlipFlop_0.Qbar EN 0.03748f
C2711 D_FlipFlop_1.nPRE a_41413_54751# 0.05925f
C2712 D_FlipFlop_1.3-input-nand_2.C a_45856_48405# 0.04443f
C2713 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout EN 0.08727f
C2714 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.08462f
C2715 a_13751_54751# VDD 0.02521f
C2716 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.Nand_Gate_1.Vout 0.1541f
C2717 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C EN 0.07565f
C2718 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.30156f
C2719 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.10915f
C2720 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout a_23593_59439# 0.04995f
C2721 a_41413_59439# VDD 0.01186f
C2722 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout a_30721_59439# 0.01335f
C2723 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B EN 0.33743f
C2724 a_28007_61411# EN 0.07048f
C2725 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_3.Qbar 0.07122f
C2726 a_34285_55365# a_34285_54751# 0.05935f
C2727 a_49391_60797# CLK 0.06211f
C2728 And_Gate_6.Nand_Gate_0.Vout a_40815_52049# 0.05964f
C2729 a_30721_58825# VDD 0.02521f
C2730 a_24443_59439# a_24443_58825# 0.05935f
C2731 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C CLK 0.20012f
C2732 Nand_Gate_2.A a_9337_60797# 0.10368f
C2733 D_FlipFlop_2.3-input-nand_1.Vout Q6 0.02179f
C2734 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.10915f
C2735 a_41168_48405# a_41782_48405# 0.05935f
C2736 a_20879_59439# VDD 0.05686f
C2737 Ring_Counter_0.D_FlipFlop_16.Q a_12901_60797# 0.01768f
C2738 And_Gate_4.A CLK 1.52489f
C2739 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.25966f
C2740 a_38699_60797# Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.05964f
C2741 a_10187_58825# VDD 0.02578f
C2742 a_13751_58825# Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.04443f
C2743 a_10187_54751# VDD 0.02521f
C2744 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_1.Vout 0.08671f
C2745 a_10808_48405# VDD 0.02521f
C2746 a_12901_59439# EN 0.045f
C2747 D_FlipFlop_2.3-input-nand_2.Vout a_34992_48405# 0.04443f
C2748 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout VDD 2.07898f
C2749 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout VDD 2.8343f
C2750 Nand_Gate_0.A a_5773_55365# 0.01335f
C2751 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C a_31571_56723# 0.04443f
C2752 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C a_23593_58825# 0.04443f
C2753 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.01202f
C2754 a_n7004_52049# VDD 0.02521f
C2755 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout a_31571_58825# 0.04444f
C2756 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B 0.02535f
C2757 a_29690_51119# a_30304_51119# 0.05935f
C2758 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout EN 0.08727f
C2759 D_FlipFlop_2.CLK a_34992_48405# 0.02953f
C2760 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout VDD 2.29929f
C2761 CDAC_v3_0.OUT m3_3428_9615# 1.25228f
C2762 a_17315_59439# Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 0.01335f
C2763 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.15413f
C2764 a_6623_54751# VDD 0.02521f
C2765 Ring_Counter_0.D_FlipFlop_16.Q a_37849_60797# 0.01768f
C2766 D_FlipFlop_1.3-input-nand_2.Vout Q7 0.01585f
C2767 D_FlipFlop_7.3-input-nand_1.B D_FlipFlop_7.3-input-nand_1.Vout 0.08641f
C2768 a_n505_59439# CLK 0.03166f
C2769 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_4.Z 5.93382f
C2770 CDAC_v3_0.switch_8.Z CDAC_v3_0.switch_6.Z 0.19987f
C2771 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_7.Z 0.06747f
C2772 And_Gate_0.Nand_Gate_0.Vout VDD 1.42724f
C2773 D_FlipFlop_6.3-input-nand_2.Vout a_2046_51119# 0.04443f
C2774 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C VDD 3.50703f
C2775 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 1.09973f
C2776 a_16854_51119# a_17468_51119# 0.05935f
C2777 D_FlipFlop_3.Inverter_1.Vout a_28332_48405# 0.04995f
C2778 Nand_Gate_0.A a_2209_55365# 0.05925f
C2779 a_6623_61411# Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.01335f
C2780 a_30721_55365# a_30721_54751# 0.05935f
C2781 D_FlipFlop_3.CLK D_FlipFlop_3.3-input-nand_1.Vout 0.67419f
C2782 CDAC_v3_0.switch_2.Z VDD 1.09756f
C2783 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.25966f
C2784 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout VDD 2.72531f
C2785 D_FlipFlop_2.nPRE EN 0.79742f
C2786 a_38699_56723# Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.05964f
C2787 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.30048f
C2788 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD 1.89599f
C2789 Nand_Gate_5.A Nand_Gate_7.A 0.04584f
C2790 a_35430_45397# Q7 0.46416f
C2791 a_5773_61411# VDD 0.08862f
C2792 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout EN 0.61998f
C2793 D_FlipFlop_1.CLK D_FlipFlop_1.3-input-nand_2.Vout 0.1192f
C2794 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_n505_54751# 0.04444f
C2795 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout 0.01202f
C2796 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_7.Qbar 0.11657f
C2797 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_n1355_54751# 0.04444f
C2798 D_FlipFlop_4.3-input-nand_1.B VDD 1.3477f
C2799 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.09856f
C2800 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout a_5773_58825# 0.04444f
C2801 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD 1.48403f
C2802 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.16431f
C2803 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B CLK 0.08407f
C2804 a_23644_48405# a_24258_48405# 0.05935f
C2805 a_3059_54751# VDD 0.02521f
C2806 D_FlipFlop_7.3-input-nand_2.Vout VDD 2.67043f
C2807 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B EN 0.3979f
C2808 And_Gate_1.A D_FlipFlop_6.CLK 0.06897f
C2809 D_FlipFlop_2.3-input-nand_1.Vout a_34992_48405# 0.04444f
C2810 a_n4919_59439# VDD 0.01186f
C2811 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B CLK 0.08407f
C2812 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B a_31571_61411# 0.04995f
C2813 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout a_2209_58825# 0.05964f
C2814 D_FlipFlop_1.nPRE a_40815_52049# 0.02193f
C2815 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout VDD 2.72531f
C2816 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B 0.02535f
C2817 D_FlipFlop_1.3-input-nand_2.Vout a_45856_51119# 0.04443f
C2818 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD 1.89599f
C2819 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B a_20879_61411# 0.04995f
C2820 a_30721_61411# VDD 0.08862f
C2821 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B a_42263_60797# 0.04443f
C2822 a_23644_51119# D_FlipFlop_3.3-input-nand_0.Vout 0.01335f
C2823 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_1.Vout 0.08671f
C2824 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.25936f
C2825 a_n505_54751# VDD 0.02521f
C2826 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.Vout 1.01753f
C2827 Nand_Gate_3.A a_27157_54751# 0.06359f
C2828 D_FlipFlop_5.Qbar VDD 1.96371f
C2829 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.06955f
C2830 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B CLK 0.08407f
C2831 Nand_Gate_1.A a_n1355_55365# 0.01335f
C2832 a_27157_55365# a_27157_54751# 0.05935f
C2833 And_Gate_3.A a_19282_52049# 0.05964f
C2834 a_34285_56723# VDD 0.02521f
C2835 Nand_Gate_5.A a_37849_58825# 0.05925f
C2836 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.08582f
C2837 a_50544_51119# VDD 0.02521f
C2838 a_55976_48405# EN 0.04443f
C2839 And_Gate_5.A And_Gate_5.Nand_Gate_0.Vout 0.24482f
C2840 a_29690_48405# VDD 0.01186f
C2841 D_FlipFlop_4.3-input-nand_2.C VDD 2.67765f
C2842 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.0646f
C2843 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.06462f
C2844 Nand_Gate_7.A And_Gate_7.A 0.11778f
C2845 Ring_Counter_0.D_FlipFlop_16.Q a_n1355_61411# 0.01252f
C2846 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.1143f
C2847 a_31571_61411# Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.01335f
C2848 a_n4069_54751# VDD 0.02521f
C2849 D_FlipFlop_5.nPRE a_19282_52049# 0.04597f
C2850 a_6120_48405# a_6734_48405# 0.05935f
C2851 Nand_Gate_3.A a_23593_54751# 0.05925f
C2852 D_FlipFlop_3.CLK D_FlipFlop_3.3-input-nand_1.B 0.06986f
C2853 D_FlipFlop_5.3-input-nand_1.Vout a_14882_48405# 0.01335f
C2854 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.07084f
C2855 Nand_Gate_1.A a_n4919_55365# 0.0598f
C2856 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B CLK 0.08407f
C2857 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.17551f
C2858 a_n1355_59439# a_n1355_58825# 0.05935f
C2859 Ring_Counter_0.D_FlipFlop_16.Q CLK 7.36469f
C2860 a_15710_45397# Q2 0.47258f
C2861 And_Gate_3.A VDD 1.34057f
C2862 D_FlipFlop_4.Qbar a_12166_48405# 0.01335f
C2863 D_FlipFlop_7.3-input-nand_1.Vout a_n9432_48405# 0.04543f
C2864 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B 0.02535f
C2865 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout a_37849_56723# 0.04443f
C2866 Nand_Gate_5.A And_Gate_6.A 0.1048f
C2867 D_FlipFlop_4.CLK a_6734_48405# 0.04443f
C2868 a_49577_52049# CLK 0.04479f
C2869 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.0646f
C2870 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.06462f
C2871 a_n7633_54751# VDD 0.02521f
C2872 Ring_Counter_0.D_FlipFlop_16.Q a_23593_61411# 0.01252f
C2873 And_Gate_5.Nand_Gate_0.Vout a_32053_52049# 0.05964f
C2874 D_FlipFlop_0.3-input-nand_2.C a_54618_48405# 0.04443f
C2875 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_6623_55365# 0.04995f
C2876 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout 0.06837f
C2877 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_31571_54751# 0.04444f
C2878 D_FlipFlop_5.nPRE VDD 7.38458f
C2879 D_FlipFlop_5.nPRE Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.1091f
C2880 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_5773_55365# 0.04995f
C2881 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_30721_54751# 0.04444f
C2882 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.01202f
C2883 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout EN 0.08727f
C2884 a_23593_55365# a_23593_54751# 0.05935f
C2885 a_n505_61411# a_n505_60797# 0.05935f
C2886 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B CLK 0.08407f
C2887 a_n4069_60797# VDD 0.02865f
C2888 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout a_n1355_60797# 0.05964f
C2889 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.01262f
C2890 a_39066_48405# Q5 0.05747f
C2891 Nand_Gate_7.A Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.29165f
C2892 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B VDD 1.71455f
C2893 D_FlipFlop_2.Inverter_1.Vout VDD 1.70303f
C2894 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C a_n7633_56723# 0.04443f
C2895 a_10187_56723# VDD 0.02578f
C2896 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout a_41413_58825# 0.04444f
C2897 a_n5358_48405# VDD 0.01186f
C2898 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.26069f
C2899 Nand_Gate_1.A a_n4919_61411# 0.04995f
C2900 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.01162f
C2901 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B VDD 1.71455f
C2902 Nand_Gate_4.A And_Gate_5.A 0.08451f
C2903 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.01262f
C2904 D_FlipFlop_3.CLK D_FlipFlop_3.3-input-nand_2.C 0.19377f
C2905 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.29165f
C2906 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout EN 0.61231f
C2907 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Qbar 0.06863f
C2908 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B a_6623_61411# 0.04995f
C2909 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.25864f
C2910 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout VDD 2.29929f
C2911 a_n4919_60797# CLK 0.06211f
C2912 a_n11404_48405# a_n10790_48405# 0.05935f
C2913 D_FlipFlop_4.nPRE VDD 7.59422f
C2914 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout 0.15416f
C2915 D_FlipFlop_1.3-input-nand_2.Vout a_43754_48405# 0.04443f
C2916 Ring_Counter_0.D_FlipFlop_16.Q a_48541_61411# 0.01252f
C2917 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.25966f
C2918 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.1143f
C2919 a_45827_58825# Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.05964f
C2920 a_20879_60797# VDD 0.02865f
C2921 D_FlipFlop_2.nPRE a_34285_56723# 0.05925f
C2922 a_9337_61411# a_9337_60797# 0.05935f
C2923 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout EN 0.78583f
C2924 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.3-input-nand_2.Vout 0.0846f
C2925 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.10034f
C2926 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.01194f
C2927 D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.43587f
C2928 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.01194f
C2929 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.16917f
C2930 Nand_Gate_3.A And_Gate_4.A 0.07694f
C2931 a_47828_48405# VDD 0.02521f
C2932 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout 0.06955f
C2933 a_51902_51119# VDD 0.01186f
C2934 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout 0.26069f
C2935 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C 0.01323f
C2936 D_FlipFlop_4.3-input-nand_0.Vout VDD 1.74442f
C2937 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout CLK 0.12427f
C2938 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout EN 0.09223f
C2939 D_FlipFlop_6.nPRE VDD 7.57772f
C2940 D_FlipFlop_6.CLK CLK 0.07954f
C2941 a_20029_55365# a_20029_54751# 0.05935f
C2942 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout EN 0.96763f
C2943 a_n1355_61411# EN 0.02636f
C2944 D_FlipFlop_2.Inverter_1.Vout a_37094_48405# 0.04995f
C2945 a_20029_60797# CLK 0.06211f
C2946 VDD Q1 3.68472f
C2947 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Qbar 0.06863f
C2948 D_FlipFlop_2.Nand_Gate_1.Vout a_38452_48405# 0.04995f
C2949 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C EN 0.07565f
C2950 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout a_41413_59439# 0.01335f
C2951 a_24443_61411# a_24443_60797# 0.05935f
C2952 a_45827_60797# VDD 0.02865f
C2953 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout a_23593_60797# 0.05964f
C2954 D_FlipFlop_1.nPRE a_42263_54751# 0.05987f
C2955 EN CLK 3.62392f
C2956 D_FlipFlop_0.CLK EN 0.70896f
C2957 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C 0.07084f
C2958 a_52105_58825# VDD 0.02865f
C2959 a_35135_59439# a_35135_58825# 0.05935f
C2960 D_FlipFlop_6.nPRE Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout 0.06837f
C2961 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.04109f
C2962 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C CLK 0.19664f
C2963 D_FlipFlop_4.nPRE a_12901_59439# 0.05925f
C2964 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout a_24443_59439# 0.04543f
C2965 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.3-input-nand_2.C 0.06863f
C2966 D_FlipFlop_7.nPRE VDD 7.70785f
C2967 a_42263_59439# VDD 0.05686f
C2968 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout 0.25855f
C2969 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.08674f
C2970 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout EN 0.09223f
C2971 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout a_3059_56723# 0.04995f
C2972 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_38699_55365# 0.04995f
C2973 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout EN 0.96763f
C2974 a_31571_58825# VDD 0.02578f
C2975 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_37849_55365# 0.04995f
C2976 a_23593_61411# EN 0.02636f
C2977 a_24443_58825# Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.04443f
C2978 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.25966f
C2979 a_44977_60797# CLK 0.06211f
C2980 a_34285_59439# EN 0.045f
C2981 Ring_Counter_0.D_FlipFlop_0.Qbar a_52105_54751# 0.04443f
C2982 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout VDD 2.8343f
C2983 D_FlipFlop_4.nPRE a_12166_51119# 0.04443f
C2984 Ring_Counter_0.D_FlipFlop_16.Q a_13751_60797# 0.01768f
C2985 D_FlipFlop_2.nPRE D_FlipFlop_2.Inverter_1.Vout 0.07033f
C2986 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.15413f
C2987 And_Gate_2.A a_10520_52049# 0.05964f
C2988 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C a_34285_58825# 0.04443f
C2989 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B 0.29684f
C2990 a_12780_48405# VDD 0.02521f
C2991 a_16465_55365# a_16465_54751# 0.05935f
C2992 D_FlipFlop_3.nPRE a_25616_51119# 0.045f
C2993 a_34285_61411# a_34285_60797# 0.05935f
C2994 a_28007_59439# Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 0.01335f
C2995 D_FlipFlop_3.nPRE a_27157_58825# 0.05925f
C2996 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.08462f
C2997 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD 1.48403f
C2998 D_FlipFlop_6.CLK D_FlipFlop_6.3-input-nand_2.Vout 0.1192f
C2999 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout a_n1355_59439# 0.04995f
C3000 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout 0.06935f
C3001 a_48541_55365# EN 0.04443f
C3002 D_FlipFlop_3.CLK D_FlipFlop_3.3-input-nand_0.Vout 0.25957f
C3003 D_FlipFlop_7.Qbar a_n4744_51119# 0.04443f
C3004 a_20879_59439# CLK 0.03223f
C3005 a_1758_52049# VDD 0.02521f
C3006 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout EN 0.78583f
C3007 a_49391_55365# a_49391_54751# 0.05935f
C3008 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout EN 0.08617f
C3009 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C 1.09565f
C3010 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.16431f
C3011 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C VDD 3.50621f
C3012 a_48541_61411# EN 0.0434f
C3013 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout EN 0.08727f
C3014 a_10187_58825# CLK 0.03f
C3015 a_n11404_51119# a_n10790_51119# 0.05935f
C3016 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout a_n1355_56723# 0.04443f
C3017 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout 0.25855f
C3018 D_FlipFlop_7.Nand_Gate_1.Vout a_n6716_48405# 0.05964f
C3019 Ring_Counter_0.D_FlipFlop_16.Q a_38699_60797# 0.01768f
C3020 CDAC_v3_0.switch_0.Z CDAC_v3_0.switch_6.Z 2.4235f
C3021 CDAC_v3_0.switch_2.Z CDAC_v3_0.switch_7.Z 0.0599f
C3022 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout CLK 0.12427f
C3023 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_5.Z 21.0253f
C3024 D_FlipFlop_6.nPRE a_n670_51119# 0.045f
C3025 a_49391_61411# a_49391_60797# 0.05935f
C3026 Nand_Gate_5.A a_37849_61411# 0.04995f
C3027 a_17468_51119# D_FlipFlop_5.3-input-nand_2.Vout 0.05964f
C3028 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout a_48541_60797# 0.05964f
C3029 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.06734f
C3030 a_21542_51119# VDD 0.02521f
C3031 CDAC_v3_0.switch_3.Z VDD 1.07516f
C3032 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.01194f
C3033 a_44977_55365# EN 0.04443f
C3034 And_Gate_4.Nand_Gate_0.Vout a_23291_52049# 0.05964f
C3035 a_6623_61411# VDD 0.04448f
C3036 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout CLK 0.20785f
C3037 D_FlipFlop_5.Qbar a_20928_48405# 0.01335f
C3038 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout EN 0.61231f
C3039 Ring_Counter_0.D_FlipFlop_1.Qbar a_48541_54751# 0.04443f
C3040 a_8706_51119# VDD 0.02521f
C3041 D_FlipFlop_3.nPRE a_27157_61411# 0.04995f
C3042 a_16465_59439# VDD 0.01186f
C3043 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout a_6623_58825# 0.04444f
C3044 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout 0.30046f
C3045 And_Gate_0.Nand_Gate_0.Vout CLK 0.47616f
C3046 a_16465_56723# VDD 0.02521f
C3047 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout a_12901_58825# 0.05964f
C3048 a_5773_58825# VDD 0.02521f
C3049 Nand_Gate_5.A Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.12285f
C3050 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C CLK 0.19664f
C3051 a_12901_55365# a_12901_54751# 0.05935f
C3052 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout 0.01202f
C3053 D_FlipFlop_2.Qbar a_39066_51119# 0.04443f
C3054 D_FlipFlop_1.nPRE D_FlipFlop_1.Nand_Gate_0.Vout 0.5831f
C3055 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout CLK 0.7779f
C3056 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_16465_56723# 0.05964f
C3057 a_n4069_59439# VDD 0.05686f
C3058 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout CLK 0.36346f
C3059 D_FlipFlop_4.nPRE a_12901_60797# 0.10368f
C3060 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C3061 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.08582f
C3062 D_FlipFlop_6.CLK Q0 0.01146f
C3063 a_41413_55365# EN 0.04443f
C3064 a_32406_51119# a_33020_51119# 0.05935f
C3065 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C3066 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout CLK 0.23546f
C3067 a_45827_55365# a_45827_54751# 0.05935f
C3068 D_FlipFlop_7.3-input-nand_1.B a_n10790_48405# 0.04443f
C3069 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.04107f
C3070 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_8.Qbar 0.07122f
C3071 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.08582f
C3072 D_FlipFlop_3.3-input-nand_2.C a_26230_51119# 0.04443f
C3073 a_n4069_56723# Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.05964f
C3074 a_31571_61411# VDD 0.04448f
C3075 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout a_16465_61411# 0.01335f
C3076 D_FlipFlop_7.CLK VDD 2.17721f
C3077 D_FlipFlop_6.nPRE And_Gate_1.A 0.36235f
C3078 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C 0.08674f
C3079 D_FlipFlop_0.3-input-nand_2.Vout a_52516_48405# 0.04443f
C3080 a_37849_55365# EN 0.04443f
C3081 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout VDD 2.07898f
C3082 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout CLK 0.7779f
C3083 a_n505_58825# Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C 0.05964f
C3084 a_32406_48405# VDD 0.01186f
C3085 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK 0.36346f
C3086 Ring_Counter_0.D_FlipFlop_2.Qbar a_44977_54751# 0.04443f
C3087 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.04109f
C3088 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.01194f
C3089 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C 0.01194f
C3090 Ring_Counter_0.D_FlipFlop_16.Q a_n505_61411# 0.01252f
C3091 Nand_Gate_2.A a_9337_56723# 0.05925f
C3092 a_9337_59439# a_9337_58825# 0.05935f
C3093 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.01194f
C3094 D_FlipFlop_1.3-input-nand_1.Vout a_41168_48405# 0.01335f
C3095 a_21542_48405# Q3 0.06021f
C3096 a_9337_55365# a_9337_54751# 0.05935f
C3097 D_FlipFlop_7.nPRE And_Gate_1.A 0.02188f
C3098 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.08462f
C3099 a_n7633_56723# VDD 0.02578f
C3100 D_FlipFlop_5.nPRE a_14882_51119# 0.034f
C3101 Nand_Gate_3.A a_24443_54751# 0.05987f
C3102 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.06734f
C3103 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout a_34285_59439# 0.04995f
C3104 D_FlipFlop_7.Nand_Gate_0.Vout a_n4744_51119# 0.04444f
C3105 D_FlipFlop_0.CLK a_50544_51119# 0.04443f
C3106 D_FlipFlop_5.3-input-nand_1.Vout a_16854_48405# 0.04543f
C3107 D_FlipFlop_1.CLK a_43140_48405# 0.02953f
C3108 a_34285_55365# EN 0.04443f
C3109 D_FlipFlop_1.Inverter_1.Vout a_45856_48405# 0.04995f
C3110 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_9.Qbar 1.27948f
C3111 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.21777f
C3112 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C a_20879_56723# 0.04443f
C3113 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout a_20029_56723# 0.04443f
C3114 a_42263_55365# a_42263_54751# 0.05935f
C3115 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout 0.30046f
C3116 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout a_n4919_59439# 0.01335f
C3117 D_FlipFlop_4.CLK a_8706_48405# 0.02953f
C3118 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout VDD 2.09665f
C3119 Ring_Counter_0.D_FlipFlop_16.Q a_24443_61411# 0.01252f
C3120 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.15413f
C3121 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_12.Qbar 0.11657f
C3122 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.04107f
C3123 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout a_28007_56723# 0.04995f
C3124 a_n505_60797# Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.05964f
C3125 And_Gate_3.A CLK 1.58585f
C3126 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout a_41413_61411# 0.01335f
C3127 And_Gate_5.A D_FlipFlop_2.CLK 0.06897f
C3128 a_30721_55365# EN 0.04443f
C3129 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout EN 0.08727f
C3130 Nand_Gate_6.A Ring_Counter_0.D_FlipFlop_10.Qbar 0.11806f
C3131 And_Gate_1.A a_1758_52049# 0.05964f
C3132 Ring_Counter_0.D_FlipFlop_3.Qbar a_41413_54751# 0.04443f
C3133 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout a_42263_58825# 0.04444f
C3134 Nand_Gate_4.A a_34285_54751# 0.06359f
C3135 a_n2642_48405# VDD 0.01186f
C3136 D_FlipFlop_2.Nand_Gate_0.Vout a_39066_51119# 0.04444f
C3137 D_FlipFlop_2.3-input-nand_2.C Q7 0.0189f
C3138 D_FlipFlop_1.nPRE EN 0.79742f
C3139 D_FlipFlop_5.nPRE CLK 0.9416f
C3140 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.16431f
C3141 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C 0.01323f
C3142 a_5773_55365# a_5773_54751# 0.05935f
C3143 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout a_34285_56723# 0.04443f
C3144 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout 0.26069f
C3145 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.08582f
C3146 a_n4069_60797# CLK 0.06211f
C3147 Nand_Gate_3.A EN 0.79742f
C3148 Ring_Counter_0.D_FlipFlop_16.Q a_49391_61411# 0.01252f
C3149 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout 0.06935f
C3150 a_27157_55365# EN 0.04443f
C3151 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B CLK 0.08407f
C3152 CDAC_v3_0.switch_2.Z Q0 0.02452f
C3153 D_FlipFlop_3.3-input-nand_0.Vout a_26230_51119# 0.04444f
C3154 a_37094_51119# VDD 0.02521f
C3155 D_FlipFlop_4.nPRE a_12901_56723# 0.05925f
C3156 a_38699_55365# a_38699_54751# 0.05935f
C3157 D_FlipFlop_7.Qbar VDD 1.96371f
C3158 Nand_Gate_4.A a_30721_54751# 0.05925f
C3159 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B CLK 0.08407f
C3160 a_11766_45397# CDAC_v3_0.switch_0.Z 0.27828f
C3161 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.16917f
C3162 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout a_2209_56723# 0.04443f
C3163 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout a_42263_56723# 0.04995f
C3164 a_16465_60797# VDD 0.02521f
C3165 D_FlipFlop_2.nPRE a_32406_48405# 0.0452f
C3166 a_24258_51119# VDD 0.02521f
C3167 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_41413_56723# 0.05964f
C3168 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout a_16465_58825# 0.04444f
C3169 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout CLK 0.20785f
C3170 D_FlipFlop_1.nPRE a_41413_59439# 0.05925f
C3171 D_FlipFlop_4.nPRE CLK 0.7408f
C3172 a_50544_48405# VDD 0.02521f
C3173 D_FlipFlop_7.nPRE Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.20928f
C3174 D_FlipFlop_0.3-input-nand_2.Vout VDD 2.77268f
C3175 And_Gate_3.Nand_Gate_0.Vout a_14529_52049# 0.05964f
C3176 CDAC_v3_0.switch_0.Z Q7 0.02962f
C3177 a_23593_55365# EN 0.04443f
C3178 a_n505_61411# EN 0.07048f
C3179 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout a_52105_59439# 0.01335f
C3180 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.01162f
C3181 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.Qbar 1.26888f
C3182 a_20879_60797# CLK 0.06211f
C3183 a_20879_56723# Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.05964f
C3184 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout a_48541_56723# 0.04443f
C3185 Ring_Counter_0.D_FlipFlop_4.Qbar a_37849_54751# 0.04443f
C3186 a_45827_59439# a_45827_58825# 0.05935f
C3187 D_FlipFlop_3.Qbar a_29690_48405# 0.01335f
C3188 D_FlipFlop_5.nPRE D_FlipFlop_5.3-input-nand_1.B 0.27142f
C3189 a_24443_60797# Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.05964f
C3190 a_2209_55365# a_2209_54751# 0.05935f
C3191 a_41413_60797# VDD 0.02521f
C3192 D_FlipFlop_4.Inverter_1.Vout a_10808_51119# 0.04443f
C3193 D_FlipFlop_6.nPRE CLK 0.70812f
C3194 a_35135_58825# Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.04443f
C3195 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.06955f
C3196 a_20029_55365# EN 0.04443f
C3197 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout VDD 2.8343f
C3198 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout 0.04109f
C3199 D_FlipFlop_7.nPRE a_n1355_61411# 0.04995f
C3200 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.10034f
C3201 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_12.Qbar 0.118f
C3202 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_13751_54751# 0.04444f
C3203 a_35135_55365# a_35135_54751# 0.05935f
C3204 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout Ring_Counter_0.D_FlipFlop_3.Qbar 0.11657f
C3205 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_12901_54751# 0.04444f
C3206 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.Inverter_1.Vout 0.06895f
C3207 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C a_44977_58825# 0.04443f
C3208 a_24443_61411# EN 0.07048f
C3209 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout VDD 1.78952f
C3210 a_45827_60797# CLK 0.06211f
C3211 D_FlipFlop_6.3-input-nand_1.B a_n2028_48405# 0.04443f
C3212 a_42263_56723# VDD 0.02578f
C3213 a_38699_59439# Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C 0.01335f
C3214 a_43140_48405# a_43754_48405# 0.05935f
C3215 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout a_27157_56723# 0.04443f
C3216 D_FlipFlop_4.Inverter_1.Vout VDD 1.70303f
C3217 Ring_Counter_0.D_FlipFlop_16.Q a_9337_60797# 0.01768f
C3218 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.30156f
C3219 D_FlipFlop_7.nPRE CLK 0.73874f
C3220 a_42263_59439# CLK 0.03166f
C3221 a_15496_48405# VDD 0.02521f
C3222 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout EN 0.61231f
C3223 D_FlipFlop_3.nPRE D_FlipFlop_3.3-input-nand_2.Vout 0.76528f
C3224 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout EN 0.78583f
C3225 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C 0.07084f
C3226 a_16465_55365# EN 0.04443f
C3227 a_n7633_61411# Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.01335f
C3228 a_2046_51119# D_FlipFlop_6.Nand_Gate_0.Vout 0.05964f
C3229 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C 1.09973f
C3230 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C VDD 3.50703f
C3231 a_31571_58825# CLK 0.03f
C3232 Q5 Q7 0.14098f
C3233 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout a_n505_59439# 0.04543f
C3234 Ring_Counter_0.D_FlipFlop_5.Qbar a_34285_54751# 0.04443f
C3235 a_n1355_56723# VDD 0.02521f
C3236 a_49391_55365# EN 0.04443f
C3237 D_FlipFlop_5.nPRE D_FlipFlop_5.3-input-nand_2.C 0.05823f
C3238 D_FlipFlop_3.nPRE VDD 7.35688f
C3239 D_FlipFlop_0.Inverter_1.Vout a_54618_51119# 0.04443f
C3240 a_10520_52049# VDD 0.02521f
C3241 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout CLK 0.12757f
C3242 D_FlipFlop_5.Nand_Gate_1.Vout a_19570_48405# 0.05964f
C3243 a_49391_54751# Ring_Counter_0.D_FlipFlop_0.Qbar 0.06113f
C3244 a_n1355_55365# a_n1355_54751# 0.05935f
C3245 a_49391_61411# EN 0.04073f
C3246 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.Nand_Gate_0.Vout 0.16429f
C3247 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout EN 0.08727f
C3248 a_n10790_51119# D_FlipFlop_7.3-input-nand_0.Vout 0.05964f
C3249 a_25616_51119# D_FlipFlop_3.3-input-nand_2.Vout 0.01335f
C3250 D_FlipFlop_7.Nand_Gate_1.Vout a_n4744_48405# 0.04444f
C3251 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.Inverter_1.Vout 0.26069f
C3252 a_38452_51119# VDD 0.01186f
C3253 And_Gate_2.A VDD 1.33707f
C3254 CDAC_v3_0.switch_2.Z CDAC_v3_0.switch_6.Z 2.49453f
C3255 CDAC_v3_0.switch_3.Z CDAC_v3_0.switch_7.Z 0.89198f
C3256 CDAC_v3_0.switch_8.Z CDAC_v3_0.OUT 5.0664f
C3257 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C EN 0.07565f
C3258 D_FlipFlop_6.nPRE D_FlipFlop_6.3-input-nand_2.Vout 0.76528f
C3259 Ring_Counter_0.D_FlipFlop_16.Q a_34285_60797# 0.01768f
C3260 D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.43587f
C3261 a_12901_55365# EN 0.04443f
C3262 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B VDD 1.71455f
C3263 a_37849_59439# VDD 0.01186f
C3264 a_49391_60797# Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout 0.05964f
C3265 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_13.Qbar 1.27148f
C3266 a_25616_51119# VDD 0.01186f
C3267 a_31571_55365# a_31571_54751# 0.05935f
C3268 CDAC_v3_0.switch_4.Z VDD 1.07378f
C3269 D_FlipFlop_0.Inverter_1.Vout a_54618_48405# 0.04995f
C3270 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.30156f
C3271 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout a_23593_58825# 0.05964f
C3272 a_27157_58825# VDD 0.02521f
C3273 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C CLK 0.26982f
C3274 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout VDD 2.72531f
C3275 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout a_52105_58825# 0.04444f
C3276 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD 1.89599f
C3277 a_2209_61411# VDD 0.08862f
C3278 a_17315_59439# VDD 0.05686f
C3279 D_FlipFlop_3.nPRE Q4 0.03683f
C3280 a_45856_51119# D_FlipFlop_1.Nand_Gate_0.Vout 0.05964f
C3281 And_Gate_0.A a_n7004_52049# 0.05964f
C3282 a_25616_48405# a_26230_48405# 0.05935f
C3283 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout VDD 2.07898f
C3284 a_6623_58825# VDD 0.02578f
C3285 Nand_Gate_5.A a_37849_56723# 0.05925f
C3286 a_9337_59439# EN 0.045f
C3287 a_9337_55365# EN 0.04443f
C3288 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout 0.01202f
C3289 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.01202f
C3290 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout VDD 2.8343f
C3291 D_FlipFlop_1.Qbar D_FlipFlop_1.Nand_Gate_1.Vout 0.11654f
C3292 D_FlipFlop_3.CLK D_FlipFlop_3.Inverter_1.Vout 0.20785f
C3293 Nand_Gate_0.A Ring_Counter_0.D_FlipFlop_14.Qbar 0.1225f
C3294 Ring_Counter_0.D_FlipFlop_6.Qbar a_30721_54751# 0.04443f
C3295 D_FlipFlop_0.Nand_Gate_1.Vout EN 0.61318f
C3296 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.Nand_Gate_0.Vout 0.16429f
C3297 a_4018_48405# Q1 0.05747f
C3298 And_Gate_0.A And_Gate_0.Nand_Gate_0.Vout 0.34057f
C3299 a_33020_51119# D_FlipFlop_2.3-input-nand_0.Vout 0.05964f
C3300 Ring_Counter_0.D_FlipFlop_16.Q a_n4919_55365# 0.01335f
C3301 Nand_Gate_1.A a_n4919_58825# 0.05925f
C3302 CDAC_v3_0.switch_4.Z Q4 0.17526f
C3303 a_45827_54751# Ring_Counter_0.D_FlipFlop_1.Qbar 0.06113f
C3304 a_17315_61411# Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.01335f
C3305 a_n4919_55365# a_n4919_54751# 0.05935f
C3306 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout 0.26069f
C3307 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_20879_55365# 0.04995f
C3308 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout VDD 2.72531f
C3309 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_45827_54751# 0.04444f
C3310 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_20029_55365# 0.04995f
C3311 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD 1.89599f
C3312 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_44977_54751# 0.04444f
C3313 D_FlipFlop_4.CLK a_6734_51119# 0.04443f
C3314 a_27157_61411# VDD 0.08862f
C3315 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout 0.3011f
C3316 a_10187_58825# Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.05964f
C3317 a_n4069_59439# CLK 0.03166f
C3318 a_45827_56723# Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.05964f
C3319 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B a_n7633_60797# 0.04443f
C3320 a_5773_55365# EN 0.04443f
C3321 D_FlipFlop_6.nPRE Q0 0.01264f
C3322 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.01194f
C3323 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C VDD 3.42554f
C3324 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C 0.01194f
C3325 a_28007_55365# a_28007_54751# 0.05935f
C3326 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C a_49391_56723# 0.04443f
C3327 Q0 Q1 2.27848f
C3328 a_20029_59439# a_20029_58825# 0.05935f
C3329 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.48403f
C3330 a_34378_48405# VDD 0.01186f
C3331 And_Gate_2.Nand_Gate_0.Vout a_5767_52049# 0.05964f
C3332 D_FlipFlop_7.CLK CLK 0.07954f
C3333 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.0646f
C3334 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.06462f
C3335 D_FlipFlop_6.Nand_Gate_0.Vout a_3404_51119# 0.04543f
C3336 Ring_Counter_0.D_FlipFlop_16.Q a_n4919_61411# 0.01252f
C3337 EN Q7 0.06332f
C3338 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.15413f
C3339 Nand_Gate_2.A Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.16911f
C3340 D_FlipFlop_1.3-input-nand_1.Vout a_43140_48405# 0.04543f
C3341 Nand_Gate_6.A a_16465_61411# 0.04995f
C3342 a_8092_48405# a_8706_48405# 0.05935f
C3343 D_FlipFlop_5.nPRE Nand_Gate_3.A 0.04143f
C3344 a_2209_55365# EN 0.04443f
C3345 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout a_35135_59439# 0.04543f
C3346 D_FlipFlop_5.nPRE D_FlipFlop_5.3-input-nand_0.Vout 0.94459f
C3347 a_52105_61411# VDD 0.09807f
C3348 D_FlipFlop_7.nPRE Q0 0.03683f
C3349 D_FlipFlop_1.nPRE Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B 0.02535f
C3350 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout a_5773_59439# 0.01335f
C3351 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout VDD 2.29925f
C3352 D_FlipFlop_2.nPRE a_38452_51119# 0.04443f
C3353 Ring_Counter_0.D_FlipFlop_7.Qbar a_27157_54751# 0.04443f
C3354 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.Qbar 1.27567f
C3355 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C 0.08674f
C3356 D_FlipFlop_7.3-input-nand_2.C a_n8818_48405# 0.05964f
C3357 a_n505_59439# a_n505_58825# 0.05935f
C3358 D_FlipFlop_7.3-input-nand_0.Vout a_n9432_51119# 0.04543f
C3359 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B 0.29684f
C3360 a_42263_54751# Ring_Counter_0.D_FlipFlop_2.Qbar 0.06113f
C3361 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout EN 0.08727f
C3362 D_FlipFlop_2.Qbar a_38452_48405# 0.01335f
C3363 a_n4744_51119# VDD 0.02521f
C3364 Nand_Gate_3.A Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B 0.02535f
C3365 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.16431f
C3366 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.0646f
C3367 D_FlipFlop_4.Qbar D_FlipFlop_4.Nand_Gate_1.Vout 0.11654f
C3368 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.06462f
C3369 a_48541_56723# VDD 0.02521f
C3370 a_n1355_55365# EN 0.04443f
C3371 Ring_Counter_0.D_FlipFlop_16.Q a_20029_61411# 0.01252f
C3372 D_FlipFlop_5.CLK D_FlipFlop_5.3-input-nand_1.Vout 0.67419f
C3373 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B VDD 1.71455f
C3374 D_FlipFlop_5.nPRE a_23593_55365# 0.01335f
C3375 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.08462f
C3376 a_24443_55365# a_24443_54751# 0.05935f
C3377 a_42263_61411# Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.01335f
C3378 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.Qbar 0.14288f
C3379 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout a_9337_59439# 0.04995f
C3380 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C a_n1355_58825# 0.04443f
C3381 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout EN 0.08727f
C3382 D_FlipFlop_1.Nand_Gate_0.Vout a_47214_51119# 0.04543f
C3383 a_n7633_60797# VDD 0.03137f
C3384 a_n4919_61411# a_n4919_60797# 0.05935f
C3385 a_n670_48405# VDD 0.01186f
C3386 a_n7633_59439# Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C 0.01335f
C3387 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.01262f
C3388 D_FlipFlop_4.3-input-nand_1.B a_6734_48405# 0.04443f
C3389 Nand_Gate_1.A Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.29165f
C3390 D_FlipFlop_0.3-input-nand_1.Vout EN 0.95784f
C3391 D_FlipFlop_2.3-input-nand_0.Vout a_34378_51119# 0.04543f
C3392 a_n4919_55365# EN 0.04443f
C3393 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_13.Qbar 0.07122f
C3394 D_FlipFlop_5.nPRE a_20029_55365# 0.05925f
C3395 a_n9432_48405# a_n8818_48405# 0.05935f
C3396 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B VDD 1.71455f
C3397 Ring_Counter_0.D_FlipFlop_8.Qbar a_23593_54751# 0.04443f
C3398 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout 0.06685f
C3399 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout a_52105_55365# 0.04995f
C3400 Ring_Counter_0.D_FlipFlop_16.Q Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.06658f
C3401 CDAC_v3_0.switch_5.Z m3_3428_33935# 1.89962f
C3402 D_FlipFlop_6.3-input-nand_1.Vout a_n2028_48405# 0.05964f
C3403 Ring_Counter_0.D_FlipFlop_16.Q a_44977_61411# 0.01252f
C3404 a_41168_51119# VDD 0.01186f
C3405 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.30156f
C3406 a_38699_54751# Ring_Counter_0.D_FlipFlop_3.Qbar 0.06113f
C3407 D_FlipFlop_4.nPRE Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.17364f
C3408 Nand_Gate_4.A a_31571_54751# 0.05987f
C3409 a_11766_45397# CDAC_v3_0.switch_2.Z 0.01245f
C3410 CDAC_v3_0.switch_0.Z a_15710_45397# 0.02206f
C3411 a_10187_61411# a_10187_60797# 0.05935f
C3412 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.06935f
C3413 D_FlipFlop_2.nPRE Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.20928f
C3414 a_17315_60797# VDD 0.02865f
C3415 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout a_9337_60797# 0.05964f
C3416 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout a_17315_58825# 0.04444f
C3417 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.01202f
C3418 a_52516_48405# VDD 0.02521f
C3419 Nand_Gate_4.A Ring_Counter_0.D_FlipFlop_16.Q 0.19783f
C3420 a_20879_55365# a_20879_54751# 0.05935f
C3421 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout 0.01202f
C3422 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B a_24443_61411# 0.04995f
C3423 a_24443_56723# VDD 0.02578f
C3424 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B VDD 1.71455f
C3425 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout EN 0.09223f
C3426 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout EN 0.96763f
C3427 And_Gate_3.Nand_Gate_0.Vout D_FlipFlop_5.CLK 0.25559f
C3428 a_n4919_61411# EN 0.02636f
C3429 a_3404_51119# a_4018_51119# 0.05935f
C3430 Vin GND 0.55041f
C3431 Q7 GND 7.80174f
C3432 Q6 GND 4.72225f
C3433 Q5 GND 6.21717f
C3434 Q4 GND 6.62305f
C3435 Q3 GND 5.64729f
C3436 Q2 GND 6.13248f
C3437 Q1 GND 6.43323f
C3438 Q0 GND 7.96605f
C3439 CLK GND 9.42962f
C3440 EN GND -34.32108f
C3441 Vbias GND 29.5259f
C3442 VDD GND 2.05091p
C3443 m3_3428_4751# GND 5.74304f $ **FLOATING
C3444 m3_3428_9615# GND 5.74304f $ **FLOATING
C3445 m3_3428_33935# GND 5.74323f $ **FLOATING
C3446 m3_3428_38799# GND 5.74323f $ **FLOATING
C3447 CDAC_v3_0.OUT GND 0.29318p
C3448 CDAC_v3_0.switch_6.Z GND 0.24278p
C3449 a_35430_45397# GND 2.17508f
C3450 CDAC_v3_0.switch_7.Z GND 0.17577p
C3451 a_31486_45397# GND 2.17477f
C3452 CDAC_v3_0.switch_5.Z GND 77.37109f
C3453 a_27542_45397# GND 2.17494f
C3454 CDAC_v3_0.switch_4.Z GND 52.97243f
C3455 a_23598_45397# GND 2.17493f
C3456 CDAC_v3_0.switch_3.Z GND 29.2262f
C3457 a_19654_45397# GND 2.17406f
C3458 CDAC_v3_0.switch_2.Z GND 17.21227f
C3459 a_15710_45397# GND 2.18883f
C3460 CDAC_v3_0.switch_0.Z GND 23.77117f
C3461 a_11766_45397# GND 2.17383f
C3462 CDAC_v3_0.switch_8.Z GND 10.86813f
C3463 a_7822_45397# GND 2.17355f
C3464 a_56590_48405# GND 0.25913f
C3465 a_55976_48405# GND 0.3185f
C3466 a_54618_48405# GND 0.3185f
C3467 a_52516_48405# GND 0.25914f
C3468 a_51902_48405# GND 0.3185f
C3469 a_50544_48405# GND 0.25914f
C3470 a_49930_48405# GND 0.3185f
C3471 a_47828_48405# GND 0.25913f
C3472 a_47214_48405# GND 0.3185f
C3473 a_45856_48405# GND 0.3185f
C3474 a_43754_48405# GND 0.25914f
C3475 a_43140_48405# GND 0.3185f
C3476 a_41782_48405# GND 0.25914f
C3477 a_41168_48405# GND 0.3198f
C3478 a_39066_48405# GND 0.25913f
C3479 a_38452_48405# GND 0.3185f
C3480 a_37094_48405# GND 0.3185f
C3481 a_34992_48405# GND 0.25914f
C3482 a_34378_48405# GND 0.3185f
C3483 a_33020_48405# GND 0.25914f
C3484 a_32406_48405# GND 0.3198f
C3485 a_30304_48405# GND 0.25913f
C3486 a_29690_48405# GND 0.3185f
C3487 a_28332_48405# GND 0.3185f
C3488 a_26230_48405# GND 0.25914f
C3489 a_25616_48405# GND 0.3185f
C3490 a_24258_48405# GND 0.25914f
C3491 a_23644_48405# GND 0.3198f
C3492 a_21542_48405# GND 0.25913f
C3493 a_20928_48405# GND 0.3185f
C3494 a_19570_48405# GND 0.3185f
C3495 a_17468_48405# GND 0.25914f
C3496 a_16854_48405# GND 0.3185f
C3497 a_15496_48405# GND 0.25914f
C3498 a_14882_48405# GND 0.3198f
C3499 a_12780_48405# GND 0.25913f
C3500 a_12166_48405# GND 0.3185f
C3501 a_10808_48405# GND 0.3185f
C3502 a_8706_48405# GND 0.25914f
C3503 a_8092_48405# GND 0.3185f
C3504 a_6734_48405# GND 0.25914f
C3505 a_6120_48405# GND 0.3198f
C3506 a_4018_48405# GND 0.25913f
C3507 a_3404_48405# GND 0.3185f
C3508 a_2046_48405# GND 0.3185f
C3509 a_n56_48405# GND 0.25914f
C3510 a_n670_48405# GND 0.3185f
C3511 a_n2028_48405# GND 0.25914f
C3512 a_n2642_48405# GND 0.3198f
C3513 a_n4744_48405# GND 0.25913f
C3514 a_n5358_48405# GND 0.3185f
C3515 a_n6716_48405# GND 0.3185f
C3516 a_n8818_48405# GND 0.25914f
C3517 a_n9432_48405# GND 0.3185f
C3518 a_n10790_48405# GND 0.25914f
C3519 a_n11404_48405# GND 0.3198f
C3520 D_FlipFlop_0.Nand_Gate_1.Vout GND 1.60762f
C3521 D_FlipFlop_0.3-input-nand_1.Vout GND 1.49358f
C3522 D_FlipFlop_1.Nand_Gate_1.Vout GND 1.5862f
C3523 D_FlipFlop_1.3-input-nand_1.Vout GND 1.49358f
C3524 D_FlipFlop_2.Nand_Gate_1.Vout GND 1.5862f
C3525 D_FlipFlop_2.3-input-nand_1.Vout GND 1.49358f
C3526 D_FlipFlop_3.Nand_Gate_1.Vout GND 1.5862f
C3527 D_FlipFlop_3.3-input-nand_1.Vout GND 1.49358f
C3528 D_FlipFlop_5.Nand_Gate_1.Vout GND 1.58593f
C3529 D_FlipFlop_5.3-input-nand_1.Vout GND 1.49307f
C3530 D_FlipFlop_4.Nand_Gate_1.Vout GND 1.58458f
C3531 D_FlipFlop_4.3-input-nand_1.Vout GND 1.49155f
C3532 D_FlipFlop_6.Nand_Gate_1.Vout GND 1.5862f
C3533 D_FlipFlop_6.3-input-nand_1.Vout GND 1.49358f
C3534 D_FlipFlop_7.Nand_Gate_1.Vout GND 1.5862f
C3535 D_FlipFlop_7.3-input-nand_1.Vout GND 1.49359f
C3536 a_56590_51119# GND 0.26272f
C3537 a_55976_51119# GND 0.31973f
C3538 D_FlipFlop_0.Qbar GND 1.76012f
C3539 D_FlipFlop_0.Nand_Gate_0.Vout GND 1.63403f
C3540 a_54618_51119# GND 0.3185f
C3541 D_FlipFlop_0.Inverter_1.Vout GND 2.74535f
C3542 D_FlipFlop_0.3-input-nand_2.Vout GND 2.1715f
C3543 a_52516_51119# GND 0.25913f
C3544 a_51902_51119# GND 0.3185f
C3545 D_FlipFlop_0.3-input-nand_2.C GND 2.16692f
C3546 D_FlipFlop_0.3-input-nand_0.Vout GND 1.63339f
C3547 a_50544_51119# GND 0.25914f
C3548 a_49930_51119# GND 0.3185f
C3549 D_FlipFlop_0.3-input-nand_1.B GND 1.68849f
C3550 a_47828_51119# GND 0.26317f
C3551 a_47214_51119# GND 0.31983f
C3552 D_FlipFlop_1.Qbar GND 1.62513f
C3553 D_FlipFlop_1.Nand_Gate_0.Vout GND 1.43997f
C3554 a_45856_51119# GND 0.3185f
C3555 D_FlipFlop_1.Inverter_1.Vout GND 2.74508f
C3556 D_FlipFlop_1.3-input-nand_2.Vout GND 2.19529f
C3557 a_43754_51119# GND 0.25913f
C3558 a_43140_51119# GND 0.3185f
C3559 D_FlipFlop_1.3-input-nand_2.C GND 2.20192f
C3560 D_FlipFlop_1.3-input-nand_0.Vout GND 1.45964f
C3561 a_41782_51119# GND 0.25914f
C3562 a_41168_51119# GND 0.3185f
C3563 D_FlipFlop_1.3-input-nand_1.B GND 1.85749f
C3564 a_39066_51119# GND 0.26317f
C3565 a_38452_51119# GND 0.31983f
C3566 D_FlipFlop_2.Qbar GND 1.62554f
C3567 D_FlipFlop_2.Nand_Gate_0.Vout GND 1.43997f
C3568 a_37094_51119# GND 0.3185f
C3569 D_FlipFlop_2.Inverter_1.Vout GND 2.74508f
C3570 D_FlipFlop_2.3-input-nand_2.Vout GND 2.19475f
C3571 a_34992_51119# GND 0.25913f
C3572 a_34378_51119# GND 0.3185f
C3573 D_FlipFlop_2.3-input-nand_2.C GND 2.20068f
C3574 D_FlipFlop_2.3-input-nand_0.Vout GND 1.45964f
C3575 a_33020_51119# GND 0.25914f
C3576 a_32406_51119# GND 0.3185f
C3577 D_FlipFlop_2.3-input-nand_1.B GND 1.85546f
C3578 a_30304_51119# GND 0.26317f
C3579 a_29690_51119# GND 0.31983f
C3580 D_FlipFlop_3.Qbar GND 1.62554f
C3581 D_FlipFlop_3.Nand_Gate_0.Vout GND 1.43997f
C3582 a_28332_51119# GND 0.3185f
C3583 D_FlipFlop_3.Inverter_1.Vout GND 2.74454f
C3584 D_FlipFlop_3.3-input-nand_2.Vout GND 2.19529f
C3585 a_26230_51119# GND 0.25913f
C3586 a_25616_51119# GND 0.3185f
C3587 D_FlipFlop_3.3-input-nand_2.C GND 2.20138f
C3588 D_FlipFlop_3.3-input-nand_0.Vout GND 1.45964f
C3589 a_24258_51119# GND 0.25914f
C3590 a_23644_51119# GND 0.3185f
C3591 D_FlipFlop_3.3-input-nand_1.B GND 1.85695f
C3592 a_21542_51119# GND 0.26317f
C3593 a_20928_51119# GND 0.31983f
C3594 D_FlipFlop_5.Qbar GND 1.62554f
C3595 D_FlipFlop_5.Nand_Gate_0.Vout GND 1.43997f
C3596 a_19570_51119# GND 0.3185f
C3597 D_FlipFlop_5.Inverter_1.Vout GND 2.74454f
C3598 D_FlipFlop_5.3-input-nand_2.Vout GND 2.19529f
C3599 a_17468_51119# GND 0.25913f
C3600 a_16854_51119# GND 0.3185f
C3601 D_FlipFlop_5.3-input-nand_2.C GND 2.20165f
C3602 D_FlipFlop_5.3-input-nand_0.Vout GND 1.45964f
C3603 a_15496_51119# GND 0.25914f
C3604 a_14882_51119# GND 0.3185f
C3605 D_FlipFlop_5.3-input-nand_1.B GND 1.85746f
C3606 a_12780_51119# GND 0.26317f
C3607 a_12166_51119# GND 0.31983f
C3608 D_FlipFlop_4.Qbar GND 1.62554f
C3609 D_FlipFlop_4.Nand_Gate_0.Vout GND 1.43997f
C3610 a_10808_51119# GND 0.3185f
C3611 D_FlipFlop_4.Inverter_1.Vout GND 2.74508f
C3612 D_FlipFlop_4.3-input-nand_2.Vout GND 2.19326f
C3613 a_8706_51119# GND 0.25913f
C3614 a_8092_51119# GND 0.3185f
C3615 D_FlipFlop_4.3-input-nand_2.C GND 2.20192f
C3616 D_FlipFlop_4.3-input-nand_0.Vout GND 1.45964f
C3617 a_6734_51119# GND 0.25914f
C3618 a_6120_51119# GND 0.3185f
C3619 D_FlipFlop_4.3-input-nand_1.B GND 1.85749f
C3620 a_4018_51119# GND 0.26317f
C3621 a_3404_51119# GND 0.31983f
C3622 D_FlipFlop_6.Qbar GND 1.62554f
C3623 D_FlipFlop_6.Nand_Gate_0.Vout GND 1.43997f
C3624 a_2046_51119# GND 0.3185f
C3625 D_FlipFlop_6.Inverter_1.Vout GND 2.74508f
C3626 D_FlipFlop_6.3-input-nand_2.Vout GND 2.19529f
C3627 a_n56_51119# GND 0.25913f
C3628 a_n670_51119# GND 0.3185f
C3629 D_FlipFlop_6.3-input-nand_2.C GND 2.20192f
C3630 D_FlipFlop_6.3-input-nand_0.Vout GND 1.45964f
C3631 a_n2028_51119# GND 0.25914f
C3632 a_n2642_51119# GND 0.3185f
C3633 D_FlipFlop_6.3-input-nand_1.B GND 1.85749f
C3634 a_n4744_51119# GND 0.26317f
C3635 a_n5358_51119# GND 0.31983f
C3636 D_FlipFlop_7.Qbar GND 1.62554f
C3637 D_FlipFlop_7.Nand_Gate_0.Vout GND 1.43997f
C3638 a_n6716_51119# GND 0.3185f
C3639 D_FlipFlop_7.Inverter_1.Vout GND 2.74508f
C3640 D_FlipFlop_7.3-input-nand_2.Vout GND 2.19529f
C3641 a_n8818_51119# GND 0.25913f
C3642 a_n9432_51119# GND 0.3185f
C3643 D_FlipFlop_7.3-input-nand_2.C GND 2.20192f
C3644 D_FlipFlop_7.3-input-nand_0.Vout GND 1.45965f
C3645 a_n10790_51119# GND 0.25914f
C3646 a_n11404_51119# GND 0.3185f
C3647 D_FlipFlop_7.3-input-nand_1.B GND 1.90098f
C3648 a_54330_52049# GND 0.3185f
C3649 a_49577_52049# GND 0.3185f
C3650 a_45568_52049# GND 0.3185f
C3651 a_40815_52049# GND 0.3185f
C3652 a_36806_52049# GND 0.3185f
C3653 a_32053_52049# GND 0.3185f
C3654 a_28044_52049# GND 0.3185f
C3655 a_23291_52049# GND 0.3185f
C3656 a_19282_52049# GND 0.3185f
C3657 a_14529_52049# GND 0.3185f
C3658 a_10520_52049# GND 0.3185f
C3659 a_5767_52049# GND 0.3185f
C3660 a_1758_52049# GND 0.3185f
C3661 a_n2995_52049# GND 0.3185f
C3662 a_n7004_52049# GND 0.3185f
C3663 a_n11757_52049# GND 0.3185f
C3664 D_FlipFlop_0.CLK GND 4.2308f
C3665 And_Gate_7.Nand_Gate_0.Vout GND 1.68958f
C3666 And_Gate_7.A GND 3.26532f
C3667 D_FlipFlop_1.CLK GND 4.36804f
C3668 And_Gate_6.Nand_Gate_0.Vout GND 1.68434f
C3669 And_Gate_6.A GND 2.71982f
C3670 D_FlipFlop_2.CLK GND 4.366f
C3671 And_Gate_5.Nand_Gate_0.Vout GND 1.68476f
C3672 And_Gate_5.A GND 2.71197f
C3673 D_FlipFlop_3.CLK GND 4.36698f
C3674 And_Gate_4.Nand_Gate_0.Vout GND 1.69006f
C3675 And_Gate_4.A GND 2.7221f
C3676 D_FlipFlop_5.CLK GND 4.36642f
C3677 And_Gate_3.Nand_Gate_0.Vout GND 1.67767f
C3678 And_Gate_3.A GND 2.71472f
C3679 D_FlipFlop_4.CLK GND 4.36804f
C3680 And_Gate_2.Nand_Gate_0.Vout GND 1.6879f
C3681 And_Gate_2.A GND 2.72006f
C3682 D_FlipFlop_6.CLK GND 4.36804f
C3683 And_Gate_1.Nand_Gate_0.Vout GND 1.6768f
C3684 And_Gate_1.A GND 2.71843f
C3685 D_FlipFlop_7.CLK GND 4.36804f
C3686 And_Gate_0.Nand_Gate_0.Vout GND 1.70549f
C3687 And_Gate_0.A GND 2.71443f
C3688 a_52105_54751# GND 0.25913f
C3689 a_52105_55365# GND 0.3185f
C3690 Ring_Counter_0.D_FlipFlop_0.Qbar GND 1.52381f
C3691 a_49391_54751# GND 0.25913f
C3692 a_49391_55365# GND 0.3185f
C3693 a_48541_54751# GND 0.25913f
C3694 a_48541_55365# GND 0.3185f
C3695 Ring_Counter_0.D_FlipFlop_1.Qbar GND 1.55944f
C3696 a_45827_54751# GND 0.25913f
C3697 a_45827_55365# GND 0.3185f
C3698 a_44977_54751# GND 0.25913f
C3699 a_44977_55365# GND 0.3185f
C3700 Ring_Counter_0.D_FlipFlop_2.Qbar GND 1.55879f
C3701 a_42263_54751# GND 0.25913f
C3702 a_42263_55365# GND 0.3185f
C3703 a_41413_54751# GND 0.25913f
C3704 a_41413_55365# GND 0.3185f
C3705 Ring_Counter_0.D_FlipFlop_3.Qbar GND 1.53573f
C3706 a_38699_54751# GND 0.25913f
C3707 a_38699_55365# GND 0.3185f
C3708 a_37849_54751# GND 0.25913f
C3709 a_37849_55365# GND 0.3185f
C3710 Ring_Counter_0.D_FlipFlop_4.Qbar GND 1.53567f
C3711 a_35135_54751# GND 0.25913f
C3712 a_35135_55365# GND 0.3185f
C3713 a_34285_54751# GND 0.25913f
C3714 a_34285_55365# GND 0.3185f
C3715 Ring_Counter_0.D_FlipFlop_5.Qbar GND 1.53431f
C3716 a_31571_54751# GND 0.25913f
C3717 a_31571_55365# GND 0.3185f
C3718 a_30721_54751# GND 0.25913f
C3719 a_30721_55365# GND 0.3185f
C3720 Ring_Counter_0.D_FlipFlop_6.Qbar GND 1.55551f
C3721 a_28007_54751# GND 0.25913f
C3722 a_28007_55365# GND 0.3185f
C3723 a_27157_54751# GND 0.25913f
C3724 a_27157_55365# GND 0.3185f
C3725 Ring_Counter_0.D_FlipFlop_7.Qbar GND 1.5594f
C3726 a_24443_54751# GND 0.25913f
C3727 a_24443_55365# GND 0.3185f
C3728 a_23593_54751# GND 0.25913f
C3729 a_23593_55365# GND 0.3185f
C3730 Ring_Counter_0.D_FlipFlop_8.Qbar GND 1.53783f
C3731 a_20879_54751# GND 0.25913f
C3732 a_20879_55365# GND 0.3185f
C3733 a_20029_54751# GND 0.25913f
C3734 a_20029_55365# GND 0.3185f
C3735 Ring_Counter_0.D_FlipFlop_9.Qbar GND 1.55166f
C3736 a_17315_54751# GND 0.25913f
C3737 a_17315_55365# GND 0.3185f
C3738 a_16465_54751# GND 0.25913f
C3739 a_16465_55365# GND 0.3185f
C3740 Ring_Counter_0.D_FlipFlop_10.Qbar GND 1.53418f
C3741 a_13751_54751# GND 0.25913f
C3742 a_13751_55365# GND 0.3185f
C3743 a_12901_54751# GND 0.25913f
C3744 a_12901_55365# GND 0.3185f
C3745 Ring_Counter_0.D_FlipFlop_11.Qbar GND 1.53684f
C3746 a_10187_54751# GND 0.25913f
C3747 a_10187_55365# GND 0.3185f
C3748 a_9337_54751# GND 0.25913f
C3749 a_9337_55365# GND 0.3185f
C3750 Ring_Counter_0.D_FlipFlop_12.Qbar GND 1.55944f
C3751 a_6623_54751# GND 0.25913f
C3752 a_6623_55365# GND 0.3185f
C3753 a_5773_54751# GND 0.25913f
C3754 a_5773_55365# GND 0.3185f
C3755 Ring_Counter_0.D_FlipFlop_13.Qbar GND 1.55797f
C3756 a_3059_54751# GND 0.25913f
C3757 a_3059_55365# GND 0.3185f
C3758 a_2209_54751# GND 0.25913f
C3759 a_2209_55365# GND 0.3185f
C3760 Ring_Counter_0.D_FlipFlop_14.Qbar GND 1.53527f
C3761 a_n505_54751# GND 0.25913f
C3762 a_n505_55365# GND 0.3185f
C3763 a_n1355_54751# GND 0.25913f
C3764 a_n1355_55365# GND 0.3185f
C3765 Ring_Counter_0.D_FlipFlop_15.Qbar GND 1.53393f
C3766 a_n4069_54751# GND 0.25913f
C3767 a_n4069_55365# GND 0.3185f
C3768 a_n4919_54751# GND 0.25913f
C3769 a_n4919_55365# GND 0.3185f
C3770 Ring_Counter_0.D_FlipFlop_16.Qbar GND 1.5991f
C3771 a_n7633_54751# GND 0.25913f
C3772 a_n7633_55365# GND 0.3185f
C3773 a_52105_56723# GND 0.3185f
C3774 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout GND 1.47014f
C3775 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_1.Vout GND 1.52315f
C3776 a_49391_56723# GND 0.3185f
C3777 a_48541_56723# GND 0.3185f
C3778 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_0.Vout GND 1.50487f
C3779 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout GND 1.39179f
C3780 a_45827_56723# GND 0.3185f
C3781 a_44977_56723# GND 0.3185f
C3782 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_0.Vout GND 1.50487f
C3783 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout GND 1.39179f
C3784 a_42263_56723# GND 0.3185f
C3785 a_41413_56723# GND 0.3185f
C3786 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_0.Vout GND 1.50487f
C3787 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout GND 1.39179f
C3788 a_38699_56723# GND 0.3185f
C3789 a_37849_56723# GND 0.3185f
C3790 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_0.Vout GND 1.50487f
C3791 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout GND 1.39179f
C3792 a_35135_56723# GND 0.3185f
C3793 a_34285_56723# GND 0.3185f
C3794 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_0.Vout GND 1.50487f
C3795 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout GND 1.39179f
C3796 a_31571_56723# GND 0.3185f
C3797 a_30721_56723# GND 0.3185f
C3798 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_0.Vout GND 1.50487f
C3799 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout GND 1.39179f
C3800 a_28007_56723# GND 0.3185f
C3801 a_27157_56723# GND 0.3185f
C3802 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_0.Vout GND 1.50487f
C3803 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout GND 1.39179f
C3804 a_24443_56723# GND 0.3185f
C3805 a_23593_56723# GND 0.3185f
C3806 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_0.Vout GND 1.50487f
C3807 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout GND 1.39179f
C3808 a_20879_56723# GND 0.3185f
C3809 a_20029_56723# GND 0.3185f
C3810 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_0.Vout GND 1.50487f
C3811 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout GND 1.39179f
C3812 a_17315_56723# GND 0.3185f
C3813 a_16465_56723# GND 0.3185f
C3814 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_0.Vout GND 1.50487f
C3815 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout GND 1.39179f
C3816 a_13751_56723# GND 0.3185f
C3817 a_12901_56723# GND 0.3185f
C3818 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_0.Vout GND 1.50487f
C3819 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout GND 1.39179f
C3820 a_10187_56723# GND 0.3185f
C3821 a_9337_56723# GND 0.3185f
C3822 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_0.Vout GND 1.50487f
C3823 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout GND 1.39179f
C3824 a_6623_56723# GND 0.3185f
C3825 a_5773_56723# GND 0.3185f
C3826 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_0.Vout GND 1.50487f
C3827 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout GND 1.39179f
C3828 a_3059_56723# GND 0.3185f
C3829 a_2209_56723# GND 0.3185f
C3830 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_0.Vout GND 1.50487f
C3831 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout GND 1.39179f
C3832 a_n505_56723# GND 0.3185f
C3833 a_n1355_56723# GND 0.3185f
C3834 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_0.Vout GND 1.50487f
C3835 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout GND 1.39179f
C3836 a_n4069_56723# GND 0.3185f
C3837 a_n4919_56723# GND 0.3185f
C3838 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_0.Vout GND 1.48635f
C3839 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout GND 1.46375f
C3840 a_n7633_56723# GND 0.3185f
C3841 Ring_Counter_0.D_FlipFlop_0.Inverter_1.Vout GND 2.61957f
C3842 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout GND 2.54791f
C3843 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout GND 2.54791f
C3844 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout GND 2.54791f
C3845 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout GND 2.54791f
C3846 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout GND 2.54791f
C3847 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout GND 2.54791f
C3848 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout GND 2.54791f
C3849 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout GND 2.54791f
C3850 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout GND 2.54509f
C3851 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout GND 2.54791f
C3852 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout GND 2.54791f
C3853 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout GND 2.54791f
C3854 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout GND 2.54791f
C3855 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout GND 2.54791f
C3856 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout GND 2.54791f
C3857 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout GND 2.632f
C3858 a_52105_58825# GND 0.25913f
C3859 a_52105_59439# GND 0.3185f
C3860 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C GND 2.41442f
C3861 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout GND 2.56749f
C3862 a_49391_58825# GND 0.25914f
C3863 a_49391_59439# GND 0.3185f
C3864 a_48541_58825# GND 0.25913f
C3865 a_48541_59439# GND 0.3185f
C3866 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C GND 2.36687f
C3867 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout GND 2.56429f
C3868 a_45827_58825# GND 0.25914f
C3869 a_45827_59439# GND 0.3185f
C3870 a_44977_58825# GND 0.25913f
C3871 a_44977_59439# GND 0.3185f
C3872 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C GND 2.36687f
C3873 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout GND 2.56429f
C3874 a_42263_58825# GND 0.25914f
C3875 a_42263_59439# GND 0.3185f
C3876 a_41413_58825# GND 0.25913f
C3877 a_41413_59439# GND 0.3185f
C3878 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C GND 2.36687f
C3879 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout GND 2.56429f
C3880 a_38699_58825# GND 0.25914f
C3881 a_38699_59439# GND 0.3185f
C3882 a_37849_58825# GND 0.25913f
C3883 a_37849_59439# GND 0.3185f
C3884 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C GND 2.36687f
C3885 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout GND 2.56429f
C3886 a_35135_58825# GND 0.25914f
C3887 a_35135_59439# GND 0.3185f
C3888 a_34285_58825# GND 0.25913f
C3889 a_34285_59439# GND 0.3185f
C3890 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C GND 2.36687f
C3891 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout GND 2.56429f
C3892 a_31571_58825# GND 0.25914f
C3893 a_31571_59439# GND 0.3185f
C3894 a_30721_58825# GND 0.25913f
C3895 a_30721_59439# GND 0.3185f
C3896 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C GND 2.36687f
C3897 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout GND 2.56429f
C3898 a_28007_58825# GND 0.25914f
C3899 a_28007_59439# GND 0.3185f
C3900 a_27157_58825# GND 0.25913f
C3901 a_27157_59439# GND 0.3185f
C3902 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C GND 2.36687f
C3903 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout GND 2.56429f
C3904 a_24443_58825# GND 0.25914f
C3905 a_24443_59439# GND 0.3185f
C3906 a_23593_58825# GND 0.25913f
C3907 a_23593_59439# GND 0.3185f
C3908 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C GND 2.36687f
C3909 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout GND 2.56429f
C3910 a_20879_58825# GND 0.25914f
C3911 a_20879_59439# GND 0.3185f
C3912 a_20029_58825# GND 0.25913f
C3913 a_20029_59439# GND 0.3185f
C3914 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C GND 2.36335f
C3915 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout GND 2.55948f
C3916 a_17315_58825# GND 0.25914f
C3917 a_17315_59439# GND 0.3185f
C3918 a_16465_58825# GND 0.25913f
C3919 a_16465_59439# GND 0.3185f
C3920 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C GND 2.36687f
C3921 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout GND 2.56429f
C3922 a_13751_58825# GND 0.25914f
C3923 a_13751_59439# GND 0.3185f
C3924 a_12901_58825# GND 0.25913f
C3925 a_12901_59439# GND 0.3185f
C3926 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C GND 2.36687f
C3927 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout GND 2.56429f
C3928 a_10187_58825# GND 0.25914f
C3929 a_10187_59439# GND 0.3185f
C3930 a_9337_58825# GND 0.25913f
C3931 a_9337_59439# GND 0.3185f
C3932 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C GND 2.36687f
C3933 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout GND 2.56429f
C3934 a_6623_58825# GND 0.25914f
C3935 a_6623_59439# GND 0.3185f
C3936 a_5773_58825# GND 0.25913f
C3937 a_5773_59439# GND 0.3185f
C3938 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C GND 2.36687f
C3939 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout GND 2.56429f
C3940 a_3059_58825# GND 0.25914f
C3941 a_3059_59439# GND 0.3185f
C3942 a_2209_58825# GND 0.25913f
C3943 a_2209_59439# GND 0.3185f
C3944 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C GND 2.36687f
C3945 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout GND 2.56429f
C3946 a_n505_58825# GND 0.25914f
C3947 a_n505_59439# GND 0.3185f
C3948 a_n1355_58825# GND 0.25913f
C3949 a_n1355_59439# GND 0.3185f
C3950 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C GND 2.36687f
C3951 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout GND 2.56429f
C3952 a_n4069_58825# GND 0.25914f
C3953 a_n4069_59439# GND 0.3185f
C3954 a_n4919_58825# GND 0.25913f
C3955 a_n4919_59439# GND 0.3185f
C3956 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C GND 2.38184f
C3957 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout GND 2.57457f
C3958 a_n7633_58825# GND 0.25914f
C3959 a_n7633_59439# GND 0.3185f
C3960 a_52105_60797# GND 0.25914f
C3961 a_52105_61411# GND 0.31934f
C3962 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout GND 1.45832f
C3963 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.Vout GND 1.4841f
C3964 a_49391_60797# GND 0.25914f
C3965 a_49391_61411# GND 0.3185f
C3966 a_48541_60797# GND 0.25914f
C3967 a_48541_61411# GND 0.3185f
C3968 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.Vout GND 1.52089f
C3969 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout GND 1.33275f
C3970 a_45827_60797# GND 0.25914f
C3971 a_45827_61411# GND 0.3185f
C3972 a_44977_60797# GND 0.25914f
C3973 a_44977_61411# GND 0.3185f
C3974 Ring_Counter_0.D_FlipFlop_2.3-input-nand_0.Vout GND 1.52144f
C3975 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout GND 1.33275f
C3976 a_42263_60797# GND 0.25914f
C3977 a_42263_61411# GND 0.3185f
C3978 a_41413_60797# GND 0.25914f
C3979 a_41413_61411# GND 0.3185f
C3980 Ring_Counter_0.D_FlipFlop_3.3-input-nand_0.Vout GND 1.52144f
C3981 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout GND 1.33275f
C3982 a_38699_60797# GND 0.25914f
C3983 a_38699_61411# GND 0.3185f
C3984 a_37849_60797# GND 0.25914f
C3985 a_37849_61411# GND 0.3185f
C3986 Ring_Counter_0.D_FlipFlop_4.3-input-nand_0.Vout GND 1.52144f
C3987 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout GND 1.33275f
C3988 a_35135_60797# GND 0.25914f
C3989 a_35135_61411# GND 0.3185f
C3990 a_34285_60797# GND 0.25914f
C3991 a_34285_61411# GND 0.3185f
C3992 Ring_Counter_0.D_FlipFlop_5.3-input-nand_0.Vout GND 1.52144f
C3993 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout GND 1.33275f
C3994 a_31571_60797# GND 0.25914f
C3995 a_31571_61411# GND 0.3185f
C3996 a_30721_60797# GND 0.25914f
C3997 a_30721_61411# GND 0.3185f
C3998 Ring_Counter_0.D_FlipFlop_6.3-input-nand_0.Vout GND 1.52144f
C3999 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout GND 1.33275f
C4000 a_28007_60797# GND 0.25914f
C4001 a_28007_61411# GND 0.3185f
C4002 a_27157_60797# GND 0.25914f
C4003 a_27157_61411# GND 0.3185f
C4004 Ring_Counter_0.D_FlipFlop_7.3-input-nand_0.Vout GND 1.52144f
C4005 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout GND 1.33275f
C4006 a_24443_60797# GND 0.25914f
C4007 a_24443_61411# GND 0.3185f
C4008 a_23593_60797# GND 0.25914f
C4009 a_23593_61411# GND 0.3185f
C4010 Ring_Counter_0.D_FlipFlop_8.3-input-nand_0.Vout GND 1.52144f
C4011 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout GND 1.33275f
C4012 a_20879_60797# GND 0.25914f
C4013 a_20879_61411# GND 0.3185f
C4014 a_20029_60797# GND 0.25914f
C4015 a_20029_61411# GND 0.3185f
C4016 Ring_Counter_0.D_FlipFlop_9.3-input-nand_0.Vout GND 1.52144f
C4017 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout GND 1.33275f
C4018 a_17315_60797# GND 0.25914f
C4019 a_17315_61411# GND 0.3185f
C4020 a_16465_60797# GND 0.25914f
C4021 a_16465_61411# GND 0.3185f
C4022 Ring_Counter_0.D_FlipFlop_10.3-input-nand_0.Vout GND 1.52144f
C4023 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout GND 1.33275f
C4024 a_13751_60797# GND 0.25914f
C4025 a_13751_61411# GND 0.3185f
C4026 a_12901_60797# GND 0.25914f
C4027 a_12901_61411# GND 0.3185f
C4028 Ring_Counter_0.D_FlipFlop_11.3-input-nand_0.Vout GND 1.52144f
C4029 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout GND 1.33275f
C4030 a_10187_60797# GND 0.25914f
C4031 a_10187_61411# GND 0.3185f
C4032 a_9337_60797# GND 0.25914f
C4033 a_9337_61411# GND 0.3185f
C4034 Ring_Counter_0.D_FlipFlop_12.3-input-nand_0.Vout GND 1.52144f
C4035 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout GND 1.33275f
C4036 a_6623_60797# GND 0.25914f
C4037 a_6623_61411# GND 0.3185f
C4038 a_5773_60797# GND 0.25914f
C4039 a_5773_61411# GND 0.3185f
C4040 Ring_Counter_0.D_FlipFlop_13.3-input-nand_0.Vout GND 1.52144f
C4041 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout GND 1.33275f
C4042 a_3059_60797# GND 0.25914f
C4043 a_3059_61411# GND 0.3185f
C4044 a_2209_60797# GND 0.25914f
C4045 a_2209_61411# GND 0.3185f
C4046 Ring_Counter_0.D_FlipFlop_14.3-input-nand_0.Vout GND 1.52144f
C4047 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout GND 1.33275f
C4048 a_n505_60797# GND 0.25914f
C4049 a_n505_61411# GND 0.3185f
C4050 a_n1355_60797# GND 0.25914f
C4051 a_n1355_61411# GND 0.3185f
C4052 Ring_Counter_0.D_FlipFlop_15.3-input-nand_0.Vout GND 1.52144f
C4053 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout GND 1.33275f
C4054 a_n4069_60797# GND 0.25914f
C4055 a_n4069_61411# GND 0.3185f
C4056 a_n4919_60797# GND 0.25914f
C4057 a_n4919_61411# GND 0.3185f
C4058 Ring_Counter_0.D_FlipFlop_16.3-input-nand_0.Vout GND 1.52144f
C4059 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout GND 1.34224f
C4060 a_n7633_60797# GND 0.25914f
C4061 a_n7633_61411# GND 0.31975f
C4062 Ring_Counter_0.D_FlipFlop_0.3-input-nand_1.B GND 1.86477f
C4063 Ring_Counter_0.D_FlipFlop_16.Q GND 6.94307f
C4064 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.B GND 1.86492f
C4065 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.B GND 1.86504f
C4066 Nand_Gate_7.A GND 10.32324f
C4067 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.B GND 1.86504f
C4068 D_FlipFlop_1.nPRE GND 12.79961f
C4069 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.B GND 1.86504f
C4070 Nand_Gate_5.A GND 9.78145f
C4071 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.B GND 1.86504f
C4072 D_FlipFlop_2.nPRE GND 12.71656f
C4073 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.B GND 1.86504f
C4074 Nand_Gate_4.A GND 9.20569f
C4075 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.B GND 1.86504f
C4076 D_FlipFlop_3.nPRE GND 13.04615f
C4077 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.B GND 1.86504f
C4078 Nand_Gate_3.A GND 8.91418f
C4079 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.B GND 1.86504f
C4080 D_FlipFlop_5.nPRE GND 13.8624f
C4081 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.B GND 1.86504f
C4082 Nand_Gate_6.A GND 8.44478f
C4083 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.B GND 1.86504f
C4084 D_FlipFlop_4.nPRE GND 14.35231f
C4085 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.B GND 1.86504f
C4086 Nand_Gate_2.A GND 8.19601f
C4087 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.B GND 1.86504f
C4088 D_FlipFlop_6.nPRE GND 14.21687f
C4089 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.B GND 1.86504f
C4090 Nand_Gate_0.A GND 8.57607f
C4091 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.B GND 1.86504f
C4092 D_FlipFlop_7.nPRE GND 14.7645f
C4093 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.B GND 1.88159f
C4094 Nand_Gate_1.A GND 8.72453f
C4095 a_50454_10637.t2 GND 0.70901f
C4096 a_50454_10637.t4 GND 0.66541f
C4097 a_50454_10637.t3 GND 1.2388f
C4098 a_50454_10637.n0 GND 0.6901f
C4099 a_50454_10637.t1 GND 1.2388f
C4100 a_50454_10637.n1 GND 0.3967f
C4101 a_50454_10637.n2 GND 0.44526f
C4102 a_50454_10637.t0 GND 2.81593f
C4103 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 GND 0.07411f
C4104 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 GND 0.16107f
C4105 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 GND 0.08416f
C4106 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 GND 0.29566f
C4107 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 GND 0.14335f
C4108 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 GND 0.56804f
C4109 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 GND 0.1051f
C4110 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 GND 0.06271f
C4111 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 GND 0.15391f
C4112 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 GND 0.15391f
C4113 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 GND 0.07722f
C4114 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 GND 0.07866f
C4115 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 GND 0.07705f
C4116 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 GND 0.43817f
C4117 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 GND 0.286f
C4118 Ring_Counter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 GND 0.09223f
C4119 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 GND 0.07411f
C4120 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 GND 0.16107f
C4121 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 GND 0.08416f
C4122 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 GND 0.29566f
C4123 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 GND 0.14335f
C4124 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 GND 0.56804f
C4125 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 GND 0.1051f
C4126 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 GND 0.06271f
C4127 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 GND 0.15391f
C4128 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 GND 0.15391f
C4129 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 GND 0.07722f
C4130 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 GND 0.07866f
C4131 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 GND 0.07705f
C4132 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 GND 0.43817f
C4133 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 GND 0.286f
C4134 Ring_Counter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 GND 0.09223f
C4135 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 GND 0.07411f
C4136 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 GND 0.16107f
C4137 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 GND 0.08416f
C4138 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 GND 0.29566f
C4139 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 GND 0.14335f
C4140 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 GND 0.56804f
C4141 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 GND 0.1051f
C4142 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 GND 0.06271f
C4143 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 GND 0.15391f
C4144 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 GND 0.15391f
C4145 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 GND 0.07722f
C4146 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 GND 0.07866f
C4147 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 GND 0.07705f
C4148 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 GND 0.43817f
C4149 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 GND 0.286f
C4150 Ring_Counter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 GND 0.09223f
C4151 D_FlipFlop_5.3-input-nand_2.C.t7 GND 0.3425f
C4152 D_FlipFlop_5.3-input-nand_2.C.n0 GND 0.3551f
C4153 D_FlipFlop_5.3-input-nand_2.C.n1 GND 0.03842f
C4154 D_FlipFlop_5.3-input-nand_2.C.t2 GND 0.04469f
C4155 D_FlipFlop_5.3-input-nand_2.C.n2 GND 0.04327f
C4156 D_FlipFlop_5.3-input-nand_2.C.n3 GND 0.09193f
C4157 D_FlipFlop_5.3-input-nand_2.C.t5 GND 0.17806f
C4158 D_FlipFlop_5.3-input-nand_2.C.t6 GND 0.34248f
C4159 D_FlipFlop_5.3-input-nand_2.C.n4 GND 0.10005f
C4160 D_FlipFlop_5.3-input-nand_2.C.n5 GND 0.04279f
C4161 D_FlipFlop_5.3-input-nand_2.C.n6 GND 0.079f
C4162 D_FlipFlop_5.3-input-nand_2.C.n7 GND 0.13677f
C4163 D_FlipFlop_5.3-input-nand_2.C.n8 GND 0.10181f
C4164 D_FlipFlop_5.3-input-nand_2.C.n9 GND 0.04823f
C4165 D_FlipFlop_5.3-input-nand_2.C.n10 GND 0.124f
C4166 D_FlipFlop_5.3-input-nand_2.C.t3 GND 0.04742f
C4167 D_FlipFlop_5.3-input-nand_2.C.t0 GND 0.04645f
C4168 D_FlipFlop_5.3-input-nand_2.C.n11 GND 0.26418f
C4169 D_FlipFlop_5.3-input-nand_2.C.n12 GND 0.08722f
C4170 D_FlipFlop_5.3-input-nand_2.C.t1 GND 0.04645f
C4171 D_FlipFlop_5.3-input-nand_2.C.n13 GND 0.293f
C4172 D_FlipFlop_5.3-input-nand_2.C.t4 GND 0.17045f
C4173 D_FlipFlop_5.3-input-nand_2.C.n14 GND 0.05129f
C4174 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t1 GND 0.05f
C4175 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n0 GND 0.10867f
C4176 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n1 GND 0.05678f
C4177 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t3 GND 0.38491f
C4178 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n2 GND 0.16589f
C4179 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t5 GND 0.30131f
C4180 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t2 GND 0.30153f
C4181 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n3 GND 0.09671f
C4182 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t4 GND 0.38323f
C4183 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n4 GND 0.0709f
C4184 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n5 GND 0.04231f
C4185 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n6 GND 0.10383f
C4186 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n7 GND 0.10383f
C4187 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.t0 GND 0.05284f
C4188 Ring_Counter_0.D_FlipFlop_11.Inverter_1.Vout.n8 GND 0.17757f
C4189 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 GND 0.07411f
C4190 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 GND 0.16107f
C4191 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 GND 0.08416f
C4192 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 GND 0.29566f
C4193 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 GND 0.14335f
C4194 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 GND 0.56804f
C4195 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 GND 0.1051f
C4196 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 GND 0.06271f
C4197 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 GND 0.15391f
C4198 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 GND 0.15391f
C4199 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 GND 0.07722f
C4200 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 GND 0.07866f
C4201 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 GND 0.07705f
C4202 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 GND 0.43817f
C4203 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 GND 0.286f
C4204 Ring_Counter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 GND 0.09223f
C4205 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 GND 0.07411f
C4206 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 GND 0.16107f
C4207 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 GND 0.08416f
C4208 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 GND 0.29566f
C4209 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 GND 0.14335f
C4210 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 GND 0.56804f
C4211 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 GND 0.1051f
C4212 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 GND 0.06271f
C4213 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 GND 0.15391f
C4214 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 GND 0.15391f
C4215 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 GND 0.07722f
C4216 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 GND 0.07866f
C4217 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 GND 0.07705f
C4218 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 GND 0.43817f
C4219 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 GND 0.286f
C4220 Ring_Counter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 GND 0.09223f
C4221 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 GND 0.07411f
C4222 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 GND 0.16107f
C4223 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 GND 0.08416f
C4224 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 GND 0.29566f
C4225 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 GND 0.14335f
C4226 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 GND 0.56804f
C4227 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 GND 0.1051f
C4228 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 GND 0.06271f
C4229 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 GND 0.15391f
C4230 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 GND 0.15391f
C4231 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 GND 0.07722f
C4232 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 GND 0.07866f
C4233 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 GND 0.07705f
C4234 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 GND 0.43817f
C4235 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 GND 0.286f
C4236 Ring_Counter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 GND 0.09223f
C4237 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 GND 0.07411f
C4238 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 GND 0.16107f
C4239 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 GND 0.08416f
C4240 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 GND 0.29566f
C4241 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 GND 0.14335f
C4242 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 GND 0.56804f
C4243 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 GND 0.1051f
C4244 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 GND 0.06271f
C4245 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 GND 0.15391f
C4246 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 GND 0.15391f
C4247 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 GND 0.07722f
C4248 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 GND 0.07866f
C4249 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 GND 0.07705f
C4250 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 GND 0.43817f
C4251 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 GND 0.286f
C4252 Ring_Counter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 GND 0.09223f
C4253 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 GND 0.07411f
C4254 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 GND 0.16107f
C4255 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 GND 0.08416f
C4256 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 GND 0.29566f
C4257 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 GND 0.14335f
C4258 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 GND 0.56804f
C4259 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 GND 0.1051f
C4260 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 GND 0.06271f
C4261 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 GND 0.15391f
C4262 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 GND 0.15391f
C4263 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 GND 0.07722f
C4264 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 GND 0.07866f
C4265 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 GND 0.07705f
C4266 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 GND 0.43817f
C4267 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 GND 0.286f
C4268 Ring_Counter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 GND 0.09223f
C4269 CDAC_v3_0.switch_4.Z.t1 GND 0.06525f
C4270 CDAC_v3_0.switch_4.Z.t2 GND 0.06525f
C4271 CDAC_v3_0.switch_4.Z.n0 GND 0.23436f
C4272 CDAC_v3_0.switch_4.Z.n1 GND 0.72258f
C4273 CDAC_v3_0.switch_4.Z.n2 GND 0.06761f
C4274 CDAC_v3_0.switch_4.Z.t14 GND 8.56099f
C4275 CDAC_v3_0.switch_4.Z.t18 GND 8.56099f
C4276 CDAC_v3_0.switch_4.Z.t7 GND 8.56099f
C4277 CDAC_v3_0.switch_4.Z.t10 GND 10.7681f
C4278 CDAC_v3_0.switch_4.Z.n3 GND 2.72934f
C4279 CDAC_v3_0.switch_4.Z.n4 GND 2.6404f
C4280 CDAC_v3_0.switch_4.Z.n5 GND 3.02056f
C4281 CDAC_v3_0.switch_4.Z.t16 GND 8.56099f
C4282 CDAC_v3_0.switch_4.Z.t19 GND 8.56099f
C4283 CDAC_v3_0.switch_4.Z.t8 GND 8.56099f
C4284 CDAC_v3_0.switch_4.Z.t12 GND 10.5936f
C4285 CDAC_v3_0.switch_4.Z.n6 GND 2.72231f
C4286 CDAC_v3_0.switch_4.Z.n7 GND 2.6404f
C4287 CDAC_v3_0.switch_4.Z.n8 GND 2.94179f
C4288 CDAC_v3_0.switch_4.Z.n9 GND 2.61915f
C4289 CDAC_v3_0.switch_4.Z.t5 GND 8.56099f
C4290 CDAC_v3_0.switch_4.Z.t4 GND 8.56099f
C4291 CDAC_v3_0.switch_4.Z.t6 GND 8.56099f
C4292 CDAC_v3_0.switch_4.Z.t9 GND 11.3609f
C4293 CDAC_v3_0.switch_4.Z.n10 GND 2.75323f
C4294 CDAC_v3_0.switch_4.Z.n11 GND 2.6404f
C4295 CDAC_v3_0.switch_4.Z.n12 GND 2.48992f
C4296 CDAC_v3_0.switch_4.Z.n13 GND 1.39753f
C4297 CDAC_v3_0.switch_4.Z.t13 GND 8.56099f
C4298 CDAC_v3_0.switch_4.Z.t11 GND 8.56099f
C4299 CDAC_v3_0.switch_4.Z.t15 GND 8.56099f
C4300 CDAC_v3_0.switch_4.Z.t17 GND 11.1864f
C4301 CDAC_v3_0.switch_4.Z.n14 GND 2.7462f
C4302 CDAC_v3_0.switch_4.Z.n15 GND 2.6404f
C4303 CDAC_v3_0.switch_4.Z.n16 GND 2.59534f
C4304 CDAC_v3_0.switch_4.Z.n17 GND 7.6393f
C4305 CDAC_v3_0.switch_4.Z.n18 GND 4.1383f
C4306 CDAC_v3_0.switch_4.Z.n19 GND 0.02147f
C4307 CDAC_v3_0.switch_4.Z.t0 GND 0.0632f
C4308 CDAC_v3_0.switch_4.Z.n20 GND 0.13877f
C4309 CDAC_v3_0.switch_4.Z.t3 GND 0.06307f
C4310 D_FlipFlop_7.3-input-nand_2.C.t1 GND 0.04469f
C4311 D_FlipFlop_7.3-input-nand_2.C.n0 GND 0.04327f
C4312 D_FlipFlop_7.3-input-nand_2.C.n1 GND 0.09193f
C4313 D_FlipFlop_7.3-input-nand_2.C.t6 GND 0.17806f
C4314 D_FlipFlop_7.3-input-nand_2.C.t7 GND 0.34248f
C4315 D_FlipFlop_7.3-input-nand_2.C.n2 GND 0.10005f
C4316 D_FlipFlop_7.3-input-nand_2.C.n3 GND 0.04279f
C4317 D_FlipFlop_7.3-input-nand_2.C.n4 GND 0.079f
C4318 D_FlipFlop_7.3-input-nand_2.C.n5 GND 0.13677f
C4319 D_FlipFlop_7.3-input-nand_2.C.n6 GND 0.10181f
C4320 D_FlipFlop_7.3-input-nand_2.C.n7 GND 0.04823f
C4321 D_FlipFlop_7.3-input-nand_2.C.t5 GND 0.3425f
C4322 D_FlipFlop_7.3-input-nand_2.C.n8 GND 0.3551f
C4323 D_FlipFlop_7.3-input-nand_2.C.n9 GND 0.03842f
C4324 D_FlipFlop_7.3-input-nand_2.C.n10 GND 0.05129f
C4325 D_FlipFlop_7.3-input-nand_2.C.t4 GND 0.17045f
C4326 D_FlipFlop_7.3-input-nand_2.C.t0 GND 0.04645f
C4327 D_FlipFlop_7.3-input-nand_2.C.n11 GND 0.293f
C4328 D_FlipFlop_7.3-input-nand_2.C.t3 GND 0.04742f
C4329 D_FlipFlop_7.3-input-nand_2.C.t2 GND 0.04645f
C4330 D_FlipFlop_7.3-input-nand_2.C.n12 GND 0.26418f
C4331 D_FlipFlop_7.3-input-nand_2.C.n13 GND 0.08722f
C4332 D_FlipFlop_7.3-input-nand_2.C.n14 GND 0.124f
C4333 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 GND 0.06443f
C4334 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 GND 0.14002f
C4335 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 GND 0.07316f
C4336 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 GND 0.25702f
C4337 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 GND 0.12462f
C4338 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 GND 0.4938f
C4339 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 GND 0.09136f
C4340 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 GND 0.05451f
C4341 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 GND 0.13379f
C4342 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 GND 0.13379f
C4343 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 GND 0.06713f
C4344 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 GND 0.07989f
C4345 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 GND 0.43786f
C4346 Ring_Counter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 GND 0.08018f
C4347 Q4.t3 GND 0.03196f
C4348 Q4.n0 GND 0.15671f
C4349 Q4.n1 GND 0.03572f
C4350 Q4.t0 GND 0.03392f
C4351 Q4.t1 GND 0.03323f
C4352 Q4.n2 GND 0.18898f
C4353 Q4.n3 GND 0.06166f
C4354 Q4.t2 GND 0.03323f
C4355 Q4.n4 GND 0.05119f
C4356 Q4.n5 GND 0.09064f
C4357 Q4.n6 GND 0.03575f
C4358 Q4.t9 GND 0.24499f
C4359 Q4.n7 GND 0.07157f
C4360 Q4.n8 GND 0.03105f
C4361 Q4.n9 GND 0.13653f
C4362 Q4.t6 GND 0.11394f
C4363 Q4.n10 GND 0.29918f
C4364 Q4.n11 GND 0.88845f
C4365 Q4.t8 GND 0.12746f
C4366 Q4.t5 GND 0.24611f
C4367 Q4.n12 GND 0.1827f
C4368 Q4.n13 GND 0.03381f
C4369 Q4.t7 GND 0.12746f
C4370 Q4.t4 GND 0.24611f
C4371 Q4.n14 GND 0.18156f
C4372 Q4.n15 GND 0.03642f
C4373 Q4.n16 GND 0.07573f
C4374 Q4.n17 GND 0.39779f
C4375 D_FlipFlop_7.3-input-nand_2.Vout.t7 GND 0.34247f
C4376 D_FlipFlop_7.3-input-nand_2.Vout.n0 GND 0.10005f
C4377 D_FlipFlop_7.3-input-nand_2.Vout.n1 GND 0.04341f
C4378 D_FlipFlop_7.3-input-nand_2.Vout.t3 GND 0.04467f
C4379 D_FlipFlop_7.3-input-nand_2.Vout.n2 GND 0.21241f
C4380 D_FlipFlop_7.3-input-nand_2.Vout.n3 GND 0.04823f
C4381 D_FlipFlop_7.3-input-nand_2.Vout.t4 GND 0.34248f
C4382 D_FlipFlop_7.3-input-nand_2.Vout.n4 GND 0.35447f
C4383 D_FlipFlop_7.3-input-nand_2.Vout.t6 GND 0.17806f
C4384 D_FlipFlop_7.3-input-nand_2.Vout.n5 GND 0.17459f
C4385 D_FlipFlop_7.3-input-nand_2.Vout.n6 GND 0.1018f
C4386 D_FlipFlop_7.3-input-nand_2.Vout.n7 GND 0.01283f
C4387 D_FlipFlop_7.3-input-nand_2.Vout.n8 GND 0.01019f
C4388 D_FlipFlop_7.3-input-nand_2.Vout.t1 GND 0.04742f
C4389 D_FlipFlop_7.3-input-nand_2.Vout.t0 GND 0.04645f
C4390 D_FlipFlop_7.3-input-nand_2.Vout.n9 GND 0.26417f
C4391 D_FlipFlop_7.3-input-nand_2.Vout.n10 GND 0.0862f
C4392 D_FlipFlop_7.3-input-nand_2.Vout.t2 GND 0.04645f
C4393 D_FlipFlop_7.3-input-nand_2.Vout.n11 GND 0.29241f
C4394 D_FlipFlop_7.3-input-nand_2.Vout.t5 GND 0.17113f
C4395 D_FlipFlop_7.3-input-nand_2.Vout.n12 GND 0.19086f
C4396 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 GND 0.07411f
C4397 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 GND 0.16107f
C4398 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 GND 0.08416f
C4399 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 GND 0.29566f
C4400 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 GND 0.14335f
C4401 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 GND 0.56804f
C4402 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 GND 0.1051f
C4403 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 GND 0.06271f
C4404 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 GND 0.15391f
C4405 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 GND 0.15391f
C4406 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 GND 0.07722f
C4407 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 GND 0.07866f
C4408 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 GND 0.07705f
C4409 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 GND 0.43817f
C4410 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 GND 0.286f
C4411 Ring_Counter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 GND 0.09223f
C4412 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 GND 0.07411f
C4413 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 GND 0.16107f
C4414 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 GND 0.08416f
C4415 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 GND 0.29566f
C4416 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 GND 0.14335f
C4417 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 GND 0.56804f
C4418 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 GND 0.1051f
C4419 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 GND 0.06271f
C4420 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 GND 0.15391f
C4421 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 GND 0.15391f
C4422 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 GND 0.07722f
C4423 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 GND 0.07866f
C4424 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 GND 0.07705f
C4425 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 GND 0.43817f
C4426 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 GND 0.286f
C4427 Ring_Counter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 GND 0.09223f
C4428 Nand_Gate_5.A.t2 GND 0.05077f
C4429 Nand_Gate_5.A.t10 GND 0.36044f
C4430 Nand_Gate_5.A.n0 GND 0.1053f
C4431 Nand_Gate_5.A.n1 GND 0.04569f
C4432 Nand_Gate_5.A.n2 GND 0.20088f
C4433 Nand_Gate_5.A.t7 GND 0.22562f
C4434 Nand_Gate_5.A.t11 GND 0.1874f
C4435 Nand_Gate_5.A.n3 GND 0.04909f
C4436 Nand_Gate_5.A.n4 GND 0.04503f
C4437 Nand_Gate_5.A.t6 GND 0.36093f
C4438 Nand_Gate_5.A.n5 GND 0.10827f
C4439 Nand_Gate_5.A.t4 GND 0.1874f
C4440 Nand_Gate_5.A.n6 GND 0.04909f
C4441 Nand_Gate_5.A.n7 GND 0.04503f
C4442 Nand_Gate_5.A.n8 GND 0.11393f
C4443 Nand_Gate_5.A.n9 GND 0.11393f
C4444 Nand_Gate_5.A.n10 GND 0.10827f
C4445 Nand_Gate_5.A.t9 GND 0.46089f
C4446 Nand_Gate_5.A.n11 GND 0.11304f
C4447 Nand_Gate_5.A.n12 GND 1.66069f
C4448 Nand_Gate_5.A.n13 GND 0.22898f
C4449 Nand_Gate_5.A.t5 GND 0.36044f
C4450 Nand_Gate_5.A.n14 GND 0.15699f
C4451 Nand_Gate_5.A.t8 GND 0.16824f
C4452 Nand_Gate_5.A.n15 GND 0.10982f
C4453 Nand_Gate_5.A.n16 GND 0.05259f
C4454 Nand_Gate_5.A.n17 GND 0.13335f
C4455 Nand_Gate_5.A.t1 GND 0.04889f
C4456 Nand_Gate_5.A.n18 GND 0.07531f
C4457 Nand_Gate_5.A.t3 GND 0.04991f
C4458 Nand_Gate_5.A.t0 GND 0.04889f
C4459 Nand_Gate_5.A.n19 GND 0.27804f
C4460 Nand_Gate_5.A.n20 GND 0.09072f
C4461 Nand_Gate_5.A.n21 GND 0.18266f
C4462 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 GND 0.06443f
C4463 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 GND 0.14002f
C4464 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 GND 0.07316f
C4465 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 GND 0.25702f
C4466 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 GND 0.12462f
C4467 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 GND 0.4938f
C4468 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 GND 0.09136f
C4469 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 GND 0.05451f
C4470 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 GND 0.13379f
C4471 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 GND 0.13379f
C4472 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 GND 0.06713f
C4473 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 GND 0.07989f
C4474 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 GND 0.43786f
C4475 Ring_Counter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 GND 0.08018f
C4476 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t1 GND 0.05f
C4477 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n0 GND 0.10867f
C4478 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n1 GND 0.05678f
C4479 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t4 GND 0.38491f
C4480 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n2 GND 0.16589f
C4481 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t5 GND 0.30131f
C4482 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t3 GND 0.30153f
C4483 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n3 GND 0.09671f
C4484 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t2 GND 0.38323f
C4485 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n4 GND 0.0709f
C4486 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n5 GND 0.04231f
C4487 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n6 GND 0.10383f
C4488 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n7 GND 0.10383f
C4489 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.t0 GND 0.05284f
C4490 Ring_Counter_0.D_FlipFlop_1.Inverter_1.Vout.n8 GND 0.17757f
C4491 Ring_Counter_0.D_FlipFlop_4.Qbar.t5 GND 0.41161f
C4492 Ring_Counter_0.D_FlipFlop_4.Qbar.n0 GND 0.1774f
C4493 Ring_Counter_0.D_FlipFlop_4.Qbar.t4 GND 0.18986f
C4494 Ring_Counter_0.D_FlipFlop_4.Qbar.n1 GND 0.23199f
C4495 Ring_Counter_0.D_FlipFlop_4.Qbar.n2 GND 0.05991f
C4496 Ring_Counter_0.D_FlipFlop_4.Qbar.t1 GND 0.05347f
C4497 Ring_Counter_0.D_FlipFlop_4.Qbar.n3 GND 0.15403f
C4498 Ring_Counter_0.D_FlipFlop_4.Qbar.t2 GND 0.05675f
C4499 Ring_Counter_0.D_FlipFlop_4.Qbar.t3 GND 0.05559f
C4500 Ring_Counter_0.D_FlipFlop_4.Qbar.n4 GND 0.31612f
C4501 Ring_Counter_0.D_FlipFlop_4.Qbar.n5 GND 0.16106f
C4502 Ring_Counter_0.D_FlipFlop_4.Qbar.t0 GND 0.05559f
C4503 Ring_Counter_0.D_FlipFlop_4.Qbar.n6 GND 0.09627f
C4504 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t1 GND 0.05f
C4505 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n0 GND 0.10867f
C4506 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n1 GND 0.05678f
C4507 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t4 GND 0.38491f
C4508 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n2 GND 0.16589f
C4509 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t2 GND 0.30131f
C4510 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t3 GND 0.30153f
C4511 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n3 GND 0.09671f
C4512 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t5 GND 0.38323f
C4513 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n4 GND 0.0709f
C4514 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n5 GND 0.04231f
C4515 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n6 GND 0.10383f
C4516 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n7 GND 0.10383f
C4517 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.t0 GND 0.05284f
C4518 Ring_Counter_0.D_FlipFlop_5.Inverter_1.Vout.n8 GND 0.17757f
C4519 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 GND 0.06443f
C4520 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 GND 0.14002f
C4521 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 GND 0.07316f
C4522 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 GND 0.25702f
C4523 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 GND 0.12462f
C4524 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 GND 0.4938f
C4525 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 GND 0.09136f
C4526 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 GND 0.05451f
C4527 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 GND 0.13379f
C4528 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 GND 0.13379f
C4529 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 GND 0.06713f
C4530 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 GND 0.07989f
C4531 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 GND 0.43786f
C4532 Ring_Counter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 GND 0.08018f
C4533 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 GND 0.06443f
C4534 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 GND 0.14002f
C4535 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 GND 0.07316f
C4536 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 GND 0.25702f
C4537 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 GND 0.12462f
C4538 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 GND 0.4938f
C4539 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 GND 0.09136f
C4540 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 GND 0.05451f
C4541 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 GND 0.13379f
C4542 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 GND 0.13379f
C4543 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 GND 0.06713f
C4544 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 GND 0.07989f
C4545 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 GND 0.43786f
C4546 Ring_Counter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 GND 0.08018f
C4547 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t3 GND 0.05969f
C4548 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n0 GND 0.15363f
C4549 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n1 GND 0.12493f
C4550 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t6 GND 0.23786f
C4551 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t4 GND 0.4575f
C4552 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n2 GND 0.10854f
C4553 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n3 GND 0.10766f
C4554 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n4 GND 0.1827f
C4555 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n5 GND 0.136f
C4556 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t7 GND 0.4595f
C4557 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n6 GND 0.19804f
C4558 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t5 GND 0.22769f
C4559 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t2 GND 0.06205f
C4560 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n7 GND 0.3914f
C4561 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t0 GND 0.06335f
C4562 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.t1 GND 0.06205f
C4563 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n8 GND 0.3529f
C4564 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n9 GND 0.12232f
C4565 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.C.n10 GND 0.07613f
C4566 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t1 GND 0.05f
C4567 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n0 GND 0.10867f
C4568 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n1 GND 0.05678f
C4569 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t5 GND 0.38491f
C4570 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n2 GND 0.16589f
C4571 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t3 GND 0.30131f
C4572 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t2 GND 0.30153f
C4573 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n3 GND 0.09671f
C4574 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t4 GND 0.38323f
C4575 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n4 GND 0.0709f
C4576 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n5 GND 0.04231f
C4577 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n6 GND 0.10383f
C4578 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n7 GND 0.10383f
C4579 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.t0 GND 0.05284f
C4580 Ring_Counter_0.D_FlipFlop_15.Inverter_1.Vout.n8 GND 0.17757f
C4581 D_FlipFlop_5.3-input-nand_2.Vout.t6 GND 0.34247f
C4582 D_FlipFlop_5.3-input-nand_2.Vout.n0 GND 0.10005f
C4583 D_FlipFlop_5.3-input-nand_2.Vout.n1 GND 0.04341f
C4584 D_FlipFlop_5.3-input-nand_2.Vout.n2 GND 0.19086f
C4585 D_FlipFlop_5.3-input-nand_2.Vout.t5 GND 0.17113f
C4586 D_FlipFlop_5.3-input-nand_2.Vout.t2 GND 0.04645f
C4587 D_FlipFlop_5.3-input-nand_2.Vout.n3 GND 0.29241f
C4588 D_FlipFlop_5.3-input-nand_2.Vout.t1 GND 0.04742f
C4589 D_FlipFlop_5.3-input-nand_2.Vout.t3 GND 0.04645f
C4590 D_FlipFlop_5.3-input-nand_2.Vout.n4 GND 0.26417f
C4591 D_FlipFlop_5.3-input-nand_2.Vout.n5 GND 0.0862f
C4592 D_FlipFlop_5.3-input-nand_2.Vout.n6 GND 0.01019f
C4593 D_FlipFlop_5.3-input-nand_2.Vout.n7 GND 0.01283f
C4594 D_FlipFlop_5.3-input-nand_2.Vout.t4 GND 0.34248f
C4595 D_FlipFlop_5.3-input-nand_2.Vout.n8 GND 0.35447f
C4596 D_FlipFlop_5.3-input-nand_2.Vout.t7 GND 0.17806f
C4597 D_FlipFlop_5.3-input-nand_2.Vout.n9 GND 0.17459f
C4598 D_FlipFlop_5.3-input-nand_2.Vout.n10 GND 0.1018f
C4599 D_FlipFlop_5.3-input-nand_2.Vout.n11 GND 0.04823f
C4600 D_FlipFlop_5.3-input-nand_2.Vout.t0 GND 0.04467f
C4601 D_FlipFlop_5.3-input-nand_2.Vout.n12 GND 0.21241f
C4602 D_FlipFlop_3.3-input-nand_2.C.t7 GND 0.3425f
C4603 D_FlipFlop_3.3-input-nand_2.C.n0 GND 0.3551f
C4604 D_FlipFlop_3.3-input-nand_2.C.n1 GND 0.03842f
C4605 D_FlipFlop_3.3-input-nand_2.C.t3 GND 0.04469f
C4606 D_FlipFlop_3.3-input-nand_2.C.n2 GND 0.04327f
C4607 D_FlipFlop_3.3-input-nand_2.C.n3 GND 0.09193f
C4608 D_FlipFlop_3.3-input-nand_2.C.t5 GND 0.17806f
C4609 D_FlipFlop_3.3-input-nand_2.C.t6 GND 0.34248f
C4610 D_FlipFlop_3.3-input-nand_2.C.n4 GND 0.10005f
C4611 D_FlipFlop_3.3-input-nand_2.C.n5 GND 0.04279f
C4612 D_FlipFlop_3.3-input-nand_2.C.n6 GND 0.079f
C4613 D_FlipFlop_3.3-input-nand_2.C.n7 GND 0.13677f
C4614 D_FlipFlop_3.3-input-nand_2.C.n8 GND 0.10181f
C4615 D_FlipFlop_3.3-input-nand_2.C.n9 GND 0.04823f
C4616 D_FlipFlop_3.3-input-nand_2.C.n10 GND 0.124f
C4617 D_FlipFlop_3.3-input-nand_2.C.t1 GND 0.04742f
C4618 D_FlipFlop_3.3-input-nand_2.C.t0 GND 0.04645f
C4619 D_FlipFlop_3.3-input-nand_2.C.n11 GND 0.26418f
C4620 D_FlipFlop_3.3-input-nand_2.C.n12 GND 0.08722f
C4621 D_FlipFlop_3.3-input-nand_2.C.t2 GND 0.04645f
C4622 D_FlipFlop_3.3-input-nand_2.C.n13 GND 0.293f
C4623 D_FlipFlop_3.3-input-nand_2.C.t4 GND 0.17045f
C4624 D_FlipFlop_3.3-input-nand_2.C.n14 GND 0.05129f
C4625 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 GND 0.07411f
C4626 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 GND 0.16107f
C4627 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 GND 0.08416f
C4628 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 GND 0.29566f
C4629 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 GND 0.14335f
C4630 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 GND 0.56804f
C4631 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 GND 0.1051f
C4632 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 GND 0.06271f
C4633 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 GND 0.15391f
C4634 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 GND 0.15391f
C4635 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 GND 0.07722f
C4636 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 GND 0.07866f
C4637 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 GND 0.07705f
C4638 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 GND 0.43817f
C4639 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 GND 0.286f
C4640 Ring_Counter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 GND 0.09223f
C4641 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 GND 0.05215f
C4642 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 GND 0.18008f
C4643 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 GND 0.37825f
C4644 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 GND 0.19588f
C4645 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 GND 0.28346f
C4646 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 GND 0.11199f
C4647 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 GND 0.01587f
C4648 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 GND 0.37675f
C4649 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 GND 0.16409f
C4650 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 GND 0.18888f
C4651 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 GND 0.0511f
C4652 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 GND 0.32168f
C4653 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 GND 0.05217f
C4654 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 GND 0.0511f
C4655 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 GND 0.29061f
C4656 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 GND 0.09483f
C4657 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 GND 0.01203f
C4658 D_FlipFlop_3.3-input-nand_2.Vout.t5 GND 0.34247f
C4659 D_FlipFlop_3.3-input-nand_2.Vout.n0 GND 0.10005f
C4660 D_FlipFlop_3.3-input-nand_2.Vout.n1 GND 0.04341f
C4661 D_FlipFlop_3.3-input-nand_2.Vout.t3 GND 0.04467f
C4662 D_FlipFlop_3.3-input-nand_2.Vout.n2 GND 0.21241f
C4663 D_FlipFlop_3.3-input-nand_2.Vout.n3 GND 0.04823f
C4664 D_FlipFlop_3.3-input-nand_2.Vout.t7 GND 0.34248f
C4665 D_FlipFlop_3.3-input-nand_2.Vout.n4 GND 0.35447f
C4666 D_FlipFlop_3.3-input-nand_2.Vout.t6 GND 0.17806f
C4667 D_FlipFlop_3.3-input-nand_2.Vout.n5 GND 0.17459f
C4668 D_FlipFlop_3.3-input-nand_2.Vout.n6 GND 0.1018f
C4669 D_FlipFlop_3.3-input-nand_2.Vout.n7 GND 0.01283f
C4670 D_FlipFlop_3.3-input-nand_2.Vout.n8 GND 0.01019f
C4671 D_FlipFlop_3.3-input-nand_2.Vout.t1 GND 0.04742f
C4672 D_FlipFlop_3.3-input-nand_2.Vout.t0 GND 0.04645f
C4673 D_FlipFlop_3.3-input-nand_2.Vout.n9 GND 0.26417f
C4674 D_FlipFlop_3.3-input-nand_2.Vout.n10 GND 0.0862f
C4675 D_FlipFlop_3.3-input-nand_2.Vout.t2 GND 0.04645f
C4676 D_FlipFlop_3.3-input-nand_2.Vout.n11 GND 0.29241f
C4677 D_FlipFlop_3.3-input-nand_2.Vout.t4 GND 0.17113f
C4678 D_FlipFlop_3.3-input-nand_2.Vout.n12 GND 0.19086f
C4679 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t1 GND 0.05f
C4680 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n0 GND 0.10867f
C4681 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n1 GND 0.05678f
C4682 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t4 GND 0.38491f
C4683 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n2 GND 0.16589f
C4684 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t2 GND 0.30131f
C4685 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t3 GND 0.30153f
C4686 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n3 GND 0.09671f
C4687 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t5 GND 0.38323f
C4688 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n4 GND 0.0709f
C4689 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n5 GND 0.04231f
C4690 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n6 GND 0.10383f
C4691 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n7 GND 0.10383f
C4692 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.t0 GND 0.05284f
C4693 Ring_Counter_0.D_FlipFlop_7.Inverter_1.Vout.n8 GND 0.17757f
C4694 Q3.t1 GND 0.03635f
C4695 Q3.n0 GND 0.17828f
C4696 Q3.n1 GND 0.04063f
C4697 Q3.t2 GND 0.03859f
C4698 Q3.t3 GND 0.0378f
C4699 Q3.n2 GND 0.21499f
C4700 Q3.n3 GND 0.07015f
C4701 Q3.t0 GND 0.0378f
C4702 Q3.n4 GND 0.05823f
C4703 Q3.n5 GND 0.10311f
C4704 Q3.n6 GND 0.04067f
C4705 Q3.t5 GND 0.27871f
C4706 Q3.n7 GND 0.08142f
C4707 Q3.n8 GND 0.03533f
C4708 Q3.n9 GND 0.15533f
C4709 Q3.t9 GND 0.12962f
C4710 Q3.n10 GND 0.35398f
C4711 Q3.n11 GND 0.27121f
C4712 Q3.t8 GND 0.145f
C4713 Q3.t4 GND 0.27998f
C4714 Q3.n12 GND 0.20785f
C4715 Q3.n13 GND 0.03846f
C4716 Q3.t7 GND 0.145f
C4717 Q3.t6 GND 0.27998f
C4718 Q3.n14 GND 0.20655f
C4719 Q3.n15 GND 0.04143f
C4720 Q3.n16 GND 0.07978f
C4721 Q3.n17 GND 0.09791f
C4722 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 GND 0.07411f
C4723 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 GND 0.16107f
C4724 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 GND 0.08416f
C4725 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 GND 0.29566f
C4726 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 GND 0.14335f
C4727 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 GND 0.56804f
C4728 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 GND 0.1051f
C4729 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 GND 0.06271f
C4730 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 GND 0.15391f
C4731 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 GND 0.15391f
C4732 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 GND 0.07722f
C4733 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 GND 0.07866f
C4734 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 GND 0.07705f
C4735 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 GND 0.43817f
C4736 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 GND 0.286f
C4737 Ring_Counter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 GND 0.09223f
C4738 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t3 GND 0.06145f
C4739 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n0 GND 0.15815f
C4740 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n1 GND 0.12861f
C4741 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t5 GND 0.24486f
C4742 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t4 GND 0.47095f
C4743 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n2 GND 0.11174f
C4744 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n3 GND 0.11082f
C4745 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n4 GND 0.18808f
C4746 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n5 GND 0.14f
C4747 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t7 GND 0.47302f
C4748 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n6 GND 0.20386f
C4749 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t6 GND 0.23439f
C4750 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t2 GND 0.06388f
C4751 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n7 GND 0.40291f
C4752 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t0 GND 0.06521f
C4753 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.t1 GND 0.06388f
C4754 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n8 GND 0.36328f
C4755 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n9 GND 0.12591f
C4756 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.C.n10 GND 0.07837f
C4757 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t1 GND 0.05f
C4758 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n0 GND 0.10867f
C4759 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n1 GND 0.05678f
C4760 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t5 GND 0.38491f
C4761 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n2 GND 0.16589f
C4762 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t2 GND 0.30131f
C4763 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t4 GND 0.30153f
C4764 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n3 GND 0.09671f
C4765 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t3 GND 0.38323f
C4766 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n4 GND 0.0709f
C4767 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n5 GND 0.04231f
C4768 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n6 GND 0.10383f
C4769 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n7 GND 0.10383f
C4770 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.t0 GND 0.05284f
C4771 Ring_Counter_0.D_FlipFlop_16.Inverter_1.Vout.n8 GND 0.17757f
C4772 Q2.t7 GND 0.13741f
C4773 Q2.t5 GND 0.26533f
C4774 Q2.n0 GND 0.19697f
C4775 Q2.n1 GND 0.03645f
C4776 Q2.t8 GND 0.13741f
C4777 Q2.t4 GND 0.26533f
C4778 Q2.n2 GND 0.19574f
C4779 Q2.n3 GND 0.03926f
C4780 Q2.n4 GND 0.06963f
C4781 Q2.n5 GND 0.62922f
C4782 Q2.t1 GND 0.03445f
C4783 Q2.n6 GND 0.16895f
C4784 Q2.n7 GND 0.0385f
C4785 Q2.t2 GND 0.03657f
C4786 Q2.t3 GND 0.03582f
C4787 Q2.n8 GND 0.20374f
C4788 Q2.n9 GND 0.06648f
C4789 Q2.t0 GND 0.03582f
C4790 Q2.n10 GND 0.05519f
C4791 Q2.n11 GND 0.09771f
C4792 Q2.n12 GND 0.03854f
C4793 Q2.t9 GND 0.26412f
C4794 Q2.n13 GND 0.07716f
C4795 Q2.n14 GND 0.03348f
C4796 Q2.n15 GND 0.1472f
C4797 Q2.t6 GND 0.12284f
C4798 Q2.n16 GND 0.34819f
C4799 Q2.n17 GND 0.23438f
C4800 D_FlipFlop_1.3-input-nand_2.Vout.t5 GND 0.34247f
C4801 D_FlipFlop_1.3-input-nand_2.Vout.n0 GND 0.10005f
C4802 D_FlipFlop_1.3-input-nand_2.Vout.n1 GND 0.04341f
C4803 D_FlipFlop_1.3-input-nand_2.Vout.t1 GND 0.04467f
C4804 D_FlipFlop_1.3-input-nand_2.Vout.n2 GND 0.21241f
C4805 D_FlipFlop_1.3-input-nand_2.Vout.n3 GND 0.04823f
C4806 D_FlipFlop_1.3-input-nand_2.Vout.t6 GND 0.34248f
C4807 D_FlipFlop_1.3-input-nand_2.Vout.n4 GND 0.35447f
C4808 D_FlipFlop_1.3-input-nand_2.Vout.t7 GND 0.17806f
C4809 D_FlipFlop_1.3-input-nand_2.Vout.n5 GND 0.17459f
C4810 D_FlipFlop_1.3-input-nand_2.Vout.n6 GND 0.1018f
C4811 D_FlipFlop_1.3-input-nand_2.Vout.n7 GND 0.01283f
C4812 D_FlipFlop_1.3-input-nand_2.Vout.n8 GND 0.01019f
C4813 D_FlipFlop_1.3-input-nand_2.Vout.t2 GND 0.04742f
C4814 D_FlipFlop_1.3-input-nand_2.Vout.t3 GND 0.04645f
C4815 D_FlipFlop_1.3-input-nand_2.Vout.n9 GND 0.26417f
C4816 D_FlipFlop_1.3-input-nand_2.Vout.n10 GND 0.0862f
C4817 D_FlipFlop_1.3-input-nand_2.Vout.t0 GND 0.04645f
C4818 D_FlipFlop_1.3-input-nand_2.Vout.n11 GND 0.29241f
C4819 D_FlipFlop_1.3-input-nand_2.Vout.t4 GND 0.17113f
C4820 D_FlipFlop_1.3-input-nand_2.Vout.n12 GND 0.19086f
C4821 D_FlipFlop_1.3-input-nand_2.C.t1 GND 0.04469f
C4822 D_FlipFlop_1.3-input-nand_2.C.n0 GND 0.04327f
C4823 D_FlipFlop_1.3-input-nand_2.C.n1 GND 0.09193f
C4824 D_FlipFlop_1.3-input-nand_2.C.t5 GND 0.17806f
C4825 D_FlipFlop_1.3-input-nand_2.C.t7 GND 0.34248f
C4826 D_FlipFlop_1.3-input-nand_2.C.n2 GND 0.10005f
C4827 D_FlipFlop_1.3-input-nand_2.C.n3 GND 0.04279f
C4828 D_FlipFlop_1.3-input-nand_2.C.n4 GND 0.079f
C4829 D_FlipFlop_1.3-input-nand_2.C.n5 GND 0.13677f
C4830 D_FlipFlop_1.3-input-nand_2.C.n6 GND 0.10181f
C4831 D_FlipFlop_1.3-input-nand_2.C.n7 GND 0.04823f
C4832 D_FlipFlop_1.3-input-nand_2.C.t6 GND 0.3425f
C4833 D_FlipFlop_1.3-input-nand_2.C.n8 GND 0.3551f
C4834 D_FlipFlop_1.3-input-nand_2.C.n9 GND 0.03842f
C4835 D_FlipFlop_1.3-input-nand_2.C.n10 GND 0.05129f
C4836 D_FlipFlop_1.3-input-nand_2.C.t4 GND 0.17045f
C4837 D_FlipFlop_1.3-input-nand_2.C.t0 GND 0.04645f
C4838 D_FlipFlop_1.3-input-nand_2.C.n11 GND 0.293f
C4839 D_FlipFlop_1.3-input-nand_2.C.t3 GND 0.04742f
C4840 D_FlipFlop_1.3-input-nand_2.C.t2 GND 0.04645f
C4841 D_FlipFlop_1.3-input-nand_2.C.n12 GND 0.26418f
C4842 D_FlipFlop_1.3-input-nand_2.C.n13 GND 0.08722f
C4843 D_FlipFlop_1.3-input-nand_2.C.n14 GND 0.124f
C4844 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t2 GND 0.06145f
C4845 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n0 GND 0.15815f
C4846 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n1 GND 0.12861f
C4847 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t7 GND 0.24486f
C4848 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t4 GND 0.47095f
C4849 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n2 GND 0.11174f
C4850 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n3 GND 0.11082f
C4851 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n4 GND 0.18808f
C4852 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n5 GND 0.14f
C4853 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t5 GND 0.47302f
C4854 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n6 GND 0.20386f
C4855 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t6 GND 0.23439f
C4856 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t3 GND 0.06388f
C4857 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n7 GND 0.40291f
C4858 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t0 GND 0.06521f
C4859 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.t1 GND 0.06388f
C4860 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n8 GND 0.36328f
C4861 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n9 GND 0.12591f
C4862 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.C.n10 GND 0.07837f
C4863 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t3 GND 0.06145f
C4864 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n0 GND 0.15815f
C4865 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n1 GND 0.12861f
C4866 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t5 GND 0.24486f
C4867 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t7 GND 0.47095f
C4868 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n2 GND 0.11174f
C4869 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n3 GND 0.11082f
C4870 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n4 GND 0.18808f
C4871 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n5 GND 0.14f
C4872 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t6 GND 0.47302f
C4873 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n6 GND 0.20386f
C4874 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t4 GND 0.23439f
C4875 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t2 GND 0.06388f
C4876 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n7 GND 0.40291f
C4877 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t1 GND 0.06521f
C4878 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.t0 GND 0.06388f
C4879 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n8 GND 0.36328f
C4880 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n9 GND 0.12591f
C4881 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.C.n10 GND 0.07837f
C4882 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 GND 0.06443f
C4883 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 GND 0.14002f
C4884 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 GND 0.07316f
C4885 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 GND 0.25702f
C4886 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 GND 0.12462f
C4887 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 GND 0.4938f
C4888 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 GND 0.09136f
C4889 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 GND 0.05451f
C4890 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 GND 0.13379f
C4891 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 GND 0.13379f
C4892 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 GND 0.06713f
C4893 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 GND 0.07989f
C4894 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 GND 0.43786f
C4895 Ring_Counter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 GND 0.08018f
C4896 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t1 GND 0.06145f
C4897 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n0 GND 0.15815f
C4898 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n1 GND 0.12861f
C4899 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t4 GND 0.24486f
C4900 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t6 GND 0.47095f
C4901 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n2 GND 0.11174f
C4902 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n3 GND 0.11082f
C4903 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n4 GND 0.18808f
C4904 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n5 GND 0.14f
C4905 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t7 GND 0.47302f
C4906 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n6 GND 0.20386f
C4907 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t5 GND 0.23439f
C4908 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t3 GND 0.06388f
C4909 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n7 GND 0.40291f
C4910 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t0 GND 0.06521f
C4911 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.t2 GND 0.06388f
C4912 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n8 GND 0.36328f
C4913 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n9 GND 0.12591f
C4914 Ring_Counter_0.D_FlipFlop_8.3-input-nand_2.C.n10 GND 0.07837f
C4915 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 GND 0.05215f
C4916 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 GND 0.18008f
C4917 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 GND 0.37825f
C4918 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 GND 0.19588f
C4919 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 GND 0.28346f
C4920 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 GND 0.11199f
C4921 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 GND 0.01587f
C4922 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 GND 0.37675f
C4923 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 GND 0.16409f
C4924 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 GND 0.18888f
C4925 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 GND 0.0511f
C4926 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 GND 0.32168f
C4927 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 GND 0.05217f
C4928 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 GND 0.0511f
C4929 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 GND 0.29061f
C4930 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 GND 0.09483f
C4931 Ring_Counter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 GND 0.01203f
C4932 Ring_Counter_0.D_FlipFlop_16.Q.t3 GND 0.10344f
C4933 Ring_Counter_0.D_FlipFlop_16.Q.t8 GND 0.7344f
C4934 Ring_Counter_0.D_FlipFlop_16.Q.n0 GND 0.31987f
C4935 Ring_Counter_0.D_FlipFlop_16.Q.t9 GND 0.34281f
C4936 Ring_Counter_0.D_FlipFlop_16.Q.n1 GND 0.03889f
C4937 Ring_Counter_0.D_FlipFlop_16.Q.n2 GND 0.0855f
C4938 Ring_Counter_0.D_FlipFlop_16.Q.t7 GND 0.7354f
C4939 Ring_Counter_0.D_FlipFlop_16.Q.n3 GND 0.22061f
C4940 Ring_Counter_0.D_FlipFlop_16.Q.t6 GND 0.38183f
C4941 Ring_Counter_0.D_FlipFlop_16.Q.n4 GND 0.10003f
C4942 Ring_Counter_0.D_FlipFlop_16.Q.n5 GND 0.09174f
C4943 Ring_Counter_0.D_FlipFlop_16.Q.n6 GND 0.11063f
C4944 Ring_Counter_0.D_FlipFlop_16.Q.t4 GND 0.7354f
C4945 Ring_Counter_0.D_FlipFlop_16.Q.n7 GND 0.22061f
C4946 Ring_Counter_0.D_FlipFlop_16.Q.t5 GND 0.38183f
C4947 Ring_Counter_0.D_FlipFlop_16.Q.n8 GND 0.10003f
C4948 Ring_Counter_0.D_FlipFlop_16.Q.n9 GND 0.09174f
C4949 Ring_Counter_0.D_FlipFlop_16.Q.n10 GND 0.01324f
C4950 Ring_Counter_0.D_FlipFlop_16.Q.n11 GND 15.259f
C4951 Ring_Counter_0.D_FlipFlop_16.Q.n12 GND 9.67439f
C4952 Ring_Counter_0.D_FlipFlop_16.Q.n13 GND 0.11314f
C4953 Ring_Counter_0.D_FlipFlop_16.Q.n14 GND 0.22205f
C4954 Ring_Counter_0.D_FlipFlop_16.Q.t2 GND 0.09961f
C4955 Ring_Counter_0.D_FlipFlop_16.Q.n15 GND 0.15345f
C4956 Ring_Counter_0.D_FlipFlop_16.Q.t1 GND 0.1017f
C4957 Ring_Counter_0.D_FlipFlop_16.Q.t0 GND 0.09961f
C4958 Ring_Counter_0.D_FlipFlop_16.Q.n16 GND 0.5665f
C4959 Ring_Counter_0.D_FlipFlop_16.Q.n17 GND 0.18485f
C4960 Ring_Counter_0.D_FlipFlop_16.Q.n18 GND 0.37218f
C4961 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 GND 0.37675f
C4962 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 GND 0.16409f
C4963 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 GND 0.18888f
C4964 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 GND 0.0511f
C4965 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 GND 0.32168f
C4966 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 GND 0.05217f
C4967 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 GND 0.0511f
C4968 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 GND 0.29061f
C4969 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 GND 0.09483f
C4970 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 GND 0.01203f
C4971 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 GND 0.01587f
C4972 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 GND 0.37825f
C4973 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 GND 0.19588f
C4974 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 GND 0.28346f
C4975 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 GND 0.11199f
C4976 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 GND 0.05215f
C4977 Ring_Counter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 GND 0.18008f
C4978 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t1 GND 0.06616f
C4979 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n0 GND 0.21243f
C4980 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t4 GND 0.49448f
C4981 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n1 GND 0.14833f
C4982 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t3 GND 0.25674f
C4983 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n2 GND 0.06726f
C4984 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n3 GND 0.06169f
C4985 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n4 GND 0.13379f
C4986 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n5 GND 0.13379f
C4987 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n6 GND 0.08249f
C4988 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t0 GND 0.06713f
C4989 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.t2 GND 0.07989f
C4990 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n7 GND 0.40234f
C4991 Ring_Counter_0.D_FlipFlop_0.Nand_Gate_0.Vout.n8 GND 0.04156f
C4992 D_FlipFlop_6.3-input-nand_2.C.t1 GND 0.04469f
C4993 D_FlipFlop_6.3-input-nand_2.C.n0 GND 0.04327f
C4994 D_FlipFlop_6.3-input-nand_2.C.n1 GND 0.09193f
C4995 D_FlipFlop_6.3-input-nand_2.C.t4 GND 0.17806f
C4996 D_FlipFlop_6.3-input-nand_2.C.t6 GND 0.34248f
C4997 D_FlipFlop_6.3-input-nand_2.C.n2 GND 0.10005f
C4998 D_FlipFlop_6.3-input-nand_2.C.n3 GND 0.04279f
C4999 D_FlipFlop_6.3-input-nand_2.C.n4 GND 0.079f
C5000 D_FlipFlop_6.3-input-nand_2.C.n5 GND 0.13677f
C5001 D_FlipFlop_6.3-input-nand_2.C.n6 GND 0.10181f
C5002 D_FlipFlop_6.3-input-nand_2.C.n7 GND 0.04823f
C5003 D_FlipFlop_6.3-input-nand_2.C.t5 GND 0.3425f
C5004 D_FlipFlop_6.3-input-nand_2.C.n8 GND 0.3551f
C5005 D_FlipFlop_6.3-input-nand_2.C.n9 GND 0.03842f
C5006 D_FlipFlop_6.3-input-nand_2.C.n10 GND 0.05129f
C5007 D_FlipFlop_6.3-input-nand_2.C.t7 GND 0.17045f
C5008 D_FlipFlop_6.3-input-nand_2.C.t0 GND 0.04645f
C5009 D_FlipFlop_6.3-input-nand_2.C.n11 GND 0.293f
C5010 D_FlipFlop_6.3-input-nand_2.C.t2 GND 0.04742f
C5011 D_FlipFlop_6.3-input-nand_2.C.t3 GND 0.04645f
C5012 D_FlipFlop_6.3-input-nand_2.C.n12 GND 0.26418f
C5013 D_FlipFlop_6.3-input-nand_2.C.n13 GND 0.08722f
C5014 D_FlipFlop_6.3-input-nand_2.C.n14 GND 0.124f
C5015 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 GND 0.06443f
C5016 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 GND 0.14002f
C5017 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 GND 0.07316f
C5018 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 GND 0.25702f
C5019 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 GND 0.12462f
C5020 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 GND 0.4938f
C5021 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 GND 0.09136f
C5022 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 GND 0.05451f
C5023 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 GND 0.13379f
C5024 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 GND 0.13379f
C5025 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 GND 0.06713f
C5026 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 GND 0.07989f
C5027 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 GND 0.43786f
C5028 Ring_Counter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 GND 0.08018f
C5029 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t1 GND 0.05f
C5030 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n0 GND 0.10867f
C5031 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n1 GND 0.05678f
C5032 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t4 GND 0.38491f
C5033 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n2 GND 0.16589f
C5034 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t5 GND 0.30131f
C5035 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t3 GND 0.30153f
C5036 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n3 GND 0.09671f
C5037 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t2 GND 0.38323f
C5038 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n4 GND 0.0709f
C5039 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n5 GND 0.04231f
C5040 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n6 GND 0.10383f
C5041 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n7 GND 0.10383f
C5042 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.t0 GND 0.05284f
C5043 Ring_Counter_0.D_FlipFlop_8.Inverter_1.Vout.n8 GND 0.17757f
C5044 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t2 GND 0.06145f
C5045 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n0 GND 0.15815f
C5046 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n1 GND 0.12861f
C5047 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t5 GND 0.24486f
C5048 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t4 GND 0.47095f
C5049 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n2 GND 0.11174f
C5050 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n3 GND 0.11082f
C5051 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n4 GND 0.18808f
C5052 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n5 GND 0.14f
C5053 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t6 GND 0.47302f
C5054 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n6 GND 0.20386f
C5055 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t7 GND 0.23439f
C5056 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t1 GND 0.06388f
C5057 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n7 GND 0.40291f
C5058 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t0 GND 0.06521f
C5059 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.t3 GND 0.06388f
C5060 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n8 GND 0.36328f
C5061 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n9 GND 0.12591f
C5062 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.C.n10 GND 0.07837f
C5063 Nand_Gate_7.A.t2 GND 0.04841f
C5064 Nand_Gate_7.A.t8 GND 0.3437f
C5065 Nand_Gate_7.A.n0 GND 0.1004f
C5066 Nand_Gate_7.A.n1 GND 0.04356f
C5067 Nand_Gate_7.A.n2 GND 0.19155f
C5068 Nand_Gate_7.A.t7 GND 0.23519f
C5069 Nand_Gate_7.A.t11 GND 0.1787f
C5070 Nand_Gate_7.A.n3 GND 0.04681f
C5071 Nand_Gate_7.A.n4 GND 0.04294f
C5072 Nand_Gate_7.A.t6 GND 0.34417f
C5073 Nand_Gate_7.A.n5 GND 0.10324f
C5074 Nand_Gate_7.A.t4 GND 0.1787f
C5075 Nand_Gate_7.A.n6 GND 0.04681f
C5076 Nand_Gate_7.A.n7 GND 0.04294f
C5077 Nand_Gate_7.A.n8 GND 0.10864f
C5078 Nand_Gate_7.A.n9 GND 0.10864f
C5079 Nand_Gate_7.A.n10 GND 0.10324f
C5080 Nand_Gate_7.A.t10 GND 0.43948f
C5081 Nand_Gate_7.A.n11 GND 0.10779f
C5082 Nand_Gate_7.A.n12 GND 1.89329f
C5083 Nand_Gate_7.A.n13 GND 0.21834f
C5084 Nand_Gate_7.A.t9 GND 0.3437f
C5085 Nand_Gate_7.A.n14 GND 0.1497f
C5086 Nand_Gate_7.A.t5 GND 0.16042f
C5087 Nand_Gate_7.A.n15 GND 0.10472f
C5088 Nand_Gate_7.A.n16 GND 0.05015f
C5089 Nand_Gate_7.A.n17 GND 0.12716f
C5090 Nand_Gate_7.A.t3 GND 0.04662f
C5091 Nand_Gate_7.A.n18 GND 0.07181f
C5092 Nand_Gate_7.A.t1 GND 0.04759f
C5093 Nand_Gate_7.A.t0 GND 0.04662f
C5094 Nand_Gate_7.A.n19 GND 0.26512f
C5095 Nand_Gate_7.A.n20 GND 0.08651f
C5096 Nand_Gate_7.A.n21 GND 0.17418f
C5097 Ring_Counter_0.D_FlipFlop_11.Qbar.t2 GND 0.05347f
C5098 Ring_Counter_0.D_FlipFlop_11.Qbar.t4 GND 0.41161f
C5099 Ring_Counter_0.D_FlipFlop_11.Qbar.n0 GND 0.1774f
C5100 Ring_Counter_0.D_FlipFlop_11.Qbar.t5 GND 0.18986f
C5101 Ring_Counter_0.D_FlipFlop_11.Qbar.n1 GND 0.23199f
C5102 Ring_Counter_0.D_FlipFlop_11.Qbar.n2 GND 0.05991f
C5103 Ring_Counter_0.D_FlipFlop_11.Qbar.t1 GND 0.05559f
C5104 Ring_Counter_0.D_FlipFlop_11.Qbar.n3 GND 0.09627f
C5105 Ring_Counter_0.D_FlipFlop_11.Qbar.t0 GND 0.05675f
C5106 Ring_Counter_0.D_FlipFlop_11.Qbar.t3 GND 0.05559f
C5107 Ring_Counter_0.D_FlipFlop_11.Qbar.n4 GND 0.31612f
C5108 Ring_Counter_0.D_FlipFlop_11.Qbar.n5 GND 0.16106f
C5109 Ring_Counter_0.D_FlipFlop_11.Qbar.n6 GND 0.15403f
C5110 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 GND 0.06713f
C5111 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 GND 0.07989f
C5112 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 GND 0.43786f
C5113 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 GND 0.08018f
C5114 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 GND 0.25702f
C5115 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 GND 0.12462f
C5116 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 GND 0.4938f
C5117 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 GND 0.09136f
C5118 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 GND 0.05451f
C5119 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 GND 0.13379f
C5120 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 GND 0.13379f
C5121 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 GND 0.07316f
C5122 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 GND 0.06443f
C5123 Ring_Counter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 GND 0.14002f
C5124 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 GND 0.06443f
C5125 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 GND 0.14002f
C5126 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 GND 0.07316f
C5127 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 GND 0.25702f
C5128 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 GND 0.12462f
C5129 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 GND 0.4938f
C5130 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 GND 0.09136f
C5131 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 GND 0.05451f
C5132 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 GND 0.13379f
C5133 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 GND 0.13379f
C5134 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 GND 0.06713f
C5135 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 GND 0.07989f
C5136 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 GND 0.43786f
C5137 Ring_Counter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 GND 0.08018f
C5138 Nand_Gate_4.A.t2 GND 0.05206f
C5139 Nand_Gate_4.A.t7 GND 0.36961f
C5140 Nand_Gate_4.A.n0 GND 0.10797f
C5141 Nand_Gate_4.A.n1 GND 0.04685f
C5142 Nand_Gate_4.A.n2 GND 0.20599f
C5143 Nand_Gate_4.A.t6 GND 0.21736f
C5144 Nand_Gate_4.A.t10 GND 0.19217f
C5145 Nand_Gate_4.A.n3 GND 0.05034f
C5146 Nand_Gate_4.A.n4 GND 0.04617f
C5147 Nand_Gate_4.A.t9 GND 0.37011f
C5148 Nand_Gate_4.A.n5 GND 0.11103f
C5149 Nand_Gate_4.A.t5 GND 0.19217f
C5150 Nand_Gate_4.A.n6 GND 0.05034f
C5151 Nand_Gate_4.A.n7 GND 0.04617f
C5152 Nand_Gate_4.A.n8 GND 0.11683f
C5153 Nand_Gate_4.A.n9 GND 0.11683f
C5154 Nand_Gate_4.A.n10 GND 0.11103f
C5155 Nand_Gate_4.A.t11 GND 0.47261f
C5156 Nand_Gate_4.A.n11 GND 0.11592f
C5157 Nand_Gate_4.A.n12 GND 1.43638f
C5158 Nand_Gate_4.A.n13 GND 0.2348f
C5159 Nand_Gate_4.A.t8 GND 0.36961f
C5160 Nand_Gate_4.A.n14 GND 0.16099f
C5161 Nand_Gate_4.A.t4 GND 0.17251f
C5162 Nand_Gate_4.A.n15 GND 0.11261f
C5163 Nand_Gate_4.A.n16 GND 0.05393f
C5164 Nand_Gate_4.A.n17 GND 0.13674f
C5165 Nand_Gate_4.A.t1 GND 0.05013f
C5166 Nand_Gate_4.A.n18 GND 0.07723f
C5167 Nand_Gate_4.A.t3 GND 0.05118f
C5168 Nand_Gate_4.A.t0 GND 0.05013f
C5169 Nand_Gate_4.A.n19 GND 0.28511f
C5170 Nand_Gate_4.A.n20 GND 0.09303f
C5171 Nand_Gate_4.A.n21 GND 0.18731f
C5172 Ring_Counter_0.D_FlipFlop_5.Qbar.t5 GND 0.41161f
C5173 Ring_Counter_0.D_FlipFlop_5.Qbar.n0 GND 0.1774f
C5174 Ring_Counter_0.D_FlipFlop_5.Qbar.t4 GND 0.18986f
C5175 Ring_Counter_0.D_FlipFlop_5.Qbar.n1 GND 0.23199f
C5176 Ring_Counter_0.D_FlipFlop_5.Qbar.n2 GND 0.05991f
C5177 Ring_Counter_0.D_FlipFlop_5.Qbar.t2 GND 0.05559f
C5178 Ring_Counter_0.D_FlipFlop_5.Qbar.n3 GND 0.09627f
C5179 Ring_Counter_0.D_FlipFlop_5.Qbar.t3 GND 0.05675f
C5180 Ring_Counter_0.D_FlipFlop_5.Qbar.t1 GND 0.05559f
C5181 Ring_Counter_0.D_FlipFlop_5.Qbar.n4 GND 0.31612f
C5182 Ring_Counter_0.D_FlipFlop_5.Qbar.n5 GND 0.16106f
C5183 Ring_Counter_0.D_FlipFlop_5.Qbar.t0 GND 0.05347f
C5184 Ring_Counter_0.D_FlipFlop_5.Qbar.n6 GND 0.15403f
C5185 Nand_Gate_2.A.t1 GND 0.0374f
C5186 Nand_Gate_2.A.t11 GND 0.26554f
C5187 Nand_Gate_2.A.n0 GND 0.07757f
C5188 Nand_Gate_2.A.n1 GND 0.03366f
C5189 Nand_Gate_2.A.n2 GND 0.14799f
C5190 Nand_Gate_2.A.t10 GND 0.12312f
C5191 Nand_Gate_2.A.t8 GND 0.13806f
C5192 Nand_Gate_2.A.n3 GND 0.03617f
C5193 Nand_Gate_2.A.n4 GND 0.03317f
C5194 Nand_Gate_2.A.t5 GND 0.2659f
C5195 Nand_Gate_2.A.n5 GND 0.07976f
C5196 Nand_Gate_2.A.t4 GND 0.13806f
C5197 Nand_Gate_2.A.n6 GND 0.03617f
C5198 Nand_Gate_2.A.n7 GND 0.03317f
C5199 Nand_Gate_2.A.n8 GND 0.08394f
C5200 Nand_Gate_2.A.n9 GND 0.08394f
C5201 Nand_Gate_2.A.n10 GND 0.07976f
C5202 Nand_Gate_2.A.t7 GND 0.33953f
C5203 Nand_Gate_2.A.n11 GND 0.09029f
C5204 Nand_Gate_2.A.n12 GND 0.33595f
C5205 Nand_Gate_2.A.n13 GND 0.16168f
C5206 Nand_Gate_2.A.t6 GND 0.26554f
C5207 Nand_Gate_2.A.n14 GND 0.11566f
C5208 Nand_Gate_2.A.t9 GND 0.12394f
C5209 Nand_Gate_2.A.n15 GND 0.0809f
C5210 Nand_Gate_2.A.n16 GND 0.03875f
C5211 Nand_Gate_2.A.n17 GND 0.09824f
C5212 Nand_Gate_2.A.t2 GND 0.03602f
C5213 Nand_Gate_2.A.n18 GND 0.05548f
C5214 Nand_Gate_2.A.t3 GND 0.03677f
C5215 Nand_Gate_2.A.t0 GND 0.03602f
C5216 Nand_Gate_2.A.n19 GND 0.20483f
C5217 Nand_Gate_2.A.n20 GND 0.06684f
C5218 Nand_Gate_2.A.n21 GND 0.13457f
C5219 CDAC_v3_0.switch_2.Z.t6 GND 0.08313f
C5220 CDAC_v3_0.switch_2.Z.t1 GND 0.08296f
C5221 CDAC_v3_0.switch_2.Z.n0 GND 0.18251f
C5222 CDAC_v3_0.switch_2.Z.n1 GND 0.02824f
C5223 CDAC_v3_0.switch_2.Z.t3 GND 11.2597f
C5224 CDAC_v3_0.switch_2.Z.t5 GND 11.2597f
C5225 CDAC_v3_0.switch_2.Z.t2 GND 12.1819f
C5226 CDAC_v3_0.switch_2.Z.n2 GND 5.82928f
C5227 CDAC_v3_0.switch_2.Z.t4 GND 11.5599f
C5228 CDAC_v3_0.switch_2.Z.n3 GND 4.98503f
C5229 CDAC_v3_0.switch_2.Z.n4 GND 8.7732f
C5230 CDAC_v3_0.switch_2.Z.n5 GND 5.96162f
C5231 CDAC_v3_0.switch_2.Z.n6 GND 0.08892f
C5232 CDAC_v3_0.switch_2.Z.t7 GND 0.08582f
C5233 CDAC_v3_0.switch_2.Z.t0 GND 0.08582f
C5234 CDAC_v3_0.switch_2.Z.n7 GND 0.30824f
C5235 CDAC_v3_0.switch_2.Z.n8 GND 0.95036f
C5236 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 GND 0.06443f
C5237 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 GND 0.14002f
C5238 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 GND 0.07316f
C5239 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 GND 0.25702f
C5240 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 GND 0.12462f
C5241 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 GND 0.4938f
C5242 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 GND 0.09136f
C5243 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 GND 0.05451f
C5244 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 GND 0.13379f
C5245 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 GND 0.13379f
C5246 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 GND 0.06713f
C5247 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 GND 0.07989f
C5248 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 GND 0.43786f
C5249 Ring_Counter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 GND 0.08018f
C5250 CDAC_v3_0.switch_0.Z.t1 GND 0.08228f
C5251 CDAC_v3_0.switch_0.Z.t4 GND 0.08228f
C5252 CDAC_v3_0.switch_0.Z.n0 GND 0.29554f
C5253 CDAC_v3_0.switch_0.Z.n1 GND 0.9112f
C5254 CDAC_v3_0.switch_0.Z.n2 GND 0.08525f
C5255 CDAC_v3_0.switch_0.Z.t2 GND 10.7957f
C5256 CDAC_v3_0.switch_0.Z.t3 GND 10.9185f
C5257 CDAC_v3_0.switch_0.Z.n3 GND 15.6517f
C5258 CDAC_v3_0.switch_0.Z.n4 GND 9.79336f
C5259 CDAC_v3_0.switch_0.Z.n5 GND 0.02708f
C5260 CDAC_v3_0.switch_0.Z.t0 GND 0.0797f
C5261 CDAC_v3_0.switch_0.Z.n6 GND 0.17499f
C5262 CDAC_v3_0.switch_0.Z.t5 GND 0.07954f
C5263 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 GND 0.37675f
C5264 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 GND 0.16409f
C5265 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 GND 0.18888f
C5266 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 GND 0.0511f
C5267 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 GND 0.32168f
C5268 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 GND 0.05217f
C5269 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 GND 0.0511f
C5270 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 GND 0.29061f
C5271 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 GND 0.09483f
C5272 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 GND 0.01203f
C5273 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 GND 0.01587f
C5274 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 GND 0.37825f
C5275 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 GND 0.19588f
C5276 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 GND 0.28346f
C5277 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 GND 0.11199f
C5278 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 GND 0.05215f
C5279 Ring_Counter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 GND 0.18008f
C5280 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 GND 0.05215f
C5281 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 GND 0.18008f
C5282 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 GND 0.37825f
C5283 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 GND 0.19588f
C5284 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 GND 0.28346f
C5285 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 GND 0.11199f
C5286 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 GND 0.01587f
C5287 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 GND 0.37675f
C5288 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 GND 0.16409f
C5289 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 GND 0.18888f
C5290 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 GND 0.0511f
C5291 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 GND 0.32168f
C5292 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 GND 0.05217f
C5293 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 GND 0.0511f
C5294 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 GND 0.29061f
C5295 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 GND 0.09483f
C5296 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 GND 0.01203f
C5297 D_FlipFlop_6.3-input-nand_2.Vout.t7 GND 0.34247f
C5298 D_FlipFlop_6.3-input-nand_2.Vout.n0 GND 0.10005f
C5299 D_FlipFlop_6.3-input-nand_2.Vout.n1 GND 0.04341f
C5300 D_FlipFlop_6.3-input-nand_2.Vout.t1 GND 0.04467f
C5301 D_FlipFlop_6.3-input-nand_2.Vout.n2 GND 0.21241f
C5302 D_FlipFlop_6.3-input-nand_2.Vout.n3 GND 0.04823f
C5303 D_FlipFlop_6.3-input-nand_2.Vout.t6 GND 0.34248f
C5304 D_FlipFlop_6.3-input-nand_2.Vout.n4 GND 0.35447f
C5305 D_FlipFlop_6.3-input-nand_2.Vout.t4 GND 0.17806f
C5306 D_FlipFlop_6.3-input-nand_2.Vout.n5 GND 0.17459f
C5307 D_FlipFlop_6.3-input-nand_2.Vout.n6 GND 0.1018f
C5308 D_FlipFlop_6.3-input-nand_2.Vout.n7 GND 0.01283f
C5309 D_FlipFlop_6.3-input-nand_2.Vout.n8 GND 0.01019f
C5310 D_FlipFlop_6.3-input-nand_2.Vout.t3 GND 0.04742f
C5311 D_FlipFlop_6.3-input-nand_2.Vout.t0 GND 0.04645f
C5312 D_FlipFlop_6.3-input-nand_2.Vout.n9 GND 0.26417f
C5313 D_FlipFlop_6.3-input-nand_2.Vout.n10 GND 0.0862f
C5314 D_FlipFlop_6.3-input-nand_2.Vout.t2 GND 0.04645f
C5315 D_FlipFlop_6.3-input-nand_2.Vout.n11 GND 0.29241f
C5316 D_FlipFlop_6.3-input-nand_2.Vout.t5 GND 0.17113f
C5317 D_FlipFlop_6.3-input-nand_2.Vout.n12 GND 0.19086f
C5318 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 GND 0.06443f
C5319 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 GND 0.14002f
C5320 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 GND 0.07316f
C5321 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 GND 0.25702f
C5322 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 GND 0.12462f
C5323 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 GND 0.4938f
C5324 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 GND 0.09136f
C5325 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 GND 0.05451f
C5326 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 GND 0.13379f
C5327 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 GND 0.13379f
C5328 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 GND 0.06713f
C5329 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 GND 0.07989f
C5330 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 GND 0.43786f
C5331 Ring_Counter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 GND 0.08018f
C5332 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t1 GND 0.05f
C5333 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n0 GND 0.10867f
C5334 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n1 GND 0.05678f
C5335 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t5 GND 0.38491f
C5336 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n2 GND 0.16589f
C5337 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t3 GND 0.30131f
C5338 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t4 GND 0.30153f
C5339 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n3 GND 0.09671f
C5340 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t2 GND 0.38323f
C5341 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n4 GND 0.0709f
C5342 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n5 GND 0.04231f
C5343 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n6 GND 0.10383f
C5344 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n7 GND 0.10383f
C5345 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.t0 GND 0.05284f
C5346 Ring_Counter_0.D_FlipFlop_13.Inverter_1.Vout.n8 GND 0.17757f
C5347 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t1 GND 0.06145f
C5348 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n0 GND 0.15815f
C5349 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n1 GND 0.12861f
C5350 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t7 GND 0.24486f
C5351 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t4 GND 0.47095f
C5352 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n2 GND 0.11174f
C5353 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n3 GND 0.11082f
C5354 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n4 GND 0.18808f
C5355 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n5 GND 0.14f
C5356 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t6 GND 0.47302f
C5357 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n6 GND 0.20386f
C5358 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t5 GND 0.23439f
C5359 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t2 GND 0.06388f
C5360 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n7 GND 0.40291f
C5361 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t0 GND 0.06521f
C5362 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.t3 GND 0.06388f
C5363 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n8 GND 0.36328f
C5364 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n9 GND 0.12591f
C5365 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.C.n10 GND 0.07837f
C5366 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 GND 0.05215f
C5367 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 GND 0.18008f
C5368 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 GND 0.37825f
C5369 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 GND 0.19588f
C5370 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 GND 0.28346f
C5371 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 GND 0.11199f
C5372 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 GND 0.01587f
C5373 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 GND 0.37675f
C5374 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 GND 0.16409f
C5375 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 GND 0.18888f
C5376 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 GND 0.0511f
C5377 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 GND 0.32168f
C5378 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 GND 0.05217f
C5379 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 GND 0.0511f
C5380 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 GND 0.29061f
C5381 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 GND 0.09483f
C5382 Ring_Counter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 GND 0.01203f
C5383 D_FlipFlop_4.3-input-nand_2.Vout.t6 GND 0.34247f
C5384 D_FlipFlop_4.3-input-nand_2.Vout.n0 GND 0.10005f
C5385 D_FlipFlop_4.3-input-nand_2.Vout.n1 GND 0.04341f
C5386 D_FlipFlop_4.3-input-nand_2.Vout.t1 GND 0.04467f
C5387 D_FlipFlop_4.3-input-nand_2.Vout.n2 GND 0.21241f
C5388 D_FlipFlop_4.3-input-nand_2.Vout.n3 GND 0.04823f
C5389 D_FlipFlop_4.3-input-nand_2.Vout.t5 GND 0.34248f
C5390 D_FlipFlop_4.3-input-nand_2.Vout.n4 GND 0.35447f
C5391 D_FlipFlop_4.3-input-nand_2.Vout.t7 GND 0.17806f
C5392 D_FlipFlop_4.3-input-nand_2.Vout.n5 GND 0.17459f
C5393 D_FlipFlop_4.3-input-nand_2.Vout.n6 GND 0.1018f
C5394 D_FlipFlop_4.3-input-nand_2.Vout.n7 GND 0.01283f
C5395 D_FlipFlop_4.3-input-nand_2.Vout.n8 GND 0.01019f
C5396 D_FlipFlop_4.3-input-nand_2.Vout.t2 GND 0.04742f
C5397 D_FlipFlop_4.3-input-nand_2.Vout.t3 GND 0.04645f
C5398 D_FlipFlop_4.3-input-nand_2.Vout.n9 GND 0.26417f
C5399 D_FlipFlop_4.3-input-nand_2.Vout.n10 GND 0.0862f
C5400 D_FlipFlop_4.3-input-nand_2.Vout.t0 GND 0.04645f
C5401 D_FlipFlop_4.3-input-nand_2.Vout.n11 GND 0.29241f
C5402 D_FlipFlop_4.3-input-nand_2.Vout.t4 GND 0.17113f
C5403 D_FlipFlop_4.3-input-nand_2.Vout.n12 GND 0.19086f
C5404 D_FlipFlop_4.3-input-nand_2.C.t1 GND 0.04469f
C5405 D_FlipFlop_4.3-input-nand_2.C.n0 GND 0.04327f
C5406 D_FlipFlop_4.3-input-nand_2.C.n1 GND 0.09193f
C5407 D_FlipFlop_4.3-input-nand_2.C.t5 GND 0.17806f
C5408 D_FlipFlop_4.3-input-nand_2.C.t7 GND 0.34248f
C5409 D_FlipFlop_4.3-input-nand_2.C.n2 GND 0.10005f
C5410 D_FlipFlop_4.3-input-nand_2.C.n3 GND 0.04279f
C5411 D_FlipFlop_4.3-input-nand_2.C.n4 GND 0.079f
C5412 D_FlipFlop_4.3-input-nand_2.C.n5 GND 0.13677f
C5413 D_FlipFlop_4.3-input-nand_2.C.n6 GND 0.10181f
C5414 D_FlipFlop_4.3-input-nand_2.C.n7 GND 0.04823f
C5415 D_FlipFlop_4.3-input-nand_2.C.t6 GND 0.3425f
C5416 D_FlipFlop_4.3-input-nand_2.C.n8 GND 0.3551f
C5417 D_FlipFlop_4.3-input-nand_2.C.n9 GND 0.03842f
C5418 D_FlipFlop_4.3-input-nand_2.C.n10 GND 0.05129f
C5419 D_FlipFlop_4.3-input-nand_2.C.t4 GND 0.17045f
C5420 D_FlipFlop_4.3-input-nand_2.C.t0 GND 0.04645f
C5421 D_FlipFlop_4.3-input-nand_2.C.n11 GND 0.293f
C5422 D_FlipFlop_4.3-input-nand_2.C.t3 GND 0.04742f
C5423 D_FlipFlop_4.3-input-nand_2.C.t2 GND 0.04645f
C5424 D_FlipFlop_4.3-input-nand_2.C.n12 GND 0.26418f
C5425 D_FlipFlop_4.3-input-nand_2.C.n13 GND 0.08722f
C5426 D_FlipFlop_4.3-input-nand_2.C.n14 GND 0.124f
C5427 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 GND 0.07411f
C5428 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 GND 0.16107f
C5429 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 GND 0.08416f
C5430 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 GND 0.29566f
C5431 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 GND 0.14335f
C5432 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 GND 0.56804f
C5433 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 GND 0.1051f
C5434 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 GND 0.06271f
C5435 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 GND 0.15391f
C5436 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 GND 0.15391f
C5437 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 GND 0.07722f
C5438 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 GND 0.07866f
C5439 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 GND 0.07705f
C5440 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 GND 0.43817f
C5441 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 GND 0.286f
C5442 Ring_Counter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 GND 0.09223f
C5443 Q1.t8 GND 0.19299f
C5444 Q1.t6 GND 0.37263f
C5445 Q1.n0 GND 0.27664f
C5446 Q1.n1 GND 0.05119f
C5447 Q1.t9 GND 0.19299f
C5448 Q1.t4 GND 0.37263f
C5449 Q1.n2 GND 0.27491f
C5450 Q1.n3 GND 0.05514f
C5451 Q1.n4 GND 0.08945f
C5452 Q1.n5 GND 1.85817f
C5453 Q1.t1 GND 0.04838f
C5454 Q1.n6 GND 0.23728f
C5455 Q1.n7 GND 0.05408f
C5456 Q1.t2 GND 0.05137f
C5457 Q1.t3 GND 0.05031f
C5458 Q1.n8 GND 0.28614f
C5459 Q1.n9 GND 0.09337f
C5460 Q1.t0 GND 0.05031f
C5461 Q1.n10 GND 0.0775f
C5462 Q1.n11 GND 0.13724f
C5463 Q1.n12 GND 0.05413f
C5464 Q1.t7 GND 0.37094f
C5465 Q1.n13 GND 0.10836f
C5466 Q1.n14 GND 0.04702f
C5467 Q1.n15 GND 0.20673f
C5468 Q1.t5 GND 0.17252f
C5469 Q1.n16 GND 0.50673f
C5470 Q1.n17 GND 0.80118f
C5471 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 GND 0.05215f
C5472 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 GND 0.18008f
C5473 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 GND 0.37825f
C5474 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 GND 0.19588f
C5475 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 GND 0.28346f
C5476 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 GND 0.11199f
C5477 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 GND 0.01587f
C5478 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 GND 0.37675f
C5479 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 GND 0.16409f
C5480 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 GND 0.18888f
C5481 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 GND 0.0511f
C5482 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 GND 0.32168f
C5483 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 GND 0.05217f
C5484 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 GND 0.0511f
C5485 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 GND 0.29061f
C5486 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 GND 0.09483f
C5487 Ring_Counter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 GND 0.01203f
C5488 Ring_Counter_0.D_FlipFlop_8.Qbar.t2 GND 0.05347f
C5489 Ring_Counter_0.D_FlipFlop_8.Qbar.t4 GND 0.41161f
C5490 Ring_Counter_0.D_FlipFlop_8.Qbar.n0 GND 0.1774f
C5491 Ring_Counter_0.D_FlipFlop_8.Qbar.t5 GND 0.18986f
C5492 Ring_Counter_0.D_FlipFlop_8.Qbar.n1 GND 0.23199f
C5493 Ring_Counter_0.D_FlipFlop_8.Qbar.n2 GND 0.05991f
C5494 Ring_Counter_0.D_FlipFlop_8.Qbar.t1 GND 0.05559f
C5495 Ring_Counter_0.D_FlipFlop_8.Qbar.n3 GND 0.09627f
C5496 Ring_Counter_0.D_FlipFlop_8.Qbar.t0 GND 0.05675f
C5497 Ring_Counter_0.D_FlipFlop_8.Qbar.t3 GND 0.05559f
C5498 Ring_Counter_0.D_FlipFlop_8.Qbar.n4 GND 0.31612f
C5499 Ring_Counter_0.D_FlipFlop_8.Qbar.n5 GND 0.16106f
C5500 Ring_Counter_0.D_FlipFlop_8.Qbar.n6 GND 0.15403f
C5501 D_FlipFlop_5.nPRE.t13 GND 0.23587f
C5502 D_FlipFlop_5.nPRE.n0 GND 0.0689f
C5503 D_FlipFlop_5.nPRE.n1 GND 0.0299f
C5504 D_FlipFlop_5.nPRE.n2 GND 0.13145f
C5505 D_FlipFlop_5.nPRE.t10 GND 0.1097f
C5506 D_FlipFlop_5.nPRE.n3 GND 0.06295f
C5507 D_FlipFlop_5.nPRE.n4 GND 0.13342f
C5508 D_FlipFlop_5.nPRE.t14 GND 0.23588f
C5509 D_FlipFlop_5.nPRE.n5 GND 0.23754f
C5510 D_FlipFlop_5.nPRE.n6 GND 0.02534f
C5511 D_FlipFlop_5.nPRE.t6 GND 0.12263f
C5512 D_FlipFlop_5.nPRE.n7 GND 0.03533f
C5513 D_FlipFlop_5.nPRE.n9 GND 0.01466f
C5514 D_FlipFlop_5.nPRE.n10 GND 0.14628f
C5515 D_FlipFlop_5.nPRE.t7 GND 0.23588f
C5516 D_FlipFlop_5.nPRE.n11 GND 0.23754f
C5517 D_FlipFlop_5.nPRE.n12 GND 0.02534f
C5518 D_FlipFlop_5.nPRE.t12 GND 0.12263f
C5519 D_FlipFlop_5.nPRE.n13 GND 0.03533f
C5520 D_FlipFlop_5.nPRE.n15 GND 0.01466f
C5521 D_FlipFlop_5.nPRE.n17 GND 0.37966f
C5522 D_FlipFlop_5.nPRE.n18 GND 0.48265f
C5523 D_FlipFlop_5.nPRE.t5 GND 0.23587f
C5524 D_FlipFlop_5.nPRE.n19 GND 0.0689f
C5525 D_FlipFlop_5.nPRE.n20 GND 0.0299f
C5526 D_FlipFlop_5.nPRE.n21 GND 0.13145f
C5527 D_FlipFlop_5.nPRE.t15 GND 0.11092f
C5528 D_FlipFlop_5.nPRE.n22 GND 0.84704f
C5529 D_FlipFlop_5.nPRE.t11 GND 0.12263f
C5530 D_FlipFlop_5.nPRE.n23 GND 0.03213f
C5531 D_FlipFlop_5.nPRE.n24 GND 0.02947f
C5532 D_FlipFlop_5.nPRE.t8 GND 0.23619f
C5533 D_FlipFlop_5.nPRE.n25 GND 0.07085f
C5534 D_FlipFlop_5.nPRE.t16 GND 0.12263f
C5535 D_FlipFlop_5.nPRE.n26 GND 0.03213f
C5536 D_FlipFlop_5.nPRE.n27 GND 0.02947f
C5537 D_FlipFlop_5.nPRE.n28 GND 0.07456f
C5538 D_FlipFlop_5.nPRE.n29 GND 0.07456f
C5539 D_FlipFlop_5.nPRE.n30 GND 0.07085f
C5540 D_FlipFlop_5.nPRE.t17 GND 0.3016f
C5541 D_FlipFlop_5.nPRE.n31 GND 0.07397f
C5542 D_FlipFlop_5.nPRE.n32 GND 0.257f
C5543 D_FlipFlop_5.nPRE.n33 GND 0.14984f
C5544 D_FlipFlop_5.nPRE.t9 GND 0.23587f
C5545 D_FlipFlop_5.nPRE.n34 GND 0.10273f
C5546 D_FlipFlop_5.nPRE.t4 GND 0.11009f
C5547 D_FlipFlop_5.nPRE.n35 GND 0.07186f
C5548 D_FlipFlop_5.nPRE.n36 GND 0.03442f
C5549 D_FlipFlop_5.nPRE.n37 GND 0.08726f
C5550 D_FlipFlop_5.nPRE.t1 GND 0.03199f
C5551 D_FlipFlop_5.nPRE.n38 GND 0.04928f
C5552 D_FlipFlop_5.nPRE.t2 GND 0.03266f
C5553 D_FlipFlop_5.nPRE.t3 GND 0.03199f
C5554 D_FlipFlop_5.nPRE.n39 GND 0.18194f
C5555 D_FlipFlop_5.nPRE.n40 GND 0.05937f
C5556 D_FlipFlop_5.nPRE.t0 GND 0.03322f
C5557 D_FlipFlop_5.nPRE.n41 GND 0.11953f
C5558 D_FlipFlop_1.CLK.t1 GND 0.02954f
C5559 D_FlipFlop_1.CLK.t6 GND 0.22695f
C5560 D_FlipFlop_1.CLK.t5 GND 0.118f
C5561 D_FlipFlop_1.CLK.n0 GND 0.12444f
C5562 D_FlipFlop_1.CLK.t7 GND 0.22695f
C5563 D_FlipFlop_1.CLK.n1 GND 0.2009f
C5564 D_FlipFlop_1.CLK.n2 GND 0.20145f
C5565 D_FlipFlop_1.CLK.n3 GND 0.12607f
C5566 D_FlipFlop_1.CLK.t3 GND 0.10447f
C5567 D_FlipFlop_1.CLK.n4 GND 0.02736f
C5568 D_FlipFlop_1.CLK.n5 GND 0.10371f
C5569 D_FlipFlop_1.CLK.t2 GND 0.10446f
C5570 D_FlipFlop_1.CLK.n6 GND 0.03399f
C5571 D_FlipFlop_1.CLK.n7 GND 0.02546f
C5572 D_FlipFlop_1.CLK.n8 GND 0.23531f
C5573 D_FlipFlop_1.CLK.t4 GND 0.21911f
C5574 D_FlipFlop_1.CLK.n9 GND 0.16025f
C5575 D_FlipFlop_1.CLK.n11 GND 0.03049f
C5576 D_FlipFlop_1.CLK.t0 GND 0.03086f
C5577 D_FlipFlop_1.CLK.n12 GND 0.19695f
C5578 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 GND 0.06393f
C5579 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 GND 0.07609f
C5580 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 GND 0.41701f
C5581 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 GND 0.07636f
C5582 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 GND 0.24478f
C5583 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 GND 0.11868f
C5584 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 GND 0.47029f
C5585 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 GND 0.08701f
C5586 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 GND 0.05192f
C5587 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 GND 0.12742f
C5588 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 GND 0.12742f
C5589 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 GND 0.06968f
C5590 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 GND 0.06136f
C5591 Ring_Counter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 GND 0.13336f
C5592 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t1 GND 0.05f
C5593 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n0 GND 0.10867f
C5594 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n1 GND 0.05678f
C5595 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t4 GND 0.38491f
C5596 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n2 GND 0.16589f
C5597 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t2 GND 0.30131f
C5598 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t3 GND 0.30153f
C5599 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n3 GND 0.09671f
C5600 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t5 GND 0.38323f
C5601 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n4 GND 0.0709f
C5602 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n5 GND 0.04231f
C5603 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n6 GND 0.10383f
C5604 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n7 GND 0.10383f
C5605 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.t0 GND 0.05284f
C5606 Ring_Counter_0.D_FlipFlop_10.Inverter_1.Vout.n8 GND 0.17757f
C5607 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t3 GND 0.06145f
C5608 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n0 GND 0.15815f
C5609 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n1 GND 0.12861f
C5610 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t5 GND 0.24486f
C5611 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t4 GND 0.47095f
C5612 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n2 GND 0.11174f
C5613 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n3 GND 0.11082f
C5614 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n4 GND 0.18808f
C5615 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n5 GND 0.14f
C5616 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t7 GND 0.47302f
C5617 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n6 GND 0.20386f
C5618 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t6 GND 0.23439f
C5619 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t2 GND 0.06388f
C5620 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n7 GND 0.40291f
C5621 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t0 GND 0.06521f
C5622 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.t1 GND 0.06388f
C5623 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n8 GND 0.36328f
C5624 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n9 GND 0.12591f
C5625 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.C.n10 GND 0.07837f
C5626 Ring_Counter_0.D_FlipFlop_14.Qbar.t2 GND 0.05347f
C5627 Ring_Counter_0.D_FlipFlop_14.Qbar.t5 GND 0.41161f
C5628 Ring_Counter_0.D_FlipFlop_14.Qbar.n0 GND 0.1774f
C5629 Ring_Counter_0.D_FlipFlop_14.Qbar.t4 GND 0.18986f
C5630 Ring_Counter_0.D_FlipFlop_14.Qbar.n1 GND 0.23199f
C5631 Ring_Counter_0.D_FlipFlop_14.Qbar.n2 GND 0.05991f
C5632 Ring_Counter_0.D_FlipFlop_14.Qbar.t1 GND 0.05559f
C5633 Ring_Counter_0.D_FlipFlop_14.Qbar.n3 GND 0.09627f
C5634 Ring_Counter_0.D_FlipFlop_14.Qbar.t0 GND 0.05675f
C5635 Ring_Counter_0.D_FlipFlop_14.Qbar.t3 GND 0.05559f
C5636 Ring_Counter_0.D_FlipFlop_14.Qbar.n4 GND 0.31612f
C5637 Ring_Counter_0.D_FlipFlop_14.Qbar.n5 GND 0.16106f
C5638 Ring_Counter_0.D_FlipFlop_14.Qbar.n6 GND 0.15403f
C5639 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 GND 0.06443f
C5640 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 GND 0.14002f
C5641 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 GND 0.07316f
C5642 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 GND 0.25702f
C5643 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 GND 0.12462f
C5644 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 GND 0.4938f
C5645 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 GND 0.09136f
C5646 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 GND 0.05451f
C5647 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 GND 0.13379f
C5648 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 GND 0.13379f
C5649 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 GND 0.06713f
C5650 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 GND 0.07989f
C5651 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 GND 0.43786f
C5652 Ring_Counter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 GND 0.08018f
C5653 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t1 GND 0.05f
C5654 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n0 GND 0.10867f
C5655 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n1 GND 0.05678f
C5656 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t5 GND 0.38491f
C5657 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n2 GND 0.16589f
C5658 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t3 GND 0.30131f
C5659 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t4 GND 0.30153f
C5660 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n3 GND 0.09671f
C5661 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t2 GND 0.38323f
C5662 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n4 GND 0.0709f
C5663 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n5 GND 0.04231f
C5664 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n6 GND 0.10383f
C5665 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n7 GND 0.10383f
C5666 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.t0 GND 0.05284f
C5667 Ring_Counter_0.D_FlipFlop_2.Inverter_1.Vout.n8 GND 0.17757f
C5668 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t1 GND 0.05f
C5669 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n0 GND 0.10867f
C5670 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n1 GND 0.05678f
C5671 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t2 GND 0.38491f
C5672 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n2 GND 0.16589f
C5673 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t3 GND 0.30131f
C5674 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t4 GND 0.30153f
C5675 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n3 GND 0.09671f
C5676 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t5 GND 0.38323f
C5677 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n4 GND 0.0709f
C5678 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n5 GND 0.04231f
C5679 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n6 GND 0.10383f
C5680 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n7 GND 0.10383f
C5681 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.t0 GND 0.05284f
C5682 Ring_Counter_0.D_FlipFlop_9.Inverter_1.Vout.n8 GND 0.17757f
C5683 Vbias.n0 GND 0.01479f
C5684 Vbias.n1 GND 0.13893f
C5685 Vbias.n2 GND 0.25311f
C5686 Vbias.n3 GND 0.14762f
C5687 Vbias.n4 GND 0.25311f
C5688 Vbias.t0 GND 6.30217f
C5689 Vbias.n5 GND 0.33942f
C5690 Vbias.n6 GND 0.33942f
C5691 Vbias.n7 GND 0.1981f
C5692 Vbias.t5 GND 2.77483f
C5693 Vbias.n8 GND 0.42554f
C5694 Vbias.n9 GND 0.42554f
C5695 Vbias.n10 GND 0.24851f
C5696 Vbias.n11 GND 0.23241f
C5697 Vbias.n12 GND 0.20147f
C5698 Vbias.n13 GND 1.60658f
C5699 Vbias.n14 GND 1.63343f
C5700 Vbias.n15 GND 1.63343f
C5701 Vbias.n16 GND 38.8269f
C5702 Vbias.n17 GND 22.6984f
C5703 Vbias.t4 GND 16.0295f
C5704 Vbias.n19 GND 53.2088f
C5705 Vbias.t2 GND 6.30217f
C5706 Vbias.n20 GND 0.42554f
C5707 Vbias.n21 GND 0.42554f
C5708 Vbias.n22 GND 6.18459f
C5709 Vbias.n23 GND 0.41774f
C5710 Vbias.n24 GND 6.18459f
C5711 Vbias.n25 GND 0.33942f
C5712 Vbias.n26 GND 0.33218f
C5713 Vbias.n27 GND 6.18459f
C5714 Vbias.n28 GND 0.33218f
C5715 Vbias.n29 GND 0.1956f
C5716 Vbias.n30 GND 0.1981f
C5717 Vbias.n31 GND 0.1956f
C5718 Vbias.n32 GND 0.1981f
C5719 Vbias.n33 GND 0.33942f
C5720 Vbias.t9 GND 2.77483f
C5721 Vbias.n34 GND 6.18459f
C5722 Vbias.n35 GND 0.41774f
C5723 Vbias.n36 GND 0.23241f
C5724 Vbias.n37 GND 0.24851f
C5725 Vbias.n38 GND 0.29298f
C5726 Vbias.n39 GND 0.23882f
C5727 Vbias.n40 GND 0.41774f
C5728 Vbias.n41 GND 31.3933f
C5729 Vbias.n42 GND 41.0582f
C5730 Vbias.n43 GND 1.6303f
C5731 Vbias.n44 GND 1.60658f
C5732 Vbias.n45 GND 2.44638f
C5733 Vbias.n46 GND 0.17898f
C5734 Vbias.t3 GND 1.28685f
C5735 Vbias.t8 GND 0.55493f
C5736 Vbias.t1 GND 4.61738f
C5737 Vbias.n47 GND 1.06251f
C5738 Vbias.n48 GND 0.39372f
C5739 Vbias.t6 GND 1.27472f
C5740 Vbias.n49 GND 0.43846f
C5741 Vbias.n50 GND 0.48485f
C5742 Vbias.n51 GND 0.13953f
C5743 Vbias.n52 GND 0.26027f
C5744 Vbias.n53 GND 0.04006f
C5745 Vbias.n54 GND 0.0337f
C5746 Vbias.n55 GND 0.20147f
C5747 Vbias.n56 GND 0.29298f
C5748 Vbias.n57 GND 0.23882f
C5749 Vbias.n58 GND 0.41774f
C5750 Vbias.n59 GND 6.18459f
C5751 Vbias.n60 GND 6.18459f
C5752 Vbias.n61 GND 0.33218f
C5753 Vbias.n62 GND 0.1956f
C5754 Vbias.n63 GND 0.1981f
C5755 Vbias.n64 GND 0.1956f
C5756 Vbias.n65 GND 0.33218f
C5757 Vbias.n66 GND 20.1293f
C5758 Vbias.n67 GND 0.24682f
C5759 Vbias.n68 GND 20.1293f
C5760 Vbias.t7 GND 19.8588f
C5761 Vbias.n70 GND 31.017f
C5762 Vbias.n71 GND 0.13893f
C5763 Vbias.n72 GND 0.33383f
C5764 Vbias.n73 GND 0.06481f
C5765 Vbias.n74 GND 0.13569f
C5766 a_51773_21431.t2 GND 1.19983f
C5767 a_51773_21431.t1 GND 2.30305f
C5768 a_51773_21431.n0 GND 2.49728f
C5769 a_51773_21431.t0 GND 1.19983f
C5770 a_50502_29172.t1 GND 2.8982f
C5771 a_50502_29172.t3 GND 2.72029f
C5772 a_50502_29172.t2 GND 4.52607f
C5773 a_50502_29172.n0 GND 1.99489f
C5774 a_50502_29172.n1 GND 1.6646f
C5775 a_50502_29172.t0 GND 0.89595f
C5776 Nand_Gate_0.A.t1 GND 0.0354f
C5777 Nand_Gate_0.A.t8 GND 0.25136f
C5778 Nand_Gate_0.A.n0 GND 0.07343f
C5779 Nand_Gate_0.A.n1 GND 0.03186f
C5780 Nand_Gate_0.A.n2 GND 0.14008f
C5781 Nand_Gate_0.A.t7 GND 0.12766f
C5782 Nand_Gate_0.A.t6 GND 0.13069f
C5783 Nand_Gate_0.A.n3 GND 0.03424f
C5784 Nand_Gate_0.A.n4 GND 0.0314f
C5785 Nand_Gate_0.A.t11 GND 0.2517f
C5786 Nand_Gate_0.A.n5 GND 0.0755f
C5787 Nand_Gate_0.A.t9 GND 0.13069f
C5788 Nand_Gate_0.A.n6 GND 0.03424f
C5789 Nand_Gate_0.A.n7 GND 0.0314f
C5790 Nand_Gate_0.A.n8 GND 0.07945f
C5791 Nand_Gate_0.A.n9 GND 0.07945f
C5792 Nand_Gate_0.A.n10 GND 0.0755f
C5793 Nand_Gate_0.A.t4 GND 0.3214f
C5794 Nand_Gate_0.A.n11 GND 0.07883f
C5795 Nand_Gate_0.A.n12 GND 0.53654f
C5796 Nand_Gate_0.A.n13 GND 0.15968f
C5797 Nand_Gate_0.A.t10 GND 0.25136f
C5798 Nand_Gate_0.A.n14 GND 0.10948f
C5799 Nand_Gate_0.A.t5 GND 0.11732f
C5800 Nand_Gate_0.A.n15 GND 0.07658f
C5801 Nand_Gate_0.A.n16 GND 0.03668f
C5802 Nand_Gate_0.A.n17 GND 0.09299f
C5803 Nand_Gate_0.A.t0 GND 0.03409f
C5804 Nand_Gate_0.A.n18 GND 0.05252f
C5805 Nand_Gate_0.A.t2 GND 0.03481f
C5806 Nand_Gate_0.A.t3 GND 0.03409f
C5807 Nand_Gate_0.A.n19 GND 0.19389f
C5808 Nand_Gate_0.A.n20 GND 0.06327f
C5809 Nand_Gate_0.A.n21 GND 0.12738f
C5810 D_FlipFlop_0.3-input-nand_2.C.t7 GND 0.3425f
C5811 D_FlipFlop_0.3-input-nand_2.C.n0 GND 0.3551f
C5812 D_FlipFlop_0.3-input-nand_2.C.n1 GND 0.03842f
C5813 D_FlipFlop_0.3-input-nand_2.C.t3 GND 0.04469f
C5814 D_FlipFlop_0.3-input-nand_2.C.n2 GND 0.04327f
C5815 D_FlipFlop_0.3-input-nand_2.C.n3 GND 0.09193f
C5816 D_FlipFlop_0.3-input-nand_2.C.t5 GND 0.17806f
C5817 D_FlipFlop_0.3-input-nand_2.C.t6 GND 0.34248f
C5818 D_FlipFlop_0.3-input-nand_2.C.n4 GND 0.10005f
C5819 D_FlipFlop_0.3-input-nand_2.C.n5 GND 0.04279f
C5820 D_FlipFlop_0.3-input-nand_2.C.n6 GND 0.079f
C5821 D_FlipFlop_0.3-input-nand_2.C.n7 GND 0.13677f
C5822 D_FlipFlop_0.3-input-nand_2.C.n8 GND 0.10181f
C5823 D_FlipFlop_0.3-input-nand_2.C.n9 GND 0.04823f
C5824 D_FlipFlop_0.3-input-nand_2.C.n10 GND 0.124f
C5825 D_FlipFlop_0.3-input-nand_2.C.t1 GND 0.04742f
C5826 D_FlipFlop_0.3-input-nand_2.C.t0 GND 0.04645f
C5827 D_FlipFlop_0.3-input-nand_2.C.n11 GND 0.26418f
C5828 D_FlipFlop_0.3-input-nand_2.C.n12 GND 0.08722f
C5829 D_FlipFlop_0.3-input-nand_2.C.t2 GND 0.04645f
C5830 D_FlipFlop_0.3-input-nand_2.C.n13 GND 0.293f
C5831 D_FlipFlop_0.3-input-nand_2.C.t4 GND 0.17045f
C5832 D_FlipFlop_0.3-input-nand_2.C.n14 GND 0.05129f
C5833 D_FlipFlop_6.nPRE.t2 GND 0.03228f
C5834 D_FlipFlop_6.nPRE.t16 GND 0.22918f
C5835 D_FlipFlop_6.nPRE.n0 GND 0.06695f
C5836 D_FlipFlop_6.nPRE.n1 GND 0.02905f
C5837 D_FlipFlop_6.nPRE.n2 GND 0.12772f
C5838 D_FlipFlop_6.nPRE.t14 GND 0.10659f
C5839 D_FlipFlop_6.nPRE.n3 GND 0.06116f
C5840 D_FlipFlop_6.nPRE.n4 GND 0.12963f
C5841 D_FlipFlop_6.nPRE.t17 GND 0.22919f
C5842 D_FlipFlop_6.nPRE.n5 GND 0.2308f
C5843 D_FlipFlop_6.nPRE.n6 GND 0.02462f
C5844 D_FlipFlop_6.nPRE.t5 GND 0.11915f
C5845 D_FlipFlop_6.nPRE.n7 GND 0.03432f
C5846 D_FlipFlop_6.nPRE.n9 GND 0.01425f
C5847 D_FlipFlop_6.nPRE.n10 GND 0.14213f
C5848 D_FlipFlop_6.nPRE.t6 GND 0.22919f
C5849 D_FlipFlop_6.nPRE.n11 GND 0.2308f
C5850 D_FlipFlop_6.nPRE.n12 GND 0.02462f
C5851 D_FlipFlop_6.nPRE.t11 GND 0.11915f
C5852 D_FlipFlop_6.nPRE.n13 GND 0.03432f
C5853 D_FlipFlop_6.nPRE.n15 GND 0.01425f
C5854 D_FlipFlop_6.nPRE.n17 GND 0.36888f
C5855 D_FlipFlop_6.nPRE.n18 GND 0.47983f
C5856 D_FlipFlop_6.nPRE.t10 GND 0.22918f
C5857 D_FlipFlop_6.nPRE.n19 GND 0.06695f
C5858 D_FlipFlop_6.nPRE.n20 GND 0.02905f
C5859 D_FlipFlop_6.nPRE.n21 GND 0.12772f
C5860 D_FlipFlop_6.nPRE.t9 GND 0.10813f
C5861 D_FlipFlop_6.nPRE.n22 GND 1.09701f
C5862 D_FlipFlop_6.nPRE.t15 GND 0.11915f
C5863 D_FlipFlop_6.nPRE.n23 GND 0.03121f
C5864 D_FlipFlop_6.nPRE.n24 GND 0.02863f
C5865 D_FlipFlop_6.nPRE.t7 GND 0.22949f
C5866 D_FlipFlop_6.nPRE.n25 GND 0.06884f
C5867 D_FlipFlop_6.nPRE.t4 GND 0.11915f
C5868 D_FlipFlop_6.nPRE.n26 GND 0.03121f
C5869 D_FlipFlop_6.nPRE.n27 GND 0.02863f
C5870 D_FlipFlop_6.nPRE.n28 GND 0.07244f
C5871 D_FlipFlop_6.nPRE.n29 GND 0.07244f
C5872 D_FlipFlop_6.nPRE.n30 GND 0.06884f
C5873 D_FlipFlop_6.nPRE.t13 GND 0.29304f
C5874 D_FlipFlop_6.nPRE.n31 GND 0.07187f
C5875 D_FlipFlop_6.nPRE.n32 GND 0.37446f
C5876 D_FlipFlop_6.nPRE.n33 GND 0.14559f
C5877 D_FlipFlop_6.nPRE.t12 GND 0.22918f
C5878 D_FlipFlop_6.nPRE.n34 GND 0.09982f
C5879 D_FlipFlop_6.nPRE.t8 GND 0.10697f
C5880 D_FlipFlop_6.nPRE.n35 GND 0.06983f
C5881 D_FlipFlop_6.nPRE.n36 GND 0.03344f
C5882 D_FlipFlop_6.nPRE.n37 GND 0.08479f
C5883 D_FlipFlop_6.nPRE.t1 GND 0.03109f
C5884 D_FlipFlop_6.nPRE.n38 GND 0.04788f
C5885 D_FlipFlop_6.nPRE.t3 GND 0.03173f
C5886 D_FlipFlop_6.nPRE.t0 GND 0.03109f
C5887 D_FlipFlop_6.nPRE.n39 GND 0.17678f
C5888 D_FlipFlop_6.nPRE.n40 GND 0.05768f
C5889 D_FlipFlop_6.nPRE.n41 GND 0.11614f
C5890 Q7.t1 GND 0.05851f
C5891 Q7.n0 GND 0.28696f
C5892 Q7.n1 GND 0.0654f
C5893 Q7.t2 GND 0.06212f
C5894 Q7.t3 GND 0.06085f
C5895 Q7.n2 GND 0.34604f
C5896 Q7.n3 GND 0.11291f
C5897 Q7.t0 GND 0.06085f
C5898 Q7.n4 GND 0.09373f
C5899 Q7.n5 GND 0.16597f
C5900 Q7.n6 GND 0.06546f
C5901 Q7.t8 GND 0.4486f
C5902 Q7.n7 GND 0.13105f
C5903 Q7.n8 GND 0.05686f
C5904 Q7.n9 GND 0.25001f
C5905 Q7.t4 GND 0.20863f
C5906 Q7.n10 GND 0.48035f
C5907 Q7.n11 GND 5.19948f
C5908 Q7.t9 GND 0.23339f
C5909 Q7.t7 GND 0.45064f
C5910 Q7.n12 GND 0.33455f
C5911 Q7.n13 GND 0.0619f
C5912 Q7.t5 GND 0.23339f
C5913 Q7.t6 GND 0.45064f
C5914 Q7.n14 GND 0.33246f
C5915 Q7.n15 GND 0.06668f
C5916 Q7.n16 GND 0.16987f
C5917 Q7.n17 GND 2.44085f
C5918 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 GND 0.05215f
C5919 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 GND 0.18008f
C5920 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 GND 0.37825f
C5921 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 GND 0.19588f
C5922 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 GND 0.28346f
C5923 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 GND 0.11199f
C5924 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 GND 0.01587f
C5925 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 GND 0.37675f
C5926 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 GND 0.16409f
C5927 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 GND 0.18888f
C5928 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 GND 0.0511f
C5929 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 GND 0.32168f
C5930 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 GND 0.05217f
C5931 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 GND 0.0511f
C5932 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 GND 0.29061f
C5933 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 GND 0.09483f
C5934 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 GND 0.01203f
C5935 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t3 GND 0.06145f
C5936 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n0 GND 0.15815f
C5937 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n1 GND 0.12861f
C5938 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t5 GND 0.24486f
C5939 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t6 GND 0.47095f
C5940 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n2 GND 0.11174f
C5941 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n3 GND 0.11082f
C5942 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n4 GND 0.18808f
C5943 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n5 GND 0.14f
C5944 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t7 GND 0.47302f
C5945 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n6 GND 0.20386f
C5946 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t4 GND 0.23439f
C5947 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t1 GND 0.06388f
C5948 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n7 GND 0.40291f
C5949 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t0 GND 0.06521f
C5950 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.t2 GND 0.06388f
C5951 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n8 GND 0.36328f
C5952 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n9 GND 0.12591f
C5953 Ring_Counter_0.D_FlipFlop_6.3-input-nand_2.C.n10 GND 0.07837f
C5954 D_FlipFlop_3.CLK.t1 GND 0.02954f
C5955 D_FlipFlop_3.CLK.t5 GND 0.22695f
C5956 D_FlipFlop_3.CLK.t2 GND 0.118f
C5957 D_FlipFlop_3.CLK.n0 GND 0.12444f
C5958 D_FlipFlop_3.CLK.t6 GND 0.22695f
C5959 D_FlipFlop_3.CLK.n1 GND 0.2009f
C5960 D_FlipFlop_3.CLK.n2 GND 0.20145f
C5961 D_FlipFlop_3.CLK.n3 GND 0.12607f
C5962 D_FlipFlop_3.CLK.t4 GND 0.10447f
C5963 D_FlipFlop_3.CLK.n4 GND 0.02736f
C5964 D_FlipFlop_3.CLK.n5 GND 0.10371f
C5965 D_FlipFlop_3.CLK.t3 GND 0.10446f
C5966 D_FlipFlop_3.CLK.n6 GND 0.03399f
C5967 D_FlipFlop_3.CLK.n7 GND 0.02546f
C5968 D_FlipFlop_3.CLK.n8 GND 0.23531f
C5969 D_FlipFlop_3.CLK.t7 GND 0.21911f
C5970 D_FlipFlop_3.CLK.n9 GND 0.16025f
C5971 D_FlipFlop_3.CLK.n11 GND 0.03049f
C5972 D_FlipFlop_3.CLK.t0 GND 0.03086f
C5973 D_FlipFlop_3.CLK.n12 GND 0.19695f
C5974 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t2 GND 0.06145f
C5975 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n0 GND 0.15815f
C5976 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n1 GND 0.12861f
C5977 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t7 GND 0.24486f
C5978 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t6 GND 0.47095f
C5979 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n2 GND 0.11174f
C5980 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n3 GND 0.11082f
C5981 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n4 GND 0.18808f
C5982 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n5 GND 0.14f
C5983 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t5 GND 0.47302f
C5984 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n6 GND 0.20386f
C5985 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t4 GND 0.23439f
C5986 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t1 GND 0.06388f
C5987 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n7 GND 0.40291f
C5988 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t0 GND 0.06521f
C5989 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.t3 GND 0.06388f
C5990 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n8 GND 0.36328f
C5991 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n9 GND 0.12591f
C5992 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.C.n10 GND 0.07837f
C5993 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 GND 0.37675f
C5994 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 GND 0.16409f
C5995 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 GND 0.18888f
C5996 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 GND 0.0511f
C5997 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 GND 0.32168f
C5998 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 GND 0.05217f
C5999 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 GND 0.0511f
C6000 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 GND 0.29061f
C6001 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 GND 0.09483f
C6002 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 GND 0.01203f
C6003 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 GND 0.01587f
C6004 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 GND 0.37825f
C6005 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 GND 0.19588f
C6006 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 GND 0.28346f
C6007 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 GND 0.11199f
C6008 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 GND 0.05215f
C6009 Ring_Counter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 GND 0.18008f
C6010 Q5.t3 GND 0.05543f
C6011 Q5.n0 GND 0.27185f
C6012 Q5.n1 GND 0.06196f
C6013 Q5.t0 GND 0.05885f
C6014 Q5.t1 GND 0.05764f
C6015 Q5.n2 GND 0.32782f
C6016 Q5.n3 GND 0.10697f
C6017 Q5.t2 GND 0.05764f
C6018 Q5.n4 GND 0.0888f
C6019 Q5.n5 GND 0.15723f
C6020 Q5.n6 GND 0.06201f
C6021 Q5.t8 GND 0.42498f
C6022 Q5.n7 GND 0.12415f
C6023 Q5.n8 GND 0.05387f
C6024 Q5.n9 GND 0.23685f
C6025 Q5.t7 GND 0.19765f
C6026 Q5.n10 GND 0.49797f
C6027 Q5.n11 GND 2.66911f
C6028 Q5.t6 GND 0.22111f
C6029 Q5.t4 GND 0.42692f
C6030 Q5.n12 GND 0.31694f
C6031 Q5.n13 GND 0.05865f
C6032 Q5.t9 GND 0.22111f
C6033 Q5.t5 GND 0.42692f
C6034 Q5.n14 GND 0.31496f
C6035 Q5.n15 GND 0.06317f
C6036 Q5.n16 GND 0.14115f
C6037 Q5.n17 GND 1.23083f
C6038 Ring_Counter_0.D_FlipFlop_3.Qbar.t1 GND 0.05347f
C6039 Ring_Counter_0.D_FlipFlop_3.Qbar.t5 GND 0.41161f
C6040 Ring_Counter_0.D_FlipFlop_3.Qbar.n0 GND 0.1774f
C6041 Ring_Counter_0.D_FlipFlop_3.Qbar.t4 GND 0.18986f
C6042 Ring_Counter_0.D_FlipFlop_3.Qbar.n1 GND 0.23199f
C6043 Ring_Counter_0.D_FlipFlop_3.Qbar.n2 GND 0.05991f
C6044 Ring_Counter_0.D_FlipFlop_3.Qbar.t3 GND 0.05559f
C6045 Ring_Counter_0.D_FlipFlop_3.Qbar.n3 GND 0.09627f
C6046 Ring_Counter_0.D_FlipFlop_3.Qbar.t0 GND 0.05675f
C6047 Ring_Counter_0.D_FlipFlop_3.Qbar.t2 GND 0.05559f
C6048 Ring_Counter_0.D_FlipFlop_3.Qbar.n4 GND 0.31612f
C6049 Ring_Counter_0.D_FlipFlop_3.Qbar.n5 GND 0.16106f
C6050 Ring_Counter_0.D_FlipFlop_3.Qbar.n6 GND 0.15403f
C6051 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 GND 0.06443f
C6052 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 GND 0.14002f
C6053 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 GND 0.07316f
C6054 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 GND 0.25702f
C6055 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 GND 0.12462f
C6056 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 GND 0.4938f
C6057 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 GND 0.09136f
C6058 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 GND 0.05451f
C6059 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 GND 0.13379f
C6060 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 GND 0.13379f
C6061 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 GND 0.06713f
C6062 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 GND 0.07989f
C6063 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 GND 0.43786f
C6064 Ring_Counter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 GND 0.08018f
C6065 Q6.t1 GND 0.0885f
C6066 Q6.n0 GND 0.434f
C6067 Q6.n1 GND 0.09891f
C6068 Q6.t2 GND 0.09395f
C6069 Q6.t3 GND 0.09203f
C6070 Q6.n2 GND 0.52335f
C6071 Q6.n3 GND 0.17077f
C6072 Q6.t0 GND 0.09203f
C6073 Q6.n4 GND 0.14176f
C6074 Q6.n5 GND 0.25101f
C6075 Q6.n6 GND 0.099f
C6076 Q6.t6 GND 0.67847f
C6077 Q6.n7 GND 0.1982f
C6078 Q6.n8 GND 0.086f
C6079 Q6.n9 GND 0.37811f
C6080 Q6.t4 GND 0.31554f
C6081 Q6.n10 GND 0.76097f
C6082 Q6.n11 GND 6.0622f
C6083 Q6.t9 GND 0.35299f
C6084 Q6.t7 GND 0.68156f
C6085 Q6.n12 GND 0.50598f
C6086 Q6.n13 GND 0.09362f
C6087 Q6.t8 GND 0.35299f
C6088 Q6.t5 GND 0.68156f
C6089 Q6.n14 GND 0.50282f
C6090 Q6.n15 GND 0.10085f
C6091 Q6.n16 GND 0.24107f
C6092 Q6.n17 GND 2.82827f
C6093 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 GND 0.07411f
C6094 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 GND 0.16107f
C6095 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 GND 0.08416f
C6096 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 GND 0.29566f
C6097 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 GND 0.14335f
C6098 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 GND 0.56804f
C6099 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 GND 0.1051f
C6100 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 GND 0.06271f
C6101 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 GND 0.15391f
C6102 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 GND 0.15391f
C6103 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 GND 0.07722f
C6104 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 GND 0.07866f
C6105 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 GND 0.07705f
C6106 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 GND 0.43817f
C6107 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 GND 0.286f
C6108 Ring_Counter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 GND 0.09223f
C6109 D_FlipFlop_0.3-input-nand_2.Vout.t5 GND 0.35515f
C6110 D_FlipFlop_0.3-input-nand_2.Vout.n0 GND 0.10375f
C6111 D_FlipFlop_0.3-input-nand_2.Vout.n1 GND 0.04502f
C6112 D_FlipFlop_0.3-input-nand_2.Vout.t1 GND 0.04632f
C6113 D_FlipFlop_0.3-input-nand_2.Vout.n2 GND 0.22028f
C6114 D_FlipFlop_0.3-input-nand_2.Vout.n3 GND 0.05002f
C6115 D_FlipFlop_0.3-input-nand_2.Vout.t7 GND 0.35517f
C6116 D_FlipFlop_0.3-input-nand_2.Vout.n4 GND 0.36759f
C6117 D_FlipFlop_0.3-input-nand_2.Vout.t6 GND 0.18465f
C6118 D_FlipFlop_0.3-input-nand_2.Vout.n5 GND 0.18106f
C6119 D_FlipFlop_0.3-input-nand_2.Vout.n6 GND 0.10557f
C6120 D_FlipFlop_0.3-input-nand_2.Vout.n7 GND 0.01331f
C6121 D_FlipFlop_0.3-input-nand_2.Vout.n8 GND 0.01057f
C6122 D_FlipFlop_0.3-input-nand_2.Vout.t2 GND 0.04918f
C6123 D_FlipFlop_0.3-input-nand_2.Vout.t3 GND 0.04817f
C6124 D_FlipFlop_0.3-input-nand_2.Vout.n9 GND 0.27396f
C6125 D_FlipFlop_0.3-input-nand_2.Vout.n10 GND 0.08939f
C6126 D_FlipFlop_0.3-input-nand_2.Vout.t0 GND 0.04817f
C6127 D_FlipFlop_0.3-input-nand_2.Vout.n11 GND 0.30324f
C6128 D_FlipFlop_0.3-input-nand_2.Vout.t4 GND 0.17747f
C6129 D_FlipFlop_0.3-input-nand_2.Vout.n12 GND 0.19793f
C6130 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 GND 0.05215f
C6131 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 GND 0.18008f
C6132 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 GND 0.37825f
C6133 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 GND 0.19588f
C6134 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 GND 0.28346f
C6135 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 GND 0.11199f
C6136 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 GND 0.01587f
C6137 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 GND 0.37675f
C6138 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 GND 0.16409f
C6139 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 GND 0.18888f
C6140 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 GND 0.0511f
C6141 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 GND 0.32168f
C6142 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 GND 0.05217f
C6143 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 GND 0.0511f
C6144 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 GND 0.29061f
C6145 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 GND 0.09483f
C6146 Ring_Counter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 GND 0.01203f
C6147 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 GND 0.05215f
C6148 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 GND 0.18008f
C6149 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 GND 0.37825f
C6150 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 GND 0.19588f
C6151 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 GND 0.28346f
C6152 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 GND 0.11199f
C6153 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 GND 0.01587f
C6154 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 GND 0.37675f
C6155 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 GND 0.16409f
C6156 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 GND 0.18888f
C6157 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 GND 0.0511f
C6158 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 GND 0.32168f
C6159 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 GND 0.05217f
C6160 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 GND 0.0511f
C6161 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 GND 0.29061f
C6162 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 GND 0.09483f
C6163 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 GND 0.01203f
C6164 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t1 GND 0.06145f
C6165 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n0 GND 0.15815f
C6166 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n1 GND 0.12861f
C6167 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t7 GND 0.24486f
C6168 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t6 GND 0.47095f
C6169 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n2 GND 0.11174f
C6170 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n3 GND 0.11082f
C6171 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n4 GND 0.18808f
C6172 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n5 GND 0.14f
C6173 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t5 GND 0.47302f
C6174 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n6 GND 0.20386f
C6175 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t4 GND 0.23439f
C6176 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t3 GND 0.06388f
C6177 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n7 GND 0.40291f
C6178 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t0 GND 0.06521f
C6179 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.t2 GND 0.06388f
C6180 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n8 GND 0.36328f
C6181 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n9 GND 0.12591f
C6182 Ring_Counter_0.D_FlipFlop_2.3-input-nand_2.C.n10 GND 0.07837f
C6183 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t3 GND 0.06145f
C6184 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n0 GND 0.15815f
C6185 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n1 GND 0.12861f
C6186 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t6 GND 0.24486f
C6187 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t4 GND 0.47095f
C6188 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n2 GND 0.11174f
C6189 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n3 GND 0.11082f
C6190 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n4 GND 0.18808f
C6191 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n5 GND 0.14f
C6192 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t7 GND 0.47302f
C6193 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n6 GND 0.20386f
C6194 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t5 GND 0.23439f
C6195 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t2 GND 0.06388f
C6196 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n7 GND 0.40291f
C6197 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t1 GND 0.06521f
C6198 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.t0 GND 0.06388f
C6199 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n8 GND 0.36328f
C6200 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n9 GND 0.12591f
C6201 Ring_Counter_0.D_FlipFlop_15.3-input-nand_2.C.n10 GND 0.07837f
C6202 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 GND 0.07411f
C6203 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 GND 0.16107f
C6204 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 GND 0.08416f
C6205 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 GND 0.29566f
C6206 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 GND 0.14335f
C6207 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 GND 0.56804f
C6208 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 GND 0.1051f
C6209 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 GND 0.06271f
C6210 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 GND 0.15391f
C6211 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 GND 0.15391f
C6212 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 GND 0.07722f
C6213 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 GND 0.07866f
C6214 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 GND 0.07705f
C6215 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 GND 0.43817f
C6216 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 GND 0.286f
C6217 Ring_Counter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 GND 0.09223f
C6218 D_FlipFlop_7.CLK.t1 GND 0.02954f
C6219 D_FlipFlop_7.CLK.t5 GND 0.22695f
C6220 D_FlipFlop_7.CLK.t7 GND 0.118f
C6221 D_FlipFlop_7.CLK.n0 GND 0.12444f
C6222 D_FlipFlop_7.CLK.t2 GND 0.22695f
C6223 D_FlipFlop_7.CLK.n1 GND 0.2009f
C6224 D_FlipFlop_7.CLK.n2 GND 0.20145f
C6225 D_FlipFlop_7.CLK.n3 GND 0.12607f
C6226 D_FlipFlop_7.CLK.t4 GND 0.10447f
C6227 D_FlipFlop_7.CLK.n4 GND 0.02736f
C6228 D_FlipFlop_7.CLK.n5 GND 0.10371f
C6229 D_FlipFlop_7.CLK.t3 GND 0.10446f
C6230 D_FlipFlop_7.CLK.n6 GND 0.03399f
C6231 D_FlipFlop_7.CLK.n7 GND 0.02546f
C6232 D_FlipFlop_7.CLK.n8 GND 0.23531f
C6233 D_FlipFlop_7.CLK.t6 GND 0.21911f
C6234 D_FlipFlop_7.CLK.n9 GND 0.16025f
C6235 D_FlipFlop_7.CLK.n11 GND 0.03049f
C6236 D_FlipFlop_7.CLK.t0 GND 0.03086f
C6237 D_FlipFlop_7.CLK.n12 GND 0.19695f
C6238 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t4 GND 0.47302f
C6239 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n0 GND 0.20386f
C6240 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t7 GND 0.23439f
C6241 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t1 GND 0.06388f
C6242 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n1 GND 0.40291f
C6243 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t2 GND 0.06521f
C6244 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t3 GND 0.06388f
C6245 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n2 GND 0.36328f
C6246 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n3 GND 0.12591f
C6247 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n4 GND 0.07837f
C6248 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t6 GND 0.24486f
C6249 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t5 GND 0.47095f
C6250 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n5 GND 0.11174f
C6251 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n6 GND 0.11082f
C6252 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n7 GND 0.18808f
C6253 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n8 GND 0.14f
C6254 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n9 GND 0.12861f
C6255 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.t0 GND 0.06145f
C6256 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.C.n10 GND 0.15815f
C6257 D_FlipFlop_1.nPRE.t1 GND 0.04604f
C6258 D_FlipFlop_1.nPRE.t17 GND 0.3269f
C6259 D_FlipFlop_1.nPRE.n0 GND 0.0955f
C6260 D_FlipFlop_1.nPRE.n1 GND 0.04144f
C6261 D_FlipFlop_1.nPRE.n2 GND 0.18219f
C6262 D_FlipFlop_1.nPRE.t16 GND 0.15673f
C6263 D_FlipFlop_1.nPRE.t15 GND 0.3269f
C6264 D_FlipFlop_1.nPRE.n3 GND 0.0955f
C6265 D_FlipFlop_1.nPRE.n4 GND 0.04144f
C6266 D_FlipFlop_1.nPRE.n5 GND 0.18219f
C6267 D_FlipFlop_1.nPRE.t12 GND 0.15203f
C6268 D_FlipFlop_1.nPRE.n6 GND 0.08724f
C6269 D_FlipFlop_1.nPRE.n7 GND 0.18491f
C6270 D_FlipFlop_1.nPRE.t9 GND 0.32692f
C6271 D_FlipFlop_1.nPRE.n8 GND 0.32922f
C6272 D_FlipFlop_1.nPRE.n9 GND 0.03512f
C6273 D_FlipFlop_1.nPRE.t14 GND 0.16996f
C6274 D_FlipFlop_1.nPRE.n10 GND 0.04896f
C6275 D_FlipFlop_1.nPRE.n11 GND 0.01304f
C6276 D_FlipFlop_1.nPRE.n12 GND 0.02032f
C6277 D_FlipFlop_1.nPRE.n13 GND 0.20274f
C6278 D_FlipFlop_1.nPRE.t5 GND 0.32692f
C6279 D_FlipFlop_1.nPRE.n14 GND 0.32922f
C6280 D_FlipFlop_1.nPRE.n15 GND 0.03512f
C6281 D_FlipFlop_1.nPRE.t13 GND 0.16996f
C6282 D_FlipFlop_1.nPRE.n16 GND 0.04896f
C6283 D_FlipFlop_1.nPRE.n17 GND 0.01304f
C6284 D_FlipFlop_1.nPRE.n18 GND 0.02032f
C6285 D_FlipFlop_1.nPRE.n20 GND 0.52619f
C6286 D_FlipFlop_1.nPRE.n21 GND 0.54528f
C6287 D_FlipFlop_1.nPRE.n22 GND 0.91254f
C6288 D_FlipFlop_1.nPRE.t6 GND 0.16996f
C6289 D_FlipFlop_1.nPRE.n23 GND 0.04453f
C6290 D_FlipFlop_1.nPRE.n24 GND 0.04084f
C6291 D_FlipFlop_1.nPRE.t11 GND 0.32735f
C6292 D_FlipFlop_1.nPRE.n25 GND 0.0982f
C6293 D_FlipFlop_1.nPRE.t8 GND 0.16996f
C6294 D_FlipFlop_1.nPRE.n26 GND 0.04453f
C6295 D_FlipFlop_1.nPRE.n27 GND 0.04084f
C6296 D_FlipFlop_1.nPRE.n28 GND 0.10333f
C6297 D_FlipFlop_1.nPRE.n29 GND 0.10333f
C6298 D_FlipFlop_1.nPRE.n30 GND 0.0982f
C6299 D_FlipFlop_1.nPRE.t4 GND 0.418f
C6300 D_FlipFlop_1.nPRE.n31 GND 0.10252f
C6301 D_FlipFlop_1.nPRE.n32 GND 0.28221f
C6302 D_FlipFlop_1.nPRE.n33 GND 0.20767f
C6303 D_FlipFlop_1.nPRE.t10 GND 0.3269f
C6304 D_FlipFlop_1.nPRE.n34 GND 0.14238f
C6305 D_FlipFlop_1.nPRE.t7 GND 0.15258f
C6306 D_FlipFlop_1.nPRE.n35 GND 0.0996f
C6307 D_FlipFlop_1.nPRE.n36 GND 0.0477f
C6308 D_FlipFlop_1.nPRE.n37 GND 0.12094f
C6309 D_FlipFlop_1.nPRE.t0 GND 0.04434f
C6310 D_FlipFlop_1.nPRE.n38 GND 0.0683f
C6311 D_FlipFlop_1.nPRE.t2 GND 0.04527f
C6312 D_FlipFlop_1.nPRE.t3 GND 0.04434f
C6313 D_FlipFlop_1.nPRE.n39 GND 0.25216f
C6314 D_FlipFlop_1.nPRE.n40 GND 0.08228f
C6315 D_FlipFlop_1.nPRE.n41 GND 0.16567f
C6316 Nand_Gate_3.A.t2 GND 0.05065f
C6317 Nand_Gate_3.A.t10 GND 0.3596f
C6318 Nand_Gate_3.A.n0 GND 0.10505f
C6319 Nand_Gate_3.A.n1 GND 0.04558f
C6320 Nand_Gate_3.A.n2 GND 0.20041f
C6321 Nand_Gate_3.A.t9 GND 0.19713f
C6322 Nand_Gate_3.A.t4 GND 0.18696f
C6323 Nand_Gate_3.A.n3 GND 0.04898f
C6324 Nand_Gate_3.A.n4 GND 0.04492f
C6325 Nand_Gate_3.A.t5 GND 0.36008f
C6326 Nand_Gate_3.A.n5 GND 0.10802f
C6327 Nand_Gate_3.A.t7 GND 0.18696f
C6328 Nand_Gate_3.A.n6 GND 0.04898f
C6329 Nand_Gate_3.A.n7 GND 0.04492f
C6330 Nand_Gate_3.A.n8 GND 0.11367f
C6331 Nand_Gate_3.A.n9 GND 0.11367f
C6332 Nand_Gate_3.A.n10 GND 0.10802f
C6333 Nand_Gate_3.A.t11 GND 0.4598f
C6334 Nand_Gate_3.A.n11 GND 0.11278f
C6335 Nand_Gate_3.A.n12 GND 1.10144f
C6336 Nand_Gate_3.A.n13 GND 0.22844f
C6337 Nand_Gate_3.A.t8 GND 0.3596f
C6338 Nand_Gate_3.A.n14 GND 0.15662f
C6339 Nand_Gate_3.A.t6 GND 0.16784f
C6340 Nand_Gate_3.A.n15 GND 0.10956f
C6341 Nand_Gate_3.A.n16 GND 0.05247f
C6342 Nand_Gate_3.A.n17 GND 0.13304f
C6343 Nand_Gate_3.A.t1 GND 0.04878f
C6344 Nand_Gate_3.A.n18 GND 0.07513f
C6345 Nand_Gate_3.A.t3 GND 0.04979f
C6346 Nand_Gate_3.A.t0 GND 0.04878f
C6347 Nand_Gate_3.A.n19 GND 0.27738f
C6348 Nand_Gate_3.A.n20 GND 0.09051f
C6349 Nand_Gate_3.A.n21 GND 0.18223f
C6350 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t1 GND 0.05f
C6351 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n0 GND 0.10867f
C6352 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n1 GND 0.05678f
C6353 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t3 GND 0.38491f
C6354 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n2 GND 0.16589f
C6355 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t2 GND 0.30131f
C6356 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t4 GND 0.30153f
C6357 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n3 GND 0.09671f
C6358 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t5 GND 0.38323f
C6359 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n4 GND 0.0709f
C6360 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n5 GND 0.04231f
C6361 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n6 GND 0.10383f
C6362 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n7 GND 0.10383f
C6363 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.t0 GND 0.05284f
C6364 Ring_Counter_0.D_FlipFlop_3.Inverter_1.Vout.n8 GND 0.17757f
C6365 D_FlipFlop_7.nPRE.t4 GND 0.22672f
C6366 D_FlipFlop_7.nPRE.n0 GND 0.06623f
C6367 D_FlipFlop_7.nPRE.n1 GND 0.02874f
C6368 D_FlipFlop_7.nPRE.n2 GND 0.12635f
C6369 D_FlipFlop_7.nPRE.t10 GND 0.10544f
C6370 D_FlipFlop_7.nPRE.n3 GND 0.06051f
C6371 D_FlipFlop_7.nPRE.n4 GND 0.12825f
C6372 D_FlipFlop_7.nPRE.t5 GND 0.22673f
C6373 D_FlipFlop_7.nPRE.n5 GND 0.22833f
C6374 D_FlipFlop_7.nPRE.n6 GND 0.02435f
C6375 D_FlipFlop_7.nPRE.t12 GND 0.11788f
C6376 D_FlipFlop_7.nPRE.n7 GND 0.03396f
C6377 D_FlipFlop_7.nPRE.n9 GND 0.01409f
C6378 D_FlipFlop_7.nPRE.n10 GND 0.14061f
C6379 D_FlipFlop_7.nPRE.t11 GND 0.22673f
C6380 D_FlipFlop_7.nPRE.n11 GND 0.22833f
C6381 D_FlipFlop_7.nPRE.n12 GND 0.02435f
C6382 D_FlipFlop_7.nPRE.t15 GND 0.11788f
C6383 D_FlipFlop_7.nPRE.n13 GND 0.03396f
C6384 D_FlipFlop_7.nPRE.n15 GND 0.01409f
C6385 D_FlipFlop_7.nPRE.n17 GND 0.36493f
C6386 D_FlipFlop_7.nPRE.n18 GND 0.46392f
C6387 D_FlipFlop_7.nPRE.t14 GND 0.22672f
C6388 D_FlipFlop_7.nPRE.n19 GND 0.06623f
C6389 D_FlipFlop_7.nPRE.n20 GND 0.02874f
C6390 D_FlipFlop_7.nPRE.n21 GND 0.12635f
C6391 D_FlipFlop_7.nPRE.t6 GND 0.10661f
C6392 D_FlipFlop_7.nPRE.n22 GND 1.18619f
C6393 D_FlipFlop_7.nPRE.t8 GND 0.11788f
C6394 D_FlipFlop_7.nPRE.n23 GND 0.03088f
C6395 D_FlipFlop_7.nPRE.n24 GND 0.02832f
C6396 D_FlipFlop_7.nPRE.t16 GND 0.22703f
C6397 D_FlipFlop_7.nPRE.n25 GND 0.0681f
C6398 D_FlipFlop_7.nPRE.t13 GND 0.11788f
C6399 D_FlipFlop_7.nPRE.n26 GND 0.03088f
C6400 D_FlipFlop_7.nPRE.n27 GND 0.02832f
C6401 D_FlipFlop_7.nPRE.n28 GND 0.07167f
C6402 D_FlipFlop_7.nPRE.n29 GND 0.07167f
C6403 D_FlipFlop_7.nPRE.n30 GND 0.0681f
C6404 D_FlipFlop_7.nPRE.t9 GND 0.2899f
C6405 D_FlipFlop_7.nPRE.n31 GND 0.0711f
C6406 D_FlipFlop_7.nPRE.n32 GND 0.46206f
C6407 D_FlipFlop_7.nPRE.n33 GND 0.14403f
C6408 D_FlipFlop_7.nPRE.t17 GND 0.22672f
C6409 D_FlipFlop_7.nPRE.n34 GND 0.09875f
C6410 D_FlipFlop_7.nPRE.t7 GND 0.10582f
C6411 D_FlipFlop_7.nPRE.n35 GND 0.06908f
C6412 D_FlipFlop_7.nPRE.n36 GND 0.03308f
C6413 D_FlipFlop_7.nPRE.n37 GND 0.08388f
C6414 D_FlipFlop_7.nPRE.t3 GND 0.03075f
C6415 D_FlipFlop_7.nPRE.n38 GND 0.04737f
C6416 D_FlipFlop_7.nPRE.t2 GND 0.03139f
C6417 D_FlipFlop_7.nPRE.t1 GND 0.03075f
C6418 D_FlipFlop_7.nPRE.n39 GND 0.17489f
C6419 D_FlipFlop_7.nPRE.n40 GND 0.05707f
C6420 D_FlipFlop_7.nPRE.t0 GND 0.03193f
C6421 D_FlipFlop_7.nPRE.n41 GND 0.1149f
C6422 D_FlipFlop_2.3-input-nand_2.C.t7 GND 0.3425f
C6423 D_FlipFlop_2.3-input-nand_2.C.n0 GND 0.3551f
C6424 D_FlipFlop_2.3-input-nand_2.C.n1 GND 0.03842f
C6425 D_FlipFlop_2.3-input-nand_2.C.t3 GND 0.04469f
C6426 D_FlipFlop_2.3-input-nand_2.C.n2 GND 0.04327f
C6427 D_FlipFlop_2.3-input-nand_2.C.n3 GND 0.09193f
C6428 D_FlipFlop_2.3-input-nand_2.C.t4 GND 0.17806f
C6429 D_FlipFlop_2.3-input-nand_2.C.t6 GND 0.34248f
C6430 D_FlipFlop_2.3-input-nand_2.C.n4 GND 0.10005f
C6431 D_FlipFlop_2.3-input-nand_2.C.n5 GND 0.04279f
C6432 D_FlipFlop_2.3-input-nand_2.C.n6 GND 0.079f
C6433 D_FlipFlop_2.3-input-nand_2.C.n7 GND 0.13677f
C6434 D_FlipFlop_2.3-input-nand_2.C.n8 GND 0.10181f
C6435 D_FlipFlop_2.3-input-nand_2.C.n9 GND 0.04823f
C6436 D_FlipFlop_2.3-input-nand_2.C.n10 GND 0.124f
C6437 D_FlipFlop_2.3-input-nand_2.C.t1 GND 0.04742f
C6438 D_FlipFlop_2.3-input-nand_2.C.t0 GND 0.04645f
C6439 D_FlipFlop_2.3-input-nand_2.C.n11 GND 0.26418f
C6440 D_FlipFlop_2.3-input-nand_2.C.n12 GND 0.08722f
C6441 D_FlipFlop_2.3-input-nand_2.C.t2 GND 0.04645f
C6442 D_FlipFlop_2.3-input-nand_2.C.n13 GND 0.293f
C6443 D_FlipFlop_2.3-input-nand_2.C.t5 GND 0.17045f
C6444 D_FlipFlop_2.3-input-nand_2.C.n14 GND 0.05129f
C6445 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t2 GND 0.07892f
C6446 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n0 GND 0.25342f
C6447 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t4 GND 0.58988f
C6448 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n1 GND 0.17695f
C6449 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t5 GND 0.30628f
C6450 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n2 GND 0.08023f
C6451 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n3 GND 0.07359f
C6452 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n4 GND 0.15961f
C6453 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n5 GND 0.15961f
C6454 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n6 GND 0.0984f
C6455 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t1 GND 0.08008f
C6456 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t3 GND 0.08157f
C6457 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.t0 GND 0.0799f
C6458 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n7 GND 0.4544f
C6459 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n8 GND 0.25422f
C6460 Ring_Counter_0.D_FlipFlop_0.3-input-nand_0.Vout.n9 GND 0.04958f
C6461 Ring_Counter_0.D_FlipFlop_10.Qbar.t3 GND 0.05347f
C6462 Ring_Counter_0.D_FlipFlop_10.Qbar.t4 GND 0.41161f
C6463 Ring_Counter_0.D_FlipFlop_10.Qbar.n0 GND 0.1774f
C6464 Ring_Counter_0.D_FlipFlop_10.Qbar.t5 GND 0.18986f
C6465 Ring_Counter_0.D_FlipFlop_10.Qbar.n1 GND 0.23199f
C6466 Ring_Counter_0.D_FlipFlop_10.Qbar.n2 GND 0.05991f
C6467 Ring_Counter_0.D_FlipFlop_10.Qbar.t2 GND 0.05559f
C6468 Ring_Counter_0.D_FlipFlop_10.Qbar.n3 GND 0.09627f
C6469 Ring_Counter_0.D_FlipFlop_10.Qbar.t1 GND 0.05675f
C6470 Ring_Counter_0.D_FlipFlop_10.Qbar.t0 GND 0.05559f
C6471 Ring_Counter_0.D_FlipFlop_10.Qbar.n4 GND 0.31612f
C6472 Ring_Counter_0.D_FlipFlop_10.Qbar.n5 GND 0.16106f
C6473 Ring_Counter_0.D_FlipFlop_10.Qbar.n6 GND 0.15403f
C6474 D_FlipFlop_4.nPRE.t14 GND 0.23576f
C6475 D_FlipFlop_4.nPRE.n0 GND 0.06887f
C6476 D_FlipFlop_4.nPRE.n1 GND 0.02988f
C6477 D_FlipFlop_4.nPRE.n2 GND 0.13139f
C6478 D_FlipFlop_4.nPRE.t12 GND 0.10965f
C6479 D_FlipFlop_4.nPRE.n3 GND 0.06292f
C6480 D_FlipFlop_4.nPRE.n4 GND 0.13336f
C6481 D_FlipFlop_4.nPRE.t8 GND 0.23577f
C6482 D_FlipFlop_4.nPRE.n5 GND 0.23743f
C6483 D_FlipFlop_4.nPRE.n6 GND 0.02533f
C6484 D_FlipFlop_4.nPRE.t13 GND 0.12258f
C6485 D_FlipFlop_4.nPRE.n7 GND 0.03531f
C6486 D_FlipFlop_4.nPRE.n9 GND 0.01466f
C6487 D_FlipFlop_4.nPRE.n10 GND 0.14621f
C6488 D_FlipFlop_4.nPRE.t5 GND 0.23577f
C6489 D_FlipFlop_4.nPRE.n11 GND 0.23743f
C6490 D_FlipFlop_4.nPRE.n12 GND 0.02533f
C6491 D_FlipFlop_4.nPRE.t7 GND 0.12258f
C6492 D_FlipFlop_4.nPRE.n13 GND 0.03531f
C6493 D_FlipFlop_4.nPRE.n15 GND 0.01466f
C6494 D_FlipFlop_4.nPRE.n17 GND 0.37948f
C6495 D_FlipFlop_4.nPRE.n18 GND 0.48242f
C6496 D_FlipFlop_4.nPRE.t17 GND 0.23576f
C6497 D_FlipFlop_4.nPRE.n19 GND 0.06887f
C6498 D_FlipFlop_4.nPRE.n20 GND 0.02988f
C6499 D_FlipFlop_4.nPRE.n21 GND 0.13139f
C6500 D_FlipFlop_4.nPRE.t16 GND 0.11086f
C6501 D_FlipFlop_4.nPRE.n22 GND 0.98523f
C6502 D_FlipFlop_4.nPRE.t6 GND 0.12258f
C6503 D_FlipFlop_4.nPRE.n23 GND 0.03211f
C6504 D_FlipFlop_4.nPRE.n24 GND 0.02945f
C6505 D_FlipFlop_4.nPRE.t10 GND 0.23608f
C6506 D_FlipFlop_4.nPRE.n25 GND 0.07082f
C6507 D_FlipFlop_4.nPRE.t11 GND 0.12258f
C6508 D_FlipFlop_4.nPRE.n26 GND 0.03211f
C6509 D_FlipFlop_4.nPRE.n27 GND 0.02945f
C6510 D_FlipFlop_4.nPRE.n28 GND 0.07452f
C6511 D_FlipFlop_4.nPRE.n29 GND 0.07452f
C6512 D_FlipFlop_4.nPRE.n30 GND 0.07082f
C6513 D_FlipFlop_4.nPRE.t15 GND 0.30146f
C6514 D_FlipFlop_4.nPRE.n31 GND 0.07394f
C6515 D_FlipFlop_4.nPRE.n32 GND 0.32177f
C6516 D_FlipFlop_4.nPRE.n33 GND 0.14977f
C6517 D_FlipFlop_4.nPRE.t9 GND 0.23576f
C6518 D_FlipFlop_4.nPRE.n34 GND 0.10269f
C6519 D_FlipFlop_4.nPRE.t4 GND 0.11004f
C6520 D_FlipFlop_4.nPRE.n35 GND 0.07183f
C6521 D_FlipFlop_4.nPRE.n36 GND 0.0344f
C6522 D_FlipFlop_4.nPRE.n37 GND 0.08722f
C6523 D_FlipFlop_4.nPRE.t3 GND 0.03198f
C6524 D_FlipFlop_4.nPRE.n38 GND 0.04926f
C6525 D_FlipFlop_4.nPRE.t2 GND 0.03265f
C6526 D_FlipFlop_4.nPRE.t1 GND 0.03198f
C6527 D_FlipFlop_4.nPRE.n39 GND 0.18186f
C6528 D_FlipFlop_4.nPRE.n40 GND 0.05934f
C6529 D_FlipFlop_4.nPRE.t0 GND 0.03321f
C6530 D_FlipFlop_4.nPRE.n41 GND 0.11948f
C6531 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t1 GND 0.05f
C6532 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n0 GND 0.10867f
C6533 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n1 GND 0.05678f
C6534 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t2 GND 0.38491f
C6535 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n2 GND 0.16589f
C6536 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t4 GND 0.30131f
C6537 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t3 GND 0.30153f
C6538 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n3 GND 0.09671f
C6539 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t5 GND 0.38323f
C6540 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n4 GND 0.0709f
C6541 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n5 GND 0.04231f
C6542 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n6 GND 0.10383f
C6543 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n7 GND 0.10383f
C6544 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.t0 GND 0.05284f
C6545 Ring_Counter_0.D_FlipFlop_6.Inverter_1.Vout.n8 GND 0.17757f
C6546 CDAC_v3_0.switch_3.Z.t10 GND 0.07175f
C6547 CDAC_v3_0.switch_3.Z.t1 GND 0.07161f
C6548 CDAC_v3_0.switch_3.Z.n0 GND 0.15754f
C6549 CDAC_v3_0.switch_3.Z.n1 GND 0.02438f
C6550 CDAC_v3_0.switch_3.Z.t7 GND 9.71895f
C6551 CDAC_v3_0.switch_3.Z.t6 GND 9.71895f
C6552 CDAC_v3_0.switch_3.Z.t2 GND 9.71895f
C6553 CDAC_v3_0.switch_3.Z.t3 GND 11.5516f
C6554 CDAC_v3_0.switch_3.Z.n2 GND 3.07139f
C6555 CDAC_v3_0.switch_3.Z.n3 GND 2.99755f
C6556 CDAC_v3_0.switch_3.Z.n4 GND 5.21574f
C6557 CDAC_v3_0.switch_3.Z.t5 GND 9.71895f
C6558 CDAC_v3_0.switch_3.Z.t4 GND 9.71895f
C6559 CDAC_v3_0.switch_3.Z.t9 GND 9.71895f
C6560 CDAC_v3_0.switch_3.Z.t8 GND 13.3724f
C6561 CDAC_v3_0.switch_3.Z.n5 GND 3.14477f
C6562 CDAC_v3_0.switch_3.Z.n6 GND 2.99755f
C6563 CDAC_v3_0.switch_3.Z.n7 GND 2.55083f
C6564 CDAC_v3_0.switch_3.Z.n8 GND 11.5649f
C6565 CDAC_v3_0.switch_3.Z.n9 GND 4.49259f
C6566 CDAC_v3_0.switch_3.Z.n10 GND 0.07675f
C6567 CDAC_v3_0.switch_3.Z.t11 GND 0.07408f
C6568 CDAC_v3_0.switch_3.Z.t0 GND 0.07408f
C6569 CDAC_v3_0.switch_3.Z.n11 GND 0.26607f
C6570 CDAC_v3_0.switch_3.Z.n12 GND 0.82032f
C6571 D_FlipFlop_2.nPRE.t1 GND 0.04588f
C6572 D_FlipFlop_2.nPRE.t13 GND 0.32577f
C6573 D_FlipFlop_2.nPRE.n0 GND 0.09517f
C6574 D_FlipFlop_2.nPRE.n1 GND 0.04129f
C6575 D_FlipFlop_2.nPRE.n2 GND 0.18156f
C6576 D_FlipFlop_2.nPRE.t17 GND 0.15404f
C6577 D_FlipFlop_2.nPRE.t9 GND 0.32577f
C6578 D_FlipFlop_2.nPRE.n3 GND 0.09517f
C6579 D_FlipFlop_2.nPRE.n4 GND 0.04129f
C6580 D_FlipFlop_2.nPRE.n5 GND 0.18156f
C6581 D_FlipFlop_2.nPRE.t14 GND 0.15151f
C6582 D_FlipFlop_2.nPRE.n6 GND 0.08694f
C6583 D_FlipFlop_2.nPRE.n7 GND 0.18428f
C6584 D_FlipFlop_2.nPRE.t11 GND 0.32579f
C6585 D_FlipFlop_2.nPRE.n8 GND 0.32808f
C6586 D_FlipFlop_2.nPRE.n9 GND 0.03499f
C6587 D_FlipFlop_2.nPRE.t4 GND 0.16938f
C6588 D_FlipFlop_2.nPRE.n10 GND 0.04879f
C6589 D_FlipFlop_2.nPRE.n11 GND 0.01299f
C6590 D_FlipFlop_2.nPRE.n12 GND 0.02025f
C6591 D_FlipFlop_2.nPRE.n13 GND 0.20204f
C6592 D_FlipFlop_2.nPRE.t8 GND 0.32579f
C6593 D_FlipFlop_2.nPRE.n14 GND 0.32808f
C6594 D_FlipFlop_2.nPRE.n15 GND 0.03499f
C6595 D_FlipFlop_2.nPRE.t15 GND 0.16938f
C6596 D_FlipFlop_2.nPRE.n16 GND 0.04879f
C6597 D_FlipFlop_2.nPRE.n17 GND 0.01299f
C6598 D_FlipFlop_2.nPRE.n18 GND 0.02025f
C6599 D_FlipFlop_2.nPRE.n20 GND 0.52437f
C6600 D_FlipFlop_2.nPRE.n21 GND 0.62078f
C6601 D_FlipFlop_2.nPRE.n22 GND 0.86804f
C6602 D_FlipFlop_2.nPRE.t16 GND 0.16938f
C6603 D_FlipFlop_2.nPRE.n23 GND 0.04437f
C6604 D_FlipFlop_2.nPRE.n24 GND 0.0407f
C6605 D_FlipFlop_2.nPRE.t6 GND 0.32622f
C6606 D_FlipFlop_2.nPRE.n25 GND 0.09786f
C6607 D_FlipFlop_2.nPRE.t5 GND 0.16938f
C6608 D_FlipFlop_2.nPRE.n26 GND 0.04437f
C6609 D_FlipFlop_2.nPRE.n27 GND 0.0407f
C6610 D_FlipFlop_2.nPRE.n28 GND 0.10298f
C6611 D_FlipFlop_2.nPRE.n29 GND 0.10298f
C6612 D_FlipFlop_2.nPRE.n30 GND 0.09786f
C6613 D_FlipFlop_2.nPRE.t12 GND 0.41655f
C6614 D_FlipFlop_2.nPRE.n31 GND 0.10217f
C6615 D_FlipFlop_2.nPRE.n32 GND 0.28124f
C6616 D_FlipFlop_2.nPRE.n33 GND 0.20695f
C6617 D_FlipFlop_2.nPRE.t10 GND 0.32577f
C6618 D_FlipFlop_2.nPRE.n34 GND 0.14189f
C6619 D_FlipFlop_2.nPRE.t7 GND 0.15205f
C6620 D_FlipFlop_2.nPRE.n35 GND 0.09926f
C6621 D_FlipFlop_2.nPRE.n36 GND 0.04754f
C6622 D_FlipFlop_2.nPRE.n37 GND 0.12052f
C6623 D_FlipFlop_2.nPRE.t0 GND 0.04419f
C6624 D_FlipFlop_2.nPRE.n38 GND 0.06807f
C6625 D_FlipFlop_2.nPRE.t3 GND 0.04511f
C6626 D_FlipFlop_2.nPRE.t2 GND 0.04419f
C6627 D_FlipFlop_2.nPRE.n39 GND 0.25129f
C6628 D_FlipFlop_2.nPRE.n40 GND 0.082f
C6629 D_FlipFlop_2.nPRE.n41 GND 0.16509f
C6630 D_FlipFlop_5.CLK.t1 GND 0.02954f
C6631 D_FlipFlop_5.CLK.t6 GND 0.22695f
C6632 D_FlipFlop_5.CLK.t5 GND 0.118f
C6633 D_FlipFlop_5.CLK.n0 GND 0.12444f
C6634 D_FlipFlop_5.CLK.t7 GND 0.22695f
C6635 D_FlipFlop_5.CLK.n1 GND 0.2009f
C6636 D_FlipFlop_5.CLK.n2 GND 0.20145f
C6637 D_FlipFlop_5.CLK.n3 GND 0.12607f
C6638 D_FlipFlop_5.CLK.t4 GND 0.10447f
C6639 D_FlipFlop_5.CLK.n4 GND 0.02736f
C6640 D_FlipFlop_5.CLK.n5 GND 0.10371f
C6641 D_FlipFlop_5.CLK.t3 GND 0.10446f
C6642 D_FlipFlop_5.CLK.n6 GND 0.03399f
C6643 D_FlipFlop_5.CLK.n7 GND 0.02546f
C6644 D_FlipFlop_5.CLK.n8 GND 0.23531f
C6645 D_FlipFlop_5.CLK.t2 GND 0.21911f
C6646 D_FlipFlop_5.CLK.n9 GND 0.16025f
C6647 D_FlipFlop_5.CLK.n11 GND 0.03049f
C6648 D_FlipFlop_5.CLK.t0 GND 0.03086f
C6649 D_FlipFlop_5.CLK.n12 GND 0.19695f
C6650 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 GND 0.37675f
C6651 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 GND 0.16409f
C6652 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 GND 0.18888f
C6653 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 GND 0.0511f
C6654 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 GND 0.32168f
C6655 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 GND 0.05217f
C6656 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 GND 0.0511f
C6657 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 GND 0.29061f
C6658 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 GND 0.09483f
C6659 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 GND 0.01203f
C6660 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 GND 0.01587f
C6661 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 GND 0.37825f
C6662 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 GND 0.19588f
C6663 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 GND 0.28346f
C6664 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 GND 0.11199f
C6665 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 GND 0.05215f
C6666 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 GND 0.18008f
C6667 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t4 GND 0.47302f
C6668 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t3 GND 0.06145f
C6669 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n0 GND 0.15815f
C6670 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n1 GND 0.12861f
C6671 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t5 GND 0.24486f
C6672 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t6 GND 0.47095f
C6673 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n2 GND 0.11174f
C6674 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n3 GND 0.11082f
C6675 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n4 GND 0.18808f
C6676 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n5 GND 0.14f
C6677 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n6 GND 0.07837f
C6678 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t1 GND 0.06521f
C6679 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t2 GND 0.06388f
C6680 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n7 GND 0.36328f
C6681 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n8 GND 0.12591f
C6682 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t0 GND 0.06388f
C6683 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n9 GND 0.40291f
C6684 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.t7 GND 0.23439f
C6685 Ring_Counter_0.D_FlipFlop_13.3-input-nand_2.C.n10 GND 0.20386f
C6686 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 GND 0.37675f
C6687 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 GND 0.16409f
C6688 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 GND 0.18888f
C6689 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 GND 0.0511f
C6690 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 GND 0.32168f
C6691 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 GND 0.05217f
C6692 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 GND 0.0511f
C6693 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 GND 0.29061f
C6694 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 GND 0.09483f
C6695 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 GND 0.01203f
C6696 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 GND 0.01587f
C6697 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 GND 0.37825f
C6698 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 GND 0.19588f
C6699 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 GND 0.28346f
C6700 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 GND 0.11199f
C6701 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 GND 0.05215f
C6702 Ring_Counter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 GND 0.18008f
C6703 D_FlipFlop_3.nPRE.t3 GND 0.04395f
C6704 D_FlipFlop_3.nPRE.t13 GND 0.31207f
C6705 D_FlipFlop_3.nPRE.n0 GND 0.09117f
C6706 D_FlipFlop_3.nPRE.n1 GND 0.03956f
C6707 D_FlipFlop_3.nPRE.n2 GND 0.17392f
C6708 D_FlipFlop_3.nPRE.t12 GND 0.14514f
C6709 D_FlipFlop_3.nPRE.n3 GND 0.08328f
C6710 D_FlipFlop_3.nPRE.n4 GND 0.17653f
C6711 D_FlipFlop_3.nPRE.t8 GND 0.31209f
C6712 D_FlipFlop_3.nPRE.n5 GND 0.31429f
C6713 D_FlipFlop_3.nPRE.n6 GND 0.03352f
C6714 D_FlipFlop_3.nPRE.t10 GND 0.16226f
C6715 D_FlipFlop_3.nPRE.n7 GND 0.04674f
C6716 D_FlipFlop_3.nPRE.n8 GND 0.01245f
C6717 D_FlipFlop_3.nPRE.n9 GND 0.0194f
C6718 D_FlipFlop_3.nPRE.n10 GND 0.19354f
C6719 D_FlipFlop_3.nPRE.t6 GND 0.31209f
C6720 D_FlipFlop_3.nPRE.n11 GND 0.31429f
C6721 D_FlipFlop_3.nPRE.n12 GND 0.03352f
C6722 D_FlipFlop_3.nPRE.t9 GND 0.16226f
C6723 D_FlipFlop_3.nPRE.n13 GND 0.04674f
C6724 D_FlipFlop_3.nPRE.n14 GND 0.01245f
C6725 D_FlipFlop_3.nPRE.n15 GND 0.0194f
C6726 D_FlipFlop_3.nPRE.n17 GND 0.50232f
C6727 D_FlipFlop_3.nPRE.n18 GND 0.63858f
C6728 D_FlipFlop_3.nPRE.t17 GND 0.31207f
C6729 D_FlipFlop_3.nPRE.n19 GND 0.09117f
C6730 D_FlipFlop_3.nPRE.n20 GND 0.03956f
C6731 D_FlipFlop_3.nPRE.n21 GND 0.17392f
C6732 D_FlipFlop_3.nPRE.t16 GND 0.14671f
C6733 D_FlipFlop_3.nPRE.n22 GND 0.9087f
C6734 D_FlipFlop_3.nPRE.t15 GND 0.16226f
C6735 D_FlipFlop_3.nPRE.n23 GND 0.04251f
C6736 D_FlipFlop_3.nPRE.n24 GND 0.03898f
C6737 D_FlipFlop_3.nPRE.t7 GND 0.3125f
C6738 D_FlipFlop_3.nPRE.n25 GND 0.09374f
C6739 D_FlipFlop_3.nPRE.t4 GND 0.16226f
C6740 D_FlipFlop_3.nPRE.n26 GND 0.04251f
C6741 D_FlipFlop_3.nPRE.n27 GND 0.03898f
C6742 D_FlipFlop_3.nPRE.n28 GND 0.09865f
C6743 D_FlipFlop_3.nPRE.n29 GND 0.09865f
C6744 D_FlipFlop_3.nPRE.n30 GND 0.09374f
C6745 D_FlipFlop_3.nPRE.t14 GND 0.39904f
C6746 D_FlipFlop_3.nPRE.n31 GND 0.09787f
C6747 D_FlipFlop_3.nPRE.n32 GND 0.26129f
C6748 D_FlipFlop_3.nPRE.n33 GND 0.19825f
C6749 D_FlipFlop_3.nPRE.t11 GND 0.31207f
C6750 D_FlipFlop_3.nPRE.n34 GND 0.13593f
C6751 D_FlipFlop_3.nPRE.t5 GND 0.14566f
C6752 D_FlipFlop_3.nPRE.n35 GND 0.09508f
C6753 D_FlipFlop_3.nPRE.n36 GND 0.04554f
C6754 D_FlipFlop_3.nPRE.n37 GND 0.11546f
C6755 D_FlipFlop_3.nPRE.t2 GND 0.04233f
C6756 D_FlipFlop_3.nPRE.n38 GND 0.0652f
C6757 D_FlipFlop_3.nPRE.t1 GND 0.04321f
C6758 D_FlipFlop_3.nPRE.t0 GND 0.04233f
C6759 D_FlipFlop_3.nPRE.n39 GND 0.24073f
C6760 D_FlipFlop_3.nPRE.n40 GND 0.07855f
C6761 D_FlipFlop_3.nPRE.n41 GND 0.15815f
C6762 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 GND 0.06443f
C6763 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 GND 0.14002f
C6764 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 GND 0.07316f
C6765 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 GND 0.25702f
C6766 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 GND 0.12462f
C6767 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 GND 0.4938f
C6768 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 GND 0.09136f
C6769 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 GND 0.05451f
C6770 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 GND 0.13379f
C6771 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 GND 0.13379f
C6772 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 GND 0.06713f
C6773 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 GND 0.07989f
C6774 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 GND 0.43786f
C6775 Ring_Counter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 GND 0.08018f
C6776 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t1 GND 0.05f
C6777 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n0 GND 0.10867f
C6778 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n1 GND 0.05678f
C6779 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t5 GND 0.38491f
C6780 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n2 GND 0.16589f
C6781 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t4 GND 0.30131f
C6782 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t3 GND 0.30153f
C6783 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n3 GND 0.09671f
C6784 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t2 GND 0.38323f
C6785 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n4 GND 0.0709f
C6786 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n5 GND 0.04231f
C6787 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n6 GND 0.10383f
C6788 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n7 GND 0.10383f
C6789 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.t0 GND 0.05284f
C6790 Ring_Counter_0.D_FlipFlop_4.Inverter_1.Vout.n8 GND 0.17757f
C6791 D_FlipFlop_7.D.t9 GND 0.24193f
C6792 D_FlipFlop_0.Inverter_0.Vin GND -0.21921f
C6793 D_FlipFlop_7.D.n0 GND 0.23325f
C6794 D_FlipFlop_7.D.n1 GND 0.02599f
C6795 D_FlipFlop_7.D.t30 GND 0.24193f
C6796 D_FlipFlop_7.Inverter_0.Vin GND -0.21921f
C6797 D_FlipFlop_7.D.n2 GND 0.23325f
C6798 D_FlipFlop_7.D.n3 GND 0.02599f
C6799 D_FlipFlop_7.D.t10 GND 0.12578f
C6800 D_FlipFlop_7.D.n4 GND 0.03623f
C6801 D_FlipFlop_7.D.n5 GND 0.01553f
C6802 D_FlipFlop_7.D.n6 GND 0.02909f
C6803 D_FlipFlop_7.D.t23 GND 0.24193f
C6804 D_FlipFlop_7.3-input-nand_0.B GND -0.17613f
C6805 D_FlipFlop_7.D.n7 GND 0.23776f
C6806 D_FlipFlop_7.D.n8 GND 0.02599f
C6807 D_FlipFlop_7.D.t15 GND 0.12578f
C6808 D_FlipFlop_7.D.n9 GND 0.03623f
C6809 D_FlipFlop_7.D.n10 GND 0.01553f
C6810 D_FlipFlop_7.D.n11 GND 0.02909f
C6811 D_FlipFlop_7.D.n12 GND 0.07647f
C6812 D_FlipFlop_7.D.n13 GND 0.07647f
C6813 D_FlipFlop_7.D.n14 GND 0.01888f
C6814 D_FlipFlop_7.D.n15 GND 0.02679f
C6815 D_FlipFlop_7.D.n16 GND 0.36101f
C6816 D_FlipFlop_7.D.t5 GND 0.24193f
C6817 D_FlipFlop_6.Inverter_0.Vin GND -0.21921f
C6818 D_FlipFlop_7.D.n17 GND 0.23325f
C6819 D_FlipFlop_7.D.n18 GND 0.02599f
C6820 D_FlipFlop_7.D.t28 GND 0.12578f
C6821 D_FlipFlop_7.D.n19 GND 0.03623f
C6822 D_FlipFlop_7.D.n20 GND 0.01553f
C6823 D_FlipFlop_7.D.n21 GND 0.02909f
C6824 D_FlipFlop_7.D.t11 GND 0.24193f
C6825 D_FlipFlop_6.3-input-nand_0.B GND -0.17613f
C6826 D_FlipFlop_7.D.n22 GND 0.23776f
C6827 D_FlipFlop_7.D.n23 GND 0.02599f
C6828 D_FlipFlop_7.D.t22 GND 0.12578f
C6829 D_FlipFlop_7.D.n24 GND 0.03623f
C6830 D_FlipFlop_7.D.n25 GND 0.01553f
C6831 D_FlipFlop_7.D.n26 GND 0.02909f
C6832 D_FlipFlop_7.D.n27 GND 0.07647f
C6833 D_FlipFlop_7.D.n28 GND 0.07647f
C6834 D_FlipFlop_7.D.n29 GND 0.01888f
C6835 D_FlipFlop_7.D.n30 GND 0.02679f
C6836 D_FlipFlop_7.D.n32 GND 0.92838f
C6837 D_FlipFlop_7.D.t24 GND 0.24193f
C6838 D_FlipFlop_4.Inverter_0.Vin GND -0.21921f
C6839 D_FlipFlop_7.D.n33 GND 0.23325f
C6840 D_FlipFlop_7.D.n34 GND 0.02599f
C6841 D_FlipFlop_7.D.t33 GND 0.12578f
C6842 D_FlipFlop_7.D.n35 GND 0.03623f
C6843 D_FlipFlop_7.D.n36 GND 0.01553f
C6844 D_FlipFlop_7.D.n37 GND 0.02909f
C6845 D_FlipFlop_7.D.t31 GND 0.24193f
C6846 D_FlipFlop_4.3-input-nand_0.B GND -0.17613f
C6847 D_FlipFlop_7.D.n38 GND 0.23776f
C6848 D_FlipFlop_7.D.n39 GND 0.02599f
C6849 D_FlipFlop_7.D.t14 GND 0.12578f
C6850 D_FlipFlop_7.D.n40 GND 0.03623f
C6851 D_FlipFlop_7.D.n41 GND 0.01553f
C6852 D_FlipFlop_7.D.n42 GND 0.02909f
C6853 D_FlipFlop_7.D.n43 GND 0.07647f
C6854 D_FlipFlop_7.D.n44 GND 0.07647f
C6855 D_FlipFlop_7.D.n45 GND 0.01888f
C6856 D_FlipFlop_7.D.n46 GND 0.02679f
C6857 D_FlipFlop_7.D.n48 GND 0.86083f
C6858 D_FlipFlop_7.D.t6 GND 0.24193f
C6859 D_FlipFlop_5.Inverter_0.Vin GND -0.21921f
C6860 D_FlipFlop_7.D.n49 GND 0.23325f
C6861 D_FlipFlop_7.D.n50 GND 0.02599f
C6862 D_FlipFlop_7.D.t20 GND 0.12578f
C6863 D_FlipFlop_7.D.n51 GND 0.03623f
C6864 D_FlipFlop_7.D.n52 GND 0.01553f
C6865 D_FlipFlop_7.D.n53 GND 0.02909f
C6866 D_FlipFlop_7.D.t17 GND 0.24193f
C6867 D_FlipFlop_5.3-input-nand_0.B GND -0.17613f
C6868 D_FlipFlop_7.D.n54 GND 0.23776f
C6869 D_FlipFlop_7.D.n55 GND 0.02599f
C6870 D_FlipFlop_7.D.t12 GND 0.12578f
C6871 D_FlipFlop_7.D.n56 GND 0.03623f
C6872 D_FlipFlop_7.D.n57 GND 0.01553f
C6873 D_FlipFlop_7.D.n58 GND 0.02909f
C6874 D_FlipFlop_7.D.n59 GND 0.07647f
C6875 D_FlipFlop_7.D.n60 GND 0.07647f
C6876 D_FlipFlop_7.D.n61 GND 0.01888f
C6877 D_FlipFlop_7.D.n62 GND 0.02679f
C6878 D_FlipFlop_7.D.n64 GND 0.86083f
C6879 D_FlipFlop_7.D.t32 GND 0.24193f
C6880 D_FlipFlop_3.Inverter_0.Vin GND -0.21921f
C6881 D_FlipFlop_7.D.n65 GND 0.23325f
C6882 D_FlipFlop_7.D.n66 GND 0.02599f
C6883 D_FlipFlop_7.D.t3 GND 0.12578f
C6884 D_FlipFlop_7.D.n67 GND 0.03623f
C6885 D_FlipFlop_7.D.n68 GND 0.01553f
C6886 D_FlipFlop_7.D.n69 GND 0.02909f
C6887 D_FlipFlop_7.D.t25 GND 0.24193f
C6888 D_FlipFlop_3.3-input-nand_0.B GND -0.17613f
C6889 D_FlipFlop_7.D.n70 GND 0.23776f
C6890 D_FlipFlop_7.D.n71 GND 0.02599f
C6891 D_FlipFlop_7.D.t4 GND 0.12578f
C6892 D_FlipFlop_7.D.n72 GND 0.03623f
C6893 D_FlipFlop_7.D.n73 GND 0.01553f
C6894 D_FlipFlop_7.D.n74 GND 0.02909f
C6895 D_FlipFlop_7.D.n75 GND 0.07647f
C6896 D_FlipFlop_7.D.n76 GND 0.07647f
C6897 D_FlipFlop_7.D.n77 GND 0.01888f
C6898 D_FlipFlop_7.D.n78 GND 0.02679f
C6899 D_FlipFlop_7.D.n80 GND 0.86083f
C6900 D_FlipFlop_7.D.t13 GND 0.24193f
C6901 D_FlipFlop_2.Inverter_0.Vin GND -0.21921f
C6902 D_FlipFlop_7.D.n81 GND 0.23325f
C6903 D_FlipFlop_7.D.n82 GND 0.02599f
C6904 D_FlipFlop_7.D.t27 GND 0.12578f
C6905 D_FlipFlop_7.D.n83 GND 0.03623f
C6906 D_FlipFlop_7.D.n84 GND 0.01553f
C6907 D_FlipFlop_7.D.n85 GND 0.02909f
C6908 D_FlipFlop_7.D.t19 GND 0.24193f
C6909 D_FlipFlop_2.3-input-nand_0.B GND -0.17613f
C6910 D_FlipFlop_7.D.n86 GND 0.23776f
C6911 D_FlipFlop_7.D.n87 GND 0.02599f
C6912 D_FlipFlop_7.D.t35 GND 0.12578f
C6913 D_FlipFlop_7.D.n88 GND 0.03623f
C6914 D_FlipFlop_7.D.n89 GND 0.01553f
C6915 D_FlipFlop_7.D.n90 GND 0.02909f
C6916 D_FlipFlop_7.D.n91 GND 0.07647f
C6917 D_FlipFlop_7.D.n92 GND 0.07647f
C6918 D_FlipFlop_7.D.n93 GND 0.01888f
C6919 D_FlipFlop_7.D.n94 GND 0.02679f
C6920 D_FlipFlop_7.D.n96 GND 0.86083f
C6921 D_FlipFlop_7.D.t7 GND 0.24193f
C6922 D_FlipFlop_1.Inverter_0.Vin GND -0.21921f
C6923 D_FlipFlop_7.D.n97 GND 0.23325f
C6924 D_FlipFlop_7.D.n98 GND 0.02599f
C6925 D_FlipFlop_7.D.t21 GND 0.12578f
C6926 D_FlipFlop_7.D.n99 GND 0.03623f
C6927 D_FlipFlop_7.D.n100 GND 0.01553f
C6928 D_FlipFlop_7.D.n101 GND 0.02909f
C6929 D_FlipFlop_7.D.t34 GND 0.24193f
C6930 D_FlipFlop_1.3-input-nand_0.B GND -0.17613f
C6931 D_FlipFlop_7.D.n102 GND 0.23776f
C6932 D_FlipFlop_7.D.n103 GND 0.02599f
C6933 D_FlipFlop_7.D.t16 GND 0.12578f
C6934 D_FlipFlop_7.D.n104 GND 0.03623f
C6935 D_FlipFlop_7.D.n105 GND 0.01553f
C6936 D_FlipFlop_7.D.n106 GND 0.02909f
C6937 D_FlipFlop_7.D.n107 GND 0.07647f
C6938 D_FlipFlop_7.D.n108 GND 0.07647f
C6939 D_FlipFlop_7.D.n109 GND 0.01888f
C6940 D_FlipFlop_7.D.n110 GND 0.02679f
C6941 D_FlipFlop_7.D.n112 GND 0.92838f
C6942 D_FlipFlop_7.D.n113 GND 0.36101f
C6943 D_FlipFlop_7.D.n114 GND 0.02679f
C6944 D_FlipFlop_7.D.n115 GND 0.01888f
C6945 D_FlipFlop_7.D.t26 GND 0.24193f
C6946 D_FlipFlop_0.3-input-nand_0.B GND -0.17613f
C6947 D_FlipFlop_7.D.n116 GND 0.23776f
C6948 D_FlipFlop_7.D.n117 GND 0.02599f
C6949 D_FlipFlop_7.D.t8 GND 0.12578f
C6950 D_FlipFlop_7.D.n118 GND 0.03623f
C6951 D_FlipFlop_7.D.n119 GND 0.01553f
C6952 D_FlipFlop_7.D.n120 GND 0.02909f
C6953 D_FlipFlop_7.D.n121 GND 0.07647f
C6954 D_FlipFlop_7.D.n122 GND 0.07647f
C6955 D_FlipFlop_7.D.n123 GND 0.02909f
C6956 D_FlipFlop_7.D.n124 GND 0.01553f
C6957 D_FlipFlop_7.D.t1 GND 3.02085f
C6958 D_FlipFlop_7.D.t0 GND 0.70735f
C6959 Comparator_0.Vout GND 0.11269f
C6960 D_FlipFlop_7.D.t29 GND 0.91151f
C6961 D_FlipFlop_7.D.n125 GND 0.26608f
C6962 D_FlipFlop_7.D.n126 GND 1.88431f
C6963 D_FlipFlop_7.D.t2 GND 1.9676f
C6964 D_FlipFlop_7.D.n127 GND 2.53644f
C6965 D_FlipFlop_7.D.n128 GND 1.88054f
C6966 D_FlipFlop_7.D.n129 GND 3.37696f
C6967 D_FlipFlop_7.D.t18 GND 0.32617f
C6968 D_FlipFlop_7.D.n130 GND 0.03623f
C6969 D_FlipFlop_6.CLK.t1 GND 0.02954f
C6970 D_FlipFlop_6.CLK.t6 GND 0.22695f
C6971 D_FlipFlop_6.CLK.t5 GND 0.118f
C6972 D_FlipFlop_6.CLK.n0 GND 0.12444f
C6973 D_FlipFlop_6.CLK.t3 GND 0.22695f
C6974 D_FlipFlop_6.CLK.n1 GND 0.2009f
C6975 D_FlipFlop_6.CLK.n2 GND 0.20145f
C6976 D_FlipFlop_6.CLK.n3 GND 0.12607f
C6977 D_FlipFlop_6.CLK.t2 GND 0.10447f
C6978 D_FlipFlop_6.CLK.n4 GND 0.02736f
C6979 D_FlipFlop_6.CLK.n5 GND 0.10371f
C6980 D_FlipFlop_6.CLK.t7 GND 0.10446f
C6981 D_FlipFlop_6.CLK.n6 GND 0.03399f
C6982 D_FlipFlop_6.CLK.n7 GND 0.02546f
C6983 D_FlipFlop_6.CLK.n8 GND 0.23531f
C6984 D_FlipFlop_6.CLK.t4 GND 0.21911f
C6985 D_FlipFlop_6.CLK.n9 GND 0.16025f
C6986 D_FlipFlop_6.CLK.n11 GND 0.03049f
C6987 D_FlipFlop_6.CLK.t0 GND 0.03086f
C6988 D_FlipFlop_6.CLK.n12 GND 0.19695f
C6989 Nand_Gate_6.A.t1 GND 0.03519f
C6990 Nand_Gate_6.A.t6 GND 0.24981f
C6991 Nand_Gate_6.A.n0 GND 0.07298f
C6992 Nand_Gate_6.A.n1 GND 0.03166f
C6993 Nand_Gate_6.A.n2 GND 0.13922f
C6994 Nand_Gate_6.A.t10 GND 0.12848f
C6995 Nand_Gate_6.A.t9 GND 0.12988f
C6996 Nand_Gate_6.A.n3 GND 0.03403f
C6997 Nand_Gate_6.A.n4 GND 0.03121f
C6998 Nand_Gate_6.A.t4 GND 0.25015f
C6999 Nand_Gate_6.A.n5 GND 0.07504f
C7000 Nand_Gate_6.A.t11 GND 0.12988f
C7001 Nand_Gate_6.A.n6 GND 0.03403f
C7002 Nand_Gate_6.A.n7 GND 0.03121f
C7003 Nand_Gate_6.A.n8 GND 0.07897f
C7004 Nand_Gate_6.A.n9 GND 0.07897f
C7005 Nand_Gate_6.A.n10 GND 0.07504f
C7006 Nand_Gate_6.A.t8 GND 0.31943f
C7007 Nand_Gate_6.A.n11 GND 0.07835f
C7008 Nand_Gate_6.A.n12 GND 0.55804f
C7009 Nand_Gate_6.A.n13 GND 0.1587f
C7010 Nand_Gate_6.A.t7 GND 0.24981f
C7011 Nand_Gate_6.A.n14 GND 0.10881f
C7012 Nand_Gate_6.A.t5 GND 0.1166f
C7013 Nand_Gate_6.A.n15 GND 0.07611f
C7014 Nand_Gate_6.A.n16 GND 0.03645f
C7015 Nand_Gate_6.A.n17 GND 0.09242f
C7016 Nand_Gate_6.A.t0 GND 0.03388f
C7017 Nand_Gate_6.A.n18 GND 0.0522f
C7018 Nand_Gate_6.A.t3 GND 0.03459f
C7019 Nand_Gate_6.A.t2 GND 0.03388f
C7020 Nand_Gate_6.A.n19 GND 0.1927f
C7021 Nand_Gate_6.A.n20 GND 0.06288f
C7022 Nand_Gate_6.A.n21 GND 0.1266f
C7023 a_51632_31172.t2 GND 1.56705f
C7024 a_51632_31172.t3 GND 2.25506f
C7025 a_51632_31172.t1 GND 2.25426f
C7026 a_51632_31172.n0 GND 1.45916f
C7027 a_51632_31172.n1 GND 0.92425f
C7028 a_51632_31172.t0 GND 0.74021f
C7029 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t2 GND 0.06145f
C7030 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n0 GND 0.15815f
C7031 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n1 GND 0.12861f
C7032 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t6 GND 0.24486f
C7033 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t7 GND 0.47095f
C7034 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n2 GND 0.11174f
C7035 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n3 GND 0.11082f
C7036 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n4 GND 0.18808f
C7037 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n5 GND 0.14f
C7038 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t4 GND 0.47302f
C7039 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n6 GND 0.20386f
C7040 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t5 GND 0.23439f
C7041 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t3 GND 0.06388f
C7042 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n7 GND 0.40291f
C7043 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t0 GND 0.06521f
C7044 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.t1 GND 0.06388f
C7045 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n8 GND 0.36328f
C7046 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n9 GND 0.12591f
C7047 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.C.n10 GND 0.07837f
C7048 D_FlipFlop_2.CLK.t1 GND 0.02954f
C7049 D_FlipFlop_2.CLK.t2 GND 0.22695f
C7050 D_FlipFlop_2.CLK.t4 GND 0.118f
C7051 D_FlipFlop_2.CLK.n0 GND 0.12444f
C7052 D_FlipFlop_2.CLK.t7 GND 0.22695f
C7053 D_FlipFlop_2.CLK.n1 GND 0.2009f
C7054 D_FlipFlop_2.CLK.n2 GND 0.20145f
C7055 D_FlipFlop_2.CLK.n3 GND 0.12607f
C7056 D_FlipFlop_2.CLK.t6 GND 0.10447f
C7057 D_FlipFlop_2.CLK.n4 GND 0.02736f
C7058 D_FlipFlop_2.CLK.n5 GND 0.10371f
C7059 D_FlipFlop_2.CLK.t5 GND 0.10446f
C7060 D_FlipFlop_2.CLK.n6 GND 0.03399f
C7061 D_FlipFlop_2.CLK.n7 GND 0.02546f
C7062 D_FlipFlop_2.CLK.n8 GND 0.23531f
C7063 D_FlipFlop_2.CLK.t3 GND 0.21911f
C7064 D_FlipFlop_2.CLK.n9 GND 0.16025f
C7065 D_FlipFlop_2.CLK.n11 GND 0.03049f
C7066 D_FlipFlop_2.CLK.t0 GND 0.03086f
C7067 D_FlipFlop_2.CLK.n12 GND 0.19695f
C7068 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 GND 0.05029f
C7069 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 GND 0.17365f
C7070 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 GND 0.36474f
C7071 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 GND 0.18889f
C7072 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 GND 0.27334f
C7073 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 GND 0.10799f
C7074 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 GND 0.0153f
C7075 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 GND 0.36329f
C7076 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 GND 0.15823f
C7077 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 GND 0.18214f
C7078 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 GND 0.04928f
C7079 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 GND 0.31019f
C7080 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 GND 0.05031f
C7081 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 GND 0.04928f
C7082 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 GND 0.28023f
C7083 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 GND 0.09144f
C7084 Ring_Counter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 GND 0.0116f
C7085 CDAC_v3_0.switch_5.Z.t1 GND 0.05033f
C7086 CDAC_v3_0.switch_5.Z.t2 GND 0.05033f
C7087 CDAC_v3_0.switch_5.Z.n0 GND 0.18079f
C7088 CDAC_v3_0.switch_5.Z.n1 GND 0.55739f
C7089 CDAC_v3_0.switch_5.Z.n2 GND 0.05215f
C7090 CDAC_v3_0.switch_5.Z.t33 GND 6.60385f
C7091 CDAC_v3_0.switch_5.Z.t25 GND 6.60385f
C7092 CDAC_v3_0.switch_5.Z.t20 GND 6.60385f
C7093 CDAC_v3_0.switch_5.Z.t5 GND 6.60385f
C7094 CDAC_v3_0.switch_5.Z.t8 GND 6.60385f
C7095 CDAC_v3_0.switch_5.Z.t31 GND 6.60385f
C7096 CDAC_v3_0.switch_5.Z.t12 GND 6.60385f
C7097 CDAC_v3_0.switch_5.Z.t34 GND 7.23284f
C7098 CDAC_v3_0.switch_5.Z.n3 GND 1.13605f
C7099 CDAC_v3_0.switch_5.Z.n4 GND 1.08536f
C7100 CDAC_v3_0.switch_5.Z.n5 GND 1.08536f
C7101 CDAC_v3_0.switch_5.Z.n6 GND 1.08536f
C7102 CDAC_v3_0.switch_5.Z.n7 GND 1.08536f
C7103 CDAC_v3_0.switch_5.Z.n8 GND 1.08536f
C7104 CDAC_v3_0.switch_5.Z.n9 GND 1.79745f
C7105 CDAC_v3_0.switch_5.Z.t29 GND 6.60385f
C7106 CDAC_v3_0.switch_5.Z.t11 GND 6.60385f
C7107 CDAC_v3_0.switch_5.Z.t15 GND 6.60385f
C7108 CDAC_v3_0.switch_5.Z.t9 GND 6.60385f
C7109 CDAC_v3_0.switch_5.Z.t7 GND 6.60385f
C7110 CDAC_v3_0.switch_5.Z.t13 GND 6.60385f
C7111 CDAC_v3_0.switch_5.Z.t32 GND 6.60385f
C7112 CDAC_v3_0.switch_5.Z.t22 GND 7.23284f
C7113 CDAC_v3_0.switch_5.Z.n10 GND 1.13605f
C7114 CDAC_v3_0.switch_5.Z.n11 GND 1.08536f
C7115 CDAC_v3_0.switch_5.Z.n12 GND 1.08536f
C7116 CDAC_v3_0.switch_5.Z.n13 GND 1.08536f
C7117 CDAC_v3_0.switch_5.Z.n14 GND 1.08536f
C7118 CDAC_v3_0.switch_5.Z.n15 GND 1.08536f
C7119 CDAC_v3_0.switch_5.Z.n16 GND 1.52631f
C7120 CDAC_v3_0.switch_5.Z.n17 GND 3.43598f
C7121 CDAC_v3_0.switch_5.Z.t26 GND 6.60385f
C7122 CDAC_v3_0.switch_5.Z.t27 GND 6.60385f
C7123 CDAC_v3_0.switch_5.Z.t17 GND 6.60385f
C7124 CDAC_v3_0.switch_5.Z.t19 GND 6.60385f
C7125 CDAC_v3_0.switch_5.Z.t6 GND 6.60385f
C7126 CDAC_v3_0.switch_5.Z.t14 GND 6.60385f
C7127 CDAC_v3_0.switch_5.Z.t35 GND 6.60385f
C7128 CDAC_v3_0.switch_5.Z.t16 GND 7.80268f
C7129 CDAC_v3_0.switch_5.Z.n18 GND 1.18198f
C7130 CDAC_v3_0.switch_5.Z.n19 GND 1.08536f
C7131 CDAC_v3_0.switch_5.Z.n20 GND 1.08536f
C7132 CDAC_v3_0.switch_5.Z.n21 GND 1.08536f
C7133 CDAC_v3_0.switch_5.Z.n22 GND 1.08536f
C7134 CDAC_v3_0.switch_5.Z.n23 GND 1.08536f
C7135 CDAC_v3_0.switch_5.Z.n24 GND 1.15346f
C7136 CDAC_v3_0.switch_5.Z.n25 GND 2.57703f
C7137 CDAC_v3_0.switch_5.Z.t28 GND 6.60385f
C7138 CDAC_v3_0.switch_5.Z.t30 GND 6.60385f
C7139 CDAC_v3_0.switch_5.Z.t23 GND 6.60385f
C7140 CDAC_v3_0.switch_5.Z.t24 GND 6.60385f
C7141 CDAC_v3_0.switch_5.Z.t10 GND 6.60385f
C7142 CDAC_v3_0.switch_5.Z.t18 GND 6.60385f
C7143 CDAC_v3_0.switch_5.Z.t4 GND 6.60385f
C7144 CDAC_v3_0.switch_5.Z.t21 GND 7.80268f
C7145 CDAC_v3_0.switch_5.Z.n26 GND 1.18198f
C7146 CDAC_v3_0.switch_5.Z.n27 GND 1.08536f
C7147 CDAC_v3_0.switch_5.Z.n28 GND 1.08536f
C7148 CDAC_v3_0.switch_5.Z.n29 GND 1.08536f
C7149 CDAC_v3_0.switch_5.Z.n30 GND 1.08536f
C7150 CDAC_v3_0.switch_5.Z.n31 GND 1.08536f
C7151 CDAC_v3_0.switch_5.Z.n32 GND 1.15346f
C7152 CDAC_v3_0.switch_5.Z.n33 GND 4.04925f
C7153 CDAC_v3_0.switch_5.Z.n34 GND 1.68696f
C7154 CDAC_v3_0.switch_5.Z.n35 GND 0.01656f
C7155 CDAC_v3_0.switch_5.Z.t0 GND 0.04875f
C7156 CDAC_v3_0.switch_5.Z.n36 GND 0.10705f
C7157 CDAC_v3_0.switch_5.Z.t3 GND 0.04865f
C7158 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 GND 0.06443f
C7159 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 GND 0.14002f
C7160 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 GND 0.07316f
C7161 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 GND 0.25702f
C7162 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 GND 0.12462f
C7163 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 GND 0.4938f
C7164 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 GND 0.09136f
C7165 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 GND 0.05451f
C7166 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 GND 0.13379f
C7167 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 GND 0.13379f
C7168 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 GND 0.06713f
C7169 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 GND 0.07989f
C7170 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 GND 0.43786f
C7171 Ring_Counter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 GND 0.08018f
C7172 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 GND 0.06443f
C7173 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 GND 0.14002f
C7174 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 GND 0.07316f
C7175 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 GND 0.25702f
C7176 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 GND 0.12462f
C7177 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 GND 0.4938f
C7178 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 GND 0.09136f
C7179 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 GND 0.05451f
C7180 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 GND 0.13379f
C7181 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 GND 0.13379f
C7182 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 GND 0.06713f
C7183 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 GND 0.07989f
C7184 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 GND 0.43786f
C7185 Ring_Counter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 GND 0.08018f
C7186 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t1 GND 0.05f
C7187 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n0 GND 0.10867f
C7188 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n1 GND 0.05678f
C7189 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t5 GND 0.38491f
C7190 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n2 GND 0.16589f
C7191 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t3 GND 0.30131f
C7192 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t4 GND 0.30153f
C7193 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n3 GND 0.09671f
C7194 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t2 GND 0.38323f
C7195 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n4 GND 0.0709f
C7196 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n5 GND 0.04231f
C7197 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n6 GND 0.10383f
C7198 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n7 GND 0.10383f
C7199 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.t0 GND 0.05284f
C7200 Ring_Counter_0.D_FlipFlop_12.Inverter_1.Vout.n8 GND 0.17757f
C7201 FFCLR.t3 GND 0.06306f
C7202 Nand_Gate_7.B GND -0.12174f
C7203 FFCLR.t35 GND 0.44775f
C7204 FFCLR.n0 GND 0.1308f
C7205 FFCLR.n1 GND 0.05675f
C7206 FFCLR.n2 GND 0.24953f
C7207 FFCLR.t32 GND 0.22375f
C7208 D_FlipFlop_0.3-input-nand_1.A GND -0.12174f
C7209 FFCLR.t4 GND 0.44775f
C7210 FFCLR.n3 GND 0.1308f
C7211 FFCLR.n4 GND 0.05675f
C7212 FFCLR.n5 GND 0.24953f
C7213 FFCLR.t54 GND 0.20824f
C7214 D_FlipFlop_0.nPRE GND -0.07257f
C7215 FFCLR.n6 GND 0.03766f
C7216 FFCLR.n7 GND 0.08143f
C7217 FFCLR.t26 GND 0.44777f
C7218 D_FlipFlop_7.3-input-nand_0.A GND -0.2662f
C7219 FFCLR.n8 GND 0.46425f
C7220 FFCLR.n9 GND 0.05023f
C7221 FFCLR.n10 GND 0.06706f
C7222 FFCLR.t25 GND 0.20914f
C7223 D_FlipFlop_7.nCLR GND -0.24492f
C7224 FFCLR.n11 GND 0.31064f
C7225 FFCLR.n12 GND 0.12314f
C7226 FFCLR.t34 GND 0.2328f
C7227 D_FlipFlop_7.3-input-nand_5.A GND -0.20104f
C7228 FFCLR.n13 GND 0.21717f
C7229 FFCLR.n14 GND 0.0481f
C7230 FFCLR.t49 GND 0.44775f
C7231 FFCLR.n15 GND 0.1308f
C7232 FFCLR.n16 GND 0.04343f
C7233 FFCLR.n17 GND 0.07336f
C7234 FFCLR.n18 GND 0.27768f
C7235 FFCLR.t57 GND 0.2328f
C7236 D_FlipFlop_7.3-input-nand_3.A GND -0.20104f
C7237 FFCLR.n19 GND 0.21717f
C7238 FFCLR.n20 GND 0.0481f
C7239 FFCLR.t11 GND 0.44775f
C7240 FFCLR.n21 GND 0.1308f
C7241 FFCLR.n22 GND 0.04343f
C7242 FFCLR.n23 GND 0.07336f
C7243 FFCLR.n25 GND 0.7054f
C7244 FFCLR.n26 GND 0.10317f
C7245 FFCLR.n27 GND 0.219f
C7246 FFCLR.n28 GND 0.71616f
C7247 FFCLR.t18 GND 0.44777f
C7248 D_FlipFlop_6.3-input-nand_0.A GND -0.2662f
C7249 FFCLR.n29 GND 0.46425f
C7250 FFCLR.n30 GND 0.05023f
C7251 FFCLR.n31 GND 0.06706f
C7252 FFCLR.t38 GND 0.20914f
C7253 D_FlipFlop_6.nCLR GND -0.24492f
C7254 FFCLR.n32 GND 0.31064f
C7255 FFCLR.n33 GND 0.12314f
C7256 FFCLR.t10 GND 0.2328f
C7257 D_FlipFlop_6.3-input-nand_5.A GND -0.20104f
C7258 FFCLR.n34 GND 0.21717f
C7259 FFCLR.n35 GND 0.0481f
C7260 FFCLR.t33 GND 0.44775f
C7261 FFCLR.n36 GND 0.1308f
C7262 FFCLR.n37 GND 0.04343f
C7263 FFCLR.n38 GND 0.07336f
C7264 FFCLR.n39 GND 0.27768f
C7265 FFCLR.t29 GND 0.2328f
C7266 D_FlipFlop_6.3-input-nand_3.A GND -0.20104f
C7267 FFCLR.n40 GND 0.21717f
C7268 FFCLR.n41 GND 0.0481f
C7269 FFCLR.t44 GND 0.44775f
C7270 FFCLR.n42 GND 0.1308f
C7271 FFCLR.n43 GND 0.04343f
C7272 FFCLR.n44 GND 0.07336f
C7273 FFCLR.n46 GND 0.7054f
C7274 FFCLR.n47 GND 0.10317f
C7275 FFCLR.n48 GND 0.219f
C7276 FFCLR.n50 GND 1.69854f
C7277 FFCLR.t59 GND 0.44777f
C7278 D_FlipFlop_4.3-input-nand_0.A GND -0.2662f
C7279 FFCLR.n51 GND 0.46425f
C7280 FFCLR.n52 GND 0.05023f
C7281 FFCLR.n53 GND 0.06706f
C7282 FFCLR.t28 GND 0.20914f
C7283 D_FlipFlop_4.nCLR GND -0.24492f
C7284 FFCLR.n54 GND 0.31064f
C7285 FFCLR.n55 GND 0.12314f
C7286 FFCLR.t30 GND 0.2328f
C7287 D_FlipFlop_4.3-input-nand_5.A GND -0.20104f
C7288 FFCLR.n56 GND 0.21717f
C7289 FFCLR.n57 GND 0.0481f
C7290 FFCLR.t52 GND 0.44775f
C7291 FFCLR.n58 GND 0.1308f
C7292 FFCLR.n59 GND 0.04343f
C7293 FFCLR.n60 GND 0.07336f
C7294 FFCLR.n61 GND 0.27768f
C7295 FFCLR.t17 GND 0.2328f
C7296 D_FlipFlop_4.3-input-nand_3.A GND -0.20104f
C7297 FFCLR.n62 GND 0.21717f
C7298 FFCLR.n63 GND 0.0481f
C7299 FFCLR.t43 GND 0.44775f
C7300 FFCLR.n64 GND 0.1308f
C7301 FFCLR.n65 GND 0.04343f
C7302 FFCLR.n66 GND 0.07336f
C7303 FFCLR.n68 GND 0.7054f
C7304 FFCLR.n69 GND 0.10317f
C7305 FFCLR.n70 GND 0.219f
C7306 FFCLR.n72 GND 1.59688f
C7307 FFCLR.t15 GND 0.44777f
C7308 D_FlipFlop_5.3-input-nand_0.A GND -0.2662f
C7309 FFCLR.n73 GND 0.46425f
C7310 FFCLR.n74 GND 0.05023f
C7311 FFCLR.n75 GND 0.06706f
C7312 FFCLR.t42 GND 0.20914f
C7313 D_FlipFlop_5.nCLR GND -0.24492f
C7314 FFCLR.n76 GND 0.31064f
C7315 FFCLR.n77 GND 0.12314f
C7316 FFCLR.t19 GND 0.2328f
C7317 D_FlipFlop_5.3-input-nand_5.A GND -0.20104f
C7318 FFCLR.n78 GND 0.21717f
C7319 FFCLR.n79 GND 0.0481f
C7320 FFCLR.t24 GND 0.44775f
C7321 FFCLR.n80 GND 0.1308f
C7322 FFCLR.n81 GND 0.04343f
C7323 FFCLR.n82 GND 0.07336f
C7324 FFCLR.n83 GND 0.27768f
C7325 FFCLR.t50 GND 0.2328f
C7326 D_FlipFlop_5.3-input-nand_3.A GND -0.20104f
C7327 FFCLR.n84 GND 0.21717f
C7328 FFCLR.n85 GND 0.0481f
C7329 FFCLR.t53 GND 0.44775f
C7330 FFCLR.n86 GND 0.1308f
C7331 FFCLR.n87 GND 0.04343f
C7332 FFCLR.n88 GND 0.07336f
C7333 FFCLR.n90 GND 0.7054f
C7334 FFCLR.n91 GND 0.10317f
C7335 FFCLR.n92 GND 0.219f
C7336 FFCLR.n94 GND 1.59688f
C7337 FFCLR.t58 GND 0.44777f
C7338 D_FlipFlop_3.3-input-nand_0.A GND -0.2662f
C7339 FFCLR.n95 GND 0.46425f
C7340 FFCLR.n96 GND 0.05023f
C7341 FFCLR.n97 GND 0.06706f
C7342 FFCLR.t27 GND 0.20914f
C7343 D_FlipFlop_3.nCLR GND -0.24492f
C7344 FFCLR.n98 GND 0.31064f
C7345 FFCLR.n99 GND 0.12314f
C7346 FFCLR.t21 GND 0.2328f
C7347 D_FlipFlop_3.3-input-nand_5.A GND -0.20104f
C7348 FFCLR.n100 GND 0.21717f
C7349 FFCLR.n101 GND 0.0481f
C7350 FFCLR.t47 GND 0.44775f
C7351 FFCLR.n102 GND 0.1308f
C7352 FFCLR.n103 GND 0.04343f
C7353 FFCLR.n104 GND 0.07336f
C7354 FFCLR.n105 GND 0.27768f
C7355 FFCLR.t20 GND 0.2328f
C7356 D_FlipFlop_3.3-input-nand_3.A GND -0.20104f
C7357 FFCLR.n106 GND 0.21717f
C7358 FFCLR.n107 GND 0.0481f
C7359 FFCLR.t39 GND 0.44775f
C7360 FFCLR.n108 GND 0.1308f
C7361 FFCLR.n109 GND 0.04343f
C7362 FFCLR.n110 GND 0.07336f
C7363 FFCLR.n112 GND 0.7054f
C7364 FFCLR.n113 GND 0.10317f
C7365 FFCLR.n114 GND 0.219f
C7366 FFCLR.n116 GND 1.59688f
C7367 FFCLR.t48 GND 0.44777f
C7368 D_FlipFlop_2.3-input-nand_0.A GND -0.2662f
C7369 FFCLR.n117 GND 0.46425f
C7370 FFCLR.n118 GND 0.05023f
C7371 FFCLR.n119 GND 0.06706f
C7372 FFCLR.t36 GND 0.20914f
C7373 D_FlipFlop_2.nCLR GND -0.24492f
C7374 FFCLR.n120 GND 0.31064f
C7375 FFCLR.n121 GND 0.12314f
C7376 FFCLR.t9 GND 0.2328f
C7377 D_FlipFlop_2.3-input-nand_5.A GND -0.20104f
C7378 FFCLR.n122 GND 0.21717f
C7379 FFCLR.n123 GND 0.0481f
C7380 FFCLR.t16 GND 0.44775f
C7381 FFCLR.n124 GND 0.1308f
C7382 FFCLR.n125 GND 0.04343f
C7383 FFCLR.n126 GND 0.07336f
C7384 FFCLR.n127 GND 0.27768f
C7385 FFCLR.t46 GND 0.2328f
C7386 D_FlipFlop_2.3-input-nand_3.A GND -0.20104f
C7387 FFCLR.n128 GND 0.21717f
C7388 FFCLR.n129 GND 0.0481f
C7389 FFCLR.t51 GND 0.44775f
C7390 FFCLR.n130 GND 0.1308f
C7391 FFCLR.n131 GND 0.04343f
C7392 FFCLR.n132 GND 0.07336f
C7393 FFCLR.n134 GND 0.7054f
C7394 FFCLR.n135 GND 0.10317f
C7395 FFCLR.n136 GND 0.219f
C7396 FFCLR.n138 GND 1.59688f
C7397 FFCLR.t7 GND 0.44777f
C7398 D_FlipFlop_1.3-input-nand_0.A GND -0.2662f
C7399 FFCLR.n139 GND 0.46425f
C7400 FFCLR.n140 GND 0.05023f
C7401 FFCLR.n141 GND 0.06706f
C7402 FFCLR.t31 GND 0.20914f
C7403 D_FlipFlop_1.nCLR GND -0.24492f
C7404 FFCLR.n142 GND 0.31064f
C7405 FFCLR.n143 GND 0.12314f
C7406 FFCLR.t40 GND 0.2328f
C7407 D_FlipFlop_1.3-input-nand_5.A GND -0.20104f
C7408 FFCLR.n144 GND 0.21717f
C7409 FFCLR.n145 GND 0.0481f
C7410 FFCLR.t8 GND 0.44775f
C7411 FFCLR.n146 GND 0.1308f
C7412 FFCLR.n147 GND 0.04343f
C7413 FFCLR.n148 GND 0.07336f
C7414 FFCLR.n149 GND 0.27768f
C7415 FFCLR.t37 GND 0.2328f
C7416 D_FlipFlop_1.3-input-nand_3.A GND -0.20104f
C7417 FFCLR.n150 GND 0.21717f
C7418 FFCLR.n151 GND 0.0481f
C7419 FFCLR.t45 GND 0.44775f
C7420 FFCLR.n152 GND 0.1308f
C7421 FFCLR.n153 GND 0.04343f
C7422 FFCLR.n154 GND 0.07336f
C7423 FFCLR.n156 GND 0.7054f
C7424 FFCLR.n157 GND 0.10317f
C7425 FFCLR.n158 GND 0.219f
C7426 FFCLR.n160 GND 1.6827f
C7427 FFCLR.n161 GND 0.68812f
C7428 FFCLR.n162 GND 0.12314f
C7429 FFCLR.n163 GND 0.20904f
C7430 FFCLR.t56 GND 0.44777f
C7431 D_FlipFlop_0.3-input-nand_4.A GND -0.29997f
C7432 FFCLR.n164 GND 0.45092f
C7433 FFCLR.n165 GND 0.0481f
C7434 FFCLR.t12 GND 0.23279f
C7435 FFCLR.n166 GND 0.06706f
C7436 FFCLR.n167 GND 0.01786f
C7437 FFCLR.n168 GND 0.02783f
C7438 FFCLR.n169 GND 0.27768f
C7439 FFCLR.t55 GND 0.44777f
C7440 D_FlipFlop_0.3-input-nand_2.A GND -0.29997f
C7441 FFCLR.n170 GND 0.45092f
C7442 FFCLR.n171 GND 0.0481f
C7443 FFCLR.t6 GND 0.23279f
C7444 FFCLR.n172 GND 0.06706f
C7445 FFCLR.n173 GND 0.01786f
C7446 FFCLR.n174 GND 0.02783f
C7447 FFCLR.n176 GND 0.7207f
C7448 FFCLR.n177 GND 0.67869f
C7449 FFCLR.n178 GND 1.35554f
C7450 Ring_Counter_0.D_FlipFlop_1.3-input-nand_0.B GND -0.0577f
C7451 FFCLR.t5 GND 0.23279f
C7452 FFCLR.n179 GND 0.06098f
C7453 FFCLR.n180 GND 0.05593f
C7454 FFCLR.t14 GND 0.44836f
C7455 Ring_Counter_0.D_FlipFlop_1.Inverter_0.Vin GND -0.0577f
C7456 FFCLR.n181 GND 0.1345f
C7457 FFCLR.t23 GND 0.23279f
C7458 FFCLR.n182 GND 0.06098f
C7459 FFCLR.n183 GND 0.05593f
C7460 FFCLR.n184 GND 0.14153f
C7461 FFCLR.n185 GND 0.14153f
C7462 FFCLR.n186 GND 0.1345f
C7463 FFCLR.t41 GND 0.57252f
C7464 Ring_Counter_0.Q0 GND 0.37211f
C7465 FFCLR.n187 GND 0.14042f
C7466 FFCLR.n188 GND -0.01433f
C7467 FFCLR.n189 GND 0.28444f
C7468 FFCLR.t13 GND 0.44775f
C7469 FFCLR.n190 GND 0.19502f
C7470 FFCLR.t22 GND 0.20898f
C7471 FFCLR.n191 GND 0.13642f
C7472 Ring_Counter_0.D_FlipFlop_0.Q GND 0.5111f
C7473 FFCLR.n192 GND 0.06533f
C7474 FFCLR.n193 GND 0.16565f
C7475 FFCLR.t2 GND 0.06073f
C7476 FFCLR.n194 GND 0.09355f
C7477 FFCLR.t0 GND 0.062f
C7478 FFCLR.t1 GND 0.06073f
C7479 FFCLR.n195 GND 0.34538f
C7480 FFCLR.n196 GND 0.1127f
C7481 FFCLR.n197 GND 0.22691f
C7482 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t1 GND 0.05f
C7483 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n0 GND 0.10867f
C7484 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n1 GND 0.05678f
C7485 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t3 GND 0.38491f
C7486 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n2 GND 0.16589f
C7487 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t2 GND 0.30131f
C7488 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t5 GND 0.30153f
C7489 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n3 GND 0.09671f
C7490 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t4 GND 0.38323f
C7491 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n4 GND 0.0709f
C7492 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n5 GND 0.04231f
C7493 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n6 GND 0.10383f
C7494 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n7 GND 0.10383f
C7495 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.t0 GND 0.05284f
C7496 Ring_Counter_0.D_FlipFlop_14.Inverter_1.Vout.n8 GND 0.17757f
C7497 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 GND 0.07411f
C7498 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 GND 0.16107f
C7499 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 GND 0.08416f
C7500 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 GND 0.29566f
C7501 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 GND 0.14335f
C7502 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 GND 0.56804f
C7503 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 GND 0.1051f
C7504 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 GND 0.06271f
C7505 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 GND 0.15391f
C7506 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 GND 0.15391f
C7507 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 GND 0.07722f
C7508 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 GND 0.07866f
C7509 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 GND 0.07705f
C7510 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 GND 0.43817f
C7511 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 GND 0.286f
C7512 Ring_Counter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 GND 0.09223f
C7513 D_FlipFlop_0.CLK.t1 GND 0.02954f
C7514 D_FlipFlop_0.CLK.t3 GND 0.22695f
C7515 D_FlipFlop_0.CLK.t4 GND 0.118f
C7516 D_FlipFlop_0.CLK.n0 GND 0.12444f
C7517 D_FlipFlop_0.CLK.t5 GND 0.22695f
C7518 D_FlipFlop_0.CLK.n1 GND 0.2009f
C7519 D_FlipFlop_0.CLK.n2 GND 0.20145f
C7520 D_FlipFlop_0.CLK.n3 GND 0.12607f
C7521 D_FlipFlop_0.CLK.t2 GND 0.10447f
C7522 D_FlipFlop_0.CLK.n4 GND 0.02736f
C7523 D_FlipFlop_0.CLK.n5 GND 0.10371f
C7524 D_FlipFlop_0.CLK.t7 GND 0.10446f
C7525 D_FlipFlop_0.CLK.n6 GND 0.03399f
C7526 D_FlipFlop_0.CLK.n7 GND 0.02546f
C7527 D_FlipFlop_0.CLK.n8 GND 0.23531f
C7528 D_FlipFlop_0.CLK.t6 GND 0.21911f
C7529 D_FlipFlop_0.CLK.n9 GND 0.16025f
C7530 D_FlipFlop_0.CLK.n11 GND 0.03049f
C7531 D_FlipFlop_0.CLK.t0 GND 0.03086f
C7532 D_FlipFlop_0.CLK.n12 GND 0.19695f
C7533 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t1 GND 0.06145f
C7534 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n0 GND 0.15815f
C7535 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n1 GND 0.12861f
C7536 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t6 GND 0.24486f
C7537 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t5 GND 0.47095f
C7538 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n2 GND 0.11174f
C7539 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n3 GND 0.11082f
C7540 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n4 GND 0.18808f
C7541 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n5 GND 0.14f
C7542 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t4 GND 0.47302f
C7543 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n6 GND 0.20386f
C7544 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t7 GND 0.23439f
C7545 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t2 GND 0.06388f
C7546 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n7 GND 0.40291f
C7547 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t0 GND 0.06521f
C7548 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.t3 GND 0.06388f
C7549 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n8 GND 0.36328f
C7550 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n9 GND 0.12591f
C7551 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.C.n10 GND 0.07837f
C7552 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 GND 0.05215f
C7553 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 GND 0.18008f
C7554 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 GND 0.37825f
C7555 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 GND 0.19588f
C7556 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 GND 0.28346f
C7557 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 GND 0.11199f
C7558 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 GND 0.01587f
C7559 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 GND 0.37675f
C7560 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 GND 0.16409f
C7561 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 GND 0.18888f
C7562 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 GND 0.0511f
C7563 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 GND 0.32168f
C7564 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 GND 0.05217f
C7565 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 GND 0.0511f
C7566 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 GND 0.29061f
C7567 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 GND 0.09483f
C7568 Ring_Counter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 GND 0.01203f
C7569 CLK.t77 GND 0.31985f
C7570 CLK.n0 GND 0.13785f
C7571 CLK.t2 GND 0.14658f
C7572 CLK.n1 GND 0.14553f
C7573 CLK.n2 GND 0.03839f
C7574 CLK.t6 GND 0.31846f
C7575 CLK.t48 GND 0.16606f
C7576 CLK.t25 GND 0.31846f
C7577 CLK.n3 GND 0.34246f
C7578 CLK.n4 GND 0.34324f
C7579 CLK.t100 GND 0.14706f
C7580 CLK.n5 GND 0.05973f
C7581 CLK.n6 GND 5.52957f
C7582 CLK.n7 GND 4.79885f
C7583 CLK.t13 GND 0.31985f
C7584 CLK.n8 GND 0.13785f
C7585 CLK.t103 GND 0.14658f
C7586 CLK.n9 GND 0.06019f
C7587 CLK.n10 GND 0.08229f
C7588 CLK.n11 GND 0.03839f
C7589 CLK.t80 GND 0.31846f
C7590 CLK.t29 GND 0.16606f
C7591 CLK.t99 GND 0.31846f
C7592 CLK.n12 GND 0.34246f
C7593 CLK.n13 GND 0.34324f
C7594 CLK.t84 GND 0.14706f
C7595 CLK.n14 GND 0.05973f
C7596 CLK.n15 GND 5.19984f
C7597 CLK.n16 GND 4.4991f
C7598 CLK.t41 GND 0.31985f
C7599 CLK.n17 GND 0.13785f
C7600 CLK.t86 GND 0.14658f
C7601 CLK.n18 GND 0.06019f
C7602 CLK.n19 GND 0.08229f
C7603 CLK.n20 GND 0.03839f
C7604 CLK.t56 GND 0.31846f
C7605 CLK.t42 GND 0.16606f
C7606 CLK.t78 GND 0.31846f
C7607 CLK.n21 GND 0.34246f
C7608 CLK.n22 GND 0.34324f
C7609 CLK.t92 GND 0.14706f
C7610 CLK.n23 GND 0.05973f
C7611 CLK.n24 GND 4.87011f
C7612 CLK.n25 GND 4.19934f
C7613 CLK.t63 GND 0.31985f
C7614 CLK.n26 GND 0.13785f
C7615 CLK.t114 GND 0.14658f
C7616 CLK.n27 GND 0.06019f
C7617 CLK.n28 GND 0.08229f
C7618 CLK.n29 GND 0.03839f
C7619 CLK.t23 GND 0.31846f
C7620 CLK.t108 GND 0.16606f
C7621 CLK.t46 GND 0.31846f
C7622 CLK.n30 GND 0.34246f
C7623 CLK.n31 GND 0.34324f
C7624 CLK.t28 GND 0.14706f
C7625 CLK.n32 GND 0.05973f
C7626 CLK.n33 GND 4.54039f
C7627 CLK.n34 GND 3.89959f
C7628 CLK.t34 GND 0.31985f
C7629 CLK.n35 GND 0.13785f
C7630 CLK.t93 GND 0.14658f
C7631 CLK.n36 GND 0.06019f
C7632 CLK.n37 GND 0.08229f
C7633 CLK.n38 GND 0.03839f
C7634 CLK.t50 GND 0.31846f
C7635 CLK.t35 GND 0.16606f
C7636 CLK.t72 GND 0.31846f
C7637 CLK.n39 GND 0.34246f
C7638 CLK.n40 GND 0.34324f
C7639 CLK.t89 GND 0.14706f
C7640 CLK.n41 GND 0.05973f
C7641 CLK.n42 GND 4.21066f
C7642 CLK.n43 GND 3.59984f
C7643 CLK.t12 GND 0.31985f
C7644 CLK.n44 GND 0.13785f
C7645 CLK.t73 GND 0.14658f
C7646 CLK.n45 GND 0.06019f
C7647 CLK.n46 GND 0.08229f
C7648 CLK.n47 GND 0.03839f
C7649 CLK.t43 GND 0.31846f
C7650 CLK.t27 GND 0.16606f
C7651 CLK.t64 GND 0.31846f
C7652 CLK.n48 GND 0.34246f
C7653 CLK.n49 GND 0.34324f
C7654 CLK.t81 GND 0.14706f
C7655 CLK.n50 GND 0.05973f
C7656 CLK.n51 GND 3.88093f
C7657 CLK.n52 GND 3.30009f
C7658 CLK.t51 GND 0.31985f
C7659 CLK.n53 GND 0.13785f
C7660 CLK.t90 GND 0.14658f
C7661 CLK.n54 GND 0.06019f
C7662 CLK.n55 GND 0.08229f
C7663 CLK.n56 GND 0.03839f
C7664 CLK.t44 GND 0.31846f
C7665 CLK.t9 GND 0.16606f
C7666 CLK.t65 GND 0.31846f
C7667 CLK.n57 GND 0.34246f
C7668 CLK.n58 GND 0.34324f
C7669 CLK.t61 GND 0.14706f
C7670 CLK.n59 GND 0.05973f
C7671 CLK.n60 GND 3.5512f
C7672 CLK.n61 GND 3.00033f
C7673 CLK.t5 GND 0.31985f
C7674 CLK.n62 GND 0.13785f
C7675 CLK.t66 GND 0.14658f
C7676 CLK.n63 GND 0.06019f
C7677 CLK.n64 GND 0.08229f
C7678 CLK.n65 GND 0.03839f
C7679 CLK.t38 GND 0.31846f
C7680 CLK.t20 GND 0.16606f
C7681 CLK.t57 GND 0.31846f
C7682 CLK.n66 GND 0.34246f
C7683 CLK.n67 GND 0.34324f
C7684 CLK.t74 GND 0.14706f
C7685 CLK.n68 GND 0.05973f
C7686 CLK.n69 GND 3.22147f
C7687 CLK.n70 GND 2.70058f
C7688 CLK.t0 GND 0.31985f
C7689 CLK.n71 GND 0.13785f
C7690 CLK.t102 GND 0.14658f
C7691 CLK.n72 GND 0.06019f
C7692 CLK.n73 GND 0.08229f
C7693 CLK.n74 GND 0.03839f
C7694 CLK.t62 GND 0.31846f
C7695 CLK.t14 GND 0.16606f
C7696 CLK.t87 GND 0.31846f
C7697 CLK.n75 GND 0.34246f
C7698 CLK.n76 GND 0.34324f
C7699 CLK.t67 GND 0.14706f
C7700 CLK.n77 GND 0.05973f
C7701 CLK.n78 GND 2.86861f
C7702 CLK.t75 GND 0.31846f
C7703 CLK.t111 GND 0.16606f
C7704 CLK.t95 GND 0.31846f
C7705 CLK.n79 GND 0.34246f
C7706 CLK.n80 GND 0.34324f
C7707 CLK.t32 GND 0.14706f
C7708 CLK.n81 GND 0.05945f
C7709 CLK.n82 GND 0.03839f
C7710 CLK.n83 GND 0.08229f
C7711 CLK.t3 GND 0.31985f
C7712 CLK.n84 GND 0.13785f
C7713 CLK.t7 GND 0.14658f
C7714 CLK.n85 GND 0.06019f
C7715 CLK.n86 GND 0.30255f
C7716 CLK.n87 GND 0.58364f
C7717 CLK.t88 GND 0.31846f
C7718 CLK.t94 GND 0.16606f
C7719 CLK.t104 GND 0.31846f
C7720 CLK.n88 GND 0.34246f
C7721 CLK.n89 GND 0.34324f
C7722 CLK.t11 GND 0.14706f
C7723 CLK.n90 GND 0.05973f
C7724 CLK.n91 GND 0.03839f
C7725 CLK.n92 GND 0.08229f
C7726 CLK.t112 GND 0.31985f
C7727 CLK.n93 GND 0.13785f
C7728 CLK.t17 GND 0.14658f
C7729 CLK.n94 GND 0.06019f
C7730 CLK.n95 GND 0.60231f
C7731 CLK.n96 GND 0.91337f
C7732 CLK.t109 GND 0.31846f
C7733 CLK.t49 GND 0.16606f
C7734 CLK.t1 GND 0.31846f
C7735 CLK.n97 GND 0.34246f
C7736 CLK.n98 GND 0.34324f
C7737 CLK.t101 GND 0.14706f
C7738 CLK.n99 GND 0.05973f
C7739 CLK.n100 GND 0.03839f
C7740 CLK.n101 GND 0.08229f
C7741 CLK.t69 GND 0.31985f
C7742 CLK.n102 GND 0.13785f
C7743 CLK.t117 GND 0.14658f
C7744 CLK.n103 GND 0.06019f
C7745 CLK.n104 GND 0.90206f
C7746 CLK.n105 GND 1.2431f
C7747 CLK.t60 GND 0.31846f
C7748 CLK.t24 GND 0.16606f
C7749 CLK.t83 GND 0.31846f
C7750 CLK.n106 GND 0.34246f
C7751 CLK.n107 GND 0.34324f
C7752 CLK.t79 GND 0.14706f
C7753 CLK.n108 GND 0.05973f
C7754 CLK.n109 GND 0.03839f
C7755 CLK.n110 GND 0.08229f
C7756 CLK.t10 GND 0.31985f
C7757 CLK.n111 GND 0.13785f
C7758 CLK.t71 GND 0.14658f
C7759 CLK.n112 GND 0.06019f
C7760 CLK.n113 GND 1.20181f
C7761 CLK.n114 GND 1.57283f
C7762 CLK.t47 GND 0.31846f
C7763 CLK.t33 GND 0.16606f
C7764 CLK.t70 GND 0.31846f
C7765 CLK.n115 GND 0.34246f
C7766 CLK.n116 GND 0.34324f
C7767 CLK.t85 GND 0.14706f
C7768 CLK.n117 GND 0.05973f
C7769 CLK.n118 GND 0.03839f
C7770 CLK.n119 GND 0.08229f
C7771 CLK.t16 GND 0.31985f
C7772 CLK.n120 GND 0.13785f
C7773 CLK.t76 GND 0.14658f
C7774 CLK.n121 GND 0.06019f
C7775 CLK.n122 GND 1.50157f
C7776 CLK.n123 GND 1.90256f
C7777 CLK.t36 GND 0.31846f
C7778 CLK.t113 GND 0.16606f
C7779 CLK.t55 GND 0.31846f
C7780 CLK.n124 GND 0.34246f
C7781 CLK.n125 GND 0.34324f
C7782 CLK.t39 GND 0.14706f
C7783 CLK.n126 GND 0.05973f
C7784 CLK.n127 GND 0.03839f
C7785 CLK.n128 GND 0.08229f
C7786 CLK.t31 GND 0.31985f
C7787 CLK.n129 GND 0.13785f
C7788 CLK.t106 GND 0.14658f
C7789 CLK.n130 GND 0.06019f
C7790 CLK.n131 GND 1.80132f
C7791 CLK.n132 GND 2.23229f
C7792 CLK.t21 GND 0.31846f
C7793 CLK.t8 GND 0.16606f
C7794 CLK.t45 GND 0.31846f
C7795 CLK.n133 GND 0.34246f
C7796 CLK.n134 GND 0.34324f
C7797 CLK.t59 GND 0.14706f
C7798 CLK.n135 GND 0.05973f
C7799 CLK.n136 GND 0.03839f
C7800 CLK.n137 GND 0.08229f
C7801 CLK.t116 GND 0.31985f
C7802 CLK.n138 GND 0.13785f
C7803 CLK.t53 GND 0.14658f
C7804 CLK.n139 GND 0.06019f
C7805 CLK.n140 GND 2.10107f
C7806 CLK.n141 GND 2.56201f
C7807 CLK.t30 GND 0.31846f
C7808 CLK.t15 GND 0.16606f
C7809 CLK.t52 GND 0.31846f
C7810 CLK.n142 GND 0.34246f
C7811 CLK.n143 GND 0.34324f
C7812 CLK.t68 GND 0.14706f
C7813 CLK.n144 GND 0.05973f
C7814 CLK.n145 GND 0.03839f
C7815 CLK.n146 GND 0.08229f
C7816 CLK.t54 GND 0.31985f
C7817 CLK.n147 GND 0.13785f
C7818 CLK.t58 GND 0.14658f
C7819 CLK.n148 GND 0.06019f
C7820 CLK.n149 GND 2.17029f
C7821 CLK.n150 GND 0.87916f
C7822 CLK.t98 GND 0.16557f
C7823 CLK.t18 GND 0.31846f
C7824 CLK.n151 GND 0.09303f
C7825 CLK.n152 GND 0.03978f
C7826 CLK.n153 GND 0.07346f
C7827 CLK.n154 GND 0.51556f
C7828 CLK.t82 GND 0.16557f
C7829 CLK.t91 GND 0.31846f
C7830 CLK.n155 GND 0.09303f
C7831 CLK.n156 GND 0.03978f
C7832 CLK.n157 GND 0.07346f
C7833 CLK.n158 GND 0.03825f
C7834 CLK.n159 GND 1.22359f
C7835 CLK.t107 GND 0.16557f
C7836 CLK.t19 GND 0.31846f
C7837 CLK.n160 GND 0.09303f
C7838 CLK.n161 GND 0.03978f
C7839 CLK.n162 GND 0.07346f
C7840 CLK.n163 GND 0.03825f
C7841 CLK.n164 GND 1.1332f
C7842 CLK.t40 GND 0.16557f
C7843 CLK.t96 GND 0.31846f
C7844 CLK.n165 GND 0.09303f
C7845 CLK.n166 GND 0.03978f
C7846 CLK.n167 GND 0.07346f
C7847 CLK.n168 GND 0.03825f
C7848 CLK.n169 GND 0.85039f
C7849 CLK.t105 GND 0.16557f
C7850 CLK.t97 GND 0.31846f
C7851 CLK.n170 GND 0.09303f
C7852 CLK.n171 GND 0.03978f
C7853 CLK.n172 GND 0.07346f
C7854 CLK.n173 GND 0.51556f
C7855 CLK.t4 GND 0.16557f
C7856 CLK.t26 GND 0.31846f
C7857 CLK.n174 GND 0.09303f
C7858 CLK.n175 GND 0.03978f
C7859 CLK.n176 GND 0.07346f
C7860 CLK.n177 GND 0.03825f
C7861 CLK.n178 GND 1.22359f
C7862 CLK.t22 GND 0.16557f
C7863 CLK.t37 GND 0.31846f
C7864 CLK.n179 GND 0.09303f
C7865 CLK.n180 GND 0.03978f
C7866 CLK.n181 GND 0.07346f
C7867 CLK.n182 GND 0.03825f
C7868 CLK.n183 GND 1.1332f
C7869 CLK.t110 GND 0.16557f
C7870 CLK.t115 GND 0.31846f
C7871 CLK.n184 GND 0.09303f
C7872 CLK.n185 GND 0.03978f
C7873 CLK.n186 GND 0.07346f
C7874 CLK.n187 GND 0.03825f
C7875 CLK.n188 GND 0.85039f
C7876 CLK.n189 GND 0.57148f
C7877 CLK.n190 GND 0.64951f
C7878 D_FlipFlop_4.CLK.t1 GND 0.02954f
C7879 D_FlipFlop_4.CLK.t4 GND 0.22695f
C7880 D_FlipFlop_4.CLK.t5 GND 0.118f
C7881 D_FlipFlop_4.CLK.n0 GND 0.12444f
C7882 D_FlipFlop_4.CLK.t6 GND 0.22695f
C7883 D_FlipFlop_4.CLK.n1 GND 0.2009f
C7884 D_FlipFlop_4.CLK.n2 GND 0.20145f
C7885 D_FlipFlop_4.CLK.n3 GND 0.12607f
C7886 D_FlipFlop_4.CLK.t3 GND 0.10447f
C7887 D_FlipFlop_4.CLK.n4 GND 0.02736f
C7888 D_FlipFlop_4.CLK.n5 GND 0.10371f
C7889 D_FlipFlop_4.CLK.t2 GND 0.10446f
C7890 D_FlipFlop_4.CLK.n6 GND 0.03399f
C7891 D_FlipFlop_4.CLK.n7 GND 0.02546f
C7892 D_FlipFlop_4.CLK.n8 GND 0.23531f
C7893 D_FlipFlop_4.CLK.t7 GND 0.21911f
C7894 D_FlipFlop_4.CLK.n9 GND 0.16025f
C7895 D_FlipFlop_4.CLK.n11 GND 0.03049f
C7896 D_FlipFlop_4.CLK.t0 GND 0.03086f
C7897 D_FlipFlop_4.CLK.n12 GND 0.19695f
C7898 CDAC_v3_0.switch_7.Z.t66 GND 0.04192f
C7899 CDAC_v3_0.switch_7.Z.t1 GND 0.04184f
C7900 CDAC_v3_0.switch_7.Z.n0 GND 0.09205f
C7901 CDAC_v3_0.switch_7.Z.n1 GND 0.01424f
C7902 CDAC_v3_0.switch_7.Z.t63 GND 5.67859f
C7903 CDAC_v3_0.switch_7.Z.t16 GND 5.67859f
C7904 CDAC_v3_0.switch_7.Z.t35 GND 5.67859f
C7905 CDAC_v3_0.switch_7.Z.t58 GND 5.67859f
C7906 CDAC_v3_0.switch_7.Z.t10 GND 5.67859f
C7907 CDAC_v3_0.switch_7.Z.t64 GND 5.67859f
C7908 CDAC_v3_0.switch_7.Z.t50 GND 5.67859f
C7909 CDAC_v3_0.switch_7.Z.t61 GND 6.21945f
C7910 CDAC_v3_0.switch_7.Z.n2 GND 0.97688f
C7911 CDAC_v3_0.switch_7.Z.n3 GND 0.93329f
C7912 CDAC_v3_0.switch_7.Z.n4 GND 0.93329f
C7913 CDAC_v3_0.switch_7.Z.n5 GND 0.93329f
C7914 CDAC_v3_0.switch_7.Z.n6 GND 0.93329f
C7915 CDAC_v3_0.switch_7.Z.n7 GND 0.93329f
C7916 CDAC_v3_0.switch_7.Z.n8 GND 1.53271f
C7917 CDAC_v3_0.switch_7.Z.t5 GND 5.67859f
C7918 CDAC_v3_0.switch_7.Z.t20 GND 5.67859f
C7919 CDAC_v3_0.switch_7.Z.t39 GND 5.67859f
C7920 CDAC_v3_0.switch_7.Z.t65 GND 5.67859f
C7921 CDAC_v3_0.switch_7.Z.t12 GND 5.67859f
C7922 CDAC_v3_0.switch_7.Z.t7 GND 5.67859f
C7923 CDAC_v3_0.switch_7.Z.t56 GND 5.67859f
C7924 CDAC_v3_0.switch_7.Z.t2 GND 6.21945f
C7925 CDAC_v3_0.switch_7.Z.n9 GND 0.97688f
C7926 CDAC_v3_0.switch_7.Z.n10 GND 0.93329f
C7927 CDAC_v3_0.switch_7.Z.n11 GND 0.93329f
C7928 CDAC_v3_0.switch_7.Z.n12 GND 0.93329f
C7929 CDAC_v3_0.switch_7.Z.n13 GND 0.93329f
C7930 CDAC_v3_0.switch_7.Z.n14 GND 0.93329f
C7931 CDAC_v3_0.switch_7.Z.n15 GND 1.30044f
C7932 CDAC_v3_0.switch_7.Z.n16 GND 1.67932f
C7933 CDAC_v3_0.switch_7.Z.t22 GND 5.67859f
C7934 CDAC_v3_0.switch_7.Z.t47 GND 5.67859f
C7935 CDAC_v3_0.switch_7.Z.t18 GND 5.67859f
C7936 CDAC_v3_0.switch_7.Z.t51 GND 5.67859f
C7937 CDAC_v3_0.switch_7.Z.t25 GND 5.67859f
C7938 CDAC_v3_0.switch_7.Z.t23 GND 5.67859f
C7939 CDAC_v3_0.switch_7.Z.t34 GND 5.67859f
C7940 CDAC_v3_0.switch_7.Z.t31 GND 6.21945f
C7941 CDAC_v3_0.switch_7.Z.n17 GND 0.97688f
C7942 CDAC_v3_0.switch_7.Z.n18 GND 0.93329f
C7943 CDAC_v3_0.switch_7.Z.n19 GND 0.93329f
C7944 CDAC_v3_0.switch_7.Z.n20 GND 0.93329f
C7945 CDAC_v3_0.switch_7.Z.n21 GND 0.93329f
C7946 CDAC_v3_0.switch_7.Z.n22 GND 0.93329f
C7947 CDAC_v3_0.switch_7.Z.n23 GND 1.30044f
C7948 CDAC_v3_0.switch_7.Z.n24 GND 1.15755f
C7949 CDAC_v3_0.switch_7.Z.t32 GND 5.67859f
C7950 CDAC_v3_0.switch_7.Z.t53 GND 5.67859f
C7951 CDAC_v3_0.switch_7.Z.t27 GND 5.67859f
C7952 CDAC_v3_0.switch_7.Z.t62 GND 5.67859f
C7953 CDAC_v3_0.switch_7.Z.t36 GND 5.67859f
C7954 CDAC_v3_0.switch_7.Z.t33 GND 5.67859f
C7955 CDAC_v3_0.switch_7.Z.t43 GND 5.67859f
C7956 CDAC_v3_0.switch_7.Z.t41 GND 6.21945f
C7957 CDAC_v3_0.switch_7.Z.n25 GND 0.97688f
C7958 CDAC_v3_0.switch_7.Z.n26 GND 0.93329f
C7959 CDAC_v3_0.switch_7.Z.n27 GND 0.93329f
C7960 CDAC_v3_0.switch_7.Z.n28 GND 0.93329f
C7961 CDAC_v3_0.switch_7.Z.n29 GND 0.93329f
C7962 CDAC_v3_0.switch_7.Z.n30 GND 0.93329f
C7963 CDAC_v3_0.switch_7.Z.n31 GND 1.30044f
C7964 CDAC_v3_0.switch_7.Z.n32 GND 1.56661f
C7965 CDAC_v3_0.switch_7.Z.t4 GND 5.67859f
C7966 CDAC_v3_0.switch_7.Z.t15 GND 5.67859f
C7967 CDAC_v3_0.switch_7.Z.t52 GND 5.67859f
C7968 CDAC_v3_0.switch_7.Z.t26 GND 5.67859f
C7969 CDAC_v3_0.switch_7.Z.t29 GND 5.67859f
C7970 CDAC_v3_0.switch_7.Z.t59 GND 5.67859f
C7971 CDAC_v3_0.switch_7.Z.t38 GND 5.67859f
C7972 CDAC_v3_0.switch_7.Z.t8 GND 6.70945f
C7973 CDAC_v3_0.switch_7.Z.n33 GND 1.01637f
C7974 CDAC_v3_0.switch_7.Z.n34 GND 0.93329f
C7975 CDAC_v3_0.switch_7.Z.n35 GND 0.93329f
C7976 CDAC_v3_0.switch_7.Z.n36 GND 0.93329f
C7977 CDAC_v3_0.switch_7.Z.n37 GND 0.93329f
C7978 CDAC_v3_0.switch_7.Z.n38 GND 0.93329f
C7979 CDAC_v3_0.switch_7.Z.n39 GND 0.9783f
C7980 CDAC_v3_0.switch_7.Z.n40 GND 1.35926f
C7981 CDAC_v3_0.switch_7.Z.t19 GND 5.67859f
C7982 CDAC_v3_0.switch_7.Z.t37 GND 5.67859f
C7983 CDAC_v3_0.switch_7.Z.t9 GND 5.67859f
C7984 CDAC_v3_0.switch_7.Z.t46 GND 5.67859f
C7985 CDAC_v3_0.switch_7.Z.t48 GND 5.67859f
C7986 CDAC_v3_0.switch_7.Z.t13 GND 5.67859f
C7987 CDAC_v3_0.switch_7.Z.t54 GND 5.67859f
C7988 CDAC_v3_0.switch_7.Z.t28 GND 6.70945f
C7989 CDAC_v3_0.switch_7.Z.n41 GND 1.01637f
C7990 CDAC_v3_0.switch_7.Z.n42 GND 0.93329f
C7991 CDAC_v3_0.switch_7.Z.n43 GND 0.93329f
C7992 CDAC_v3_0.switch_7.Z.n44 GND 0.93329f
C7993 CDAC_v3_0.switch_7.Z.n45 GND 0.93329f
C7994 CDAC_v3_0.switch_7.Z.n46 GND 0.93329f
C7995 CDAC_v3_0.switch_7.Z.n47 GND 0.9783f
C7996 CDAC_v3_0.switch_7.Z.n48 GND 0.9502f
C7997 CDAC_v3_0.switch_7.Z.t30 GND 5.67859f
C7998 CDAC_v3_0.switch_7.Z.t45 GND 5.67859f
C7999 CDAC_v3_0.switch_7.Z.t17 GND 5.67859f
C8000 CDAC_v3_0.switch_7.Z.t55 GND 5.67859f
C8001 CDAC_v3_0.switch_7.Z.t60 GND 5.67859f
C8002 CDAC_v3_0.switch_7.Z.t24 GND 5.67859f
C8003 CDAC_v3_0.switch_7.Z.t6 GND 5.67859f
C8004 CDAC_v3_0.switch_7.Z.t40 GND 6.70945f
C8005 CDAC_v3_0.switch_7.Z.n49 GND 1.01637f
C8006 CDAC_v3_0.switch_7.Z.n50 GND 0.93329f
C8007 CDAC_v3_0.switch_7.Z.n51 GND 0.93329f
C8008 CDAC_v3_0.switch_7.Z.n52 GND 0.93329f
C8009 CDAC_v3_0.switch_7.Z.n53 GND 0.93329f
C8010 CDAC_v3_0.switch_7.Z.n54 GND 0.93329f
C8011 CDAC_v3_0.switch_7.Z.n55 GND 0.9783f
C8012 CDAC_v3_0.switch_7.Z.n56 GND 0.9502f
C8013 CDAC_v3_0.switch_7.Z.t49 GND 5.67859f
C8014 CDAC_v3_0.switch_7.Z.t3 GND 5.67859f
C8015 CDAC_v3_0.switch_7.Z.t42 GND 5.67859f
C8016 CDAC_v3_0.switch_7.Z.t11 GND 5.67859f
C8017 CDAC_v3_0.switch_7.Z.t14 GND 5.67859f
C8018 CDAC_v3_0.switch_7.Z.t44 GND 5.67859f
C8019 CDAC_v3_0.switch_7.Z.t21 GND 5.67859f
C8020 CDAC_v3_0.switch_7.Z.t57 GND 6.70945f
C8021 CDAC_v3_0.switch_7.Z.n57 GND 1.01637f
C8022 CDAC_v3_0.switch_7.Z.n58 GND 0.93329f
C8023 CDAC_v3_0.switch_7.Z.n59 GND 0.93329f
C8024 CDAC_v3_0.switch_7.Z.n60 GND 0.93329f
C8025 CDAC_v3_0.switch_7.Z.n61 GND 0.93329f
C8026 CDAC_v3_0.switch_7.Z.n62 GND 0.93329f
C8027 CDAC_v3_0.switch_7.Z.n63 GND 0.9783f
C8028 CDAC_v3_0.switch_7.Z.n64 GND 4.43744f
C8029 CDAC_v3_0.switch_7.Z.n65 GND 2.2303f
C8030 CDAC_v3_0.switch_7.Z.n66 GND 0.04484f
C8031 CDAC_v3_0.switch_7.Z.t67 GND 0.04328f
C8032 CDAC_v3_0.switch_7.Z.t0 GND 0.04328f
C8033 CDAC_v3_0.switch_7.Z.n67 GND 0.15546f
C8034 CDAC_v3_0.switch_7.Z.n68 GND 0.4793f
C8035 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 GND 0.05215f
C8036 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 GND 0.18008f
C8037 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 GND 0.37825f
C8038 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 GND 0.19588f
C8039 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 GND 0.28346f
C8040 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 GND 0.11199f
C8041 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 GND 0.01587f
C8042 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 GND 0.37675f
C8043 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 GND 0.16409f
C8044 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 GND 0.18888f
C8045 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 GND 0.0511f
C8046 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 GND 0.32168f
C8047 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 GND 0.05217f
C8048 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 GND 0.0511f
C8049 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 GND 0.29061f
C8050 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 GND 0.09483f
C8051 Ring_Counter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 GND 0.01203f
C8052 D_FlipFlop_2.3-input-nand_2.Vout.t5 GND 0.34247f
C8053 D_FlipFlop_2.3-input-nand_2.Vout.n0 GND 0.10005f
C8054 D_FlipFlop_2.3-input-nand_2.Vout.n1 GND 0.04341f
C8055 D_FlipFlop_2.3-input-nand_2.Vout.t3 GND 0.04467f
C8056 D_FlipFlop_2.3-input-nand_2.Vout.n2 GND 0.21241f
C8057 D_FlipFlop_2.3-input-nand_2.Vout.n3 GND 0.04823f
C8058 D_FlipFlop_2.3-input-nand_2.Vout.t7 GND 0.34248f
C8059 D_FlipFlop_2.3-input-nand_2.Vout.n4 GND 0.35447f
C8060 D_FlipFlop_2.3-input-nand_2.Vout.t4 GND 0.17806f
C8061 D_FlipFlop_2.3-input-nand_2.Vout.n5 GND 0.17459f
C8062 D_FlipFlop_2.3-input-nand_2.Vout.n6 GND 0.1018f
C8063 D_FlipFlop_2.3-input-nand_2.Vout.n7 GND 0.01283f
C8064 D_FlipFlop_2.3-input-nand_2.Vout.n8 GND 0.01019f
C8065 D_FlipFlop_2.3-input-nand_2.Vout.t2 GND 0.04742f
C8066 D_FlipFlop_2.3-input-nand_2.Vout.t0 GND 0.04645f
C8067 D_FlipFlop_2.3-input-nand_2.Vout.n9 GND 0.26417f
C8068 D_FlipFlop_2.3-input-nand_2.Vout.n10 GND 0.0862f
C8069 D_FlipFlop_2.3-input-nand_2.Vout.t1 GND 0.04645f
C8070 D_FlipFlop_2.3-input-nand_2.Vout.n11 GND 0.29241f
C8071 D_FlipFlop_2.3-input-nand_2.Vout.t6 GND 0.17113f
C8072 D_FlipFlop_2.3-input-nand_2.Vout.n12 GND 0.19086f
C8073 CDAC_v3_0.switch_6.Z.t2 GND 0.04156f
C8074 CDAC_v3_0.switch_6.Z.t1 GND 0.04148f
C8075 CDAC_v3_0.switch_6.Z.n0 GND 0.09126f
C8076 CDAC_v3_0.switch_6.Z.n1 GND 0.01412f
C8077 CDAC_v3_0.switch_6.Z.t30 GND 5.62981f
C8078 CDAC_v3_0.switch_6.Z.t129 GND 5.62981f
C8079 CDAC_v3_0.switch_6.Z.t118 GND 5.62981f
C8080 CDAC_v3_0.switch_6.Z.t48 GND 5.62981f
C8081 CDAC_v3_0.switch_6.Z.t53 GND 5.62981f
C8082 CDAC_v3_0.switch_6.Z.t17 GND 5.62981f
C8083 CDAC_v3_0.switch_6.Z.t95 GND 5.62981f
C8084 CDAC_v3_0.switch_6.Z.t34 GND 6.01712f
C8085 CDAC_v3_0.switch_6.Z.t88 GND 5.76479f
C8086 CDAC_v3_0.switch_6.Z.n2 GND 0.49725f
C8087 CDAC_v3_0.switch_6.Z.n3 GND 0.51837f
C8088 CDAC_v3_0.switch_6.Z.t3 GND 5.76479f
C8089 CDAC_v3_0.switch_6.Z.n4 GND 0.44889f
C8090 CDAC_v3_0.switch_6.Z.n5 GND 0.51837f
C8091 CDAC_v3_0.switch_6.Z.t40 GND 5.76479f
C8092 CDAC_v3_0.switch_6.Z.n6 GND 0.44889f
C8093 CDAC_v3_0.switch_6.Z.n7 GND 0.51837f
C8094 CDAC_v3_0.switch_6.Z.t83 GND 5.76479f
C8095 CDAC_v3_0.switch_6.Z.n8 GND 0.44889f
C8096 CDAC_v3_0.switch_6.Z.n9 GND 0.51837f
C8097 CDAC_v3_0.switch_6.Z.t119 GND 5.76479f
C8098 CDAC_v3_0.switch_6.Z.n10 GND 0.44889f
C8099 CDAC_v3_0.switch_6.Z.n11 GND 0.51837f
C8100 CDAC_v3_0.switch_6.Z.t94 GND 5.76479f
C8101 CDAC_v3_0.switch_6.Z.n12 GND 0.44889f
C8102 CDAC_v3_0.switch_6.Z.n13 GND 0.51837f
C8103 CDAC_v3_0.switch_6.Z.t72 GND 5.76479f
C8104 CDAC_v3_0.switch_6.Z.n14 GND 0.44889f
C8105 CDAC_v3_0.switch_6.Z.n15 GND 0.51837f
C8106 CDAC_v3_0.switch_6.Z.t86 GND 5.76479f
C8107 CDAC_v3_0.switch_6.Z.n16 GND 0.96449f
C8108 CDAC_v3_0.switch_6.Z.t43 GND 5.62981f
C8109 CDAC_v3_0.switch_6.Z.t4 GND 5.62981f
C8110 CDAC_v3_0.switch_6.Z.t127 GND 5.62981f
C8111 CDAC_v3_0.switch_6.Z.t54 GND 5.62981f
C8112 CDAC_v3_0.switch_6.Z.t59 GND 5.62981f
C8113 CDAC_v3_0.switch_6.Z.t29 GND 5.62981f
C8114 CDAC_v3_0.switch_6.Z.t103 GND 5.62981f
C8115 CDAC_v3_0.switch_6.Z.t46 GND 6.01712f
C8116 CDAC_v3_0.switch_6.Z.t15 GND 5.76479f
C8117 CDAC_v3_0.switch_6.Z.n17 GND 0.49725f
C8118 CDAC_v3_0.switch_6.Z.n18 GND 0.51837f
C8119 CDAC_v3_0.switch_6.Z.t65 GND 5.76479f
C8120 CDAC_v3_0.switch_6.Z.n19 GND 0.44889f
C8121 CDAC_v3_0.switch_6.Z.n20 GND 0.51837f
C8122 CDAC_v3_0.switch_6.Z.t7 GND 5.76479f
C8123 CDAC_v3_0.switch_6.Z.n21 GND 0.44889f
C8124 CDAC_v3_0.switch_6.Z.n22 GND 0.51837f
C8125 CDAC_v3_0.switch_6.Z.t73 GND 5.76479f
C8126 CDAC_v3_0.switch_6.Z.n23 GND 0.44889f
C8127 CDAC_v3_0.switch_6.Z.n24 GND 0.51837f
C8128 CDAC_v3_0.switch_6.Z.t19 GND 5.76479f
C8129 CDAC_v3_0.switch_6.Z.n25 GND 0.44889f
C8130 CDAC_v3_0.switch_6.Z.n26 GND 0.51837f
C8131 CDAC_v3_0.switch_6.Z.t16 GND 5.76479f
C8132 CDAC_v3_0.switch_6.Z.n27 GND 0.44889f
C8133 CDAC_v3_0.switch_6.Z.n28 GND 0.51837f
C8134 CDAC_v3_0.switch_6.Z.t33 GND 5.76479f
C8135 CDAC_v3_0.switch_6.Z.n29 GND 0.44889f
C8136 CDAC_v3_0.switch_6.Z.n30 GND 0.51837f
C8137 CDAC_v3_0.switch_6.Z.t31 GND 5.76479f
C8138 CDAC_v3_0.switch_6.Z.n31 GND 0.75578f
C8139 CDAC_v3_0.switch_6.Z.n32 GND 1.2746f
C8140 CDAC_v3_0.switch_6.Z.t10 GND 5.62981f
C8141 CDAC_v3_0.switch_6.Z.t66 GND 5.62981f
C8142 CDAC_v3_0.switch_6.Z.t110 GND 5.62981f
C8143 CDAC_v3_0.switch_6.Z.t57 GND 5.62981f
C8144 CDAC_v3_0.switch_6.Z.t49 GND 5.62981f
C8145 CDAC_v3_0.switch_6.Z.t97 GND 5.62981f
C8146 CDAC_v3_0.switch_6.Z.t28 GND 5.62981f
C8147 CDAC_v3_0.switch_6.Z.t124 GND 6.01712f
C8148 CDAC_v3_0.switch_6.Z.t90 GND 5.76479f
C8149 CDAC_v3_0.switch_6.Z.n33 GND 0.49725f
C8150 CDAC_v3_0.switch_6.Z.n34 GND 0.51837f
C8151 CDAC_v3_0.switch_6.Z.t13 GND 5.76479f
C8152 CDAC_v3_0.switch_6.Z.n35 GND 0.44889f
C8153 CDAC_v3_0.switch_6.Z.n36 GND 0.51837f
C8154 CDAC_v3_0.switch_6.Z.t82 GND 5.76479f
C8155 CDAC_v3_0.switch_6.Z.n37 GND 0.44889f
C8156 CDAC_v3_0.switch_6.Z.n38 GND 0.51837f
C8157 CDAC_v3_0.switch_6.Z.t25 GND 5.76479f
C8158 CDAC_v3_0.switch_6.Z.n39 GND 0.44889f
C8159 CDAC_v3_0.switch_6.Z.n40 GND 0.51837f
C8160 CDAC_v3_0.switch_6.Z.t96 GND 5.76479f
C8161 CDAC_v3_0.switch_6.Z.n41 GND 0.44889f
C8162 CDAC_v3_0.switch_6.Z.n42 GND 0.51837f
C8163 CDAC_v3_0.switch_6.Z.t91 GND 5.76479f
C8164 CDAC_v3_0.switch_6.Z.n43 GND 0.44889f
C8165 CDAC_v3_0.switch_6.Z.n44 GND 0.51837f
C8166 CDAC_v3_0.switch_6.Z.t108 GND 5.76479f
C8167 CDAC_v3_0.switch_6.Z.n45 GND 0.44889f
C8168 CDAC_v3_0.switch_6.Z.n46 GND 0.51837f
C8169 CDAC_v3_0.switch_6.Z.t107 GND 5.76479f
C8170 CDAC_v3_0.switch_6.Z.n47 GND 0.75578f
C8171 CDAC_v3_0.switch_6.Z.n48 GND 0.94156f
C8172 CDAC_v3_0.switch_6.Z.t27 GND 5.62981f
C8173 CDAC_v3_0.switch_6.Z.t77 GND 5.62981f
C8174 CDAC_v3_0.switch_6.Z.t128 GND 5.62981f
C8175 CDAC_v3_0.switch_6.Z.t69 GND 5.62981f
C8176 CDAC_v3_0.switch_6.Z.t61 GND 5.62981f
C8177 CDAC_v3_0.switch_6.Z.t113 GND 5.62981f
C8178 CDAC_v3_0.switch_6.Z.t45 GND 5.62981f
C8179 CDAC_v3_0.switch_6.Z.t11 GND 6.01712f
C8180 CDAC_v3_0.switch_6.Z.t101 GND 5.76479f
C8181 CDAC_v3_0.switch_6.Z.n49 GND 0.49725f
C8182 CDAC_v3_0.switch_6.Z.n50 GND 0.51837f
C8183 CDAC_v3_0.switch_6.Z.t21 GND 5.76479f
C8184 CDAC_v3_0.switch_6.Z.n51 GND 0.44889f
C8185 CDAC_v3_0.switch_6.Z.n52 GND 0.51837f
C8186 CDAC_v3_0.switch_6.Z.t93 GND 5.76479f
C8187 CDAC_v3_0.switch_6.Z.n53 GND 0.44889f
C8188 CDAC_v3_0.switch_6.Z.n54 GND 0.51837f
C8189 CDAC_v3_0.switch_6.Z.t38 GND 5.76479f
C8190 CDAC_v3_0.switch_6.Z.n55 GND 0.44889f
C8191 CDAC_v3_0.switch_6.Z.n56 GND 0.51837f
C8192 CDAC_v3_0.switch_6.Z.t105 GND 5.76479f
C8193 CDAC_v3_0.switch_6.Z.n57 GND 0.44889f
C8194 CDAC_v3_0.switch_6.Z.n58 GND 0.51837f
C8195 CDAC_v3_0.switch_6.Z.t102 GND 5.76479f
C8196 CDAC_v3_0.switch_6.Z.n59 GND 0.44889f
C8197 CDAC_v3_0.switch_6.Z.n60 GND 0.51837f
C8198 CDAC_v3_0.switch_6.Z.t117 GND 5.76479f
C8199 CDAC_v3_0.switch_6.Z.n61 GND 0.44889f
C8200 CDAC_v3_0.switch_6.Z.n62 GND 0.51837f
C8201 CDAC_v3_0.switch_6.Z.t115 GND 5.76479f
C8202 CDAC_v3_0.switch_6.Z.n63 GND 0.75578f
C8203 CDAC_v3_0.switch_6.Z.n64 GND 0.97258f
C8204 CDAC_v3_0.switch_6.Z.t74 GND 5.62981f
C8205 CDAC_v3_0.switch_6.Z.t75 GND 5.62981f
C8206 CDAC_v3_0.switch_6.Z.t64 GND 5.62981f
C8207 CDAC_v3_0.switch_6.Z.t67 GND 5.62981f
C8208 CDAC_v3_0.switch_6.Z.t120 GND 5.62981f
C8209 CDAC_v3_0.switch_6.Z.t58 GND 5.62981f
C8210 CDAC_v3_0.switch_6.Z.t109 GND 5.62981f
C8211 CDAC_v3_0.switch_6.Z.t63 GND 5.62981f
C8212 CDAC_v3_0.switch_6.Z.t87 GND 5.82965f
C8213 CDAC_v3_0.switch_6.Z.n65 GND 0.7112f
C8214 CDAC_v3_0.switch_6.Z.t123 GND 5.76457f
C8215 CDAC_v3_0.switch_6.Z.n66 GND 0.44859f
C8216 CDAC_v3_0.switch_6.Z.n67 GND 0.51844f
C8217 CDAC_v3_0.switch_6.Z.t70 GND 5.76457f
C8218 CDAC_v3_0.switch_6.Z.n68 GND 0.44859f
C8219 CDAC_v3_0.switch_6.Z.n69 GND 0.51844f
C8220 CDAC_v3_0.switch_6.Z.t14 GND 5.76457f
C8221 CDAC_v3_0.switch_6.Z.n70 GND 0.44859f
C8222 CDAC_v3_0.switch_6.Z.n71 GND 0.51844f
C8223 CDAC_v3_0.switch_6.Z.t22 GND 5.76457f
C8224 CDAC_v3_0.switch_6.Z.n72 GND 0.44859f
C8225 CDAC_v3_0.switch_6.Z.n73 GND 0.51844f
C8226 CDAC_v3_0.switch_6.Z.t79 GND 5.76457f
C8227 CDAC_v3_0.switch_6.Z.n74 GND 0.44859f
C8228 CDAC_v3_0.switch_6.Z.n75 GND 0.51844f
C8229 CDAC_v3_0.switch_6.Z.t39 GND 5.76457f
C8230 CDAC_v3_0.switch_6.Z.n76 GND 0.44859f
C8231 CDAC_v3_0.switch_6.Z.n77 GND 0.51844f
C8232 CDAC_v3_0.switch_6.Z.t106 GND 5.76457f
C8233 CDAC_v3_0.switch_6.Z.n78 GND 0.44859f
C8234 CDAC_v3_0.switch_6.Z.n79 GND 0.82617f
C8235 CDAC_v3_0.switch_6.Z.n80 GND 0.97306f
C8236 CDAC_v3_0.switch_6.Z.t114 GND 5.62981f
C8237 CDAC_v3_0.switch_6.Z.t116 GND 5.62981f
C8238 CDAC_v3_0.switch_6.Z.t100 GND 5.62981f
C8239 CDAC_v3_0.switch_6.Z.t104 GND 5.62981f
C8240 CDAC_v3_0.switch_6.Z.t35 GND 5.62981f
C8241 CDAC_v3_0.switch_6.Z.t92 GND 5.62981f
C8242 CDAC_v3_0.switch_6.Z.t20 GND 5.62981f
C8243 CDAC_v3_0.switch_6.Z.t99 GND 5.62981f
C8244 CDAC_v3_0.switch_6.Z.t9 GND 5.82965f
C8245 CDAC_v3_0.switch_6.Z.n81 GND 0.7112f
C8246 CDAC_v3_0.switch_6.Z.t44 GND 5.76457f
C8247 CDAC_v3_0.switch_6.Z.n82 GND 0.44859f
C8248 CDAC_v3_0.switch_6.Z.n83 GND 0.51844f
C8249 CDAC_v3_0.switch_6.Z.t112 GND 5.76457f
C8250 CDAC_v3_0.switch_6.Z.n84 GND 0.44859f
C8251 CDAC_v3_0.switch_6.Z.n85 GND 0.51844f
C8252 CDAC_v3_0.switch_6.Z.t60 GND 5.76457f
C8253 CDAC_v3_0.switch_6.Z.n86 GND 0.44859f
C8254 CDAC_v3_0.switch_6.Z.n87 GND 0.51844f
C8255 CDAC_v3_0.switch_6.Z.t68 GND 5.76457f
C8256 CDAC_v3_0.switch_6.Z.n88 GND 0.44859f
C8257 CDAC_v3_0.switch_6.Z.n89 GND 0.51844f
C8258 CDAC_v3_0.switch_6.Z.t126 GND 5.76457f
C8259 CDAC_v3_0.switch_6.Z.n90 GND 0.44859f
C8260 CDAC_v3_0.switch_6.Z.n91 GND 0.51844f
C8261 CDAC_v3_0.switch_6.Z.t76 GND 5.76457f
C8262 CDAC_v3_0.switch_6.Z.n92 GND 0.44859f
C8263 CDAC_v3_0.switch_6.Z.n93 GND 0.51844f
C8264 CDAC_v3_0.switch_6.Z.t24 GND 5.76457f
C8265 CDAC_v3_0.switch_6.Z.n94 GND 0.44859f
C8266 CDAC_v3_0.switch_6.Z.n95 GND 0.82617f
C8267 CDAC_v3_0.switch_6.Z.n96 GND 0.94204f
C8268 CDAC_v3_0.switch_6.Z.t5 GND 5.62981f
C8269 CDAC_v3_0.switch_6.Z.t6 GND 5.62981f
C8270 CDAC_v3_0.switch_6.Z.t122 GND 5.62981f
C8271 CDAC_v3_0.switch_6.Z.t125 GND 5.62981f
C8272 CDAC_v3_0.switch_6.Z.t55 GND 5.62981f
C8273 CDAC_v3_0.switch_6.Z.t111 GND 5.62981f
C8274 CDAC_v3_0.switch_6.Z.t47 GND 5.62981f
C8275 CDAC_v3_0.switch_6.Z.t121 GND 5.62981f
C8276 CDAC_v3_0.switch_6.Z.t23 GND 5.82965f
C8277 CDAC_v3_0.switch_6.Z.n97 GND 0.7112f
C8278 CDAC_v3_0.switch_6.Z.t56 GND 5.76457f
C8279 CDAC_v3_0.switch_6.Z.n98 GND 0.44859f
C8280 CDAC_v3_0.switch_6.Z.n99 GND 0.51844f
C8281 CDAC_v3_0.switch_6.Z.t130 GND 5.76457f
C8282 CDAC_v3_0.switch_6.Z.n100 GND 0.44859f
C8283 CDAC_v3_0.switch_6.Z.n101 GND 0.51844f
C8284 CDAC_v3_0.switch_6.Z.t71 GND 5.76457f
C8285 CDAC_v3_0.switch_6.Z.n102 GND 0.44859f
C8286 CDAC_v3_0.switch_6.Z.n103 GND 0.51844f
C8287 CDAC_v3_0.switch_6.Z.t80 GND 5.76457f
C8288 CDAC_v3_0.switch_6.Z.n104 GND 0.44859f
C8289 CDAC_v3_0.switch_6.Z.n105 GND 0.51844f
C8290 CDAC_v3_0.switch_6.Z.t12 GND 5.76457f
C8291 CDAC_v3_0.switch_6.Z.n106 GND 0.44859f
C8292 CDAC_v3_0.switch_6.Z.n107 GND 0.51844f
C8293 CDAC_v3_0.switch_6.Z.t89 GND 5.76457f
C8294 CDAC_v3_0.switch_6.Z.n108 GND 0.44859f
C8295 CDAC_v3_0.switch_6.Z.n109 GND 0.51844f
C8296 CDAC_v3_0.switch_6.Z.t42 GND 5.76457f
C8297 CDAC_v3_0.switch_6.Z.n110 GND 0.44859f
C8298 CDAC_v3_0.switch_6.Z.n111 GND 0.82617f
C8299 CDAC_v3_0.switch_6.Z.n112 GND 0.94204f
C8300 CDAC_v3_0.switch_6.Z.t51 GND 5.62981f
C8301 CDAC_v3_0.switch_6.Z.t52 GND 5.62981f
C8302 CDAC_v3_0.switch_6.Z.t37 GND 5.62981f
C8303 CDAC_v3_0.switch_6.Z.t41 GND 5.62981f
C8304 CDAC_v3_0.switch_6.Z.t85 GND 5.62981f
C8305 CDAC_v3_0.switch_6.Z.t26 GND 5.62981f
C8306 CDAC_v3_0.switch_6.Z.t78 GND 5.62981f
C8307 CDAC_v3_0.switch_6.Z.t36 GND 5.62981f
C8308 CDAC_v3_0.switch_6.Z.t32 GND 5.82965f
C8309 CDAC_v3_0.switch_6.Z.n113 GND 0.7112f
C8310 CDAC_v3_0.switch_6.Z.t62 GND 5.76457f
C8311 CDAC_v3_0.switch_6.Z.n114 GND 0.44859f
C8312 CDAC_v3_0.switch_6.Z.n115 GND 0.51844f
C8313 CDAC_v3_0.switch_6.Z.t8 GND 5.76457f
C8314 CDAC_v3_0.switch_6.Z.n116 GND 0.44859f
C8315 CDAC_v3_0.switch_6.Z.n117 GND 0.51844f
C8316 CDAC_v3_0.switch_6.Z.t81 GND 5.76457f
C8317 CDAC_v3_0.switch_6.Z.n118 GND 0.44859f
C8318 CDAC_v3_0.switch_6.Z.n119 GND 0.51844f
C8319 CDAC_v3_0.switch_6.Z.t84 GND 5.76457f
C8320 CDAC_v3_0.switch_6.Z.n120 GND 0.44859f
C8321 CDAC_v3_0.switch_6.Z.n121 GND 0.51844f
C8322 CDAC_v3_0.switch_6.Z.t18 GND 5.76457f
C8323 CDAC_v3_0.switch_6.Z.n122 GND 0.44859f
C8324 CDAC_v3_0.switch_6.Z.n123 GND 0.51844f
C8325 CDAC_v3_0.switch_6.Z.t98 GND 5.76457f
C8326 CDAC_v3_0.switch_6.Z.n124 GND 0.44859f
C8327 CDAC_v3_0.switch_6.Z.n125 GND 0.51844f
C8328 CDAC_v3_0.switch_6.Z.t50 GND 5.76457f
C8329 CDAC_v3_0.switch_6.Z.n126 GND 0.44859f
C8330 CDAC_v3_0.switch_6.Z.n127 GND 0.82617f
C8331 CDAC_v3_0.switch_6.Z.n128 GND 2.41061f
C8332 CDAC_v3_0.switch_6.Z.n129 GND 0.73072f
C8333 CDAC_v3_0.switch_6.Z.n130 GND 0.04446f
C8334 CDAC_v3_0.switch_6.Z.t131 GND 0.04291f
C8335 CDAC_v3_0.switch_6.Z.t0 GND 0.04291f
C8336 CDAC_v3_0.switch_6.Z.n131 GND 0.15412f
C8337 CDAC_v3_0.switch_6.Z.n132 GND 0.47518f
C8338 Nand_Gate_1.A.t2 GND 0.03449f
C8339 Nand_Gate_1.A.t5 GND 0.24485f
C8340 Nand_Gate_1.A.n0 GND 0.07153f
C8341 Nand_Gate_1.A.n1 GND 0.03103f
C8342 Nand_Gate_1.A.n2 GND 0.13646f
C8343 Nand_Gate_1.A.t7 GND 0.13313f
C8344 Nand_Gate_1.A.t6 GND 0.1273f
C8345 Nand_Gate_1.A.n3 GND 0.03335f
C8346 Nand_Gate_1.A.n4 GND 0.03059f
C8347 Nand_Gate_1.A.t4 GND 0.24518f
C8348 Nand_Gate_1.A.n5 GND 0.07355f
C8349 Nand_Gate_1.A.t8 GND 0.1273f
C8350 Nand_Gate_1.A.n6 GND 0.03335f
C8351 Nand_Gate_1.A.n7 GND 0.03059f
C8352 Nand_Gate_1.A.n8 GND 0.0774f
C8353 Nand_Gate_1.A.n9 GND 0.0774f
C8354 Nand_Gate_1.A.n10 GND 0.07355f
C8355 Nand_Gate_1.A.t9 GND 0.31308f
C8356 Nand_Gate_1.A.n11 GND 0.07679f
C8357 Nand_Gate_1.A.n12 GND 0.7252f
C8358 Nand_Gate_1.A.n13 GND 0.15555f
C8359 Nand_Gate_1.A.t11 GND 0.24485f
C8360 Nand_Gate_1.A.n14 GND 0.10664f
C8361 Nand_Gate_1.A.t10 GND 0.11428f
C8362 Nand_Gate_1.A.n15 GND 0.0746f
C8363 Nand_Gate_1.A.n16 GND 0.03573f
C8364 Nand_Gate_1.A.n17 GND 0.09059f
C8365 Nand_Gate_1.A.t1 GND 0.03321f
C8366 Nand_Gate_1.A.n18 GND 0.05116f
C8367 Nand_Gate_1.A.t0 GND 0.03391f
C8368 Nand_Gate_1.A.t3 GND 0.03321f
C8369 Nand_Gate_1.A.n19 GND 0.18887f
C8370 Nand_Gate_1.A.n20 GND 0.06163f
C8371 Nand_Gate_1.A.n21 GND 0.12408f
C8372 Ring_Counter_0.D_FlipFlop_15.Qbar.t2 GND 0.05347f
C8373 Ring_Counter_0.D_FlipFlop_15.Qbar.t4 GND 0.41161f
C8374 Ring_Counter_0.D_FlipFlop_15.Qbar.n0 GND 0.1774f
C8375 Ring_Counter_0.D_FlipFlop_15.Qbar.t5 GND 0.18986f
C8376 Ring_Counter_0.D_FlipFlop_15.Qbar.n1 GND 0.23199f
C8377 Ring_Counter_0.D_FlipFlop_15.Qbar.n2 GND 0.05991f
C8378 Ring_Counter_0.D_FlipFlop_15.Qbar.t1 GND 0.05559f
C8379 Ring_Counter_0.D_FlipFlop_15.Qbar.n3 GND 0.09627f
C8380 Ring_Counter_0.D_FlipFlop_15.Qbar.t0 GND 0.05675f
C8381 Ring_Counter_0.D_FlipFlop_15.Qbar.t3 GND 0.05559f
C8382 Ring_Counter_0.D_FlipFlop_15.Qbar.n4 GND 0.31612f
C8383 Ring_Counter_0.D_FlipFlop_15.Qbar.n5 GND 0.16106f
C8384 Ring_Counter_0.D_FlipFlop_15.Qbar.n6 GND 0.15403f
C8385 VDD.n0 GND 0.24808f
C8386 VDD.t510 GND 0.02127f
C8387 VDD.n1 GND 0.07408f
C8388 VDD.n2 GND 0.02503f
C8389 VDD.n3 GND 0.04624f
C8390 VDD.n4 GND 0.02704f
C8391 VDD.n5 GND 0.04624f
C8392 VDD.n6 GND 0.32569f
C8393 VDD.t509 GND 0.3079f
C8394 VDD.t911 GND 0.2823f
C8395 VDD.n8 GND 0.04624f
C8396 VDD.n9 GND 0.04624f
C8397 VDD.n10 GND 0.08322f
C8398 VDD.t314 GND 0.3079f
C8399 VDD.n11 GND 0.04624f
C8400 VDD.n12 GND 0.04624f
C8401 VDD.n13 GND 0.02772f
C8402 VDD.n14 GND 0.03228f
C8403 VDD.t508 GND 0.02796f
C8404 VDD.n15 GND 0.03422f
C8405 VDD.n16 GND 0.07267f
C8406 VDD.t315 GND 0.02326f
C8407 VDD.n17 GND 0.11265f
C8408 VDD.n19 GND 0.02735f
C8409 VDD.t896 GND 0.02127f
C8410 VDD.n20 GND 0.07408f
C8411 VDD.n21 GND 0.02503f
C8412 VDD.n22 GND 0.04624f
C8413 VDD.n23 GND 0.02704f
C8414 VDD.n24 GND 0.04624f
C8415 VDD.n25 GND 0.32569f
C8416 VDD.t895 GND 0.3079f
C8417 VDD.t894 GND 0.2823f
C8418 VDD.n27 GND 0.04624f
C8419 VDD.n28 GND 0.04624f
C8420 VDD.n29 GND 0.08322f
C8421 VDD.t301 GND 0.3079f
C8422 VDD.n30 GND 0.04624f
C8423 VDD.n31 GND 0.04624f
C8424 VDD.n32 GND 0.02772f
C8425 VDD.n33 GND 0.03228f
C8426 VDD.t893 GND 0.02796f
C8427 VDD.n34 GND 0.03422f
C8428 VDD.n35 GND 0.07267f
C8429 VDD.t302 GND 0.02326f
C8430 VDD.n36 GND 0.11265f
C8431 VDD.n38 GND 0.02735f
C8432 VDD.t384 GND 0.02127f
C8433 VDD.n39 GND 0.07408f
C8434 VDD.n40 GND 0.02503f
C8435 VDD.n41 GND 0.04624f
C8436 VDD.n42 GND 0.02704f
C8437 VDD.n43 GND 0.04624f
C8438 VDD.n44 GND 0.32569f
C8439 VDD.t383 GND 0.3079f
C8440 VDD.t427 GND 0.2823f
C8441 VDD.n46 GND 0.04624f
C8442 VDD.n47 GND 0.04624f
C8443 VDD.n48 GND 0.08322f
C8444 VDD.t630 GND 0.3079f
C8445 VDD.n49 GND 0.04624f
C8446 VDD.n50 GND 0.04624f
C8447 VDD.n51 GND 0.02772f
C8448 VDD.n52 GND 0.03228f
C8449 VDD.t382 GND 0.02796f
C8450 VDD.n53 GND 0.03422f
C8451 VDD.n54 GND 0.07267f
C8452 VDD.t631 GND 0.02326f
C8453 VDD.n55 GND 0.11265f
C8454 VDD.n57 GND 0.02735f
C8455 VDD.t715 GND 0.02127f
C8456 VDD.n58 GND 0.07408f
C8457 VDD.n59 GND 0.02503f
C8458 VDD.n60 GND 0.04624f
C8459 VDD.n61 GND 0.02704f
C8460 VDD.n62 GND 0.04624f
C8461 VDD.n63 GND 0.32569f
C8462 VDD.t714 GND 0.3079f
C8463 VDD.t713 GND 0.2823f
C8464 VDD.n65 GND 0.04624f
C8465 VDD.n66 GND 0.04624f
C8466 VDD.n67 GND 0.08322f
C8467 VDD.t402 GND 0.3079f
C8468 VDD.n68 GND 0.04624f
C8469 VDD.n69 GND 0.04624f
C8470 VDD.n70 GND 0.02772f
C8471 VDD.n71 GND 0.03228f
C8472 VDD.t361 GND 0.02796f
C8473 VDD.n72 GND 0.03422f
C8474 VDD.n73 GND 0.07267f
C8475 VDD.t403 GND 0.02326f
C8476 VDD.n74 GND 0.11265f
C8477 VDD.n76 GND 0.02735f
C8478 VDD.t299 GND 0.02127f
C8479 VDD.n77 GND 0.07408f
C8480 VDD.n78 GND 0.02503f
C8481 VDD.n79 GND 0.04624f
C8482 VDD.n80 GND 0.02704f
C8483 VDD.n81 GND 0.04624f
C8484 VDD.n82 GND 0.32569f
C8485 VDD.t298 GND 0.3079f
C8486 VDD.t790 GND 0.2823f
C8487 VDD.n84 GND 0.04624f
C8488 VDD.n85 GND 0.04624f
C8489 VDD.n86 GND 0.08322f
C8490 VDD.t96 GND 0.3079f
C8491 VDD.n87 GND 0.04624f
C8492 VDD.n88 GND 0.04624f
C8493 VDD.n89 GND 0.02772f
C8494 VDD.n90 GND 0.03228f
C8495 VDD.t789 GND 0.02796f
C8496 VDD.n91 GND 0.03422f
C8497 VDD.n92 GND 0.07267f
C8498 VDD.t97 GND 0.02326f
C8499 VDD.n93 GND 0.11265f
C8500 VDD.n95 GND 0.02735f
C8501 VDD.t856 GND 0.02127f
C8502 VDD.n96 GND 0.07408f
C8503 VDD.n97 GND 0.02503f
C8504 VDD.n98 GND 0.04624f
C8505 VDD.n99 GND 0.02704f
C8506 VDD.n100 GND 0.04624f
C8507 VDD.n101 GND 0.32569f
C8508 VDD.t855 GND 0.3079f
C8509 VDD.t866 GND 0.2823f
C8510 VDD.n103 GND 0.04624f
C8511 VDD.n104 GND 0.04624f
C8512 VDD.n105 GND 0.08322f
C8513 VDD.t544 GND 0.3079f
C8514 VDD.n106 GND 0.04624f
C8515 VDD.n107 GND 0.04624f
C8516 VDD.n108 GND 0.02772f
C8517 VDD.n109 GND 0.03228f
C8518 VDD.t853 GND 0.02796f
C8519 VDD.n110 GND 0.03422f
C8520 VDD.n111 GND 0.07267f
C8521 VDD.t545 GND 0.02326f
C8522 VDD.n112 GND 0.11265f
C8523 VDD.n114 GND 0.02735f
C8524 VDD.t904 GND 0.02127f
C8525 VDD.n115 GND 0.07408f
C8526 VDD.n116 GND 0.02503f
C8527 VDD.n117 GND 0.04624f
C8528 VDD.n118 GND 0.02704f
C8529 VDD.n119 GND 0.04624f
C8530 VDD.n120 GND 0.32569f
C8531 VDD.t903 GND 0.3079f
C8532 VDD.t905 GND 0.2823f
C8533 VDD.n122 GND 0.04624f
C8534 VDD.n123 GND 0.04624f
C8535 VDD.n124 GND 0.08322f
C8536 VDD.t880 GND 0.3079f
C8537 VDD.n125 GND 0.04624f
C8538 VDD.n126 GND 0.04624f
C8539 VDD.n127 GND 0.02772f
C8540 VDD.n128 GND 0.03228f
C8541 VDD.t448 GND 0.02796f
C8542 VDD.n129 GND 0.03422f
C8543 VDD.n130 GND 0.07267f
C8544 VDD.t881 GND 0.02326f
C8545 VDD.n131 GND 0.11265f
C8546 VDD.n133 GND 0.02735f
C8547 VDD.t774 GND 0.02127f
C8548 VDD.n134 GND 0.07408f
C8549 VDD.n135 GND 0.02503f
C8550 VDD.n136 GND 0.04624f
C8551 VDD.n137 GND 0.02704f
C8552 VDD.n138 GND 0.04624f
C8553 VDD.n139 GND 0.32569f
C8554 VDD.t773 GND 0.3079f
C8555 VDD.t776 GND 0.2823f
C8556 VDD.n141 GND 0.04624f
C8557 VDD.n142 GND 0.04624f
C8558 VDD.n143 GND 0.08322f
C8559 VDD.t915 GND 0.3079f
C8560 VDD.n144 GND 0.04624f
C8561 VDD.n145 GND 0.04624f
C8562 VDD.n146 GND 0.02772f
C8563 VDD.n147 GND 0.03228f
C8564 VDD.t775 GND 0.02796f
C8565 VDD.n148 GND 0.03422f
C8566 VDD.n149 GND 0.07267f
C8567 VDD.t916 GND 0.02326f
C8568 VDD.n150 GND 0.11265f
C8569 VDD.n152 GND 0.02735f
C8570 VDD.t967 GND 0.15539f
C8571 VDD.n153 GND 0.06697f
C8572 VDD.t209 GND 0.0709f
C8573 VDD.n154 GND 0.26868f
C8574 VDD.n155 GND 0.44145f
C8575 VDD.n156 GND 1.0093f
C8576 VDD.t954 GND 0.15509f
C8577 VDD.n157 GND 0.05006f
C8578 VDD.t189 GND 0.08044f
C8579 VDD.n158 GND 0.01731f
C8580 VDD.n159 GND 0.01034f
C8581 VDD.n160 GND 0.09595f
C8582 VDD.t947 GND 0.15509f
C8583 VDD.n161 GND 0.05006f
C8584 VDD.t196 GND 0.08044f
C8585 VDD.n162 GND 0.01731f
C8586 VDD.n163 GND 0.01034f
C8587 VDD.n165 GND 0.24903f
C8588 VDD.n166 GND 0.36089f
C8589 VDD.n167 GND 0.07705f
C8590 VDD.n168 GND 0.04255f
C8591 VDD.n169 GND 0.05152f
C8592 VDD.t897 GND 0.02114f
C8593 VDD.t219 GND 0.02114f
C8594 VDD.n170 GND 0.14059f
C8595 VDD.n171 GND 0.04891f
C8596 VDD.n172 GND 0.04648f
C8597 VDD.n173 GND 0.04891f
C8598 VDD.n174 GND 0.04532f
C8599 VDD.n175 GND 0.04532f
C8600 VDD.t190 GND 4.12913f
C8601 VDD.n176 GND 0.04648f
C8602 VDD.n177 GND 0.04648f
C8603 VDD.n178 GND 0.04648f
C8604 VDD.n179 GND 0.04648f
C8605 VDD.n180 GND 0.04648f
C8606 VDD.n181 GND 0.04648f
C8607 VDD.n182 GND 3.47277f
C8608 VDD.n183 GND 0.04648f
C8609 VDD.n184 GND 0.04648f
C8610 VDD.n185 GND 0.04648f
C8611 VDD.n186 GND 0.04648f
C8612 VDD.n187 GND 0.04532f
C8613 VDD.n188 GND 0.04532f
C8614 VDD.n189 GND 0.02497f
C8615 VDD.n190 GND 0.02497f
C8616 VDD.t220 GND 0.02104f
C8617 VDD.n191 GND 0.22365f
C8618 VDD.t690 GND 0.02104f
C8619 VDD.t102 GND 0.02104f
C8620 VDD.n192 GND 0.04891f
C8621 VDD.n193 GND 0.04891f
C8622 VDD.n194 GND 0.04532f
C8623 VDD.n195 GND 0.04648f
C8624 VDD.n196 GND 0.02293f
C8625 VDD.n197 GND 0.02708f
C8626 VDD.n198 GND 0.02293f
C8627 VDD.n199 GND 0.04532f
C8628 VDD.n200 GND 0.04532f
C8629 VDD.n201 GND 0.04532f
C8630 VDD.n202 GND 0.04532f
C8631 VDD.n203 GND 0.04532f
C8632 VDD.n204 GND 0.04532f
C8633 VDD.n205 GND 0.04532f
C8634 VDD.n206 GND 0.04532f
C8635 VDD.n207 GND 0.04532f
C8636 VDD.n208 GND 0.04532f
C8637 VDD.n209 GND 0.04532f
C8638 VDD.n210 GND 0.04532f
C8639 VDD.n211 GND 0.04532f
C8640 VDD.n212 GND 0.04532f
C8641 VDD.n213 GND 0.04532f
C8642 VDD.n214 GND 0.04532f
C8643 VDD.n215 GND 0.04532f
C8644 VDD.n216 GND 0.04532f
C8645 VDD.n217 GND 0.04532f
C8646 VDD.n218 GND 0.04532f
C8647 VDD.n219 GND 0.02293f
C8648 VDD.n220 GND 0.02293f
C8649 VDD.n221 GND 0.02708f
C8650 VDD.n222 GND 0.04648f
C8651 VDD.n223 GND 3.19829f
C8652 VDD.n224 GND 0.04532f
C8653 VDD.n225 GND 0.04648f
C8654 VDD.n226 GND 0.04648f
C8655 VDD.n227 GND 0.04891f
C8656 VDD.n228 GND 0.02293f
C8657 VDD.t641 GND 0.02114f
C8658 VDD.t876 GND 0.02114f
C8659 VDD.t800 GND 0.02114f
C8660 VDD.t607 GND 0.02114f
C8661 VDD.n229 GND 0.02324f
C8662 VDD.n230 GND 0.04891f
C8663 VDD.n231 GND 0.04648f
C8664 VDD.n232 GND 0.02293f
C8665 VDD.n233 GND 0.04648f
C8666 VDD.n234 GND 0.02708f
C8667 VDD.n235 GND 0.02293f
C8668 VDD.n236 GND 0.02708f
C8669 VDD.n237 GND 0.02293f
C8670 VDD.n238 GND 0.04532f
C8671 VDD.n239 GND 0.04532f
C8672 VDD.n240 GND 0.04532f
C8673 VDD.n241 GND 0.02293f
C8674 VDD.n242 GND 0.02293f
C8675 VDD.n243 GND 0.02708f
C8676 VDD.n244 GND 0.04648f
C8677 VDD.n245 GND 0.04648f
C8678 VDD.n246 GND 0.04648f
C8679 VDD.n247 GND 0.04648f
C8680 VDD.n248 GND 0.04532f
C8681 VDD.n249 GND 0.04532f
C8682 VDD.n250 GND 0.02293f
C8683 VDD.n251 GND 0.02293f
C8684 VDD.n252 GND 0.04648f
C8685 VDD.n253 GND 0.02708f
C8686 VDD.n254 GND 0.02293f
C8687 VDD.n255 GND 0.04891f
C8688 VDD.n256 GND 0.04648f
C8689 VDD.n257 GND 0.05737f
C8690 VDD.n258 GND 0.04891f
C8691 VDD.n259 GND 0.02293f
C8692 VDD.n260 GND 0.02708f
C8693 VDD.n261 GND 0.04648f
C8694 VDD.n262 GND 0.04532f
C8695 VDD.n263 GND 0.04532f
C8696 VDD.n264 GND 0.02293f
C8697 VDD.n265 GND 0.02708f
C8698 VDD.n266 GND 0.04648f
C8699 VDD.n267 GND 0.04648f
C8700 VDD.n268 GND 0.04648f
C8701 VDD.n269 GND 0.04532f
C8702 VDD.n270 GND 0.04532f
C8703 VDD.n271 GND 0.02293f
C8704 VDD.n272 GND 0.02293f
C8705 VDD.n273 GND 0.04648f
C8706 VDD.n274 GND 0.02708f
C8707 VDD.n275 GND 0.02293f
C8708 VDD.n276 GND 0.04891f
C8709 VDD.n277 GND 0.04648f
C8710 VDD.t654 GND 0.02104f
C8711 VDD.t197 GND 0.02104f
C8712 VDD.t815 GND 0.02114f
C8713 VDD.t251 GND 0.02114f
C8714 VDD.n278 GND 0.44561f
C8715 VDD.n279 GND 0.04891f
C8716 VDD.n280 GND 0.04648f
C8717 VDD.n281 GND 0.02293f
C8718 VDD.n282 GND 0.04648f
C8719 VDD.n283 GND 0.02708f
C8720 VDD.n284 GND 0.02293f
C8721 VDD.n285 GND 0.04532f
C8722 VDD.n286 GND 0.02293f
C8723 VDD.n287 GND 0.02708f
C8724 VDD.n288 GND 0.04532f
C8725 VDD.n289 GND 0.02293f
C8726 VDD.n290 GND 0.04891f
C8727 VDD.n291 GND 0.05737f
C8728 VDD.n292 GND 0.02055f
C8729 VDD.n293 GND 0.08471f
C8730 VDD.n294 GND 0.95576f
C8731 VDD.t771 GND 0.02114f
C8732 VDD.t362 GND 0.02114f
C8733 VDD.t447 GND 0.02114f
C8734 VDD.t844 GND 0.02114f
C8735 VDD.t248 GND 0.02104f
C8736 VDD.t845 GND 0.02114f
C8737 VDD.t446 GND 0.02114f
C8738 VDD.t434 GND 0.02114f
C8739 VDD.t435 GND 0.02114f
C8740 VDD.t699 GND 0.02104f
C8741 VDD.t191 GND 0.02104f
C8742 VDD.n295 GND 0.95576f
C8743 VDD.n296 GND 0.08471f
C8744 VDD.n297 GND 0.04891f
C8745 VDD.n298 GND 0.04648f
C8746 VDD.n299 GND 0.02293f
C8747 VDD.n300 GND 0.04648f
C8748 VDD.n301 GND 0.02708f
C8749 VDD.n302 GND 0.02293f
C8750 VDD.n303 GND 0.04532f
C8751 VDD.n304 GND 0.02293f
C8752 VDD.n305 GND 0.02708f
C8753 VDD.n306 GND 0.04532f
C8754 VDD.n307 GND 0.02293f
C8755 VDD.n308 GND 0.04891f
C8756 VDD.n309 GND 0.05737f
C8757 VDD.n310 GND 0.02055f
C8758 VDD.n311 GND 0.44561f
C8759 VDD.n312 GND 0.14059f
C8760 VDD.n313 GND 0.04891f
C8761 VDD.n314 GND 0.04648f
C8762 VDD.n315 GND 0.02293f
C8763 VDD.n316 GND 0.04648f
C8764 VDD.n317 GND 0.02708f
C8765 VDD.n318 GND 0.02293f
C8766 VDD.n319 GND 0.04532f
C8767 VDD.n320 GND 0.02293f
C8768 VDD.n321 GND 0.02708f
C8769 VDD.n322 GND 0.04532f
C8770 VDD.n323 GND 0.02293f
C8771 VDD.n324 GND 0.04891f
C8772 VDD.n325 GND 0.05737f
C8773 VDD.n326 GND 0.02055f
C8774 VDD.n327 GND 0.02497f
C8775 VDD.n328 GND 0.04648f
C8776 VDD.n329 GND 0.04648f
C8777 VDD.n330 GND 0.02708f
C8778 VDD.n331 GND 0.02497f
C8779 VDD.n332 GND 0.08328f
C8780 VDD.n333 GND 0.01566f
C8781 VDD.n334 GND 0.18236f
C8782 VDD.n335 GND 0.03549f
C8783 VDD.n336 GND 0.04891f
C8784 VDD.n337 GND 0.04648f
C8785 VDD.n338 GND 0.02293f
C8786 VDD.n339 GND 0.04648f
C8787 VDD.n340 GND 0.02708f
C8788 VDD.n341 GND 0.02293f
C8789 VDD.n342 GND 0.04532f
C8790 VDD.n343 GND 0.02293f
C8791 VDD.n344 GND 0.02708f
C8792 VDD.n345 GND 0.04532f
C8793 VDD.n346 GND 0.02293f
C8794 VDD.n347 GND 0.04891f
C8795 VDD.n348 GND 0.05737f
C8796 VDD.n349 GND 0.02055f
C8797 VDD.n350 GND 0.44561f
C8798 VDD.n351 GND 0.14059f
C8799 VDD.n352 GND 0.04891f
C8800 VDD.n353 GND 0.04648f
C8801 VDD.n354 GND 0.02293f
C8802 VDD.n355 GND 0.04648f
C8803 VDD.n356 GND 0.02708f
C8804 VDD.n357 GND 0.02293f
C8805 VDD.n358 GND 0.04532f
C8806 VDD.n359 GND 0.02293f
C8807 VDD.n360 GND 0.02708f
C8808 VDD.n361 GND 0.04532f
C8809 VDD.n362 GND 0.02293f
C8810 VDD.n363 GND 0.04891f
C8811 VDD.n364 GND 0.05737f
C8812 VDD.n365 GND 0.02813f
C8813 VDD.n366 GND 0.02324f
C8814 VDD.n367 GND 0.05737f
C8815 VDD.n368 GND 0.04891f
C8816 VDD.n369 GND 0.02293f
C8817 VDD.n370 GND 0.02708f
C8818 VDD.n371 GND 0.04648f
C8819 VDD.n372 GND 0.02293f
C8820 VDD.n373 GND 0.02293f
C8821 VDD.n374 GND 0.02708f
C8822 VDD.n375 GND 0.04648f
C8823 VDD.n376 GND 0.02708f
C8824 VDD.n377 GND 0.04648f
C8825 VDD.n378 GND 3.19829f
C8826 VDD.n379 GND 0.04648f
C8827 VDD.n380 GND 0.04532f
C8828 VDD.n381 GND 0.02293f
C8829 VDD.n382 GND 0.04891f
C8830 VDD.n383 GND 0.05737f
C8831 VDD.n384 GND 0.02813f
C8832 VDD.n385 GND 0.14059f
C8833 VDD.n386 GND 0.44561f
C8834 VDD.n387 GND 0.02055f
C8835 VDD.n388 GND 0.05737f
C8836 VDD.n389 GND 0.04891f
C8837 VDD.n390 GND 0.02293f
C8838 VDD.n391 GND 0.02708f
C8839 VDD.n392 GND 0.02293f
C8840 VDD.n393 GND 0.04532f
C8841 VDD.t101 GND 4.12913f
C8842 VDD.n394 GND 0.04532f
C8843 VDD.n395 GND 0.04648f
C8844 VDD.n396 GND 0.05737f
C8845 VDD.n398 GND 0.95576f
C8846 VDD.n399 GND 0.08471f
C8847 VDD.n400 GND 0.01566f
C8848 VDD.n401 GND 0.08328f
C8849 VDD.n402 GND 0.04648f
C8850 VDD.n403 GND 3.47277f
C8851 VDD.n404 GND 0.04648f
C8852 VDD.n405 GND 0.05737f
C8853 VDD.n406 GND 0.02177f
C8854 VDD.n407 GND 0.07516f
C8855 VDD.n410 GND 0.01801f
C8856 VDD.t964 GND 0.15471f
C8857 VDD.n412 GND 0.06739f
C8858 VDD.t100 GND 0.07116f
C8859 VDD.n413 GND 0.17412f
C8860 VDD.n414 GND 0.18182f
C8861 VDD.n415 GND 0.06121f
C8862 VDD.n416 GND 0.04255f
C8863 VDD.n417 GND 0.05152f
C8864 VDD.t848 GND 0.02114f
C8865 VDD.t387 GND 0.02114f
C8866 VDD.n418 GND 0.14059f
C8867 VDD.n419 GND 0.04891f
C8868 VDD.n420 GND 0.04648f
C8869 VDD.n421 GND 0.04891f
C8870 VDD.n422 GND 0.04532f
C8871 VDD.n423 GND 0.04532f
C8872 VDD.t210 GND 4.12913f
C8873 VDD.n424 GND 0.04648f
C8874 VDD.n425 GND 0.04648f
C8875 VDD.n426 GND 0.04648f
C8876 VDD.n427 GND 0.04648f
C8877 VDD.n428 GND 0.04648f
C8878 VDD.n429 GND 0.04648f
C8879 VDD.n430 GND 3.47277f
C8880 VDD.n431 GND 0.04648f
C8881 VDD.n432 GND 0.04648f
C8882 VDD.n433 GND 0.04648f
C8883 VDD.n434 GND 0.04648f
C8884 VDD.n435 GND 0.04532f
C8885 VDD.n436 GND 0.04532f
C8886 VDD.n437 GND 0.02497f
C8887 VDD.n438 GND 0.02497f
C8888 VDD.t642 GND 0.02104f
C8889 VDD.n439 GND 0.22365f
C8890 VDD.t211 GND 0.02104f
C8891 VDD.t662 GND 0.02104f
C8892 VDD.n440 GND 0.04891f
C8893 VDD.n441 GND 0.04891f
C8894 VDD.n442 GND 0.04532f
C8895 VDD.n443 GND 0.04648f
C8896 VDD.n444 GND 0.02293f
C8897 VDD.n445 GND 0.02708f
C8898 VDD.n446 GND 0.02293f
C8899 VDD.n447 GND 0.04532f
C8900 VDD.n448 GND 0.04532f
C8901 VDD.n449 GND 0.04532f
C8902 VDD.n450 GND 0.04532f
C8903 VDD.n451 GND 0.04532f
C8904 VDD.n452 GND 0.04532f
C8905 VDD.n453 GND 0.04532f
C8906 VDD.n454 GND 0.04532f
C8907 VDD.n455 GND 0.04532f
C8908 VDD.n456 GND 0.04532f
C8909 VDD.n457 GND 0.04532f
C8910 VDD.n458 GND 0.04532f
C8911 VDD.n459 GND 0.04532f
C8912 VDD.n460 GND 0.04532f
C8913 VDD.n461 GND 0.04532f
C8914 VDD.n462 GND 0.04532f
C8915 VDD.n463 GND 0.04532f
C8916 VDD.n464 GND 0.04532f
C8917 VDD.n465 GND 0.04532f
C8918 VDD.n466 GND 0.04532f
C8919 VDD.n467 GND 0.02293f
C8920 VDD.n468 GND 0.02293f
C8921 VDD.n469 GND 0.02708f
C8922 VDD.n470 GND 0.04648f
C8923 VDD.n471 GND 3.19829f
C8924 VDD.n472 GND 0.04532f
C8925 VDD.n473 GND 0.04648f
C8926 VDD.n474 GND 0.04648f
C8927 VDD.n475 GND 0.04891f
C8928 VDD.n476 GND 0.02293f
C8929 VDD.t339 GND 0.02114f
C8930 VDD.t886 GND 0.02114f
C8931 VDD.t606 GND 0.02114f
C8932 VDD.t634 GND 0.02114f
C8933 VDD.n477 GND 0.02324f
C8934 VDD.n478 GND 0.04891f
C8935 VDD.n479 GND 0.04648f
C8936 VDD.n480 GND 0.02293f
C8937 VDD.n481 GND 0.04648f
C8938 VDD.n482 GND 0.02708f
C8939 VDD.n483 GND 0.02293f
C8940 VDD.n484 GND 0.02708f
C8941 VDD.n485 GND 0.02293f
C8942 VDD.n486 GND 0.04532f
C8943 VDD.n487 GND 0.04532f
C8944 VDD.n488 GND 0.04532f
C8945 VDD.n489 GND 0.02293f
C8946 VDD.n490 GND 0.02293f
C8947 VDD.n491 GND 0.02708f
C8948 VDD.n492 GND 0.04648f
C8949 VDD.n493 GND 0.04648f
C8950 VDD.n494 GND 0.04648f
C8951 VDD.n495 GND 0.04648f
C8952 VDD.n496 GND 0.04532f
C8953 VDD.n497 GND 0.04532f
C8954 VDD.n498 GND 0.02293f
C8955 VDD.n499 GND 0.02293f
C8956 VDD.n500 GND 0.04648f
C8957 VDD.n501 GND 0.02708f
C8958 VDD.n502 GND 0.02293f
C8959 VDD.n503 GND 0.04891f
C8960 VDD.n504 GND 0.04648f
C8961 VDD.n505 GND 0.05737f
C8962 VDD.n506 GND 0.04891f
C8963 VDD.n507 GND 0.02293f
C8964 VDD.n508 GND 0.02708f
C8965 VDD.n509 GND 0.04648f
C8966 VDD.n510 GND 0.04532f
C8967 VDD.n511 GND 0.04532f
C8968 VDD.n512 GND 0.02293f
C8969 VDD.n513 GND 0.02708f
C8970 VDD.n514 GND 0.04648f
C8971 VDD.n515 GND 0.04648f
C8972 VDD.n516 GND 0.04648f
C8973 VDD.n517 GND 0.04532f
C8974 VDD.n518 GND 0.04532f
C8975 VDD.n519 GND 0.02293f
C8976 VDD.n520 GND 0.02293f
C8977 VDD.n521 GND 0.04648f
C8978 VDD.n522 GND 0.02708f
C8979 VDD.n523 GND 0.02293f
C8980 VDD.n524 GND 0.04891f
C8981 VDD.n525 GND 0.04648f
C8982 VDD.t145 GND 0.02104f
C8983 VDD.t651 GND 0.02104f
C8984 VDD.t226 GND 0.02114f
C8985 VDD.t818 GND 0.02114f
C8986 VDD.n526 GND 0.44561f
C8987 VDD.n527 GND 0.04891f
C8988 VDD.n528 GND 0.04648f
C8989 VDD.n529 GND 0.02293f
C8990 VDD.n530 GND 0.04648f
C8991 VDD.n531 GND 0.02708f
C8992 VDD.n532 GND 0.02293f
C8993 VDD.n533 GND 0.04532f
C8994 VDD.n534 GND 0.02293f
C8995 VDD.n535 GND 0.02708f
C8996 VDD.n536 GND 0.04532f
C8997 VDD.n537 GND 0.02293f
C8998 VDD.n538 GND 0.04891f
C8999 VDD.n539 GND 0.05737f
C9000 VDD.n540 GND 0.02055f
C9001 VDD.n541 GND 0.08471f
C9002 VDD.n542 GND 0.95576f
C9003 VDD.t342 GND 0.02114f
C9004 VDD.t313 GND 0.02114f
C9005 VDD.t399 GND 0.02114f
C9006 VDD.t707 GND 0.02114f
C9007 VDD.t235 GND 0.02104f
C9008 VDD.t708 GND 0.02114f
C9009 VDD.t762 GND 0.02114f
C9010 VDD.t620 GND 0.02114f
C9011 VDD.t462 GND 0.02114f
C9012 VDD.t107 GND 0.02104f
C9013 VDD.t694 GND 0.02104f
C9014 VDD.n543 GND 0.95576f
C9015 VDD.n544 GND 0.08471f
C9016 VDD.n545 GND 0.04891f
C9017 VDD.n546 GND 0.04648f
C9018 VDD.n547 GND 0.02293f
C9019 VDD.n548 GND 0.04648f
C9020 VDD.n549 GND 0.02708f
C9021 VDD.n550 GND 0.02293f
C9022 VDD.n551 GND 0.04532f
C9023 VDD.n552 GND 0.02293f
C9024 VDD.n553 GND 0.02708f
C9025 VDD.n554 GND 0.04532f
C9026 VDD.n555 GND 0.02293f
C9027 VDD.n556 GND 0.04891f
C9028 VDD.n557 GND 0.05737f
C9029 VDD.n558 GND 0.02055f
C9030 VDD.n559 GND 0.44561f
C9031 VDD.n560 GND 0.14059f
C9032 VDD.n561 GND 0.04891f
C9033 VDD.n562 GND 0.04648f
C9034 VDD.n563 GND 0.02293f
C9035 VDD.n564 GND 0.04648f
C9036 VDD.n565 GND 0.02708f
C9037 VDD.n566 GND 0.02293f
C9038 VDD.n567 GND 0.04532f
C9039 VDD.n568 GND 0.02293f
C9040 VDD.n569 GND 0.02708f
C9041 VDD.n570 GND 0.04532f
C9042 VDD.n571 GND 0.02293f
C9043 VDD.n572 GND 0.04891f
C9044 VDD.n573 GND 0.05737f
C9045 VDD.n574 GND 0.02055f
C9046 VDD.n575 GND 0.02497f
C9047 VDD.n576 GND 0.04648f
C9048 VDD.n577 GND 0.04648f
C9049 VDD.n578 GND 0.02708f
C9050 VDD.n579 GND 0.02497f
C9051 VDD.n580 GND 0.08328f
C9052 VDD.n581 GND 0.01566f
C9053 VDD.n582 GND 0.18236f
C9054 VDD.n583 GND 0.03549f
C9055 VDD.n584 GND 0.04891f
C9056 VDD.n585 GND 0.04648f
C9057 VDD.n586 GND 0.02293f
C9058 VDD.n587 GND 0.04648f
C9059 VDD.n588 GND 0.02708f
C9060 VDD.n589 GND 0.02293f
C9061 VDD.n590 GND 0.04532f
C9062 VDD.n591 GND 0.02293f
C9063 VDD.n592 GND 0.02708f
C9064 VDD.n593 GND 0.04532f
C9065 VDD.n594 GND 0.02293f
C9066 VDD.n595 GND 0.04891f
C9067 VDD.n596 GND 0.05737f
C9068 VDD.n597 GND 0.02055f
C9069 VDD.n598 GND 0.44561f
C9070 VDD.n599 GND 0.14059f
C9071 VDD.n600 GND 0.04891f
C9072 VDD.n601 GND 0.04648f
C9073 VDD.n602 GND 0.02293f
C9074 VDD.n603 GND 0.04648f
C9075 VDD.n604 GND 0.02708f
C9076 VDD.n605 GND 0.02293f
C9077 VDD.n606 GND 0.04532f
C9078 VDD.n607 GND 0.02293f
C9079 VDD.n608 GND 0.02708f
C9080 VDD.n609 GND 0.04532f
C9081 VDD.n610 GND 0.02293f
C9082 VDD.n611 GND 0.04891f
C9083 VDD.n612 GND 0.05737f
C9084 VDD.n613 GND 0.02813f
C9085 VDD.n614 GND 0.02324f
C9086 VDD.n615 GND 0.05737f
C9087 VDD.n616 GND 0.04891f
C9088 VDD.n617 GND 0.02293f
C9089 VDD.n618 GND 0.02708f
C9090 VDD.n619 GND 0.04648f
C9091 VDD.n620 GND 0.02293f
C9092 VDD.n621 GND 0.02293f
C9093 VDD.n622 GND 0.02708f
C9094 VDD.n623 GND 0.04648f
C9095 VDD.n624 GND 0.02708f
C9096 VDD.n625 GND 0.04648f
C9097 VDD.n626 GND 3.19829f
C9098 VDD.n627 GND 0.04648f
C9099 VDD.n628 GND 0.04532f
C9100 VDD.n629 GND 0.02293f
C9101 VDD.n630 GND 0.04891f
C9102 VDD.n631 GND 0.05737f
C9103 VDD.n632 GND 0.02813f
C9104 VDD.n633 GND 0.14059f
C9105 VDD.n634 GND 0.44561f
C9106 VDD.n635 GND 0.02055f
C9107 VDD.n636 GND 0.05737f
C9108 VDD.n637 GND 0.04891f
C9109 VDD.n638 GND 0.02293f
C9110 VDD.n639 GND 0.02708f
C9111 VDD.n640 GND 0.02293f
C9112 VDD.n641 GND 0.04532f
C9113 VDD.t106 GND 4.12913f
C9114 VDD.n642 GND 0.04532f
C9115 VDD.n643 GND 0.04648f
C9116 VDD.n644 GND 0.05737f
C9117 VDD.n645 GND 0.01303f
C9118 VDD.n646 GND 0.95576f
C9119 VDD.n647 GND 0.08471f
C9120 VDD.n648 GND 0.01566f
C9121 VDD.n649 GND 0.08328f
C9122 VDD.n650 GND 0.04648f
C9123 VDD.n651 GND 3.47277f
C9124 VDD.n652 GND 0.04648f
C9125 VDD.n653 GND 0.05737f
C9126 VDD.n654 GND 0.0171f
C9127 VDD.n655 GND 0.064f
C9128 VDD.n658 GND 0.06555f
C9129 VDD.n659 GND 0.03083f
C9130 VDD.t105 GND 0.08047f
C9131 VDD.n660 GND 0.03534f
C9132 VDD.t955 GND 0.15471f
C9133 VDD.n661 GND 0.03238f
C9134 VDD.n662 GND 0.02607f
C9135 VDD.n663 GND 0.09595f
C9136 VDD.t144 GND 0.08047f
C9137 VDD.n664 GND 0.03534f
C9138 VDD.t948 GND 0.15471f
C9139 VDD.n665 GND 0.03238f
C9140 VDD.n666 GND 0.02607f
C9141 VDD.n668 GND 0.24365f
C9142 VDD.n669 GND 0.03496f
C9143 VDD.n670 GND 2.50355f
C9144 VDD.n671 GND 2.18575f
C9145 VDD.t929 GND 0.15539f
C9146 VDD.n672 GND 0.06697f
C9147 VDD.t122 GND 0.07226f
C9148 VDD.n673 GND 0.05627f
C9149 VDD.n674 GND 0.05442f
C9150 VDD.n675 GND 0.04255f
C9151 VDD.n676 GND 0.05152f
C9152 VDD.t709 GND 0.02114f
C9153 VDD.t329 GND 0.02114f
C9154 VDD.n677 GND 0.14059f
C9155 VDD.n678 GND 0.04891f
C9156 VDD.n679 GND 0.04648f
C9157 VDD.n680 GND 0.04891f
C9158 VDD.n681 GND 0.04532f
C9159 VDD.n682 GND 0.04532f
C9160 VDD.t123 GND 4.12913f
C9161 VDD.n683 GND 0.04648f
C9162 VDD.n684 GND 0.04648f
C9163 VDD.n685 GND 0.04648f
C9164 VDD.n686 GND 0.04648f
C9165 VDD.n687 GND 0.04648f
C9166 VDD.n688 GND 0.04648f
C9167 VDD.n689 GND 3.47277f
C9168 VDD.n690 GND 0.04648f
C9169 VDD.n691 GND 0.04648f
C9170 VDD.n692 GND 0.04648f
C9171 VDD.n693 GND 0.04648f
C9172 VDD.n694 GND 0.04532f
C9173 VDD.n695 GND 0.04532f
C9174 VDD.n696 GND 0.02497f
C9175 VDD.n697 GND 0.02497f
C9176 VDD.t338 GND 0.02104f
C9177 VDD.n698 GND 0.22365f
C9178 VDD.t124 GND 0.02104f
C9179 VDD.t653 GND 0.02104f
C9180 VDD.n699 GND 0.04891f
C9181 VDD.n700 GND 0.04891f
C9182 VDD.n701 GND 0.04532f
C9183 VDD.n702 GND 0.04648f
C9184 VDD.n703 GND 0.02293f
C9185 VDD.n704 GND 0.02708f
C9186 VDD.n705 GND 0.02293f
C9187 VDD.n706 GND 0.04532f
C9188 VDD.n707 GND 0.04532f
C9189 VDD.n708 GND 0.04532f
C9190 VDD.n709 GND 0.04532f
C9191 VDD.n710 GND 0.04532f
C9192 VDD.n711 GND 0.04532f
C9193 VDD.n712 GND 0.04532f
C9194 VDD.n713 GND 0.04532f
C9195 VDD.n714 GND 0.04532f
C9196 VDD.n715 GND 0.04532f
C9197 VDD.n716 GND 0.04532f
C9198 VDD.n717 GND 0.04532f
C9199 VDD.n718 GND 0.04532f
C9200 VDD.n719 GND 0.04532f
C9201 VDD.n720 GND 0.04532f
C9202 VDD.n721 GND 0.04532f
C9203 VDD.n722 GND 0.04532f
C9204 VDD.n723 GND 0.04532f
C9205 VDD.n724 GND 0.04532f
C9206 VDD.n725 GND 0.04532f
C9207 VDD.n726 GND 0.02293f
C9208 VDD.n727 GND 0.02293f
C9209 VDD.n728 GND 0.02708f
C9210 VDD.n729 GND 0.04648f
C9211 VDD.n730 GND 3.19829f
C9212 VDD.n731 GND 0.04532f
C9213 VDD.n732 GND 0.04648f
C9214 VDD.n733 GND 0.04648f
C9215 VDD.n734 GND 0.04891f
C9216 VDD.n735 GND 0.02293f
C9217 VDD.t858 GND 0.02114f
C9218 VDD.t525 GND 0.02114f
C9219 VDD.t345 GND 0.02114f
C9220 VDD.t923 GND 0.02114f
C9221 VDD.n736 GND 0.02324f
C9222 VDD.n737 GND 0.04891f
C9223 VDD.n738 GND 0.04648f
C9224 VDD.n739 GND 0.02293f
C9225 VDD.n740 GND 0.04648f
C9226 VDD.n741 GND 0.02708f
C9227 VDD.n742 GND 0.02293f
C9228 VDD.n743 GND 0.02708f
C9229 VDD.n744 GND 0.02293f
C9230 VDD.n745 GND 0.04532f
C9231 VDD.n746 GND 0.04532f
C9232 VDD.n747 GND 0.04532f
C9233 VDD.n748 GND 0.02293f
C9234 VDD.n749 GND 0.02293f
C9235 VDD.n750 GND 0.02708f
C9236 VDD.n751 GND 0.04648f
C9237 VDD.n752 GND 0.04648f
C9238 VDD.n753 GND 0.04648f
C9239 VDD.n754 GND 0.04648f
C9240 VDD.n755 GND 0.04532f
C9241 VDD.n756 GND 0.04532f
C9242 VDD.n757 GND 0.02293f
C9243 VDD.n758 GND 0.02293f
C9244 VDD.n759 GND 0.04648f
C9245 VDD.n760 GND 0.02708f
C9246 VDD.n761 GND 0.02293f
C9247 VDD.n762 GND 0.04891f
C9248 VDD.n763 GND 0.04648f
C9249 VDD.n764 GND 0.05737f
C9250 VDD.n765 GND 0.04891f
C9251 VDD.n766 GND 0.02293f
C9252 VDD.n767 GND 0.02708f
C9253 VDD.n768 GND 0.04648f
C9254 VDD.n769 GND 0.04532f
C9255 VDD.n770 GND 0.04532f
C9256 VDD.n771 GND 0.02293f
C9257 VDD.n772 GND 0.02708f
C9258 VDD.n773 GND 0.04648f
C9259 VDD.n774 GND 0.04648f
C9260 VDD.n775 GND 0.04648f
C9261 VDD.n776 GND 0.04532f
C9262 VDD.n777 GND 0.04532f
C9263 VDD.n778 GND 0.02293f
C9264 VDD.n779 GND 0.02293f
C9265 VDD.n780 GND 0.04648f
C9266 VDD.n781 GND 0.02708f
C9267 VDD.n782 GND 0.02293f
C9268 VDD.n783 GND 0.04891f
C9269 VDD.n784 GND 0.04648f
C9270 VDD.t127 GND 0.02104f
C9271 VDD.t667 GND 0.02104f
C9272 VDD.t809 GND 0.02114f
C9273 VDD.t228 GND 0.02114f
C9274 VDD.n785 GND 0.44561f
C9275 VDD.n786 GND 0.04891f
C9276 VDD.n787 GND 0.04648f
C9277 VDD.n788 GND 0.02293f
C9278 VDD.n789 GND 0.04648f
C9279 VDD.n790 GND 0.02708f
C9280 VDD.n791 GND 0.02293f
C9281 VDD.n792 GND 0.04532f
C9282 VDD.n793 GND 0.02293f
C9283 VDD.n794 GND 0.02708f
C9284 VDD.n795 GND 0.04532f
C9285 VDD.n796 GND 0.02293f
C9286 VDD.n797 GND 0.04891f
C9287 VDD.n798 GND 0.05737f
C9288 VDD.n799 GND 0.02055f
C9289 VDD.n800 GND 0.08471f
C9290 VDD.n801 GND 0.95576f
C9291 VDD.t497 GND 0.02114f
C9292 VDD.t511 GND 0.02114f
C9293 VDD.t602 GND 0.02114f
C9294 VDD.t807 GND 0.02114f
C9295 VDD.t746 GND 0.02104f
C9296 VDD.t803 GND 0.02114f
C9297 VDD.t328 GND 0.02114f
C9298 VDD.t498 GND 0.02114f
C9299 VDD.t273 GND 0.02114f
C9300 VDD.t208 GND 0.02104f
C9301 VDD.t650 GND 0.02104f
C9302 VDD.n802 GND 0.95576f
C9303 VDD.n803 GND 0.08471f
C9304 VDD.n804 GND 0.04891f
C9305 VDD.n805 GND 0.04648f
C9306 VDD.n806 GND 0.02293f
C9307 VDD.n807 GND 0.04648f
C9308 VDD.n808 GND 0.02708f
C9309 VDD.n809 GND 0.02293f
C9310 VDD.n810 GND 0.04532f
C9311 VDD.n811 GND 0.02293f
C9312 VDD.n812 GND 0.02708f
C9313 VDD.n813 GND 0.04532f
C9314 VDD.n814 GND 0.02293f
C9315 VDD.n815 GND 0.04891f
C9316 VDD.n816 GND 0.05737f
C9317 VDD.n817 GND 0.02055f
C9318 VDD.n818 GND 0.44561f
C9319 VDD.n819 GND 0.14059f
C9320 VDD.n820 GND 0.04891f
C9321 VDD.n821 GND 0.04648f
C9322 VDD.n822 GND 0.02293f
C9323 VDD.n823 GND 0.04648f
C9324 VDD.n824 GND 0.02708f
C9325 VDD.n825 GND 0.02293f
C9326 VDD.n826 GND 0.04532f
C9327 VDD.n827 GND 0.02293f
C9328 VDD.n828 GND 0.02708f
C9329 VDD.n829 GND 0.04532f
C9330 VDD.n830 GND 0.02293f
C9331 VDD.n831 GND 0.04891f
C9332 VDD.n832 GND 0.05737f
C9333 VDD.n833 GND 0.02055f
C9334 VDD.n834 GND 0.02497f
C9335 VDD.n835 GND 0.04648f
C9336 VDD.n836 GND 0.04648f
C9337 VDD.n837 GND 0.02708f
C9338 VDD.n838 GND 0.02497f
C9339 VDD.n839 GND 0.08328f
C9340 VDD.n840 GND 0.01566f
C9341 VDD.n841 GND 0.18236f
C9342 VDD.n842 GND 0.03549f
C9343 VDD.n843 GND 0.04891f
C9344 VDD.n844 GND 0.04648f
C9345 VDD.n845 GND 0.02293f
C9346 VDD.n846 GND 0.04648f
C9347 VDD.n847 GND 0.02708f
C9348 VDD.n848 GND 0.02293f
C9349 VDD.n849 GND 0.04532f
C9350 VDD.n850 GND 0.02293f
C9351 VDD.n851 GND 0.02708f
C9352 VDD.n852 GND 0.04532f
C9353 VDD.n853 GND 0.02293f
C9354 VDD.n854 GND 0.04891f
C9355 VDD.n855 GND 0.05737f
C9356 VDD.n856 GND 0.02055f
C9357 VDD.n857 GND 0.44561f
C9358 VDD.n858 GND 0.14059f
C9359 VDD.n859 GND 0.04891f
C9360 VDD.n860 GND 0.04648f
C9361 VDD.n861 GND 0.02293f
C9362 VDD.n862 GND 0.04648f
C9363 VDD.n863 GND 0.02708f
C9364 VDD.n864 GND 0.02293f
C9365 VDD.n865 GND 0.04532f
C9366 VDD.n866 GND 0.02293f
C9367 VDD.n867 GND 0.02708f
C9368 VDD.n868 GND 0.04532f
C9369 VDD.n869 GND 0.02293f
C9370 VDD.n870 GND 0.04891f
C9371 VDD.n871 GND 0.05737f
C9372 VDD.n872 GND 0.02813f
C9373 VDD.n873 GND 0.02324f
C9374 VDD.n874 GND 0.05737f
C9375 VDD.n875 GND 0.04891f
C9376 VDD.n876 GND 0.02293f
C9377 VDD.n877 GND 0.02708f
C9378 VDD.n878 GND 0.04648f
C9379 VDD.n879 GND 0.02293f
C9380 VDD.n880 GND 0.02293f
C9381 VDD.n881 GND 0.02708f
C9382 VDD.n882 GND 0.04648f
C9383 VDD.n883 GND 0.02708f
C9384 VDD.n884 GND 0.04648f
C9385 VDD.n885 GND 3.19829f
C9386 VDD.n886 GND 0.04648f
C9387 VDD.n887 GND 0.04532f
C9388 VDD.n888 GND 0.02293f
C9389 VDD.n889 GND 0.04891f
C9390 VDD.n890 GND 0.05737f
C9391 VDD.n891 GND 0.02813f
C9392 VDD.n892 GND 0.14059f
C9393 VDD.n893 GND 0.44561f
C9394 VDD.n894 GND 0.02055f
C9395 VDD.n895 GND 0.05737f
C9396 VDD.n896 GND 0.04891f
C9397 VDD.n897 GND 0.02293f
C9398 VDD.n898 GND 0.02708f
C9399 VDD.n899 GND 0.02293f
C9400 VDD.n900 GND 0.04532f
C9401 VDD.t126 GND 4.12913f
C9402 VDD.n901 GND 0.04532f
C9403 VDD.n902 GND 0.04648f
C9404 VDD.n903 GND 0.05737f
C9405 VDD.n904 GND 0.01303f
C9406 VDD.n905 GND 0.95576f
C9407 VDD.n906 GND 0.08471f
C9408 VDD.n907 GND 0.01566f
C9409 VDD.n908 GND 0.08328f
C9410 VDD.n909 GND 0.04648f
C9411 VDD.n910 GND 3.47277f
C9412 VDD.n911 GND 0.04648f
C9413 VDD.n912 GND 0.05737f
C9414 VDD.n913 GND 0.0171f
C9415 VDD.n914 GND 0.064f
C9416 VDD.n917 GND 0.06555f
C9417 VDD.n918 GND 0.03083f
C9418 VDD.t207 GND 0.08047f
C9419 VDD.n919 GND 0.03534f
C9420 VDD.t949 GND 0.15471f
C9421 VDD.n920 GND 0.03238f
C9422 VDD.n921 GND 0.02607f
C9423 VDD.n922 GND 0.09595f
C9424 VDD.t125 GND 0.08047f
C9425 VDD.n923 GND 0.03534f
C9426 VDD.t933 GND 0.15471f
C9427 VDD.n924 GND 0.03238f
C9428 VDD.n925 GND 0.02607f
C9429 VDD.n927 GND 0.24365f
C9430 VDD.n928 GND 0.03496f
C9431 VDD.n929 GND 2.34336f
C9432 VDD.n930 GND 2.04012f
C9433 VDD.t943 GND 0.15539f
C9434 VDD.n931 GND 0.06697f
C9435 VDD.t201 GND 0.07226f
C9436 VDD.n932 GND 0.05627f
C9437 VDD.n933 GND 0.05442f
C9438 VDD.n934 GND 0.04255f
C9439 VDD.n935 GND 0.05152f
C9440 VDD.t80 GND 0.02114f
C9441 VDD.t857 GND 0.02114f
C9442 VDD.n936 GND 0.14059f
C9443 VDD.n937 GND 0.04891f
C9444 VDD.n938 GND 0.04648f
C9445 VDD.n939 GND 0.04891f
C9446 VDD.n940 GND 0.04532f
C9447 VDD.n941 GND 0.04532f
C9448 VDD.t12 GND 4.12913f
C9449 VDD.n942 GND 0.04648f
C9450 VDD.n943 GND 0.04648f
C9451 VDD.n944 GND 0.04648f
C9452 VDD.n945 GND 0.04648f
C9453 VDD.n946 GND 0.04648f
C9454 VDD.n947 GND 0.04648f
C9455 VDD.n948 GND 3.47277f
C9456 VDD.n949 GND 0.04648f
C9457 VDD.n950 GND 0.04648f
C9458 VDD.n951 GND 0.04648f
C9459 VDD.n952 GND 0.04648f
C9460 VDD.n953 GND 0.04532f
C9461 VDD.n954 GND 0.04532f
C9462 VDD.n955 GND 0.02497f
C9463 VDD.n956 GND 0.02497f
C9464 VDD.t859 GND 0.02104f
C9465 VDD.n957 GND 0.22365f
C9466 VDD.t202 GND 0.02104f
C9467 VDD.t684 GND 0.02104f
C9468 VDD.n958 GND 0.04891f
C9469 VDD.n959 GND 0.04891f
C9470 VDD.n960 GND 0.04532f
C9471 VDD.n961 GND 0.04648f
C9472 VDD.n962 GND 0.02293f
C9473 VDD.n963 GND 0.02708f
C9474 VDD.n964 GND 0.02293f
C9475 VDD.n965 GND 0.04532f
C9476 VDD.n966 GND 0.04532f
C9477 VDD.n967 GND 0.04532f
C9478 VDD.n968 GND 0.04532f
C9479 VDD.n969 GND 0.04532f
C9480 VDD.n970 GND 0.04532f
C9481 VDD.n971 GND 0.04532f
C9482 VDD.n972 GND 0.04532f
C9483 VDD.n973 GND 0.04532f
C9484 VDD.n974 GND 0.04532f
C9485 VDD.n975 GND 0.04532f
C9486 VDD.n976 GND 0.04532f
C9487 VDD.n977 GND 0.04532f
C9488 VDD.n978 GND 0.04532f
C9489 VDD.n979 GND 0.04532f
C9490 VDD.n980 GND 0.04532f
C9491 VDD.n981 GND 0.04532f
C9492 VDD.n982 GND 0.04532f
C9493 VDD.n983 GND 0.04532f
C9494 VDD.n984 GND 0.04532f
C9495 VDD.n985 GND 0.02293f
C9496 VDD.n986 GND 0.02293f
C9497 VDD.n987 GND 0.02708f
C9498 VDD.n988 GND 0.04648f
C9499 VDD.n989 GND 3.19829f
C9500 VDD.n990 GND 0.04532f
C9501 VDD.n991 GND 0.04648f
C9502 VDD.n992 GND 0.04648f
C9503 VDD.n993 GND 0.04891f
C9504 VDD.n994 GND 0.02293f
C9505 VDD.t749 GND 0.02114f
C9506 VDD.t50 GND 0.02114f
C9507 VDD.t52 GND 0.02114f
C9508 VDD.t67 GND 0.02114f
C9509 VDD.n995 GND 0.02324f
C9510 VDD.n996 GND 0.04891f
C9511 VDD.n997 GND 0.04648f
C9512 VDD.n998 GND 0.02293f
C9513 VDD.n999 GND 0.04648f
C9514 VDD.n1000 GND 0.02708f
C9515 VDD.n1001 GND 0.02293f
C9516 VDD.n1002 GND 0.02708f
C9517 VDD.n1003 GND 0.02293f
C9518 VDD.n1004 GND 0.04532f
C9519 VDD.n1005 GND 0.04532f
C9520 VDD.n1006 GND 0.04532f
C9521 VDD.n1007 GND 0.02293f
C9522 VDD.n1008 GND 0.02293f
C9523 VDD.n1009 GND 0.02708f
C9524 VDD.n1010 GND 0.04648f
C9525 VDD.n1011 GND 0.04648f
C9526 VDD.n1012 GND 0.04648f
C9527 VDD.n1013 GND 0.04648f
C9528 VDD.n1014 GND 0.04532f
C9529 VDD.n1015 GND 0.04532f
C9530 VDD.n1016 GND 0.02293f
C9531 VDD.n1017 GND 0.02293f
C9532 VDD.n1018 GND 0.04648f
C9533 VDD.n1019 GND 0.02708f
C9534 VDD.n1020 GND 0.02293f
C9535 VDD.n1021 GND 0.04891f
C9536 VDD.n1022 GND 0.04648f
C9537 VDD.n1023 GND 0.05737f
C9538 VDD.n1024 GND 0.04891f
C9539 VDD.n1025 GND 0.02293f
C9540 VDD.n1026 GND 0.02708f
C9541 VDD.n1027 GND 0.04648f
C9542 VDD.n1028 GND 0.04532f
C9543 VDD.n1029 GND 0.04532f
C9544 VDD.n1030 GND 0.02293f
C9545 VDD.n1031 GND 0.02708f
C9546 VDD.n1032 GND 0.04648f
C9547 VDD.n1033 GND 0.04648f
C9548 VDD.n1034 GND 0.04648f
C9549 VDD.n1035 GND 0.04532f
C9550 VDD.n1036 GND 0.04532f
C9551 VDD.n1037 GND 0.02293f
C9552 VDD.n1038 GND 0.02293f
C9553 VDD.n1039 GND 0.04648f
C9554 VDD.n1040 GND 0.02708f
C9555 VDD.n1041 GND 0.02293f
C9556 VDD.n1042 GND 0.04891f
C9557 VDD.n1043 GND 0.04648f
C9558 VDD.t186 GND 0.02104f
C9559 VDD.t698 GND 0.02104f
C9560 VDD.t234 GND 0.02114f
C9561 VDD.t832 GND 0.02114f
C9562 VDD.n1044 GND 0.44561f
C9563 VDD.n1045 GND 0.04891f
C9564 VDD.n1046 GND 0.04648f
C9565 VDD.n1047 GND 0.02293f
C9566 VDD.n1048 GND 0.04648f
C9567 VDD.n1049 GND 0.02708f
C9568 VDD.n1050 GND 0.02293f
C9569 VDD.n1051 GND 0.04532f
C9570 VDD.n1052 GND 0.02293f
C9571 VDD.n1053 GND 0.02708f
C9572 VDD.n1054 GND 0.04532f
C9573 VDD.n1055 GND 0.02293f
C9574 VDD.n1056 GND 0.04891f
C9575 VDD.n1057 GND 0.05737f
C9576 VDD.n1058 GND 0.02055f
C9577 VDD.n1059 GND 0.08471f
C9578 VDD.n1060 GND 0.95576f
C9579 VDD.t791 GND 0.02114f
C9580 VDD.t603 GND 0.02114f
C9581 VDD.t268 GND 0.02114f
C9582 VDD.t354 GND 0.02114f
C9583 VDD.t824 GND 0.02104f
C9584 VDD.t355 GND 0.02114f
C9585 VDD.t381 GND 0.02114f
C9586 VDD.t556 GND 0.02114f
C9587 VDD.t13 GND 0.02114f
C9588 VDD.t178 GND 0.02104f
C9589 VDD.t689 GND 0.02104f
C9590 VDD.n1061 GND 0.95576f
C9591 VDD.n1062 GND 0.08471f
C9592 VDD.n1063 GND 0.04891f
C9593 VDD.n1064 GND 0.04648f
C9594 VDD.n1065 GND 0.02293f
C9595 VDD.n1066 GND 0.04648f
C9596 VDD.n1067 GND 0.02708f
C9597 VDD.n1068 GND 0.02293f
C9598 VDD.n1069 GND 0.04532f
C9599 VDD.n1070 GND 0.02293f
C9600 VDD.n1071 GND 0.02708f
C9601 VDD.n1072 GND 0.04532f
C9602 VDD.n1073 GND 0.02293f
C9603 VDD.n1074 GND 0.04891f
C9604 VDD.n1075 GND 0.05737f
C9605 VDD.n1076 GND 0.02055f
C9606 VDD.n1077 GND 0.44561f
C9607 VDD.n1078 GND 0.14059f
C9608 VDD.n1079 GND 0.04891f
C9609 VDD.n1080 GND 0.04648f
C9610 VDD.n1081 GND 0.02293f
C9611 VDD.n1082 GND 0.04648f
C9612 VDD.n1083 GND 0.02708f
C9613 VDD.n1084 GND 0.02293f
C9614 VDD.n1085 GND 0.04532f
C9615 VDD.n1086 GND 0.02293f
C9616 VDD.n1087 GND 0.02708f
C9617 VDD.n1088 GND 0.04532f
C9618 VDD.n1089 GND 0.02293f
C9619 VDD.n1090 GND 0.04891f
C9620 VDD.n1091 GND 0.05737f
C9621 VDD.n1092 GND 0.02055f
C9622 VDD.n1093 GND 0.02497f
C9623 VDD.n1094 GND 0.04648f
C9624 VDD.n1095 GND 0.04648f
C9625 VDD.n1096 GND 0.02708f
C9626 VDD.n1097 GND 0.02497f
C9627 VDD.n1098 GND 0.08328f
C9628 VDD.n1099 GND 0.01566f
C9629 VDD.n1100 GND 0.18236f
C9630 VDD.n1101 GND 0.03549f
C9631 VDD.n1102 GND 0.04891f
C9632 VDD.n1103 GND 0.04648f
C9633 VDD.n1104 GND 0.02293f
C9634 VDD.n1105 GND 0.04648f
C9635 VDD.n1106 GND 0.02708f
C9636 VDD.n1107 GND 0.02293f
C9637 VDD.n1108 GND 0.04532f
C9638 VDD.n1109 GND 0.02293f
C9639 VDD.n1110 GND 0.02708f
C9640 VDD.n1111 GND 0.04532f
C9641 VDD.n1112 GND 0.02293f
C9642 VDD.n1113 GND 0.04891f
C9643 VDD.n1114 GND 0.05737f
C9644 VDD.n1115 GND 0.02055f
C9645 VDD.n1116 GND 0.44561f
C9646 VDD.n1117 GND 0.14059f
C9647 VDD.n1118 GND 0.04891f
C9648 VDD.n1119 GND 0.04648f
C9649 VDD.n1120 GND 0.02293f
C9650 VDD.n1121 GND 0.04648f
C9651 VDD.n1122 GND 0.02708f
C9652 VDD.n1123 GND 0.02293f
C9653 VDD.n1124 GND 0.04532f
C9654 VDD.n1125 GND 0.02293f
C9655 VDD.n1126 GND 0.02708f
C9656 VDD.n1127 GND 0.04532f
C9657 VDD.n1128 GND 0.02293f
C9658 VDD.n1129 GND 0.04891f
C9659 VDD.n1130 GND 0.05737f
C9660 VDD.n1131 GND 0.02813f
C9661 VDD.n1132 GND 0.02324f
C9662 VDD.n1133 GND 0.05737f
C9663 VDD.n1134 GND 0.04891f
C9664 VDD.n1135 GND 0.02293f
C9665 VDD.n1136 GND 0.02708f
C9666 VDD.n1137 GND 0.04648f
C9667 VDD.n1138 GND 0.02293f
C9668 VDD.n1139 GND 0.02293f
C9669 VDD.n1140 GND 0.02708f
C9670 VDD.n1141 GND 0.04648f
C9671 VDD.n1142 GND 0.02708f
C9672 VDD.n1143 GND 0.04648f
C9673 VDD.n1144 GND 3.19829f
C9674 VDD.n1145 GND 0.04648f
C9675 VDD.n1146 GND 0.04532f
C9676 VDD.n1147 GND 0.02293f
C9677 VDD.n1148 GND 0.04891f
C9678 VDD.n1149 GND 0.05737f
C9679 VDD.n1150 GND 0.02813f
C9680 VDD.n1151 GND 0.14059f
C9681 VDD.n1152 GND 0.44561f
C9682 VDD.n1153 GND 0.02055f
C9683 VDD.n1154 GND 0.05737f
C9684 VDD.n1155 GND 0.04891f
C9685 VDD.n1156 GND 0.02293f
C9686 VDD.n1157 GND 0.02708f
C9687 VDD.n1158 GND 0.02293f
C9688 VDD.n1159 GND 0.04532f
C9689 VDD.t51 GND 4.12913f
C9690 VDD.n1160 GND 0.04532f
C9691 VDD.n1161 GND 0.04648f
C9692 VDD.n1162 GND 0.05737f
C9693 VDD.n1163 GND 0.01303f
C9694 VDD.n1164 GND 0.95576f
C9695 VDD.n1165 GND 0.08471f
C9696 VDD.n1166 GND 0.01566f
C9697 VDD.n1167 GND 0.08328f
C9698 VDD.n1168 GND 0.04648f
C9699 VDD.n1169 GND 3.47277f
C9700 VDD.n1170 GND 0.04648f
C9701 VDD.n1171 GND 0.05737f
C9702 VDD.n1172 GND 0.0171f
C9703 VDD.n1173 GND 0.064f
C9704 VDD.n1176 GND 0.06555f
C9705 VDD.n1177 GND 0.03083f
C9706 VDD.t177 GND 0.08047f
C9707 VDD.n1178 GND 0.03534f
C9708 VDD.t930 GND 0.15471f
C9709 VDD.n1179 GND 0.03238f
C9710 VDD.n1180 GND 0.02607f
C9711 VDD.n1181 GND 0.09595f
C9712 VDD.t185 GND 0.08047f
C9713 VDD.n1182 GND 0.03534f
C9714 VDD.t970 GND 0.15471f
C9715 VDD.n1183 GND 0.03238f
C9716 VDD.n1184 GND 0.02607f
C9717 VDD.n1186 GND 0.24365f
C9718 VDD.n1187 GND 0.03496f
C9719 VDD.n1188 GND 2.18317f
C9720 VDD.n1189 GND 1.8945f
C9721 VDD.t924 GND 0.15539f
C9722 VDD.n1190 GND 0.06697f
C9723 VDD.t110 GND 0.07226f
C9724 VDD.n1191 GND 0.05627f
C9725 VDD.n1192 GND 0.05442f
C9726 VDD.n1193 GND 0.04255f
C9727 VDD.n1194 GND 0.05152f
C9728 VDD.t290 GND 0.02114f
C9729 VDD.t263 GND 0.02114f
C9730 VDD.n1195 GND 0.14059f
C9731 VDD.n1196 GND 0.04891f
C9732 VDD.n1197 GND 0.04648f
C9733 VDD.n1198 GND 0.04891f
C9734 VDD.n1199 GND 0.04532f
C9735 VDD.n1200 GND 0.04532f
C9736 VDD.t111 GND 4.12913f
C9737 VDD.n1201 GND 0.04648f
C9738 VDD.n1202 GND 0.04648f
C9739 VDD.n1203 GND 0.04648f
C9740 VDD.n1204 GND 0.04648f
C9741 VDD.n1205 GND 0.04648f
C9742 VDD.n1206 GND 0.04648f
C9743 VDD.n1207 GND 3.47277f
C9744 VDD.n1208 GND 0.04648f
C9745 VDD.n1209 GND 0.04648f
C9746 VDD.n1210 GND 0.04648f
C9747 VDD.n1211 GND 0.04648f
C9748 VDD.n1212 GND 0.04532f
C9749 VDD.n1213 GND 0.04532f
C9750 VDD.n1214 GND 0.02497f
C9751 VDD.n1215 GND 0.02497f
C9752 VDD.t370 GND 0.02104f
C9753 VDD.n1216 GND 0.22365f
C9754 VDD.t112 GND 0.02104f
C9755 VDD.t657 GND 0.02104f
C9756 VDD.n1217 GND 0.04891f
C9757 VDD.n1218 GND 0.04891f
C9758 VDD.n1219 GND 0.04532f
C9759 VDD.n1220 GND 0.04648f
C9760 VDD.n1221 GND 0.02293f
C9761 VDD.n1222 GND 0.02708f
C9762 VDD.n1223 GND 0.02293f
C9763 VDD.n1224 GND 0.04532f
C9764 VDD.n1225 GND 0.04532f
C9765 VDD.n1226 GND 0.04532f
C9766 VDD.n1227 GND 0.04532f
C9767 VDD.n1228 GND 0.04532f
C9768 VDD.n1229 GND 0.04532f
C9769 VDD.n1230 GND 0.04532f
C9770 VDD.n1231 GND 0.04532f
C9771 VDD.n1232 GND 0.04532f
C9772 VDD.n1233 GND 0.04532f
C9773 VDD.n1234 GND 0.04532f
C9774 VDD.n1235 GND 0.04532f
C9775 VDD.n1236 GND 0.04532f
C9776 VDD.n1237 GND 0.04532f
C9777 VDD.n1238 GND 0.04532f
C9778 VDD.n1239 GND 0.04532f
C9779 VDD.n1240 GND 0.04532f
C9780 VDD.n1241 GND 0.04532f
C9781 VDD.n1242 GND 0.04532f
C9782 VDD.n1243 GND 0.04532f
C9783 VDD.n1244 GND 0.02293f
C9784 VDD.n1245 GND 0.02293f
C9785 VDD.n1246 GND 0.02708f
C9786 VDD.n1247 GND 0.04648f
C9787 VDD.n1248 GND 3.19829f
C9788 VDD.n1249 GND 0.04532f
C9789 VDD.n1250 GND 0.04648f
C9790 VDD.n1251 GND 0.04648f
C9791 VDD.n1252 GND 0.04891f
C9792 VDD.n1253 GND 0.02293f
C9793 VDD.t741 GND 0.02114f
C9794 VDD.t266 GND 0.02114f
C9795 VDD.t702 GND 0.02114f
C9796 VDD.t310 GND 0.02114f
C9797 VDD.n1254 GND 0.02324f
C9798 VDD.n1255 GND 0.04891f
C9799 VDD.n1256 GND 0.04648f
C9800 VDD.n1257 GND 0.02293f
C9801 VDD.n1258 GND 0.04648f
C9802 VDD.n1259 GND 0.02708f
C9803 VDD.n1260 GND 0.02293f
C9804 VDD.n1261 GND 0.02708f
C9805 VDD.n1262 GND 0.02293f
C9806 VDD.n1263 GND 0.04532f
C9807 VDD.n1264 GND 0.04532f
C9808 VDD.n1265 GND 0.04532f
C9809 VDD.n1266 GND 0.02293f
C9810 VDD.n1267 GND 0.02293f
C9811 VDD.n1268 GND 0.02708f
C9812 VDD.n1269 GND 0.04648f
C9813 VDD.n1270 GND 0.04648f
C9814 VDD.n1271 GND 0.04648f
C9815 VDD.n1272 GND 0.04648f
C9816 VDD.n1273 GND 0.04532f
C9817 VDD.n1274 GND 0.04532f
C9818 VDD.n1275 GND 0.02293f
C9819 VDD.n1276 GND 0.02293f
C9820 VDD.n1277 GND 0.04648f
C9821 VDD.n1278 GND 0.02708f
C9822 VDD.n1279 GND 0.02293f
C9823 VDD.n1280 GND 0.04891f
C9824 VDD.n1281 GND 0.04648f
C9825 VDD.n1282 GND 0.05737f
C9826 VDD.n1283 GND 0.04891f
C9827 VDD.n1284 GND 0.02293f
C9828 VDD.n1285 GND 0.02708f
C9829 VDD.n1286 GND 0.04648f
C9830 VDD.n1287 GND 0.04532f
C9831 VDD.n1288 GND 0.04532f
C9832 VDD.n1289 GND 0.02293f
C9833 VDD.n1290 GND 0.02708f
C9834 VDD.n1291 GND 0.04648f
C9835 VDD.n1292 GND 0.04648f
C9836 VDD.n1293 GND 0.04648f
C9837 VDD.n1294 GND 0.04532f
C9838 VDD.n1295 GND 0.04532f
C9839 VDD.n1296 GND 0.02293f
C9840 VDD.n1297 GND 0.02293f
C9841 VDD.n1298 GND 0.04648f
C9842 VDD.n1299 GND 0.02708f
C9843 VDD.n1300 GND 0.02293f
C9844 VDD.n1301 GND 0.04891f
C9845 VDD.n1302 GND 0.04648f
C9846 VDD.t133 GND 0.02104f
C9847 VDD.t659 GND 0.02104f
C9848 VDD.t229 GND 0.02114f
C9849 VDD.t810 GND 0.02114f
C9850 VDD.n1303 GND 0.44561f
C9851 VDD.n1304 GND 0.04891f
C9852 VDD.n1305 GND 0.04648f
C9853 VDD.n1306 GND 0.02293f
C9854 VDD.n1307 GND 0.04648f
C9855 VDD.n1308 GND 0.02708f
C9856 VDD.n1309 GND 0.02293f
C9857 VDD.n1310 GND 0.04532f
C9858 VDD.n1311 GND 0.02293f
C9859 VDD.n1312 GND 0.02708f
C9860 VDD.n1313 GND 0.04532f
C9861 VDD.n1314 GND 0.02293f
C9862 VDD.n1315 GND 0.04891f
C9863 VDD.n1316 GND 0.05737f
C9864 VDD.n1317 GND 0.02055f
C9865 VDD.n1318 GND 0.08471f
C9866 VDD.n1319 GND 0.95576f
C9867 VDD.t918 GND 0.02114f
C9868 VDD.t798 GND 0.02114f
C9869 VDD.t593 GND 0.02114f
C9870 VDD.t841 GND 0.02114f
C9871 VDD.t238 GND 0.02104f
C9872 VDD.t54 GND 0.02114f
C9873 VDD.t320 GND 0.02114f
C9874 VDD.t514 GND 0.02114f
C9875 VDD.t516 GND 0.02114f
C9876 VDD.t99 GND 0.02104f
C9877 VDD.t700 GND 0.02104f
C9878 VDD.n1320 GND 0.95576f
C9879 VDD.n1321 GND 0.08471f
C9880 VDD.n1322 GND 0.04891f
C9881 VDD.n1323 GND 0.04648f
C9882 VDD.n1324 GND 0.02293f
C9883 VDD.n1325 GND 0.04648f
C9884 VDD.n1326 GND 0.02708f
C9885 VDD.n1327 GND 0.02293f
C9886 VDD.n1328 GND 0.04532f
C9887 VDD.n1329 GND 0.02293f
C9888 VDD.n1330 GND 0.02708f
C9889 VDD.n1331 GND 0.04532f
C9890 VDD.n1332 GND 0.02293f
C9891 VDD.n1333 GND 0.04891f
C9892 VDD.n1334 GND 0.05737f
C9893 VDD.n1335 GND 0.02055f
C9894 VDD.n1336 GND 0.44561f
C9895 VDD.n1337 GND 0.14059f
C9896 VDD.n1338 GND 0.04891f
C9897 VDD.n1339 GND 0.04648f
C9898 VDD.n1340 GND 0.02293f
C9899 VDD.n1341 GND 0.04648f
C9900 VDD.n1342 GND 0.02708f
C9901 VDD.n1343 GND 0.02293f
C9902 VDD.n1344 GND 0.04532f
C9903 VDD.n1345 GND 0.02293f
C9904 VDD.n1346 GND 0.02708f
C9905 VDD.n1347 GND 0.04532f
C9906 VDD.n1348 GND 0.02293f
C9907 VDD.n1349 GND 0.04891f
C9908 VDD.n1350 GND 0.05737f
C9909 VDD.n1351 GND 0.02055f
C9910 VDD.n1352 GND 0.02497f
C9911 VDD.n1353 GND 0.04648f
C9912 VDD.n1354 GND 0.04648f
C9913 VDD.n1355 GND 0.02708f
C9914 VDD.n1356 GND 0.02497f
C9915 VDD.n1357 GND 0.08328f
C9916 VDD.n1358 GND 0.01566f
C9917 VDD.n1359 GND 0.18236f
C9918 VDD.n1360 GND 0.03549f
C9919 VDD.n1361 GND 0.04891f
C9920 VDD.n1362 GND 0.04648f
C9921 VDD.n1363 GND 0.02293f
C9922 VDD.n1364 GND 0.04648f
C9923 VDD.n1365 GND 0.02708f
C9924 VDD.n1366 GND 0.02293f
C9925 VDD.n1367 GND 0.04532f
C9926 VDD.n1368 GND 0.02293f
C9927 VDD.n1369 GND 0.02708f
C9928 VDD.n1370 GND 0.04532f
C9929 VDD.n1371 GND 0.02293f
C9930 VDD.n1372 GND 0.04891f
C9931 VDD.n1373 GND 0.05737f
C9932 VDD.n1374 GND 0.02055f
C9933 VDD.n1375 GND 0.44561f
C9934 VDD.n1376 GND 0.14059f
C9935 VDD.n1377 GND 0.04891f
C9936 VDD.n1378 GND 0.04648f
C9937 VDD.n1379 GND 0.02293f
C9938 VDD.n1380 GND 0.04648f
C9939 VDD.n1381 GND 0.02708f
C9940 VDD.n1382 GND 0.02293f
C9941 VDD.n1383 GND 0.04532f
C9942 VDD.n1384 GND 0.02293f
C9943 VDD.n1385 GND 0.02708f
C9944 VDD.n1386 GND 0.04532f
C9945 VDD.n1387 GND 0.02293f
C9946 VDD.n1388 GND 0.04891f
C9947 VDD.n1389 GND 0.05737f
C9948 VDD.n1390 GND 0.02813f
C9949 VDD.n1391 GND 0.02324f
C9950 VDD.n1392 GND 0.05737f
C9951 VDD.n1393 GND 0.04891f
C9952 VDD.n1394 GND 0.02293f
C9953 VDD.n1395 GND 0.02708f
C9954 VDD.n1396 GND 0.04648f
C9955 VDD.n1397 GND 0.02293f
C9956 VDD.n1398 GND 0.02293f
C9957 VDD.n1399 GND 0.02708f
C9958 VDD.n1400 GND 0.04648f
C9959 VDD.n1401 GND 0.02708f
C9960 VDD.n1402 GND 0.04648f
C9961 VDD.n1403 GND 3.19829f
C9962 VDD.n1404 GND 0.04648f
C9963 VDD.n1405 GND 0.04532f
C9964 VDD.n1406 GND 0.02293f
C9965 VDD.n1407 GND 0.04891f
C9966 VDD.n1408 GND 0.05737f
C9967 VDD.n1409 GND 0.02813f
C9968 VDD.n1410 GND 0.14059f
C9969 VDD.n1411 GND 0.44561f
C9970 VDD.n1412 GND 0.02055f
C9971 VDD.n1413 GND 0.05737f
C9972 VDD.n1414 GND 0.04891f
C9973 VDD.n1415 GND 0.02293f
C9974 VDD.n1416 GND 0.02708f
C9975 VDD.n1417 GND 0.02293f
C9976 VDD.n1418 GND 0.04532f
C9977 VDD.t53 GND 4.12913f
C9978 VDD.n1419 GND 0.04532f
C9979 VDD.n1420 GND 0.04648f
C9980 VDD.n1421 GND 0.05737f
C9981 VDD.n1422 GND 0.01303f
C9982 VDD.n1423 GND 0.95576f
C9983 VDD.n1424 GND 0.08471f
C9984 VDD.n1425 GND 0.01566f
C9985 VDD.n1426 GND 0.08328f
C9986 VDD.n1427 GND 0.04648f
C9987 VDD.n1428 GND 3.47277f
C9988 VDD.n1429 GND 0.04648f
C9989 VDD.n1430 GND 0.05737f
C9990 VDD.n1431 GND 0.0171f
C9991 VDD.n1432 GND 0.064f
C9992 VDD.n1435 GND 0.06555f
C9993 VDD.n1436 GND 0.03083f
C9994 VDD.t98 GND 0.08047f
C9995 VDD.n1437 GND 0.03534f
C9996 VDD.t944 GND 0.15471f
C9997 VDD.n1438 GND 0.03238f
C9998 VDD.n1439 GND 0.02607f
C9999 VDD.n1440 GND 0.09595f
C10000 VDD.t132 GND 0.08047f
C10001 VDD.n1441 GND 0.03534f
C10002 VDD.t931 GND 0.15471f
C10003 VDD.n1442 GND 0.03238f
C10004 VDD.n1443 GND 0.02607f
C10005 VDD.n1445 GND 0.24365f
C10006 VDD.n1446 GND 0.03496f
C10007 VDD.n1447 GND 2.02298f
C10008 VDD.n1448 GND 1.74887f
C10009 VDD.t966 GND 0.15539f
C10010 VDD.n1449 GND 0.06697f
C10011 VDD.t146 GND 0.07226f
C10012 VDD.n1450 GND 0.05627f
C10013 VDD.n1451 GND 0.05442f
C10014 VDD.n1452 GND 0.04255f
C10015 VDD.n1453 GND 0.05152f
C10016 VDD.t557 GND 0.02114f
C10017 VDD.t793 GND 0.02114f
C10018 VDD.n1454 GND 0.14059f
C10019 VDD.n1455 GND 0.04891f
C10020 VDD.n1456 GND 0.04648f
C10021 VDD.n1457 GND 0.04891f
C10022 VDD.n1458 GND 0.04532f
C10023 VDD.n1459 GND 0.04532f
C10024 VDD.t147 GND 4.12913f
C10025 VDD.n1460 GND 0.04648f
C10026 VDD.n1461 GND 0.04648f
C10027 VDD.n1462 GND 0.04648f
C10028 VDD.n1463 GND 0.04648f
C10029 VDD.n1464 GND 0.04648f
C10030 VDD.n1465 GND 0.04648f
C10031 VDD.n1466 GND 3.47277f
C10032 VDD.n1467 GND 0.04648f
C10033 VDD.n1468 GND 0.04648f
C10034 VDD.n1469 GND 0.04648f
C10035 VDD.n1470 GND 0.04648f
C10036 VDD.n1471 GND 0.04532f
C10037 VDD.n1472 GND 0.04532f
C10038 VDD.n1473 GND 0.02497f
C10039 VDD.n1474 GND 0.02497f
C10040 VDD.t740 GND 0.02104f
C10041 VDD.n1475 GND 0.22365f
C10042 VDD.t148 GND 0.02104f
C10043 VDD.t663 GND 0.02104f
C10044 VDD.n1476 GND 0.04891f
C10045 VDD.n1477 GND 0.04891f
C10046 VDD.n1478 GND 0.04532f
C10047 VDD.n1479 GND 0.04648f
C10048 VDD.n1480 GND 0.02293f
C10049 VDD.n1481 GND 0.02708f
C10050 VDD.n1482 GND 0.02293f
C10051 VDD.n1483 GND 0.04532f
C10052 VDD.n1484 GND 0.04532f
C10053 VDD.n1485 GND 0.04532f
C10054 VDD.n1486 GND 0.04532f
C10055 VDD.n1487 GND 0.04532f
C10056 VDD.n1488 GND 0.04532f
C10057 VDD.n1489 GND 0.04532f
C10058 VDD.n1490 GND 0.04532f
C10059 VDD.n1491 GND 0.04532f
C10060 VDD.n1492 GND 0.04532f
C10061 VDD.n1493 GND 0.04532f
C10062 VDD.n1494 GND 0.04532f
C10063 VDD.n1495 GND 0.04532f
C10064 VDD.n1496 GND 0.04532f
C10065 VDD.n1497 GND 0.04532f
C10066 VDD.n1498 GND 0.04532f
C10067 VDD.n1499 GND 0.04532f
C10068 VDD.n1500 GND 0.04532f
C10069 VDD.n1501 GND 0.04532f
C10070 VDD.n1502 GND 0.04532f
C10071 VDD.n1503 GND 0.02293f
C10072 VDD.n1504 GND 0.02293f
C10073 VDD.n1505 GND 0.02708f
C10074 VDD.n1506 GND 0.04648f
C10075 VDD.n1507 GND 3.19829f
C10076 VDD.n1508 GND 0.04532f
C10077 VDD.n1509 GND 0.04648f
C10078 VDD.n1510 GND 0.04648f
C10079 VDD.n1511 GND 0.04891f
C10080 VDD.n1512 GND 0.02293f
C10081 VDD.t85 GND 0.02114f
C10082 VDD.t835 GND 0.02114f
C10083 VDD.t47 GND 0.02114f
C10084 VDD.t398 GND 0.02114f
C10085 VDD.n1513 GND 0.02324f
C10086 VDD.n1514 GND 0.04891f
C10087 VDD.n1515 GND 0.04648f
C10088 VDD.n1516 GND 0.02293f
C10089 VDD.n1517 GND 0.04648f
C10090 VDD.n1518 GND 0.02708f
C10091 VDD.n1519 GND 0.02293f
C10092 VDD.n1520 GND 0.02708f
C10093 VDD.n1521 GND 0.02293f
C10094 VDD.n1522 GND 0.04532f
C10095 VDD.n1523 GND 0.04532f
C10096 VDD.n1524 GND 0.04532f
C10097 VDD.n1525 GND 0.02293f
C10098 VDD.n1526 GND 0.02293f
C10099 VDD.n1527 GND 0.02708f
C10100 VDD.n1528 GND 0.04648f
C10101 VDD.n1529 GND 0.04648f
C10102 VDD.n1530 GND 0.04648f
C10103 VDD.n1531 GND 0.04648f
C10104 VDD.n1532 GND 0.04532f
C10105 VDD.n1533 GND 0.04532f
C10106 VDD.n1534 GND 0.02293f
C10107 VDD.n1535 GND 0.02293f
C10108 VDD.n1536 GND 0.04648f
C10109 VDD.n1537 GND 0.02708f
C10110 VDD.n1538 GND 0.02293f
C10111 VDD.n1539 GND 0.04891f
C10112 VDD.n1540 GND 0.04648f
C10113 VDD.n1541 GND 0.05737f
C10114 VDD.n1542 GND 0.04891f
C10115 VDD.n1543 GND 0.02293f
C10116 VDD.n1544 GND 0.02708f
C10117 VDD.n1545 GND 0.04648f
C10118 VDD.n1546 GND 0.04532f
C10119 VDD.n1547 GND 0.04532f
C10120 VDD.n1548 GND 0.02293f
C10121 VDD.n1549 GND 0.02708f
C10122 VDD.n1550 GND 0.04648f
C10123 VDD.n1551 GND 0.04648f
C10124 VDD.n1552 GND 0.04648f
C10125 VDD.n1553 GND 0.04532f
C10126 VDD.n1554 GND 0.04532f
C10127 VDD.n1555 GND 0.02293f
C10128 VDD.n1556 GND 0.02293f
C10129 VDD.n1557 GND 0.04648f
C10130 VDD.n1558 GND 0.02708f
C10131 VDD.n1559 GND 0.02293f
C10132 VDD.n1560 GND 0.04891f
C10133 VDD.n1561 GND 0.04648f
C10134 VDD.t150 GND 0.02104f
C10135 VDD.t674 GND 0.02104f
C10136 VDD.t247 GND 0.02114f
C10137 VDD.t243 GND 0.02114f
C10138 VDD.n1562 GND 0.44561f
C10139 VDD.n1563 GND 0.04891f
C10140 VDD.n1564 GND 0.04648f
C10141 VDD.n1565 GND 0.02293f
C10142 VDD.n1566 GND 0.04648f
C10143 VDD.n1567 GND 0.02708f
C10144 VDD.n1568 GND 0.02293f
C10145 VDD.n1569 GND 0.04532f
C10146 VDD.n1570 GND 0.02293f
C10147 VDD.n1571 GND 0.02708f
C10148 VDD.n1572 GND 0.04532f
C10149 VDD.n1573 GND 0.02293f
C10150 VDD.n1574 GND 0.04891f
C10151 VDD.n1575 GND 0.05737f
C10152 VDD.n1576 GND 0.02055f
C10153 VDD.n1577 GND 0.08471f
C10154 VDD.n1578 GND 0.95576f
C10155 VDD.t849 GND 0.02114f
C10156 VDD.t906 GND 0.02114f
C10157 VDD.t472 GND 0.02114f
C10158 VDD.t769 GND 0.02114f
C10159 VDD.t295 GND 0.02104f
C10160 VDD.t768 GND 0.02114f
C10161 VDD.t473 GND 0.02114f
C10162 VDD.t751 GND 0.02114f
C10163 VDD.t750 GND 0.02114f
C10164 VDD.t109 GND 0.02104f
C10165 VDD.t658 GND 0.02104f
C10166 VDD.n1579 GND 0.95576f
C10167 VDD.n1580 GND 0.08471f
C10168 VDD.n1581 GND 0.04891f
C10169 VDD.n1582 GND 0.04648f
C10170 VDD.n1583 GND 0.02293f
C10171 VDD.n1584 GND 0.04648f
C10172 VDD.n1585 GND 0.02708f
C10173 VDD.n1586 GND 0.02293f
C10174 VDD.n1587 GND 0.04532f
C10175 VDD.n1588 GND 0.02293f
C10176 VDD.n1589 GND 0.02708f
C10177 VDD.n1590 GND 0.04532f
C10178 VDD.n1591 GND 0.02293f
C10179 VDD.n1592 GND 0.04891f
C10180 VDD.n1593 GND 0.05737f
C10181 VDD.n1594 GND 0.02055f
C10182 VDD.n1595 GND 0.44561f
C10183 VDD.n1596 GND 0.14059f
C10184 VDD.n1597 GND 0.04891f
C10185 VDD.n1598 GND 0.04648f
C10186 VDD.n1599 GND 0.02293f
C10187 VDD.n1600 GND 0.04648f
C10188 VDD.n1601 GND 0.02708f
C10189 VDD.n1602 GND 0.02293f
C10190 VDD.n1603 GND 0.04532f
C10191 VDD.n1604 GND 0.02293f
C10192 VDD.n1605 GND 0.02708f
C10193 VDD.n1606 GND 0.04532f
C10194 VDD.n1607 GND 0.02293f
C10195 VDD.n1608 GND 0.04891f
C10196 VDD.n1609 GND 0.05737f
C10197 VDD.n1610 GND 0.02055f
C10198 VDD.n1611 GND 0.02497f
C10199 VDD.n1612 GND 0.04648f
C10200 VDD.n1613 GND 0.04648f
C10201 VDD.n1614 GND 0.02708f
C10202 VDD.n1615 GND 0.02497f
C10203 VDD.n1616 GND 0.08328f
C10204 VDD.n1617 GND 0.01566f
C10205 VDD.n1618 GND 0.18236f
C10206 VDD.n1619 GND 0.03549f
C10207 VDD.n1620 GND 0.04891f
C10208 VDD.n1621 GND 0.04648f
C10209 VDD.n1622 GND 0.02293f
C10210 VDD.n1623 GND 0.04648f
C10211 VDD.n1624 GND 0.02708f
C10212 VDD.n1625 GND 0.02293f
C10213 VDD.n1626 GND 0.04532f
C10214 VDD.n1627 GND 0.02293f
C10215 VDD.n1628 GND 0.02708f
C10216 VDD.n1629 GND 0.04532f
C10217 VDD.n1630 GND 0.02293f
C10218 VDD.n1631 GND 0.04891f
C10219 VDD.n1632 GND 0.05737f
C10220 VDD.n1633 GND 0.02055f
C10221 VDD.n1634 GND 0.44561f
C10222 VDD.n1635 GND 0.14059f
C10223 VDD.n1636 GND 0.04891f
C10224 VDD.n1637 GND 0.04648f
C10225 VDD.n1638 GND 0.02293f
C10226 VDD.n1639 GND 0.04648f
C10227 VDD.n1640 GND 0.02708f
C10228 VDD.n1641 GND 0.02293f
C10229 VDD.n1642 GND 0.04532f
C10230 VDD.n1643 GND 0.02293f
C10231 VDD.n1644 GND 0.02708f
C10232 VDD.n1645 GND 0.04532f
C10233 VDD.n1646 GND 0.02293f
C10234 VDD.n1647 GND 0.04891f
C10235 VDD.n1648 GND 0.05737f
C10236 VDD.n1649 GND 0.02813f
C10237 VDD.n1650 GND 0.02324f
C10238 VDD.n1651 GND 0.05737f
C10239 VDD.n1652 GND 0.04891f
C10240 VDD.n1653 GND 0.02293f
C10241 VDD.n1654 GND 0.02708f
C10242 VDD.n1655 GND 0.04648f
C10243 VDD.n1656 GND 0.02293f
C10244 VDD.n1657 GND 0.02293f
C10245 VDD.n1658 GND 0.02708f
C10246 VDD.n1659 GND 0.04648f
C10247 VDD.n1660 GND 0.02708f
C10248 VDD.n1661 GND 0.04648f
C10249 VDD.n1662 GND 3.19829f
C10250 VDD.n1663 GND 0.04648f
C10251 VDD.n1664 GND 0.04532f
C10252 VDD.n1665 GND 0.02293f
C10253 VDD.n1666 GND 0.04891f
C10254 VDD.n1667 GND 0.05737f
C10255 VDD.n1668 GND 0.02813f
C10256 VDD.n1669 GND 0.14059f
C10257 VDD.n1670 GND 0.44561f
C10258 VDD.n1671 GND 0.02055f
C10259 VDD.n1672 GND 0.05737f
C10260 VDD.n1673 GND 0.04891f
C10261 VDD.n1674 GND 0.02293f
C10262 VDD.n1675 GND 0.02708f
C10263 VDD.n1676 GND 0.02293f
C10264 VDD.n1677 GND 0.04532f
C10265 VDD.t46 GND 4.12913f
C10266 VDD.n1678 GND 0.04532f
C10267 VDD.n1679 GND 0.04648f
C10268 VDD.n1680 GND 0.05737f
C10269 VDD.n1681 GND 0.01303f
C10270 VDD.n1682 GND 0.95576f
C10271 VDD.n1683 GND 0.08471f
C10272 VDD.n1684 GND 0.01566f
C10273 VDD.n1685 GND 0.08328f
C10274 VDD.n1686 GND 0.04648f
C10275 VDD.n1687 GND 3.47277f
C10276 VDD.n1688 GND 0.04648f
C10277 VDD.n1689 GND 0.05737f
C10278 VDD.n1690 GND 0.0171f
C10279 VDD.n1691 GND 0.064f
C10280 VDD.n1694 GND 0.06555f
C10281 VDD.n1695 GND 0.03083f
C10282 VDD.t108 GND 0.08047f
C10283 VDD.n1696 GND 0.03534f
C10284 VDD.t940 GND 0.15471f
C10285 VDD.n1697 GND 0.03238f
C10286 VDD.n1698 GND 0.02607f
C10287 VDD.n1699 GND 0.09595f
C10288 VDD.t149 GND 0.08047f
C10289 VDD.n1700 GND 0.03534f
C10290 VDD.t925 GND 0.15471f
C10291 VDD.n1701 GND 0.03238f
C10292 VDD.n1702 GND 0.02607f
C10293 VDD.n1704 GND 0.24365f
C10294 VDD.n1705 GND 0.03496f
C10295 VDD.n1706 GND 1.86279f
C10296 VDD.n1707 GND 1.60325f
C10297 VDD.t935 GND 0.15539f
C10298 VDD.n1708 GND 0.06697f
C10299 VDD.t120 GND 0.07226f
C10300 VDD.n1709 GND 0.05627f
C10301 VDD.n1710 GND 0.05442f
C10302 VDD.n1711 GND 0.04255f
C10303 VDD.n1712 GND 0.05152f
C10304 VDD.t729 GND 0.02114f
C10305 VDD.t23 GND 0.02114f
C10306 VDD.n1713 GND 0.14059f
C10307 VDD.n1714 GND 0.04891f
C10308 VDD.n1715 GND 0.04648f
C10309 VDD.n1716 GND 0.04891f
C10310 VDD.n1717 GND 0.04532f
C10311 VDD.n1718 GND 0.04532f
C10312 VDD.t22 GND 4.12913f
C10313 VDD.n1719 GND 0.04648f
C10314 VDD.n1720 GND 0.04648f
C10315 VDD.n1721 GND 0.04648f
C10316 VDD.n1722 GND 0.04648f
C10317 VDD.n1723 GND 0.04648f
C10318 VDD.n1724 GND 0.04648f
C10319 VDD.n1725 GND 3.47277f
C10320 VDD.n1726 GND 0.04648f
C10321 VDD.n1727 GND 0.04648f
C10322 VDD.n1728 GND 0.04648f
C10323 VDD.n1729 GND 0.04648f
C10324 VDD.n1730 GND 0.04532f
C10325 VDD.n1731 GND 0.04532f
C10326 VDD.n1732 GND 0.02497f
C10327 VDD.n1733 GND 0.02497f
C10328 VDD.t86 GND 0.02104f
C10329 VDD.n1734 GND 0.22365f
C10330 VDD.t121 GND 0.02104f
C10331 VDD.t675 GND 0.02104f
C10332 VDD.n1735 GND 0.04891f
C10333 VDD.n1736 GND 0.04891f
C10334 VDD.n1737 GND 0.04532f
C10335 VDD.n1738 GND 0.04648f
C10336 VDD.n1739 GND 0.02293f
C10337 VDD.n1740 GND 0.02708f
C10338 VDD.n1741 GND 0.02293f
C10339 VDD.n1742 GND 0.04532f
C10340 VDD.n1743 GND 0.04532f
C10341 VDD.n1744 GND 0.04532f
C10342 VDD.n1745 GND 0.04532f
C10343 VDD.n1746 GND 0.04532f
C10344 VDD.n1747 GND 0.04532f
C10345 VDD.n1748 GND 0.04532f
C10346 VDD.n1749 GND 0.04532f
C10347 VDD.n1750 GND 0.04532f
C10348 VDD.n1751 GND 0.04532f
C10349 VDD.n1752 GND 0.04532f
C10350 VDD.n1753 GND 0.04532f
C10351 VDD.n1754 GND 0.04532f
C10352 VDD.n1755 GND 0.04532f
C10353 VDD.n1756 GND 0.04532f
C10354 VDD.n1757 GND 0.04532f
C10355 VDD.n1758 GND 0.04532f
C10356 VDD.n1759 GND 0.04532f
C10357 VDD.n1760 GND 0.04532f
C10358 VDD.n1761 GND 0.04532f
C10359 VDD.n1762 GND 0.02293f
C10360 VDD.n1763 GND 0.02293f
C10361 VDD.n1764 GND 0.02708f
C10362 VDD.n1765 GND 0.04648f
C10363 VDD.n1766 GND 3.19829f
C10364 VDD.n1767 GND 0.04532f
C10365 VDD.n1768 GND 0.04648f
C10366 VDD.n1769 GND 0.04648f
C10367 VDD.n1770 GND 0.04891f
C10368 VDD.n1771 GND 0.02293f
C10369 VDD.t711 GND 0.02114f
C10370 VDD.t907 GND 0.02114f
C10371 VDD.t360 GND 0.02114f
C10372 VDD.t491 GND 0.02114f
C10373 VDD.n1772 GND 0.02324f
C10374 VDD.n1773 GND 0.04891f
C10375 VDD.n1774 GND 0.04648f
C10376 VDD.n1775 GND 0.02293f
C10377 VDD.n1776 GND 0.04648f
C10378 VDD.n1777 GND 0.02708f
C10379 VDD.n1778 GND 0.02293f
C10380 VDD.n1779 GND 0.02708f
C10381 VDD.n1780 GND 0.02293f
C10382 VDD.n1781 GND 0.04532f
C10383 VDD.n1782 GND 0.04532f
C10384 VDD.n1783 GND 0.04532f
C10385 VDD.n1784 GND 0.02293f
C10386 VDD.n1785 GND 0.02293f
C10387 VDD.n1786 GND 0.02708f
C10388 VDD.n1787 GND 0.04648f
C10389 VDD.n1788 GND 0.04648f
C10390 VDD.n1789 GND 0.04648f
C10391 VDD.n1790 GND 0.04648f
C10392 VDD.n1791 GND 0.04532f
C10393 VDD.n1792 GND 0.04532f
C10394 VDD.n1793 GND 0.02293f
C10395 VDD.n1794 GND 0.02293f
C10396 VDD.n1795 GND 0.04648f
C10397 VDD.n1796 GND 0.02708f
C10398 VDD.n1797 GND 0.02293f
C10399 VDD.n1798 GND 0.04891f
C10400 VDD.n1799 GND 0.04648f
C10401 VDD.n1800 GND 0.05737f
C10402 VDD.n1801 GND 0.04891f
C10403 VDD.n1802 GND 0.02293f
C10404 VDD.n1803 GND 0.02708f
C10405 VDD.n1804 GND 0.04648f
C10406 VDD.n1805 GND 0.04532f
C10407 VDD.n1806 GND 0.04532f
C10408 VDD.n1807 GND 0.02293f
C10409 VDD.n1808 GND 0.02708f
C10410 VDD.n1809 GND 0.04648f
C10411 VDD.n1810 GND 0.04648f
C10412 VDD.n1811 GND 0.04648f
C10413 VDD.n1812 GND 0.04532f
C10414 VDD.n1813 GND 0.04532f
C10415 VDD.n1814 GND 0.02293f
C10416 VDD.n1815 GND 0.02293f
C10417 VDD.n1816 GND 0.04648f
C10418 VDD.n1817 GND 0.02708f
C10419 VDD.n1818 GND 0.02293f
C10420 VDD.n1819 GND 0.04891f
C10421 VDD.n1820 GND 0.04648f
C10422 VDD.t167 GND 0.02104f
C10423 VDD.t665 GND 0.02104f
C10424 VDD.t233 GND 0.02114f
C10425 VDD.t230 GND 0.02114f
C10426 VDD.n1821 GND 0.44561f
C10427 VDD.n1822 GND 0.04891f
C10428 VDD.n1823 GND 0.04648f
C10429 VDD.n1824 GND 0.02293f
C10430 VDD.n1825 GND 0.04648f
C10431 VDD.n1826 GND 0.02708f
C10432 VDD.n1827 GND 0.02293f
C10433 VDD.n1828 GND 0.04532f
C10434 VDD.n1829 GND 0.02293f
C10435 VDD.n1830 GND 0.02708f
C10436 VDD.n1831 GND 0.04532f
C10437 VDD.n1832 GND 0.02293f
C10438 VDD.n1833 GND 0.04891f
C10439 VDD.n1834 GND 0.05737f
C10440 VDD.n1835 GND 0.02055f
C10441 VDD.n1836 GND 0.08471f
C10442 VDD.n1837 GND 0.95576f
C10443 VDD.t445 GND 0.02114f
C10444 VDD.t921 GND 0.02114f
C10445 VDD.t312 GND 0.02114f
C10446 VDD.t417 GND 0.02114f
C10447 VDD.t256 GND 0.02104f
C10448 VDD.t433 GND 0.02114f
C10449 VDD.t311 GND 0.02114f
C10450 VDD.t274 GND 0.02114f
C10451 VDD.t591 GND 0.02114f
C10452 VDD.t141 GND 0.02104f
C10453 VDD.t647 GND 0.02104f
C10454 VDD.n1838 GND 0.95576f
C10455 VDD.n1839 GND 0.08471f
C10456 VDD.n1840 GND 0.04891f
C10457 VDD.n1841 GND 0.04648f
C10458 VDD.n1842 GND 0.02293f
C10459 VDD.n1843 GND 0.04648f
C10460 VDD.n1844 GND 0.02708f
C10461 VDD.n1845 GND 0.02293f
C10462 VDD.n1846 GND 0.04532f
C10463 VDD.n1847 GND 0.02293f
C10464 VDD.n1848 GND 0.02708f
C10465 VDD.n1849 GND 0.04532f
C10466 VDD.n1850 GND 0.02293f
C10467 VDD.n1851 GND 0.04891f
C10468 VDD.n1852 GND 0.05737f
C10469 VDD.n1853 GND 0.02055f
C10470 VDD.n1854 GND 0.44561f
C10471 VDD.n1855 GND 0.14059f
C10472 VDD.n1856 GND 0.04891f
C10473 VDD.n1857 GND 0.04648f
C10474 VDD.n1858 GND 0.02293f
C10475 VDD.n1859 GND 0.04648f
C10476 VDD.n1860 GND 0.02708f
C10477 VDD.n1861 GND 0.02293f
C10478 VDD.n1862 GND 0.04532f
C10479 VDD.n1863 GND 0.02293f
C10480 VDD.n1864 GND 0.02708f
C10481 VDD.n1865 GND 0.04532f
C10482 VDD.n1866 GND 0.02293f
C10483 VDD.n1867 GND 0.04891f
C10484 VDD.n1868 GND 0.05737f
C10485 VDD.n1869 GND 0.02055f
C10486 VDD.n1870 GND 0.02497f
C10487 VDD.n1871 GND 0.04648f
C10488 VDD.n1872 GND 0.04648f
C10489 VDD.n1873 GND 0.02708f
C10490 VDD.n1874 GND 0.02497f
C10491 VDD.n1875 GND 0.08328f
C10492 VDD.n1876 GND 0.01566f
C10493 VDD.n1877 GND 0.18236f
C10494 VDD.n1878 GND 0.03549f
C10495 VDD.n1879 GND 0.04891f
C10496 VDD.n1880 GND 0.04648f
C10497 VDD.n1881 GND 0.02293f
C10498 VDD.n1882 GND 0.04648f
C10499 VDD.n1883 GND 0.02708f
C10500 VDD.n1884 GND 0.02293f
C10501 VDD.n1885 GND 0.04532f
C10502 VDD.n1886 GND 0.02293f
C10503 VDD.n1887 GND 0.02708f
C10504 VDD.n1888 GND 0.04532f
C10505 VDD.n1889 GND 0.02293f
C10506 VDD.n1890 GND 0.04891f
C10507 VDD.n1891 GND 0.05737f
C10508 VDD.n1892 GND 0.02055f
C10509 VDD.n1893 GND 0.44561f
C10510 VDD.n1894 GND 0.14059f
C10511 VDD.n1895 GND 0.04891f
C10512 VDD.n1896 GND 0.04648f
C10513 VDD.n1897 GND 0.02293f
C10514 VDD.n1898 GND 0.04648f
C10515 VDD.n1899 GND 0.02708f
C10516 VDD.n1900 GND 0.02293f
C10517 VDD.n1901 GND 0.04532f
C10518 VDD.n1902 GND 0.02293f
C10519 VDD.n1903 GND 0.02708f
C10520 VDD.n1904 GND 0.04532f
C10521 VDD.n1905 GND 0.02293f
C10522 VDD.n1906 GND 0.04891f
C10523 VDD.n1907 GND 0.05737f
C10524 VDD.n1908 GND 0.02813f
C10525 VDD.n1909 GND 0.02324f
C10526 VDD.n1910 GND 0.05737f
C10527 VDD.n1911 GND 0.04891f
C10528 VDD.n1912 GND 0.02293f
C10529 VDD.n1913 GND 0.02708f
C10530 VDD.n1914 GND 0.04648f
C10531 VDD.n1915 GND 0.02293f
C10532 VDD.n1916 GND 0.02293f
C10533 VDD.n1917 GND 0.02708f
C10534 VDD.n1918 GND 0.04648f
C10535 VDD.n1919 GND 0.02708f
C10536 VDD.n1920 GND 0.04648f
C10537 VDD.n1921 GND 3.19829f
C10538 VDD.n1922 GND 0.04648f
C10539 VDD.n1923 GND 0.04532f
C10540 VDD.n1924 GND 0.02293f
C10541 VDD.n1925 GND 0.04891f
C10542 VDD.n1926 GND 0.05737f
C10543 VDD.n1927 GND 0.02813f
C10544 VDD.n1928 GND 0.14059f
C10545 VDD.n1929 GND 0.44561f
C10546 VDD.n1930 GND 0.02055f
C10547 VDD.n1931 GND 0.05737f
C10548 VDD.n1932 GND 0.04891f
C10549 VDD.n1933 GND 0.02293f
C10550 VDD.n1934 GND 0.02708f
C10551 VDD.n1935 GND 0.02293f
C10552 VDD.n1936 GND 0.04532f
C10553 VDD.t140 GND 4.12913f
C10554 VDD.n1937 GND 0.04532f
C10555 VDD.n1938 GND 0.04648f
C10556 VDD.n1939 GND 0.05737f
C10557 VDD.n1940 GND 0.01303f
C10558 VDD.n1941 GND 0.95576f
C10559 VDD.n1942 GND 0.08471f
C10560 VDD.n1943 GND 0.01566f
C10561 VDD.n1944 GND 0.08328f
C10562 VDD.n1945 GND 0.04648f
C10563 VDD.n1946 GND 3.47277f
C10564 VDD.n1947 GND 0.04648f
C10565 VDD.n1948 GND 0.05737f
C10566 VDD.n1949 GND 0.0171f
C10567 VDD.n1950 GND 0.064f
C10568 VDD.n1953 GND 0.06555f
C10569 VDD.n1954 GND 0.03083f
C10570 VDD.t139 GND 0.08047f
C10571 VDD.n1955 GND 0.03534f
C10572 VDD.t941 GND 0.15471f
C10573 VDD.n1956 GND 0.03238f
C10574 VDD.n1957 GND 0.02607f
C10575 VDD.n1958 GND 0.09595f
C10576 VDD.t166 GND 0.08047f
C10577 VDD.n1959 GND 0.03534f
C10578 VDD.t926 GND 0.15471f
C10579 VDD.n1960 GND 0.03238f
C10580 VDD.n1961 GND 0.02607f
C10581 VDD.n1963 GND 0.24365f
C10582 VDD.n1964 GND 0.03496f
C10583 VDD.n1965 GND 1.7026f
C10584 VDD.n1966 GND 1.45762f
C10585 VDD.t963 GND 0.15539f
C10586 VDD.n1967 GND 0.06697f
C10587 VDD.t155 GND 0.07226f
C10588 VDD.n1968 GND 0.05627f
C10589 VDD.n1969 GND 0.05442f
C10590 VDD.n1970 GND 0.04255f
C10591 VDD.n1971 GND 0.05152f
C10592 VDD.t217 GND 0.02114f
C10593 VDD.t367 GND 0.02114f
C10594 VDD.n1972 GND 0.14059f
C10595 VDD.n1973 GND 0.04891f
C10596 VDD.n1974 GND 0.04648f
C10597 VDD.n1975 GND 0.04891f
C10598 VDD.n1976 GND 0.04532f
C10599 VDD.n1977 GND 0.04532f
C10600 VDD.t156 GND 4.12913f
C10601 VDD.n1978 GND 0.04648f
C10602 VDD.n1979 GND 0.04648f
C10603 VDD.n1980 GND 0.04648f
C10604 VDD.n1981 GND 0.04648f
C10605 VDD.n1982 GND 0.04648f
C10606 VDD.n1983 GND 0.04648f
C10607 VDD.n1984 GND 3.47277f
C10608 VDD.n1985 GND 0.04648f
C10609 VDD.n1986 GND 0.04648f
C10610 VDD.n1987 GND 0.04648f
C10611 VDD.n1988 GND 0.04648f
C10612 VDD.n1989 GND 0.04532f
C10613 VDD.n1990 GND 0.04532f
C10614 VDD.n1991 GND 0.02497f
C10615 VDD.n1992 GND 0.02497f
C10616 VDD.t710 GND 0.02104f
C10617 VDD.n1993 GND 0.22365f
C10618 VDD.t157 GND 0.02104f
C10619 VDD.t668 GND 0.02104f
C10620 VDD.n1994 GND 0.04891f
C10621 VDD.n1995 GND 0.04891f
C10622 VDD.n1996 GND 0.04532f
C10623 VDD.n1997 GND 0.04648f
C10624 VDD.n1998 GND 0.02293f
C10625 VDD.n1999 GND 0.02708f
C10626 VDD.n2000 GND 0.02293f
C10627 VDD.n2001 GND 0.04532f
C10628 VDD.n2002 GND 0.04532f
C10629 VDD.n2003 GND 0.04532f
C10630 VDD.n2004 GND 0.04532f
C10631 VDD.n2005 GND 0.04532f
C10632 VDD.n2006 GND 0.04532f
C10633 VDD.n2007 GND 0.04532f
C10634 VDD.n2008 GND 0.04532f
C10635 VDD.n2009 GND 0.04532f
C10636 VDD.n2010 GND 0.04532f
C10637 VDD.n2011 GND 0.04532f
C10638 VDD.n2012 GND 0.04532f
C10639 VDD.n2013 GND 0.04532f
C10640 VDD.n2014 GND 0.04532f
C10641 VDD.n2015 GND 0.04532f
C10642 VDD.n2016 GND 0.04532f
C10643 VDD.n2017 GND 0.04532f
C10644 VDD.n2018 GND 0.04532f
C10645 VDD.n2019 GND 0.04532f
C10646 VDD.n2020 GND 0.04532f
C10647 VDD.n2021 GND 0.02293f
C10648 VDD.n2022 GND 0.02293f
C10649 VDD.n2023 GND 0.02708f
C10650 VDD.n2024 GND 0.04648f
C10651 VDD.n2025 GND 3.19829f
C10652 VDD.n2026 GND 0.04532f
C10653 VDD.n2027 GND 0.04648f
C10654 VDD.n2028 GND 0.04648f
C10655 VDD.n2029 GND 0.04891f
C10656 VDD.n2030 GND 0.02293f
C10657 VDD.t551 GND 0.02114f
C10658 VDD.t533 GND 0.02114f
C10659 VDD.t366 GND 0.02114f
C10660 VDD.t522 GND 0.02114f
C10661 VDD.n2031 GND 0.02324f
C10662 VDD.n2032 GND 0.04891f
C10663 VDD.n2033 GND 0.04648f
C10664 VDD.n2034 GND 0.02293f
C10665 VDD.n2035 GND 0.04648f
C10666 VDD.n2036 GND 0.02708f
C10667 VDD.n2037 GND 0.02293f
C10668 VDD.n2038 GND 0.02708f
C10669 VDD.n2039 GND 0.02293f
C10670 VDD.n2040 GND 0.04532f
C10671 VDD.n2041 GND 0.04532f
C10672 VDD.n2042 GND 0.04532f
C10673 VDD.n2043 GND 0.02293f
C10674 VDD.n2044 GND 0.02293f
C10675 VDD.n2045 GND 0.02708f
C10676 VDD.n2046 GND 0.04648f
C10677 VDD.n2047 GND 0.04648f
C10678 VDD.n2048 GND 0.04648f
C10679 VDD.n2049 GND 0.04648f
C10680 VDD.n2050 GND 0.04532f
C10681 VDD.n2051 GND 0.04532f
C10682 VDD.n2052 GND 0.02293f
C10683 VDD.n2053 GND 0.02293f
C10684 VDD.n2054 GND 0.04648f
C10685 VDD.n2055 GND 0.02708f
C10686 VDD.n2056 GND 0.02293f
C10687 VDD.n2057 GND 0.04891f
C10688 VDD.n2058 GND 0.04648f
C10689 VDD.n2059 GND 0.05737f
C10690 VDD.n2060 GND 0.04891f
C10691 VDD.n2061 GND 0.02293f
C10692 VDD.n2062 GND 0.02708f
C10693 VDD.n2063 GND 0.04648f
C10694 VDD.n2064 GND 0.04532f
C10695 VDD.n2065 GND 0.04532f
C10696 VDD.n2066 GND 0.02293f
C10697 VDD.n2067 GND 0.02708f
C10698 VDD.n2068 GND 0.04648f
C10699 VDD.n2069 GND 0.04648f
C10700 VDD.n2070 GND 0.04648f
C10701 VDD.n2071 GND 0.04532f
C10702 VDD.n2072 GND 0.04532f
C10703 VDD.n2073 GND 0.02293f
C10704 VDD.n2074 GND 0.02293f
C10705 VDD.n2075 GND 0.04648f
C10706 VDD.n2076 GND 0.02708f
C10707 VDD.n2077 GND 0.02293f
C10708 VDD.n2078 GND 0.04891f
C10709 VDD.n2079 GND 0.04648f
C10710 VDD.t159 GND 0.02104f
C10711 VDD.t678 GND 0.02104f
C10712 VDD.t244 GND 0.02114f
C10713 VDD.t321 GND 0.02114f
C10714 VDD.n2080 GND 0.44561f
C10715 VDD.n2081 GND 0.04891f
C10716 VDD.n2082 GND 0.04648f
C10717 VDD.n2083 GND 0.02293f
C10718 VDD.n2084 GND 0.04648f
C10719 VDD.n2085 GND 0.02708f
C10720 VDD.n2086 GND 0.02293f
C10721 VDD.n2087 GND 0.04532f
C10722 VDD.n2088 GND 0.02293f
C10723 VDD.n2089 GND 0.02708f
C10724 VDD.n2090 GND 0.04532f
C10725 VDD.n2091 GND 0.02293f
C10726 VDD.n2092 GND 0.04891f
C10727 VDD.n2093 GND 0.05737f
C10728 VDD.n2094 GND 0.02055f
C10729 VDD.n2095 GND 0.08471f
C10730 VDD.n2096 GND 0.95576f
C10731 VDD.t284 GND 0.02114f
C10732 VDD.t582 GND 0.02114f
C10733 VDD.t36 GND 0.02114f
C10734 VDD.t786 GND 0.02114f
C10735 VDD.t291 GND 0.02104f
C10736 VDD.t882 GND 0.02114f
C10737 VDD.t515 GND 0.02114f
C10738 VDD.t265 GND 0.02114f
C10739 VDD.t264 GND 0.02114f
C10740 VDD.t119 GND 0.02104f
C10741 VDD.t664 GND 0.02104f
C10742 VDD.n2097 GND 0.95576f
C10743 VDD.n2098 GND 0.08471f
C10744 VDD.n2099 GND 0.04891f
C10745 VDD.n2100 GND 0.04648f
C10746 VDD.n2101 GND 0.02293f
C10747 VDD.n2102 GND 0.04648f
C10748 VDD.n2103 GND 0.02708f
C10749 VDD.n2104 GND 0.02293f
C10750 VDD.n2105 GND 0.04532f
C10751 VDD.n2106 GND 0.02293f
C10752 VDD.n2107 GND 0.02708f
C10753 VDD.n2108 GND 0.04532f
C10754 VDD.n2109 GND 0.02293f
C10755 VDD.n2110 GND 0.04891f
C10756 VDD.n2111 GND 0.05737f
C10757 VDD.n2112 GND 0.02055f
C10758 VDD.n2113 GND 0.44561f
C10759 VDD.n2114 GND 0.14059f
C10760 VDD.n2115 GND 0.04891f
C10761 VDD.n2116 GND 0.04648f
C10762 VDD.n2117 GND 0.02293f
C10763 VDD.n2118 GND 0.04648f
C10764 VDD.n2119 GND 0.02708f
C10765 VDD.n2120 GND 0.02293f
C10766 VDD.n2121 GND 0.04532f
C10767 VDD.n2122 GND 0.02293f
C10768 VDD.n2123 GND 0.02708f
C10769 VDD.n2124 GND 0.04532f
C10770 VDD.n2125 GND 0.02293f
C10771 VDD.n2126 GND 0.04891f
C10772 VDD.n2127 GND 0.05737f
C10773 VDD.n2128 GND 0.02055f
C10774 VDD.n2129 GND 0.02497f
C10775 VDD.n2130 GND 0.04648f
C10776 VDD.n2131 GND 0.04648f
C10777 VDD.n2132 GND 0.02708f
C10778 VDD.n2133 GND 0.02497f
C10779 VDD.n2134 GND 0.08328f
C10780 VDD.n2135 GND 0.01566f
C10781 VDD.n2136 GND 0.18236f
C10782 VDD.n2137 GND 0.03549f
C10783 VDD.n2138 GND 0.04891f
C10784 VDD.n2139 GND 0.04648f
C10785 VDD.n2140 GND 0.02293f
C10786 VDD.n2141 GND 0.04648f
C10787 VDD.n2142 GND 0.02708f
C10788 VDD.n2143 GND 0.02293f
C10789 VDD.n2144 GND 0.04532f
C10790 VDD.n2145 GND 0.02293f
C10791 VDD.n2146 GND 0.02708f
C10792 VDD.n2147 GND 0.04532f
C10793 VDD.n2148 GND 0.02293f
C10794 VDD.n2149 GND 0.04891f
C10795 VDD.n2150 GND 0.05737f
C10796 VDD.n2151 GND 0.02055f
C10797 VDD.n2152 GND 0.44561f
C10798 VDD.n2153 GND 0.14059f
C10799 VDD.n2154 GND 0.04891f
C10800 VDD.n2155 GND 0.04648f
C10801 VDD.n2156 GND 0.02293f
C10802 VDD.n2157 GND 0.04648f
C10803 VDD.n2158 GND 0.02708f
C10804 VDD.n2159 GND 0.02293f
C10805 VDD.n2160 GND 0.04532f
C10806 VDD.n2161 GND 0.02293f
C10807 VDD.n2162 GND 0.02708f
C10808 VDD.n2163 GND 0.04532f
C10809 VDD.n2164 GND 0.02293f
C10810 VDD.n2165 GND 0.04891f
C10811 VDD.n2166 GND 0.05737f
C10812 VDD.n2167 GND 0.02813f
C10813 VDD.n2168 GND 0.02324f
C10814 VDD.n2169 GND 0.05737f
C10815 VDD.n2170 GND 0.04891f
C10816 VDD.n2171 GND 0.02293f
C10817 VDD.n2172 GND 0.02708f
C10818 VDD.n2173 GND 0.04648f
C10819 VDD.n2174 GND 0.02293f
C10820 VDD.n2175 GND 0.02293f
C10821 VDD.n2176 GND 0.02708f
C10822 VDD.n2177 GND 0.04648f
C10823 VDD.n2178 GND 0.02708f
C10824 VDD.n2179 GND 0.04648f
C10825 VDD.n2180 GND 3.19829f
C10826 VDD.n2181 GND 0.04648f
C10827 VDD.n2182 GND 0.04532f
C10828 VDD.n2183 GND 0.02293f
C10829 VDD.n2184 GND 0.04891f
C10830 VDD.n2185 GND 0.05737f
C10831 VDD.n2186 GND 0.02813f
C10832 VDD.n2187 GND 0.14059f
C10833 VDD.n2188 GND 0.44561f
C10834 VDD.n2189 GND 0.02055f
C10835 VDD.n2190 GND 0.05737f
C10836 VDD.n2191 GND 0.04891f
C10837 VDD.n2192 GND 0.02293f
C10838 VDD.n2193 GND 0.02708f
C10839 VDD.n2194 GND 0.02293f
C10840 VDD.n2195 GND 0.04532f
C10841 VDD.t35 GND 4.12913f
C10842 VDD.n2196 GND 0.04532f
C10843 VDD.n2197 GND 0.04648f
C10844 VDD.n2198 GND 0.05737f
C10845 VDD.n2199 GND 0.01303f
C10846 VDD.n2200 GND 0.95576f
C10847 VDD.n2201 GND 0.08471f
C10848 VDD.n2202 GND 0.01566f
C10849 VDD.n2203 GND 0.08328f
C10850 VDD.n2204 GND 0.04648f
C10851 VDD.n2205 GND 3.47277f
C10852 VDD.n2206 GND 0.04648f
C10853 VDD.n2207 GND 0.05737f
C10854 VDD.n2208 GND 0.0171f
C10855 VDD.n2209 GND 0.064f
C10856 VDD.n2212 GND 0.06555f
C10857 VDD.n2213 GND 0.03083f
C10858 VDD.t118 GND 0.08047f
C10859 VDD.n2214 GND 0.03534f
C10860 VDD.t936 GND 0.15471f
C10861 VDD.n2215 GND 0.03238f
C10862 VDD.n2216 GND 0.02607f
C10863 VDD.n2217 GND 0.09595f
C10864 VDD.t158 GND 0.08047f
C10865 VDD.n2218 GND 0.03534f
C10866 VDD.t973 GND 0.15471f
C10867 VDD.n2219 GND 0.03238f
C10868 VDD.n2220 GND 0.02607f
C10869 VDD.n2222 GND 0.24365f
C10870 VDD.n2223 GND 0.03496f
C10871 VDD.n2224 GND 1.54242f
C10872 VDD.n2225 GND 1.31199f
C10873 VDD.t961 GND 0.15539f
C10874 VDD.n2226 GND 0.06697f
C10875 VDD.t212 GND 0.07226f
C10876 VDD.n2227 GND 0.05627f
C10877 VDD.n2228 GND 0.05442f
C10878 VDD.n2229 GND 0.04255f
C10879 VDD.n2230 GND 0.05152f
C10880 VDD.t633 GND 0.02114f
C10881 VDD.t909 GND 0.02114f
C10882 VDD.n2231 GND 0.14059f
C10883 VDD.n2232 GND 0.04891f
C10884 VDD.n2233 GND 0.04648f
C10885 VDD.n2234 GND 0.04891f
C10886 VDD.n2235 GND 0.04532f
C10887 VDD.n2236 GND 0.04532f
C10888 VDD.t213 GND 4.12913f
C10889 VDD.n2237 GND 0.04648f
C10890 VDD.n2238 GND 0.04648f
C10891 VDD.n2239 GND 0.04648f
C10892 VDD.n2240 GND 0.04648f
C10893 VDD.n2241 GND 0.04648f
C10894 VDD.n2242 GND 0.04648f
C10895 VDD.n2243 GND 3.47277f
C10896 VDD.n2244 GND 0.04648f
C10897 VDD.n2245 GND 0.04648f
C10898 VDD.n2246 GND 0.04648f
C10899 VDD.n2247 GND 0.04648f
C10900 VDD.n2248 GND 0.04532f
C10901 VDD.n2249 GND 0.04532f
C10902 VDD.n2250 GND 0.02497f
C10903 VDD.n2251 GND 0.02497f
C10904 VDD.t552 GND 0.02104f
C10905 VDD.n2252 GND 0.22365f
C10906 VDD.t214 GND 0.02104f
C10907 VDD.t671 GND 0.02104f
C10908 VDD.n2253 GND 0.04891f
C10909 VDD.n2254 GND 0.04891f
C10910 VDD.n2255 GND 0.04532f
C10911 VDD.n2256 GND 0.04648f
C10912 VDD.n2257 GND 0.02293f
C10913 VDD.n2258 GND 0.02708f
C10914 VDD.n2259 GND 0.02293f
C10915 VDD.n2260 GND 0.04532f
C10916 VDD.n2261 GND 0.04532f
C10917 VDD.n2262 GND 0.04532f
C10918 VDD.n2263 GND 0.04532f
C10919 VDD.n2264 GND 0.04532f
C10920 VDD.n2265 GND 0.04532f
C10921 VDD.n2266 GND 0.04532f
C10922 VDD.n2267 GND 0.04532f
C10923 VDD.n2268 GND 0.04532f
C10924 VDD.n2269 GND 0.04532f
C10925 VDD.n2270 GND 0.04532f
C10926 VDD.n2271 GND 0.04532f
C10927 VDD.n2272 GND 0.04532f
C10928 VDD.n2273 GND 0.04532f
C10929 VDD.n2274 GND 0.04532f
C10930 VDD.n2275 GND 0.04532f
C10931 VDD.n2276 GND 0.04532f
C10932 VDD.n2277 GND 0.04532f
C10933 VDD.n2278 GND 0.04532f
C10934 VDD.n2279 GND 0.04532f
C10935 VDD.n2280 GND 0.02293f
C10936 VDD.n2281 GND 0.02293f
C10937 VDD.n2282 GND 0.02708f
C10938 VDD.n2283 GND 0.04648f
C10939 VDD.n2284 GND 3.19829f
C10940 VDD.n2285 GND 0.04532f
C10941 VDD.n2286 GND 0.04648f
C10942 VDD.n2287 GND 0.04648f
C10943 VDD.n2288 GND 0.04891f
C10944 VDD.n2289 GND 0.02293f
C10945 VDD.t787 GND 0.02114f
C10946 VDD.t363 GND 0.02114f
C10947 VDD.t404 GND 0.02114f
C10948 VDD.t785 GND 0.02114f
C10949 VDD.n2290 GND 0.02324f
C10950 VDD.n2291 GND 0.04891f
C10951 VDD.n2292 GND 0.04648f
C10952 VDD.n2293 GND 0.02293f
C10953 VDD.n2294 GND 0.04648f
C10954 VDD.n2295 GND 0.02708f
C10955 VDD.n2296 GND 0.02293f
C10956 VDD.n2297 GND 0.02708f
C10957 VDD.n2298 GND 0.02293f
C10958 VDD.n2299 GND 0.04532f
C10959 VDD.n2300 GND 0.04532f
C10960 VDD.n2301 GND 0.04532f
C10961 VDD.n2302 GND 0.02293f
C10962 VDD.n2303 GND 0.02293f
C10963 VDD.n2304 GND 0.02708f
C10964 VDD.n2305 GND 0.04648f
C10965 VDD.n2306 GND 0.04648f
C10966 VDD.n2307 GND 0.04648f
C10967 VDD.n2308 GND 0.04648f
C10968 VDD.n2309 GND 0.04532f
C10969 VDD.n2310 GND 0.04532f
C10970 VDD.n2311 GND 0.02293f
C10971 VDD.n2312 GND 0.02293f
C10972 VDD.n2313 GND 0.04648f
C10973 VDD.n2314 GND 0.02708f
C10974 VDD.n2315 GND 0.02293f
C10975 VDD.n2316 GND 0.04891f
C10976 VDD.n2317 GND 0.04648f
C10977 VDD.n2318 GND 0.05737f
C10978 VDD.n2319 GND 0.04891f
C10979 VDD.n2320 GND 0.02293f
C10980 VDD.n2321 GND 0.02708f
C10981 VDD.n2322 GND 0.04648f
C10982 VDD.n2323 GND 0.04532f
C10983 VDD.n2324 GND 0.04532f
C10984 VDD.n2325 GND 0.02293f
C10985 VDD.n2326 GND 0.02708f
C10986 VDD.n2327 GND 0.04648f
C10987 VDD.n2328 GND 0.04648f
C10988 VDD.n2329 GND 0.04648f
C10989 VDD.n2330 GND 0.04532f
C10990 VDD.n2331 GND 0.04532f
C10991 VDD.n2332 GND 0.02293f
C10992 VDD.n2333 GND 0.02293f
C10993 VDD.n2334 GND 0.04648f
C10994 VDD.n2335 GND 0.02708f
C10995 VDD.n2336 GND 0.02293f
C10996 VDD.n2337 GND 0.04891f
C10997 VDD.n2338 GND 0.04648f
C10998 VDD.t165 GND 0.02104f
C10999 VDD.t652 GND 0.02104f
C11000 VDD.t322 GND 0.02114f
C11001 VDD.t817 GND 0.02114f
C11002 VDD.n2339 GND 0.44561f
C11003 VDD.n2340 GND 0.04891f
C11004 VDD.n2341 GND 0.04648f
C11005 VDD.n2342 GND 0.02293f
C11006 VDD.n2343 GND 0.04648f
C11007 VDD.n2344 GND 0.02708f
C11008 VDD.n2345 GND 0.02293f
C11009 VDD.n2346 GND 0.04532f
C11010 VDD.n2347 GND 0.02293f
C11011 VDD.n2348 GND 0.02708f
C11012 VDD.n2349 GND 0.04532f
C11013 VDD.n2350 GND 0.02293f
C11014 VDD.n2351 GND 0.04891f
C11015 VDD.n2352 GND 0.05737f
C11016 VDD.n2353 GND 0.02055f
C11017 VDD.n2354 GND 0.08471f
C11018 VDD.n2355 GND 0.95576f
C11019 VDD.t616 GND 0.02114f
C11020 VDD.t920 GND 0.02114f
C11021 VDD.t723 GND 0.02114f
C11022 VDD.t868 GND 0.02114f
C11023 VDD.t240 GND 0.02104f
C11024 VDD.t867 GND 0.02114f
C11025 VDD.t334 GND 0.02114f
C11026 VDD.t30 GND 0.02114f
C11027 VDD.t218 GND 0.02114f
C11028 VDD.t131 GND 0.02104f
C11029 VDD.t696 GND 0.02104f
C11030 VDD.n2356 GND 0.95576f
C11031 VDD.n2357 GND 0.08471f
C11032 VDD.n2358 GND 0.04891f
C11033 VDD.n2359 GND 0.04648f
C11034 VDD.n2360 GND 0.02293f
C11035 VDD.n2361 GND 0.04648f
C11036 VDD.n2362 GND 0.02708f
C11037 VDD.n2363 GND 0.02293f
C11038 VDD.n2364 GND 0.04532f
C11039 VDD.n2365 GND 0.02293f
C11040 VDD.n2366 GND 0.02708f
C11041 VDD.n2367 GND 0.04532f
C11042 VDD.n2368 GND 0.02293f
C11043 VDD.n2369 GND 0.04891f
C11044 VDD.n2370 GND 0.05737f
C11045 VDD.n2371 GND 0.02055f
C11046 VDD.n2372 GND 0.44561f
C11047 VDD.n2373 GND 0.14059f
C11048 VDD.n2374 GND 0.04891f
C11049 VDD.n2375 GND 0.04648f
C11050 VDD.n2376 GND 0.02293f
C11051 VDD.n2377 GND 0.04648f
C11052 VDD.n2378 GND 0.02708f
C11053 VDD.n2379 GND 0.02293f
C11054 VDD.n2380 GND 0.04532f
C11055 VDD.n2381 GND 0.02293f
C11056 VDD.n2382 GND 0.02708f
C11057 VDD.n2383 GND 0.04532f
C11058 VDD.n2384 GND 0.02293f
C11059 VDD.n2385 GND 0.04891f
C11060 VDD.n2386 GND 0.05737f
C11061 VDD.n2387 GND 0.02055f
C11062 VDD.n2388 GND 0.02497f
C11063 VDD.n2389 GND 0.04648f
C11064 VDD.n2390 GND 0.04648f
C11065 VDD.n2391 GND 0.02708f
C11066 VDD.n2392 GND 0.02497f
C11067 VDD.n2393 GND 0.08328f
C11068 VDD.n2394 GND 0.01566f
C11069 VDD.n2395 GND 0.18236f
C11070 VDD.n2396 GND 0.03549f
C11071 VDD.n2397 GND 0.04891f
C11072 VDD.n2398 GND 0.04648f
C11073 VDD.n2399 GND 0.02293f
C11074 VDD.n2400 GND 0.04648f
C11075 VDD.n2401 GND 0.02708f
C11076 VDD.n2402 GND 0.02293f
C11077 VDD.n2403 GND 0.04532f
C11078 VDD.n2404 GND 0.02293f
C11079 VDD.n2405 GND 0.02708f
C11080 VDD.n2406 GND 0.04532f
C11081 VDD.n2407 GND 0.02293f
C11082 VDD.n2408 GND 0.04891f
C11083 VDD.n2409 GND 0.05737f
C11084 VDD.n2410 GND 0.02055f
C11085 VDD.n2411 GND 0.44561f
C11086 VDD.n2412 GND 0.14059f
C11087 VDD.n2413 GND 0.04891f
C11088 VDD.n2414 GND 0.04648f
C11089 VDD.n2415 GND 0.02293f
C11090 VDD.n2416 GND 0.04648f
C11091 VDD.n2417 GND 0.02708f
C11092 VDD.n2418 GND 0.02293f
C11093 VDD.n2419 GND 0.04532f
C11094 VDD.n2420 GND 0.02293f
C11095 VDD.n2421 GND 0.02708f
C11096 VDD.n2422 GND 0.04532f
C11097 VDD.n2423 GND 0.02293f
C11098 VDD.n2424 GND 0.04891f
C11099 VDD.n2425 GND 0.05737f
C11100 VDD.n2426 GND 0.02813f
C11101 VDD.n2427 GND 0.02324f
C11102 VDD.n2428 GND 0.05737f
C11103 VDD.n2429 GND 0.04891f
C11104 VDD.n2430 GND 0.02293f
C11105 VDD.n2431 GND 0.02708f
C11106 VDD.n2432 GND 0.04648f
C11107 VDD.n2433 GND 0.02293f
C11108 VDD.n2434 GND 0.02293f
C11109 VDD.n2435 GND 0.02708f
C11110 VDD.n2436 GND 0.04648f
C11111 VDD.n2437 GND 0.02708f
C11112 VDD.n2438 GND 0.04648f
C11113 VDD.n2439 GND 3.19829f
C11114 VDD.n2440 GND 0.04648f
C11115 VDD.n2441 GND 0.04532f
C11116 VDD.n2442 GND 0.02293f
C11117 VDD.n2443 GND 0.04891f
C11118 VDD.n2444 GND 0.05737f
C11119 VDD.n2445 GND 0.02813f
C11120 VDD.n2446 GND 0.14059f
C11121 VDD.n2447 GND 0.44561f
C11122 VDD.n2448 GND 0.02055f
C11123 VDD.n2449 GND 0.05737f
C11124 VDD.n2450 GND 0.04891f
C11125 VDD.n2451 GND 0.02293f
C11126 VDD.n2452 GND 0.02708f
C11127 VDD.n2453 GND 0.02293f
C11128 VDD.n2454 GND 0.04532f
C11129 VDD.t29 GND 4.12913f
C11130 VDD.n2455 GND 0.04532f
C11131 VDD.n2456 GND 0.04648f
C11132 VDD.n2457 GND 0.05737f
C11133 VDD.n2458 GND 0.01303f
C11134 VDD.n2459 GND 0.95576f
C11135 VDD.n2460 GND 0.08471f
C11136 VDD.n2461 GND 0.01566f
C11137 VDD.n2462 GND 0.08328f
C11138 VDD.n2463 GND 0.04648f
C11139 VDD.n2464 GND 3.47277f
C11140 VDD.n2465 GND 0.04648f
C11141 VDD.n2466 GND 0.05737f
C11142 VDD.n2467 GND 0.0171f
C11143 VDD.n2468 GND 0.064f
C11144 VDD.n2471 GND 0.06555f
C11145 VDD.n2472 GND 0.03083f
C11146 VDD.t130 GND 0.08047f
C11147 VDD.n2473 GND 0.03534f
C11148 VDD.t952 GND 0.15471f
C11149 VDD.n2474 GND 0.03238f
C11150 VDD.n2475 GND 0.02607f
C11151 VDD.n2476 GND 0.09595f
C11152 VDD.t164 GND 0.08047f
C11153 VDD.n2477 GND 0.03534f
C11154 VDD.t938 GND 0.15471f
C11155 VDD.n2478 GND 0.03238f
C11156 VDD.n2479 GND 0.02607f
C11157 VDD.n2481 GND 0.24365f
C11158 VDD.n2482 GND 0.03496f
C11159 VDD.n2483 GND 1.38223f
C11160 VDD.n2484 GND 1.16637f
C11161 VDD.t939 GND 0.15539f
C11162 VDD.n2485 GND 0.06697f
C11163 VDD.t160 GND 0.07226f
C11164 VDD.n2486 GND 0.05627f
C11165 VDD.n2487 GND 0.05442f
C11166 VDD.n2488 GND 0.04255f
C11167 VDD.n2489 GND 0.05152f
C11168 VDD.t84 GND 0.02114f
C11169 VDD.t351 GND 0.02114f
C11170 VDD.n2490 GND 0.14059f
C11171 VDD.n2491 GND 0.04891f
C11172 VDD.n2492 GND 0.04648f
C11173 VDD.n2493 GND 0.04891f
C11174 VDD.n2494 GND 0.04532f
C11175 VDD.n2495 GND 0.04532f
C11176 VDD.t72 GND 4.12913f
C11177 VDD.n2496 GND 0.04648f
C11178 VDD.n2497 GND 0.04648f
C11179 VDD.n2498 GND 0.04648f
C11180 VDD.n2499 GND 0.04648f
C11181 VDD.n2500 GND 0.04648f
C11182 VDD.n2501 GND 0.04648f
C11183 VDD.n2502 GND 3.47277f
C11184 VDD.n2503 GND 0.04648f
C11185 VDD.n2504 GND 0.04648f
C11186 VDD.n2505 GND 0.04648f
C11187 VDD.n2506 GND 0.04648f
C11188 VDD.n2507 GND 0.04532f
C11189 VDD.n2508 GND 0.04532f
C11190 VDD.n2509 GND 0.02497f
C11191 VDD.n2510 GND 0.02497f
C11192 VDD.t456 GND 0.02104f
C11193 VDD.n2511 GND 0.22365f
C11194 VDD.t161 GND 0.02104f
C11195 VDD.t672 GND 0.02104f
C11196 VDD.n2512 GND 0.04891f
C11197 VDD.n2513 GND 0.04891f
C11198 VDD.n2514 GND 0.04532f
C11199 VDD.n2515 GND 0.04648f
C11200 VDD.n2516 GND 0.02293f
C11201 VDD.n2517 GND 0.02708f
C11202 VDD.n2518 GND 0.02293f
C11203 VDD.n2519 GND 0.04532f
C11204 VDD.n2520 GND 0.04532f
C11205 VDD.n2521 GND 0.04532f
C11206 VDD.n2522 GND 0.04532f
C11207 VDD.n2523 GND 0.04532f
C11208 VDD.n2524 GND 0.04532f
C11209 VDD.n2525 GND 0.04532f
C11210 VDD.n2526 GND 0.04532f
C11211 VDD.n2527 GND 0.04532f
C11212 VDD.n2528 GND 0.04532f
C11213 VDD.n2529 GND 0.04532f
C11214 VDD.n2530 GND 0.04532f
C11215 VDD.n2531 GND 0.04532f
C11216 VDD.n2532 GND 0.04532f
C11217 VDD.n2533 GND 0.04532f
C11218 VDD.n2534 GND 0.04532f
C11219 VDD.n2535 GND 0.04532f
C11220 VDD.n2536 GND 0.04532f
C11221 VDD.n2537 GND 0.04532f
C11222 VDD.n2538 GND 0.04532f
C11223 VDD.n2539 GND 0.02293f
C11224 VDD.n2540 GND 0.02293f
C11225 VDD.n2541 GND 0.02708f
C11226 VDD.n2542 GND 0.04648f
C11227 VDD.n2543 GND 3.19829f
C11228 VDD.n2544 GND 0.04532f
C11229 VDD.n2545 GND 0.04648f
C11230 VDD.n2546 GND 0.04648f
C11231 VDD.n2547 GND 0.04891f
C11232 VDD.n2548 GND 0.02293f
C11233 VDD.t436 GND 0.02114f
C11234 VDD.t73 GND 0.02114f
C11235 VDD.t575 GND 0.02114f
C11236 VDD.t410 GND 0.02114f
C11237 VDD.n2549 GND 0.02324f
C11238 VDD.n2550 GND 0.04891f
C11239 VDD.n2551 GND 0.04648f
C11240 VDD.n2552 GND 0.02293f
C11241 VDD.n2553 GND 0.04648f
C11242 VDD.n2554 GND 0.02708f
C11243 VDD.n2555 GND 0.02293f
C11244 VDD.n2556 GND 0.02708f
C11245 VDD.n2557 GND 0.02293f
C11246 VDD.n2558 GND 0.04532f
C11247 VDD.n2559 GND 0.04532f
C11248 VDD.n2560 GND 0.04532f
C11249 VDD.n2561 GND 0.02293f
C11250 VDD.n2562 GND 0.02293f
C11251 VDD.n2563 GND 0.02708f
C11252 VDD.n2564 GND 0.04648f
C11253 VDD.n2565 GND 0.04648f
C11254 VDD.n2566 GND 0.04648f
C11255 VDD.n2567 GND 0.04648f
C11256 VDD.n2568 GND 0.04532f
C11257 VDD.n2569 GND 0.04532f
C11258 VDD.n2570 GND 0.02293f
C11259 VDD.n2571 GND 0.02293f
C11260 VDD.n2572 GND 0.04648f
C11261 VDD.n2573 GND 0.02708f
C11262 VDD.n2574 GND 0.02293f
C11263 VDD.n2575 GND 0.04891f
C11264 VDD.n2576 GND 0.04648f
C11265 VDD.n2577 GND 0.05737f
C11266 VDD.n2578 GND 0.04891f
C11267 VDD.n2579 GND 0.02293f
C11268 VDD.n2580 GND 0.02708f
C11269 VDD.n2581 GND 0.04648f
C11270 VDD.n2582 GND 0.04532f
C11271 VDD.n2583 GND 0.04532f
C11272 VDD.n2584 GND 0.02293f
C11273 VDD.n2585 GND 0.02708f
C11274 VDD.n2586 GND 0.04648f
C11275 VDD.n2587 GND 0.04648f
C11276 VDD.n2588 GND 0.04648f
C11277 VDD.n2589 GND 0.04532f
C11278 VDD.n2590 GND 0.04532f
C11279 VDD.n2591 GND 0.02293f
C11280 VDD.n2592 GND 0.02293f
C11281 VDD.n2593 GND 0.04648f
C11282 VDD.n2594 GND 0.02708f
C11283 VDD.n2595 GND 0.02293f
C11284 VDD.n2596 GND 0.04891f
C11285 VDD.n2597 GND 0.04648f
C11286 VDD.t163 GND 0.02104f
C11287 VDD.t679 GND 0.02104f
C11288 VDD.t323 GND 0.02114f
C11289 VDD.t231 GND 0.02114f
C11290 VDD.n2598 GND 0.44561f
C11291 VDD.n2599 GND 0.04891f
C11292 VDD.n2600 GND 0.04648f
C11293 VDD.n2601 GND 0.02293f
C11294 VDD.n2602 GND 0.04648f
C11295 VDD.n2603 GND 0.02708f
C11296 VDD.n2604 GND 0.02293f
C11297 VDD.n2605 GND 0.04532f
C11298 VDD.n2606 GND 0.02293f
C11299 VDD.n2607 GND 0.02708f
C11300 VDD.n2608 GND 0.04532f
C11301 VDD.n2609 GND 0.02293f
C11302 VDD.n2610 GND 0.04891f
C11303 VDD.n2611 GND 0.05737f
C11304 VDD.n2612 GND 0.02055f
C11305 VDD.n2613 GND 0.08471f
C11306 VDD.n2614 GND 0.95576f
C11307 VDD.t600 GND 0.02114f
C11308 VDD.t806 GND 0.02114f
C11309 VDD.t513 GND 0.02114f
C11310 VDD.t919 GND 0.02114f
C11311 VDD.t241 GND 0.02104f
C11312 VDD.t393 GND 0.02114f
C11313 VDD.t414 GND 0.02114f
C11314 VDD.t489 GND 0.02114f
C11315 VDD.t917 GND 0.02114f
C11316 VDD.t129 GND 0.02104f
C11317 VDD.t669 GND 0.02104f
C11318 VDD.n2615 GND 0.95576f
C11319 VDD.n2616 GND 0.08471f
C11320 VDD.n2617 GND 0.04891f
C11321 VDD.n2618 GND 0.04648f
C11322 VDD.n2619 GND 0.02293f
C11323 VDD.n2620 GND 0.04648f
C11324 VDD.n2621 GND 0.02708f
C11325 VDD.n2622 GND 0.02293f
C11326 VDD.n2623 GND 0.04532f
C11327 VDD.n2624 GND 0.02293f
C11328 VDD.n2625 GND 0.02708f
C11329 VDD.n2626 GND 0.04532f
C11330 VDD.n2627 GND 0.02293f
C11331 VDD.n2628 GND 0.04891f
C11332 VDD.n2629 GND 0.05737f
C11333 VDD.n2630 GND 0.02055f
C11334 VDD.n2631 GND 0.44561f
C11335 VDD.n2632 GND 0.14059f
C11336 VDD.n2633 GND 0.04891f
C11337 VDD.n2634 GND 0.04648f
C11338 VDD.n2635 GND 0.02293f
C11339 VDD.n2636 GND 0.04648f
C11340 VDD.n2637 GND 0.02708f
C11341 VDD.n2638 GND 0.02293f
C11342 VDD.n2639 GND 0.04532f
C11343 VDD.n2640 GND 0.02293f
C11344 VDD.n2641 GND 0.02708f
C11345 VDD.n2642 GND 0.04532f
C11346 VDD.n2643 GND 0.02293f
C11347 VDD.n2644 GND 0.04891f
C11348 VDD.n2645 GND 0.05737f
C11349 VDD.n2646 GND 0.02055f
C11350 VDD.n2647 GND 0.02497f
C11351 VDD.n2648 GND 0.04648f
C11352 VDD.n2649 GND 0.04648f
C11353 VDD.n2650 GND 0.02708f
C11354 VDD.n2651 GND 0.02497f
C11355 VDD.n2652 GND 0.08328f
C11356 VDD.n2653 GND 0.01566f
C11357 VDD.n2654 GND 0.18236f
C11358 VDD.n2655 GND 0.03549f
C11359 VDD.n2656 GND 0.04891f
C11360 VDD.n2657 GND 0.04648f
C11361 VDD.n2658 GND 0.02293f
C11362 VDD.n2659 GND 0.04648f
C11363 VDD.n2660 GND 0.02708f
C11364 VDD.n2661 GND 0.02293f
C11365 VDD.n2662 GND 0.04532f
C11366 VDD.n2663 GND 0.02293f
C11367 VDD.n2664 GND 0.02708f
C11368 VDD.n2665 GND 0.04532f
C11369 VDD.n2666 GND 0.02293f
C11370 VDD.n2667 GND 0.04891f
C11371 VDD.n2668 GND 0.05737f
C11372 VDD.n2669 GND 0.02055f
C11373 VDD.n2670 GND 0.44561f
C11374 VDD.n2671 GND 0.14059f
C11375 VDD.n2672 GND 0.04891f
C11376 VDD.n2673 GND 0.04648f
C11377 VDD.n2674 GND 0.02293f
C11378 VDD.n2675 GND 0.04648f
C11379 VDD.n2676 GND 0.02708f
C11380 VDD.n2677 GND 0.02293f
C11381 VDD.n2678 GND 0.04532f
C11382 VDD.n2679 GND 0.02293f
C11383 VDD.n2680 GND 0.02708f
C11384 VDD.n2681 GND 0.04532f
C11385 VDD.n2682 GND 0.02293f
C11386 VDD.n2683 GND 0.04891f
C11387 VDD.n2684 GND 0.05737f
C11388 VDD.n2685 GND 0.02813f
C11389 VDD.n2686 GND 0.02324f
C11390 VDD.n2687 GND 0.05737f
C11391 VDD.n2688 GND 0.04891f
C11392 VDD.n2689 GND 0.02293f
C11393 VDD.n2690 GND 0.02708f
C11394 VDD.n2691 GND 0.04648f
C11395 VDD.n2692 GND 0.02293f
C11396 VDD.n2693 GND 0.02293f
C11397 VDD.n2694 GND 0.02708f
C11398 VDD.n2695 GND 0.04648f
C11399 VDD.n2696 GND 0.02708f
C11400 VDD.n2697 GND 0.04648f
C11401 VDD.n2698 GND 3.19829f
C11402 VDD.n2699 GND 0.04648f
C11403 VDD.n2700 GND 0.04532f
C11404 VDD.n2701 GND 0.02293f
C11405 VDD.n2702 GND 0.04891f
C11406 VDD.n2703 GND 0.05737f
C11407 VDD.n2704 GND 0.02813f
C11408 VDD.n2705 GND 0.14059f
C11409 VDD.n2706 GND 0.44561f
C11410 VDD.n2707 GND 0.02055f
C11411 VDD.n2708 GND 0.05737f
C11412 VDD.n2709 GND 0.04891f
C11413 VDD.n2710 GND 0.02293f
C11414 VDD.n2711 GND 0.02708f
C11415 VDD.n2712 GND 0.02293f
C11416 VDD.n2713 GND 0.04532f
C11417 VDD.t83 GND 4.12913f
C11418 VDD.n2714 GND 0.04532f
C11419 VDD.n2715 GND 0.04648f
C11420 VDD.n2716 GND 0.05737f
C11421 VDD.n2717 GND 0.01303f
C11422 VDD.n2718 GND 0.95576f
C11423 VDD.n2719 GND 0.08471f
C11424 VDD.n2720 GND 0.01566f
C11425 VDD.n2721 GND 0.08328f
C11426 VDD.n2722 GND 0.04648f
C11427 VDD.n2723 GND 3.47277f
C11428 VDD.n2724 GND 0.04648f
C11429 VDD.n2725 GND 0.05737f
C11430 VDD.n2726 GND 0.0171f
C11431 VDD.n2727 GND 0.064f
C11432 VDD.n2730 GND 0.06555f
C11433 VDD.n2731 GND 0.03083f
C11434 VDD.t128 GND 0.08047f
C11435 VDD.n2732 GND 0.03534f
C11436 VDD.t932 GND 0.15471f
C11437 VDD.n2733 GND 0.03238f
C11438 VDD.n2734 GND 0.02607f
C11439 VDD.n2735 GND 0.09595f
C11440 VDD.t162 GND 0.08047f
C11441 VDD.n2736 GND 0.03534f
C11442 VDD.t971 GND 0.15471f
C11443 VDD.n2737 GND 0.03238f
C11444 VDD.n2738 GND 0.02607f
C11445 VDD.n2740 GND 0.24365f
C11446 VDD.n2741 GND 0.03496f
C11447 VDD.n2742 GND 1.22204f
C11448 VDD.n2743 GND 1.02074f
C11449 VDD.t959 GND 0.15539f
C11450 VDD.n2744 GND 0.06697f
C11451 VDD.t170 GND 0.07226f
C11452 VDD.n2745 GND 0.05627f
C11453 VDD.n2746 GND 0.05442f
C11454 VDD.n2747 GND 0.04255f
C11455 VDD.n2748 GND 0.05152f
C11456 VDD.t490 GND 0.02114f
C11457 VDD.t58 GND 0.02114f
C11458 VDD.n2749 GND 0.14059f
C11459 VDD.n2750 GND 0.04891f
C11460 VDD.n2751 GND 0.04648f
C11461 VDD.n2752 GND 0.04891f
C11462 VDD.n2753 GND 0.04532f
C11463 VDD.n2754 GND 0.04532f
C11464 VDD.t57 GND 4.12913f
C11465 VDD.n2755 GND 0.04648f
C11466 VDD.n2756 GND 0.04648f
C11467 VDD.n2757 GND 0.04648f
C11468 VDD.n2758 GND 0.04648f
C11469 VDD.n2759 GND 0.04648f
C11470 VDD.n2760 GND 0.04648f
C11471 VDD.n2761 GND 3.47277f
C11472 VDD.n2762 GND 0.04648f
C11473 VDD.n2763 GND 0.04648f
C11474 VDD.n2764 GND 0.04648f
C11475 VDD.n2765 GND 0.04648f
C11476 VDD.n2766 GND 0.04532f
C11477 VDD.n2767 GND 0.04532f
C11478 VDD.n2768 GND 0.02497f
C11479 VDD.n2769 GND 0.02497f
C11480 VDD.t61 GND 0.02104f
C11481 VDD.n2770 GND 0.22365f
C11482 VDD.t171 GND 0.02104f
C11483 VDD.t677 GND 0.02104f
C11484 VDD.n2771 GND 0.04891f
C11485 VDD.n2772 GND 0.04891f
C11486 VDD.n2773 GND 0.04532f
C11487 VDD.n2774 GND 0.04648f
C11488 VDD.n2775 GND 0.02293f
C11489 VDD.n2776 GND 0.02708f
C11490 VDD.n2777 GND 0.02293f
C11491 VDD.n2778 GND 0.04532f
C11492 VDD.n2779 GND 0.04532f
C11493 VDD.n2780 GND 0.04532f
C11494 VDD.n2781 GND 0.04532f
C11495 VDD.n2782 GND 0.04532f
C11496 VDD.n2783 GND 0.04532f
C11497 VDD.n2784 GND 0.04532f
C11498 VDD.n2785 GND 0.04532f
C11499 VDD.n2786 GND 0.04532f
C11500 VDD.n2787 GND 0.04532f
C11501 VDD.n2788 GND 0.04532f
C11502 VDD.n2789 GND 0.04532f
C11503 VDD.n2790 GND 0.04532f
C11504 VDD.n2791 GND 0.04532f
C11505 VDD.n2792 GND 0.04532f
C11506 VDD.n2793 GND 0.04532f
C11507 VDD.n2794 GND 0.04532f
C11508 VDD.n2795 GND 0.04532f
C11509 VDD.n2796 GND 0.04532f
C11510 VDD.n2797 GND 0.04532f
C11511 VDD.n2798 GND 0.02293f
C11512 VDD.n2799 GND 0.02293f
C11513 VDD.n2800 GND 0.02708f
C11514 VDD.n2801 GND 0.04648f
C11515 VDD.n2802 GND 3.19829f
C11516 VDD.n2803 GND 0.04532f
C11517 VDD.n2804 GND 0.04648f
C11518 VDD.n2805 GND 0.04648f
C11519 VDD.n2806 GND 0.04891f
C11520 VDD.n2807 GND 0.02293f
C11521 VDD.t588 GND 0.02114f
C11522 VDD.t706 GND 0.02114f
C11523 VDD.t11 GND 0.02114f
C11524 VDD.t587 GND 0.02114f
C11525 VDD.n2808 GND 0.02324f
C11526 VDD.n2809 GND 0.04891f
C11527 VDD.n2810 GND 0.04648f
C11528 VDD.n2811 GND 0.02293f
C11529 VDD.n2812 GND 0.04648f
C11530 VDD.n2813 GND 0.02708f
C11531 VDD.n2814 GND 0.02293f
C11532 VDD.n2815 GND 0.02708f
C11533 VDD.n2816 GND 0.02293f
C11534 VDD.n2817 GND 0.04532f
C11535 VDD.n2818 GND 0.04532f
C11536 VDD.n2819 GND 0.04532f
C11537 VDD.n2820 GND 0.02293f
C11538 VDD.n2821 GND 0.02293f
C11539 VDD.n2822 GND 0.02708f
C11540 VDD.n2823 GND 0.04648f
C11541 VDD.n2824 GND 0.04648f
C11542 VDD.n2825 GND 0.04648f
C11543 VDD.n2826 GND 0.04648f
C11544 VDD.n2827 GND 0.04532f
C11545 VDD.n2828 GND 0.04532f
C11546 VDD.n2829 GND 0.02293f
C11547 VDD.n2830 GND 0.02293f
C11548 VDD.n2831 GND 0.04648f
C11549 VDD.n2832 GND 0.02708f
C11550 VDD.n2833 GND 0.02293f
C11551 VDD.n2834 GND 0.04891f
C11552 VDD.n2835 GND 0.04648f
C11553 VDD.n2836 GND 0.05737f
C11554 VDD.n2837 GND 0.04891f
C11555 VDD.n2838 GND 0.02293f
C11556 VDD.n2839 GND 0.02708f
C11557 VDD.n2840 GND 0.04648f
C11558 VDD.n2841 GND 0.04532f
C11559 VDD.n2842 GND 0.04532f
C11560 VDD.n2843 GND 0.02293f
C11561 VDD.n2844 GND 0.02708f
C11562 VDD.n2845 GND 0.04648f
C11563 VDD.n2846 GND 0.04648f
C11564 VDD.n2847 GND 0.04648f
C11565 VDD.n2848 GND 0.04532f
C11566 VDD.n2849 GND 0.04532f
C11567 VDD.n2850 GND 0.02293f
C11568 VDD.n2851 GND 0.02293f
C11569 VDD.n2852 GND 0.04648f
C11570 VDD.n2853 GND 0.02708f
C11571 VDD.n2854 GND 0.02293f
C11572 VDD.n2855 GND 0.04891f
C11573 VDD.n2856 GND 0.04648f
C11574 VDD.t173 GND 0.02104f
C11575 VDD.t680 GND 0.02104f
C11576 VDD.t232 GND 0.02114f
C11577 VDD.t250 GND 0.02114f
C11578 VDD.n2857 GND 0.44561f
C11579 VDD.n2858 GND 0.04891f
C11580 VDD.n2859 GND 0.04648f
C11581 VDD.n2860 GND 0.02293f
C11582 VDD.n2861 GND 0.04648f
C11583 VDD.n2862 GND 0.02708f
C11584 VDD.n2863 GND 0.02293f
C11585 VDD.n2864 GND 0.04532f
C11586 VDD.n2865 GND 0.02293f
C11587 VDD.n2866 GND 0.02708f
C11588 VDD.n2867 GND 0.04532f
C11589 VDD.n2868 GND 0.02293f
C11590 VDD.n2869 GND 0.04891f
C11591 VDD.n2870 GND 0.05737f
C11592 VDD.n2871 GND 0.02055f
C11593 VDD.n2872 GND 0.08471f
C11594 VDD.n2873 GND 0.95576f
C11595 VDD.t279 GND 0.02114f
C11596 VDD.t512 GND 0.02114f
C11597 VDD.t337 GND 0.02114f
C11598 VDD.t852 GND 0.02114f
C11599 VDD.t255 GND 0.02104f
C11600 VDD.t851 GND 0.02114f
C11601 VDD.t374 GND 0.02114f
C11602 VDD.t622 GND 0.02114f
C11603 VDD.t621 GND 0.02114f
C11604 VDD.t143 GND 0.02104f
C11605 VDD.t673 GND 0.02104f
C11606 VDD.n2874 GND 0.95576f
C11607 VDD.n2875 GND 0.08471f
C11608 VDD.n2876 GND 0.04891f
C11609 VDD.n2877 GND 0.04648f
C11610 VDD.n2878 GND 0.02293f
C11611 VDD.n2879 GND 0.04648f
C11612 VDD.n2880 GND 0.02708f
C11613 VDD.n2881 GND 0.02293f
C11614 VDD.n2882 GND 0.04532f
C11615 VDD.n2883 GND 0.02293f
C11616 VDD.n2884 GND 0.02708f
C11617 VDD.n2885 GND 0.04532f
C11618 VDD.n2886 GND 0.02293f
C11619 VDD.n2887 GND 0.04891f
C11620 VDD.n2888 GND 0.05737f
C11621 VDD.n2889 GND 0.02055f
C11622 VDD.n2890 GND 0.44561f
C11623 VDD.n2891 GND 0.14059f
C11624 VDD.n2892 GND 0.04891f
C11625 VDD.n2893 GND 0.04648f
C11626 VDD.n2894 GND 0.02293f
C11627 VDD.n2895 GND 0.04648f
C11628 VDD.n2896 GND 0.02708f
C11629 VDD.n2897 GND 0.02293f
C11630 VDD.n2898 GND 0.04532f
C11631 VDD.n2899 GND 0.02293f
C11632 VDD.n2900 GND 0.02708f
C11633 VDD.n2901 GND 0.04532f
C11634 VDD.n2902 GND 0.02293f
C11635 VDD.n2903 GND 0.04891f
C11636 VDD.n2904 GND 0.05737f
C11637 VDD.n2905 GND 0.02055f
C11638 VDD.n2906 GND 0.02497f
C11639 VDD.n2907 GND 0.04648f
C11640 VDD.n2908 GND 0.04648f
C11641 VDD.n2909 GND 0.02708f
C11642 VDD.n2910 GND 0.02497f
C11643 VDD.n2911 GND 0.08328f
C11644 VDD.n2912 GND 0.01566f
C11645 VDD.n2913 GND 0.18236f
C11646 VDD.n2914 GND 0.03549f
C11647 VDD.n2915 GND 0.04891f
C11648 VDD.n2916 GND 0.04648f
C11649 VDD.n2917 GND 0.02293f
C11650 VDD.n2918 GND 0.04648f
C11651 VDD.n2919 GND 0.02708f
C11652 VDD.n2920 GND 0.02293f
C11653 VDD.n2921 GND 0.04532f
C11654 VDD.n2922 GND 0.02293f
C11655 VDD.n2923 GND 0.02708f
C11656 VDD.n2924 GND 0.04532f
C11657 VDD.n2925 GND 0.02293f
C11658 VDD.n2926 GND 0.04891f
C11659 VDD.n2927 GND 0.05737f
C11660 VDD.n2928 GND 0.02055f
C11661 VDD.n2929 GND 0.44561f
C11662 VDD.n2930 GND 0.14059f
C11663 VDD.n2931 GND 0.04891f
C11664 VDD.n2932 GND 0.04648f
C11665 VDD.n2933 GND 0.02293f
C11666 VDD.n2934 GND 0.04648f
C11667 VDD.n2935 GND 0.02708f
C11668 VDD.n2936 GND 0.02293f
C11669 VDD.n2937 GND 0.04532f
C11670 VDD.n2938 GND 0.02293f
C11671 VDD.n2939 GND 0.02708f
C11672 VDD.n2940 GND 0.04532f
C11673 VDD.n2941 GND 0.02293f
C11674 VDD.n2942 GND 0.04891f
C11675 VDD.n2943 GND 0.05737f
C11676 VDD.n2944 GND 0.02813f
C11677 VDD.n2945 GND 0.02324f
C11678 VDD.n2946 GND 0.05737f
C11679 VDD.n2947 GND 0.04891f
C11680 VDD.n2948 GND 0.02293f
C11681 VDD.n2949 GND 0.02708f
C11682 VDD.n2950 GND 0.04648f
C11683 VDD.n2951 GND 0.02293f
C11684 VDD.n2952 GND 0.02293f
C11685 VDD.n2953 GND 0.02708f
C11686 VDD.n2954 GND 0.04648f
C11687 VDD.n2955 GND 0.02708f
C11688 VDD.n2956 GND 0.04648f
C11689 VDD.n2957 GND 3.19829f
C11690 VDD.n2958 GND 0.04648f
C11691 VDD.n2959 GND 0.04532f
C11692 VDD.n2960 GND 0.02293f
C11693 VDD.n2961 GND 0.04891f
C11694 VDD.n2962 GND 0.05737f
C11695 VDD.n2963 GND 0.02813f
C11696 VDD.n2964 GND 0.14059f
C11697 VDD.n2965 GND 0.44561f
C11698 VDD.n2966 GND 0.02055f
C11699 VDD.n2967 GND 0.05737f
C11700 VDD.n2968 GND 0.04891f
C11701 VDD.n2969 GND 0.02293f
C11702 VDD.n2970 GND 0.02708f
C11703 VDD.n2971 GND 0.02293f
C11704 VDD.n2972 GND 0.04532f
C11705 VDD.t10 GND 4.12913f
C11706 VDD.n2973 GND 0.04532f
C11707 VDD.n2974 GND 0.04648f
C11708 VDD.n2975 GND 0.05737f
C11709 VDD.n2976 GND 0.01303f
C11710 VDD.n2977 GND 0.95576f
C11711 VDD.n2978 GND 0.08471f
C11712 VDD.n2979 GND 0.01566f
C11713 VDD.n2980 GND 0.08328f
C11714 VDD.n2981 GND 0.04648f
C11715 VDD.n2982 GND 3.47277f
C11716 VDD.n2983 GND 0.04648f
C11717 VDD.n2984 GND 0.05737f
C11718 VDD.n2985 GND 0.0171f
C11719 VDD.n2986 GND 0.064f
C11720 VDD.n2989 GND 0.06555f
C11721 VDD.n2990 GND 0.03083f
C11722 VDD.t142 GND 0.08047f
C11723 VDD.n2991 GND 0.03534f
C11724 VDD.t927 GND 0.15471f
C11725 VDD.n2992 GND 0.03238f
C11726 VDD.n2993 GND 0.02607f
C11727 VDD.n2994 GND 0.09595f
C11728 VDD.t172 GND 0.08047f
C11729 VDD.n2995 GND 0.03534f
C11730 VDD.t968 GND 0.15471f
C11731 VDD.n2996 GND 0.03238f
C11732 VDD.n2997 GND 0.02607f
C11733 VDD.n2999 GND 0.24365f
C11734 VDD.n3000 GND 0.03496f
C11735 VDD.n3001 GND 1.06185f
C11736 VDD.n3002 GND 0.87512f
C11737 VDD.t974 GND 0.15539f
C11738 VDD.n3003 GND 0.06697f
C11739 VDD.t205 GND 0.07226f
C11740 VDD.n3004 GND 0.05627f
C11741 VDD.n3005 GND 0.05442f
C11742 VDD.n3006 GND 0.04255f
C11743 VDD.n3007 GND 0.05152f
C11744 VDD.t56 GND 0.02114f
C11745 VDD.t589 GND 0.02114f
C11746 VDD.n3008 GND 0.14059f
C11747 VDD.n3009 GND 0.04891f
C11748 VDD.n3010 GND 0.04648f
C11749 VDD.n3011 GND 0.04891f
C11750 VDD.n3012 GND 0.04532f
C11751 VDD.n3013 GND 0.04532f
C11752 VDD.t48 GND 4.12913f
C11753 VDD.n3014 GND 0.04648f
C11754 VDD.n3015 GND 0.04648f
C11755 VDD.n3016 GND 0.04648f
C11756 VDD.n3017 GND 0.04648f
C11757 VDD.n3018 GND 0.04648f
C11758 VDD.n3019 GND 0.04648f
C11759 VDD.n3020 GND 3.47277f
C11760 VDD.n3021 GND 0.04648f
C11761 VDD.n3022 GND 0.04648f
C11762 VDD.n3023 GND 0.04648f
C11763 VDD.n3024 GND 0.04648f
C11764 VDD.n3025 GND 0.04532f
C11765 VDD.n3026 GND 0.04532f
C11766 VDD.n3027 GND 0.02497f
C11767 VDD.n3028 GND 0.02497f
C11768 VDD.t492 GND 0.02104f
C11769 VDD.n3029 GND 0.22365f
C11770 VDD.t206 GND 0.02104f
C11771 VDD.t681 GND 0.02104f
C11772 VDD.n3030 GND 0.04891f
C11773 VDD.n3031 GND 0.04891f
C11774 VDD.n3032 GND 0.04532f
C11775 VDD.n3033 GND 0.04648f
C11776 VDD.n3034 GND 0.02293f
C11777 VDD.n3035 GND 0.02708f
C11778 VDD.n3036 GND 0.02293f
C11779 VDD.n3037 GND 0.04532f
C11780 VDD.n3038 GND 0.04532f
C11781 VDD.n3039 GND 0.04532f
C11782 VDD.n3040 GND 0.04532f
C11783 VDD.n3041 GND 0.04532f
C11784 VDD.n3042 GND 0.04532f
C11785 VDD.n3043 GND 0.04532f
C11786 VDD.n3044 GND 0.04532f
C11787 VDD.n3045 GND 0.04532f
C11788 VDD.n3046 GND 0.04532f
C11789 VDD.n3047 GND 0.04532f
C11790 VDD.n3048 GND 0.04532f
C11791 VDD.n3049 GND 0.04532f
C11792 VDD.n3050 GND 0.04532f
C11793 VDD.n3051 GND 0.04532f
C11794 VDD.n3052 GND 0.04532f
C11795 VDD.n3053 GND 0.04532f
C11796 VDD.n3054 GND 0.04532f
C11797 VDD.n3055 GND 0.04532f
C11798 VDD.n3056 GND 0.04532f
C11799 VDD.n3057 GND 0.02293f
C11800 VDD.n3058 GND 0.02293f
C11801 VDD.n3059 GND 0.02708f
C11802 VDD.n3060 GND 0.04648f
C11803 VDD.n3061 GND 3.19829f
C11804 VDD.n3062 GND 0.04532f
C11805 VDD.n3063 GND 0.04648f
C11806 VDD.n3064 GND 0.04648f
C11807 VDD.n3065 GND 0.04891f
C11808 VDD.n3066 GND 0.02293f
C11809 VDD.t406 GND 0.02114f
C11810 VDD.t305 GND 0.02114f
C11811 VDD.t519 GND 0.02114f
C11812 VDD.t49 GND 0.02114f
C11813 VDD.n3067 GND 0.02324f
C11814 VDD.n3068 GND 0.04891f
C11815 VDD.n3069 GND 0.04648f
C11816 VDD.n3070 GND 0.02293f
C11817 VDD.n3071 GND 0.04648f
C11818 VDD.n3072 GND 0.02708f
C11819 VDD.n3073 GND 0.02293f
C11820 VDD.n3074 GND 0.02708f
C11821 VDD.n3075 GND 0.02293f
C11822 VDD.n3076 GND 0.04532f
C11823 VDD.n3077 GND 0.04532f
C11824 VDD.n3078 GND 0.04532f
C11825 VDD.n3079 GND 0.02293f
C11826 VDD.n3080 GND 0.02293f
C11827 VDD.n3081 GND 0.02708f
C11828 VDD.n3082 GND 0.04648f
C11829 VDD.n3083 GND 0.04648f
C11830 VDD.n3084 GND 0.04648f
C11831 VDD.n3085 GND 0.04648f
C11832 VDD.n3086 GND 0.04532f
C11833 VDD.n3087 GND 0.04532f
C11834 VDD.n3088 GND 0.02293f
C11835 VDD.n3089 GND 0.02293f
C11836 VDD.n3090 GND 0.04648f
C11837 VDD.n3091 GND 0.02708f
C11838 VDD.n3092 GND 0.02293f
C11839 VDD.n3093 GND 0.04891f
C11840 VDD.n3094 GND 0.04648f
C11841 VDD.n3095 GND 0.05737f
C11842 VDD.n3096 GND 0.04891f
C11843 VDD.n3097 GND 0.02293f
C11844 VDD.n3098 GND 0.02708f
C11845 VDD.n3099 GND 0.04648f
C11846 VDD.n3100 GND 0.04532f
C11847 VDD.n3101 GND 0.04532f
C11848 VDD.n3102 GND 0.02293f
C11849 VDD.n3103 GND 0.02708f
C11850 VDD.n3104 GND 0.04648f
C11851 VDD.n3105 GND 0.04648f
C11852 VDD.n3106 GND 0.04648f
C11853 VDD.n3107 GND 0.04532f
C11854 VDD.n3108 GND 0.04532f
C11855 VDD.n3109 GND 0.02293f
C11856 VDD.n3110 GND 0.02293f
C11857 VDD.n3111 GND 0.04648f
C11858 VDD.n3112 GND 0.02708f
C11859 VDD.n3113 GND 0.02293f
C11860 VDD.n3114 GND 0.04891f
C11861 VDD.n3115 GND 0.04648f
C11862 VDD.t180 GND 0.02104f
C11863 VDD.t648 GND 0.02104f
C11864 VDD.t743 GND 0.02114f
C11865 VDD.t821 GND 0.02114f
C11866 VDD.n3116 GND 0.44561f
C11867 VDD.n3117 GND 0.04891f
C11868 VDD.n3118 GND 0.04648f
C11869 VDD.n3119 GND 0.02293f
C11870 VDD.n3120 GND 0.04648f
C11871 VDD.n3121 GND 0.02708f
C11872 VDD.n3122 GND 0.02293f
C11873 VDD.n3123 GND 0.04532f
C11874 VDD.n3124 GND 0.02293f
C11875 VDD.n3125 GND 0.02708f
C11876 VDD.n3126 GND 0.04532f
C11877 VDD.n3127 GND 0.02293f
C11878 VDD.n3128 GND 0.04891f
C11879 VDD.n3129 GND 0.05737f
C11880 VDD.n3130 GND 0.02055f
C11881 VDD.n3131 GND 0.08471f
C11882 VDD.n3132 GND 0.95576f
C11883 VDD.t373 GND 0.02114f
C11884 VDD.t872 GND 0.02114f
C11885 VDD.t624 GND 0.02114f
C11886 VDD.t780 GND 0.02114f
C11887 VDD.t831 GND 0.02104f
C11888 VDD.t781 GND 0.02114f
C11889 VDD.t623 GND 0.02114f
C11890 VDD.t908 GND 0.02114f
C11891 VDD.t734 GND 0.02114f
C11892 VDD.t169 GND 0.02104f
C11893 VDD.t693 GND 0.02104f
C11894 VDD.n3133 GND 0.95576f
C11895 VDD.n3134 GND 0.08471f
C11896 VDD.n3135 GND 0.04891f
C11897 VDD.n3136 GND 0.04648f
C11898 VDD.n3137 GND 0.02293f
C11899 VDD.n3138 GND 0.04648f
C11900 VDD.n3139 GND 0.02708f
C11901 VDD.n3140 GND 0.02293f
C11902 VDD.n3141 GND 0.04532f
C11903 VDD.n3142 GND 0.02293f
C11904 VDD.n3143 GND 0.02708f
C11905 VDD.n3144 GND 0.04532f
C11906 VDD.n3145 GND 0.02293f
C11907 VDD.n3146 GND 0.04891f
C11908 VDD.n3147 GND 0.05737f
C11909 VDD.n3148 GND 0.02055f
C11910 VDD.n3149 GND 0.44561f
C11911 VDD.n3150 GND 0.14059f
C11912 VDD.n3151 GND 0.04891f
C11913 VDD.n3152 GND 0.04648f
C11914 VDD.n3153 GND 0.02293f
C11915 VDD.n3154 GND 0.04648f
C11916 VDD.n3155 GND 0.02708f
C11917 VDD.n3156 GND 0.02293f
C11918 VDD.n3157 GND 0.04532f
C11919 VDD.n3158 GND 0.02293f
C11920 VDD.n3159 GND 0.02708f
C11921 VDD.n3160 GND 0.04532f
C11922 VDD.n3161 GND 0.02293f
C11923 VDD.n3162 GND 0.04891f
C11924 VDD.n3163 GND 0.05737f
C11925 VDD.n3164 GND 0.02055f
C11926 VDD.n3165 GND 0.02497f
C11927 VDD.n3166 GND 0.04648f
C11928 VDD.n3167 GND 0.04648f
C11929 VDD.n3168 GND 0.02708f
C11930 VDD.n3169 GND 0.02497f
C11931 VDD.n3170 GND 0.08328f
C11932 VDD.n3171 GND 0.01566f
C11933 VDD.n3172 GND 0.18236f
C11934 VDD.n3173 GND 0.03549f
C11935 VDD.n3174 GND 0.04891f
C11936 VDD.n3175 GND 0.04648f
C11937 VDD.n3176 GND 0.02293f
C11938 VDD.n3177 GND 0.04648f
C11939 VDD.n3178 GND 0.02708f
C11940 VDD.n3179 GND 0.02293f
C11941 VDD.n3180 GND 0.04532f
C11942 VDD.n3181 GND 0.02293f
C11943 VDD.n3182 GND 0.02708f
C11944 VDD.n3183 GND 0.04532f
C11945 VDD.n3184 GND 0.02293f
C11946 VDD.n3185 GND 0.04891f
C11947 VDD.n3186 GND 0.05737f
C11948 VDD.n3187 GND 0.02055f
C11949 VDD.n3188 GND 0.44561f
C11950 VDD.n3189 GND 0.14059f
C11951 VDD.n3190 GND 0.04891f
C11952 VDD.n3191 GND 0.04648f
C11953 VDD.n3192 GND 0.02293f
C11954 VDD.n3193 GND 0.04648f
C11955 VDD.n3194 GND 0.02708f
C11956 VDD.n3195 GND 0.02293f
C11957 VDD.n3196 GND 0.04532f
C11958 VDD.n3197 GND 0.02293f
C11959 VDD.n3198 GND 0.02708f
C11960 VDD.n3199 GND 0.04532f
C11961 VDD.n3200 GND 0.02293f
C11962 VDD.n3201 GND 0.04891f
C11963 VDD.n3202 GND 0.05737f
C11964 VDD.n3203 GND 0.02813f
C11965 VDD.n3204 GND 0.02324f
C11966 VDD.n3205 GND 0.05737f
C11967 VDD.n3206 GND 0.04891f
C11968 VDD.n3207 GND 0.02293f
C11969 VDD.n3208 GND 0.02708f
C11970 VDD.n3209 GND 0.04648f
C11971 VDD.n3210 GND 0.02293f
C11972 VDD.n3211 GND 0.02293f
C11973 VDD.n3212 GND 0.02708f
C11974 VDD.n3213 GND 0.04648f
C11975 VDD.n3214 GND 0.02708f
C11976 VDD.n3215 GND 0.04648f
C11977 VDD.n3216 GND 3.19829f
C11978 VDD.n3217 GND 0.04648f
C11979 VDD.n3218 GND 0.04532f
C11980 VDD.n3219 GND 0.02293f
C11981 VDD.n3220 GND 0.04891f
C11982 VDD.n3221 GND 0.05737f
C11983 VDD.n3222 GND 0.02813f
C11984 VDD.n3223 GND 0.14059f
C11985 VDD.n3224 GND 0.44561f
C11986 VDD.n3225 GND 0.02055f
C11987 VDD.n3226 GND 0.05737f
C11988 VDD.n3227 GND 0.04891f
C11989 VDD.n3228 GND 0.02293f
C11990 VDD.n3229 GND 0.02708f
C11991 VDD.n3230 GND 0.02293f
C11992 VDD.n3231 GND 0.04532f
C11993 VDD.t55 GND 4.12913f
C11994 VDD.n3232 GND 0.04532f
C11995 VDD.n3233 GND 0.04648f
C11996 VDD.n3234 GND 0.05737f
C11997 VDD.n3235 GND 0.01303f
C11998 VDD.n3236 GND 0.95576f
C11999 VDD.n3237 GND 0.08471f
C12000 VDD.n3238 GND 0.01566f
C12001 VDD.n3239 GND 0.08328f
C12002 VDD.n3240 GND 0.04648f
C12003 VDD.n3241 GND 3.47277f
C12004 VDD.n3242 GND 0.04648f
C12005 VDD.n3243 GND 0.05737f
C12006 VDD.n3244 GND 0.0171f
C12007 VDD.n3245 GND 0.064f
C12008 VDD.n3248 GND 0.06555f
C12009 VDD.n3249 GND 0.03083f
C12010 VDD.t168 GND 0.08047f
C12011 VDD.n3250 GND 0.03534f
C12012 VDD.t934 GND 0.15471f
C12013 VDD.n3251 GND 0.03238f
C12014 VDD.n3252 GND 0.02607f
C12015 VDD.n3253 GND 0.09595f
C12016 VDD.t179 GND 0.08047f
C12017 VDD.n3254 GND 0.03534f
C12018 VDD.t972 GND 0.15471f
C12019 VDD.n3255 GND 0.03238f
C12020 VDD.n3256 GND 0.02607f
C12021 VDD.n3258 GND 0.24365f
C12022 VDD.n3259 GND 0.03496f
C12023 VDD.n3260 GND 0.90166f
C12024 VDD.n3261 GND 0.72949f
C12025 VDD.t969 GND 0.15539f
C12026 VDD.n3262 GND 0.06697f
C12027 VDD.t134 GND 0.07226f
C12028 VDD.n3263 GND 0.05627f
C12029 VDD.n3264 GND 0.05442f
C12030 VDD.n3265 GND 0.04255f
C12031 VDD.n3266 GND 0.05152f
C12032 VDD.t874 GND 0.02114f
C12033 VDD.t405 GND 0.02114f
C12034 VDD.n3267 GND 0.14059f
C12035 VDD.n3268 GND 0.04891f
C12036 VDD.n3269 GND 0.04648f
C12037 VDD.n3270 GND 0.04891f
C12038 VDD.n3271 GND 0.04532f
C12039 VDD.n3272 GND 0.04532f
C12040 VDD.t135 GND 4.12913f
C12041 VDD.n3273 GND 0.04648f
C12042 VDD.n3274 GND 0.04648f
C12043 VDD.n3275 GND 0.04648f
C12044 VDD.n3276 GND 0.04648f
C12045 VDD.n3277 GND 0.04648f
C12046 VDD.n3278 GND 0.04648f
C12047 VDD.n3279 GND 3.47277f
C12048 VDD.n3280 GND 0.04648f
C12049 VDD.n3281 GND 0.04648f
C12050 VDD.n3282 GND 0.04648f
C12051 VDD.n3283 GND 0.04648f
C12052 VDD.n3284 GND 0.04532f
C12053 VDD.n3285 GND 0.04532f
C12054 VDD.n3286 GND 0.02497f
C12055 VDD.n3287 GND 0.02497f
C12056 VDD.t802 GND 0.02104f
C12057 VDD.n3288 GND 0.22365f
C12058 VDD.t136 GND 0.02104f
C12059 VDD.t660 GND 0.02104f
C12060 VDD.n3289 GND 0.04891f
C12061 VDD.n3290 GND 0.04891f
C12062 VDD.n3291 GND 0.04532f
C12063 VDD.n3292 GND 0.04648f
C12064 VDD.n3293 GND 0.02293f
C12065 VDD.n3294 GND 0.02708f
C12066 VDD.n3295 GND 0.02293f
C12067 VDD.n3296 GND 0.04532f
C12068 VDD.n3297 GND 0.04532f
C12069 VDD.n3298 GND 0.04532f
C12070 VDD.n3299 GND 0.04532f
C12071 VDD.n3300 GND 0.04532f
C12072 VDD.n3301 GND 0.04532f
C12073 VDD.n3302 GND 0.04532f
C12074 VDD.n3303 GND 0.04532f
C12075 VDD.n3304 GND 0.04532f
C12076 VDD.n3305 GND 0.04532f
C12077 VDD.n3306 GND 0.04532f
C12078 VDD.n3307 GND 0.04532f
C12079 VDD.n3308 GND 0.04532f
C12080 VDD.n3309 GND 0.04532f
C12081 VDD.n3310 GND 0.04532f
C12082 VDD.n3311 GND 0.04532f
C12083 VDD.n3312 GND 0.04532f
C12084 VDD.n3313 GND 0.04532f
C12085 VDD.n3314 GND 0.04532f
C12086 VDD.n3315 GND 0.04532f
C12087 VDD.n3316 GND 0.02293f
C12088 VDD.n3317 GND 0.02293f
C12089 VDD.n3318 GND 0.02708f
C12090 VDD.n3319 GND 0.04648f
C12091 VDD.n3320 GND 3.19829f
C12092 VDD.n3321 GND 0.04532f
C12093 VDD.n3322 GND 0.04648f
C12094 VDD.n3323 GND 0.04648f
C12095 VDD.n3324 GND 0.04891f
C12096 VDD.n3325 GND 0.02293f
C12097 VDD.t93 GND 0.02114f
C12098 VDD.t500 GND 0.02114f
C12099 VDD.t632 GND 0.02114f
C12100 VDD.t267 GND 0.02114f
C12101 VDD.n3326 GND 0.02324f
C12102 VDD.n3327 GND 0.04891f
C12103 VDD.n3328 GND 0.04648f
C12104 VDD.n3329 GND 0.02293f
C12105 VDD.n3330 GND 0.04648f
C12106 VDD.n3331 GND 0.02708f
C12107 VDD.n3332 GND 0.02293f
C12108 VDD.n3333 GND 0.02708f
C12109 VDD.n3334 GND 0.02293f
C12110 VDD.n3335 GND 0.04532f
C12111 VDD.n3336 GND 0.04532f
C12112 VDD.n3337 GND 0.04532f
C12113 VDD.n3338 GND 0.02293f
C12114 VDD.n3339 GND 0.02293f
C12115 VDD.n3340 GND 0.02708f
C12116 VDD.n3341 GND 0.04648f
C12117 VDD.n3342 GND 0.04648f
C12118 VDD.n3343 GND 0.04648f
C12119 VDD.n3344 GND 0.04648f
C12120 VDD.n3345 GND 0.04532f
C12121 VDD.n3346 GND 0.04532f
C12122 VDD.n3347 GND 0.02293f
C12123 VDD.n3348 GND 0.02293f
C12124 VDD.n3349 GND 0.04648f
C12125 VDD.n3350 GND 0.02708f
C12126 VDD.n3351 GND 0.02293f
C12127 VDD.n3352 GND 0.04891f
C12128 VDD.n3353 GND 0.04648f
C12129 VDD.n3354 GND 0.05737f
C12130 VDD.n3355 GND 0.04891f
C12131 VDD.n3356 GND 0.02293f
C12132 VDD.n3357 GND 0.02708f
C12133 VDD.n3358 GND 0.04648f
C12134 VDD.n3359 GND 0.04532f
C12135 VDD.n3360 GND 0.04532f
C12136 VDD.n3361 GND 0.02293f
C12137 VDD.n3362 GND 0.02708f
C12138 VDD.n3363 GND 0.04648f
C12139 VDD.n3364 GND 0.04648f
C12140 VDD.n3365 GND 0.04648f
C12141 VDD.n3366 GND 0.04532f
C12142 VDD.n3367 GND 0.04532f
C12143 VDD.n3368 GND 0.02293f
C12144 VDD.n3369 GND 0.02293f
C12145 VDD.n3370 GND 0.04648f
C12146 VDD.n3371 GND 0.02708f
C12147 VDD.n3372 GND 0.02293f
C12148 VDD.n3373 GND 0.04891f
C12149 VDD.n3374 GND 0.04648f
C12150 VDD.t138 GND 0.02104f
C12151 VDD.t670 GND 0.02104f
C12152 VDD.t227 GND 0.02114f
C12153 VDD.t245 GND 0.02114f
C12154 VDD.n3375 GND 0.44561f
C12155 VDD.n3376 GND 0.04891f
C12156 VDD.n3377 GND 0.04648f
C12157 VDD.n3378 GND 0.02293f
C12158 VDD.n3379 GND 0.04648f
C12159 VDD.n3380 GND 0.02708f
C12160 VDD.n3381 GND 0.02293f
C12161 VDD.n3382 GND 0.04532f
C12162 VDD.n3383 GND 0.02293f
C12163 VDD.n3384 GND 0.02708f
C12164 VDD.n3385 GND 0.04532f
C12165 VDD.n3386 GND 0.02293f
C12166 VDD.n3387 GND 0.04891f
C12167 VDD.n3388 GND 0.05737f
C12168 VDD.n3389 GND 0.02055f
C12169 VDD.n3390 GND 0.08471f
C12170 VDD.n3391 GND 0.95576f
C12171 VDD.t850 GND 0.02114f
C12172 VDD.t608 GND 0.02114f
C12173 VDD.t463 GND 0.02114f
C12174 VDD.t861 GND 0.02114f
C12175 VDD.t237 GND 0.02104f
C12176 VDD.t860 GND 0.02114f
C12177 VDD.t464 GND 0.02114f
C12178 VDD.t521 GND 0.02114f
C12179 VDD.t520 GND 0.02114f
C12180 VDD.t104 GND 0.02104f
C12181 VDD.t655 GND 0.02104f
C12182 VDD.n3392 GND 0.95576f
C12183 VDD.n3393 GND 0.08471f
C12184 VDD.n3394 GND 0.04891f
C12185 VDD.n3395 GND 0.04648f
C12186 VDD.n3396 GND 0.02293f
C12187 VDD.n3397 GND 0.04648f
C12188 VDD.n3398 GND 0.02708f
C12189 VDD.n3399 GND 0.02293f
C12190 VDD.n3400 GND 0.04532f
C12191 VDD.n3401 GND 0.02293f
C12192 VDD.n3402 GND 0.02708f
C12193 VDD.n3403 GND 0.04532f
C12194 VDD.n3404 GND 0.02293f
C12195 VDD.n3405 GND 0.04891f
C12196 VDD.n3406 GND 0.05737f
C12197 VDD.n3407 GND 0.02055f
C12198 VDD.n3408 GND 0.44561f
C12199 VDD.n3409 GND 0.14059f
C12200 VDD.n3410 GND 0.04891f
C12201 VDD.n3411 GND 0.04648f
C12202 VDD.n3412 GND 0.02293f
C12203 VDD.n3413 GND 0.04648f
C12204 VDD.n3414 GND 0.02708f
C12205 VDD.n3415 GND 0.02293f
C12206 VDD.n3416 GND 0.04532f
C12207 VDD.n3417 GND 0.02293f
C12208 VDD.n3418 GND 0.02708f
C12209 VDD.n3419 GND 0.04532f
C12210 VDD.n3420 GND 0.02293f
C12211 VDD.n3421 GND 0.04891f
C12212 VDD.n3422 GND 0.05737f
C12213 VDD.n3423 GND 0.02055f
C12214 VDD.n3424 GND 0.02497f
C12215 VDD.n3425 GND 0.04648f
C12216 VDD.n3426 GND 0.04648f
C12217 VDD.n3427 GND 0.02708f
C12218 VDD.n3428 GND 0.02497f
C12219 VDD.n3429 GND 0.08328f
C12220 VDD.n3430 GND 0.01566f
C12221 VDD.n3431 GND 0.18236f
C12222 VDD.n3432 GND 0.03549f
C12223 VDD.n3433 GND 0.04891f
C12224 VDD.n3434 GND 0.04648f
C12225 VDD.n3435 GND 0.02293f
C12226 VDD.n3436 GND 0.04648f
C12227 VDD.n3437 GND 0.02708f
C12228 VDD.n3438 GND 0.02293f
C12229 VDD.n3439 GND 0.04532f
C12230 VDD.n3440 GND 0.02293f
C12231 VDD.n3441 GND 0.02708f
C12232 VDD.n3442 GND 0.04532f
C12233 VDD.n3443 GND 0.02293f
C12234 VDD.n3444 GND 0.04891f
C12235 VDD.n3445 GND 0.05737f
C12236 VDD.n3446 GND 0.02055f
C12237 VDD.n3447 GND 0.44561f
C12238 VDD.n3448 GND 0.14059f
C12239 VDD.n3449 GND 0.04891f
C12240 VDD.n3450 GND 0.04648f
C12241 VDD.n3451 GND 0.02293f
C12242 VDD.n3452 GND 0.04648f
C12243 VDD.n3453 GND 0.02708f
C12244 VDD.n3454 GND 0.02293f
C12245 VDD.n3455 GND 0.04532f
C12246 VDD.n3456 GND 0.02293f
C12247 VDD.n3457 GND 0.02708f
C12248 VDD.n3458 GND 0.04532f
C12249 VDD.n3459 GND 0.02293f
C12250 VDD.n3460 GND 0.04891f
C12251 VDD.n3461 GND 0.05737f
C12252 VDD.n3462 GND 0.02813f
C12253 VDD.n3463 GND 0.02324f
C12254 VDD.n3464 GND 0.05737f
C12255 VDD.n3465 GND 0.04891f
C12256 VDD.n3466 GND 0.02293f
C12257 VDD.n3467 GND 0.02708f
C12258 VDD.n3468 GND 0.04648f
C12259 VDD.n3469 GND 0.02293f
C12260 VDD.n3470 GND 0.02293f
C12261 VDD.n3471 GND 0.02708f
C12262 VDD.n3472 GND 0.04648f
C12263 VDD.n3473 GND 0.02708f
C12264 VDD.n3474 GND 0.04648f
C12265 VDD.n3475 GND 3.19829f
C12266 VDD.n3476 GND 0.04648f
C12267 VDD.n3477 GND 0.04532f
C12268 VDD.n3478 GND 0.02293f
C12269 VDD.n3479 GND 0.04891f
C12270 VDD.n3480 GND 0.05737f
C12271 VDD.n3481 GND 0.02813f
C12272 VDD.n3482 GND 0.14059f
C12273 VDD.n3483 GND 0.44561f
C12274 VDD.n3484 GND 0.02055f
C12275 VDD.n3485 GND 0.05737f
C12276 VDD.n3486 GND 0.04891f
C12277 VDD.n3487 GND 0.02293f
C12278 VDD.n3488 GND 0.02708f
C12279 VDD.n3489 GND 0.02293f
C12280 VDD.n3490 GND 0.04532f
C12281 VDD.t92 GND 4.12913f
C12282 VDD.n3491 GND 0.04532f
C12283 VDD.n3492 GND 0.04648f
C12284 VDD.n3493 GND 0.05737f
C12285 VDD.n3494 GND 0.01303f
C12286 VDD.n3495 GND 0.95576f
C12287 VDD.n3496 GND 0.08471f
C12288 VDD.n3497 GND 0.01566f
C12289 VDD.n3498 GND 0.08328f
C12290 VDD.n3499 GND 0.04648f
C12291 VDD.n3500 GND 3.47277f
C12292 VDD.n3501 GND 0.04648f
C12293 VDD.n3502 GND 0.05737f
C12294 VDD.n3503 GND 0.0171f
C12295 VDD.n3504 GND 0.064f
C12296 VDD.n3507 GND 0.06555f
C12297 VDD.n3508 GND 0.03083f
C12298 VDD.t103 GND 0.08047f
C12299 VDD.n3509 GND 0.03534f
C12300 VDD.t942 GND 0.15471f
C12301 VDD.n3510 GND 0.03238f
C12302 VDD.n3511 GND 0.02607f
C12303 VDD.n3512 GND 0.09595f
C12304 VDD.t137 GND 0.08047f
C12305 VDD.n3513 GND 0.03534f
C12306 VDD.t928 GND 0.15471f
C12307 VDD.n3514 GND 0.03238f
C12308 VDD.n3515 GND 0.02607f
C12309 VDD.n3517 GND 0.24365f
C12310 VDD.n3518 GND 0.03496f
C12311 VDD.n3519 GND 0.74147f
C12312 VDD.n3520 GND 0.58386f
C12313 VDD.t965 GND 0.15539f
C12314 VDD.n3521 GND 0.06697f
C12315 VDD.t151 GND 0.07226f
C12316 VDD.n3522 GND 0.05627f
C12317 VDD.n3523 GND 0.05442f
C12318 VDD.n3524 GND 0.04255f
C12319 VDD.n3525 GND 0.05152f
C12320 VDD.t801 GND 0.02114f
C12321 VDD.t480 GND 0.02114f
C12322 VDD.n3526 GND 0.14059f
C12323 VDD.n3527 GND 0.04891f
C12324 VDD.n3528 GND 0.04648f
C12325 VDD.n3529 GND 0.04891f
C12326 VDD.n3530 GND 0.04532f
C12327 VDD.n3531 GND 0.04532f
C12328 VDD.t24 GND 4.12913f
C12329 VDD.n3532 GND 0.04648f
C12330 VDD.n3533 GND 0.04648f
C12331 VDD.n3534 GND 0.04648f
C12332 VDD.n3535 GND 0.04648f
C12333 VDD.n3536 GND 0.04648f
C12334 VDD.n3537 GND 0.04648f
C12335 VDD.n3538 GND 3.47277f
C12336 VDD.n3539 GND 0.04648f
C12337 VDD.n3540 GND 0.04648f
C12338 VDD.n3541 GND 0.04648f
C12339 VDD.n3542 GND 0.04648f
C12340 VDD.n3543 GND 0.04532f
C12341 VDD.n3544 GND 0.04532f
C12342 VDD.n3545 GND 0.02497f
C12343 VDD.n3546 GND 0.02497f
C12344 VDD.t89 GND 0.02104f
C12345 VDD.n3547 GND 0.22365f
C12346 VDD.t152 GND 0.02104f
C12347 VDD.t666 GND 0.02104f
C12348 VDD.n3548 GND 0.04891f
C12349 VDD.n3549 GND 0.04891f
C12350 VDD.n3550 GND 0.04532f
C12351 VDD.n3551 GND 0.04648f
C12352 VDD.n3552 GND 0.02293f
C12353 VDD.n3553 GND 0.02708f
C12354 VDD.n3554 GND 0.02293f
C12355 VDD.n3555 GND 0.04532f
C12356 VDD.n3556 GND 0.04532f
C12357 VDD.n3557 GND 0.04532f
C12358 VDD.n3558 GND 0.04532f
C12359 VDD.n3559 GND 0.04532f
C12360 VDD.n3560 GND 0.04532f
C12361 VDD.n3561 GND 0.04532f
C12362 VDD.n3562 GND 0.04532f
C12363 VDD.n3563 GND 0.04532f
C12364 VDD.n3564 GND 0.04532f
C12365 VDD.n3565 GND 0.04532f
C12366 VDD.n3566 GND 0.04532f
C12367 VDD.n3567 GND 0.04532f
C12368 VDD.n3568 GND 0.04532f
C12369 VDD.n3569 GND 0.04532f
C12370 VDD.n3570 GND 0.04532f
C12371 VDD.n3571 GND 0.04532f
C12372 VDD.n3572 GND 0.04532f
C12373 VDD.n3573 GND 0.04532f
C12374 VDD.n3574 GND 0.04532f
C12375 VDD.n3575 GND 0.02293f
C12376 VDD.n3576 GND 0.02293f
C12377 VDD.n3577 GND 0.02708f
C12378 VDD.n3578 GND 0.04648f
C12379 VDD.n3579 GND 3.19829f
C12380 VDD.n3580 GND 0.04532f
C12381 VDD.n3581 GND 0.04648f
C12382 VDD.n3582 GND 0.04648f
C12383 VDD.n3583 GND 0.04891f
C12384 VDD.n3584 GND 0.02293f
C12385 VDD.t380 GND 0.02114f
C12386 VDD.t555 GND 0.02114f
C12387 VDD.t727 GND 0.02114f
C12388 VDD.t724 GND 0.02114f
C12389 VDD.n3585 GND 0.02324f
C12390 VDD.n3586 GND 0.04891f
C12391 VDD.n3587 GND 0.04648f
C12392 VDD.n3588 GND 0.02293f
C12393 VDD.n3589 GND 0.04648f
C12394 VDD.n3590 GND 0.02708f
C12395 VDD.n3591 GND 0.02293f
C12396 VDD.n3592 GND 0.02708f
C12397 VDD.n3593 GND 0.02293f
C12398 VDD.n3594 GND 0.04532f
C12399 VDD.n3595 GND 0.04532f
C12400 VDD.n3596 GND 0.04532f
C12401 VDD.n3597 GND 0.02293f
C12402 VDD.n3598 GND 0.02293f
C12403 VDD.n3599 GND 0.02708f
C12404 VDD.n3600 GND 0.04648f
C12405 VDD.n3601 GND 0.04648f
C12406 VDD.n3602 GND 0.04648f
C12407 VDD.n3603 GND 0.04648f
C12408 VDD.n3604 GND 0.04532f
C12409 VDD.n3605 GND 0.04532f
C12410 VDD.n3606 GND 0.02293f
C12411 VDD.n3607 GND 0.02293f
C12412 VDD.n3608 GND 0.04648f
C12413 VDD.n3609 GND 0.02708f
C12414 VDD.n3610 GND 0.02293f
C12415 VDD.n3611 GND 0.04891f
C12416 VDD.n3612 GND 0.04648f
C12417 VDD.n3613 GND 0.05737f
C12418 VDD.n3614 GND 0.04891f
C12419 VDD.n3615 GND 0.02293f
C12420 VDD.n3616 GND 0.02708f
C12421 VDD.n3617 GND 0.04648f
C12422 VDD.n3618 GND 0.04532f
C12423 VDD.n3619 GND 0.04532f
C12424 VDD.n3620 GND 0.02293f
C12425 VDD.n3621 GND 0.02708f
C12426 VDD.n3622 GND 0.04648f
C12427 VDD.n3623 GND 0.04648f
C12428 VDD.n3624 GND 0.04648f
C12429 VDD.n3625 GND 0.04532f
C12430 VDD.n3626 GND 0.04532f
C12431 VDD.n3627 GND 0.02293f
C12432 VDD.n3628 GND 0.02293f
C12433 VDD.n3629 GND 0.04648f
C12434 VDD.n3630 GND 0.02708f
C12435 VDD.n3631 GND 0.02293f
C12436 VDD.n3632 GND 0.04891f
C12437 VDD.n3633 GND 0.04648f
C12438 VDD.t154 GND 0.02104f
C12439 VDD.t676 GND 0.02104f
C12440 VDD.t246 GND 0.02114f
C12441 VDD.t324 GND 0.02114f
C12442 VDD.n3634 GND 0.44561f
C12443 VDD.n3635 GND 0.04891f
C12444 VDD.n3636 GND 0.04648f
C12445 VDD.n3637 GND 0.02293f
C12446 VDD.n3638 GND 0.04648f
C12447 VDD.n3639 GND 0.02708f
C12448 VDD.n3640 GND 0.02293f
C12449 VDD.n3641 GND 0.04532f
C12450 VDD.n3642 GND 0.02293f
C12451 VDD.n3643 GND 0.02708f
C12452 VDD.n3644 GND 0.04532f
C12453 VDD.n3645 GND 0.02293f
C12454 VDD.n3646 GND 0.04891f
C12455 VDD.n3647 GND 0.05737f
C12456 VDD.n3648 GND 0.02055f
C12457 VDD.n3649 GND 0.08471f
C12458 VDD.n3650 GND 0.95576f
C12459 VDD.t331 GND 0.02114f
C12460 VDD.t581 GND 0.02114f
C12461 VDD.t15 GND 0.02114f
C12462 VDD.t34 GND 0.02114f
C12463 VDD.t294 GND 0.02104f
C12464 VDD.t33 GND 0.02114f
C12465 VDD.t592 GND 0.02114f
C12466 VDD.t26 GND 0.02114f
C12467 VDD.t25 GND 0.02114f
C12468 VDD.t114 GND 0.02104f
C12469 VDD.t661 GND 0.02104f
C12470 VDD.n3651 GND 0.95576f
C12471 VDD.n3652 GND 0.08471f
C12472 VDD.n3653 GND 0.04891f
C12473 VDD.n3654 GND 0.04648f
C12474 VDD.n3655 GND 0.02293f
C12475 VDD.n3656 GND 0.04648f
C12476 VDD.n3657 GND 0.02708f
C12477 VDD.n3658 GND 0.02293f
C12478 VDD.n3659 GND 0.04532f
C12479 VDD.n3660 GND 0.02293f
C12480 VDD.n3661 GND 0.02708f
C12481 VDD.n3662 GND 0.04532f
C12482 VDD.n3663 GND 0.02293f
C12483 VDD.n3664 GND 0.04891f
C12484 VDD.n3665 GND 0.05737f
C12485 VDD.n3666 GND 0.02055f
C12486 VDD.n3667 GND 0.44561f
C12487 VDD.n3668 GND 0.14059f
C12488 VDD.n3669 GND 0.04891f
C12489 VDD.n3670 GND 0.04648f
C12490 VDD.n3671 GND 0.02293f
C12491 VDD.n3672 GND 0.04648f
C12492 VDD.n3673 GND 0.02708f
C12493 VDD.n3674 GND 0.02293f
C12494 VDD.n3675 GND 0.04532f
C12495 VDD.n3676 GND 0.02293f
C12496 VDD.n3677 GND 0.02708f
C12497 VDD.n3678 GND 0.04532f
C12498 VDD.n3679 GND 0.02293f
C12499 VDD.n3680 GND 0.04891f
C12500 VDD.n3681 GND 0.05737f
C12501 VDD.n3682 GND 0.02055f
C12502 VDD.n3683 GND 0.02497f
C12503 VDD.n3684 GND 0.04648f
C12504 VDD.n3685 GND 0.04648f
C12505 VDD.n3686 GND 0.02708f
C12506 VDD.n3687 GND 0.02497f
C12507 VDD.n3688 GND 0.08328f
C12508 VDD.n3689 GND 0.01566f
C12509 VDD.n3690 GND 0.18236f
C12510 VDD.n3691 GND 0.03549f
C12511 VDD.n3692 GND 0.04891f
C12512 VDD.n3693 GND 0.04648f
C12513 VDD.n3694 GND 0.02293f
C12514 VDD.n3695 GND 0.04648f
C12515 VDD.n3696 GND 0.02708f
C12516 VDD.n3697 GND 0.02293f
C12517 VDD.n3698 GND 0.04532f
C12518 VDD.n3699 GND 0.02293f
C12519 VDD.n3700 GND 0.02708f
C12520 VDD.n3701 GND 0.04532f
C12521 VDD.n3702 GND 0.02293f
C12522 VDD.n3703 GND 0.04891f
C12523 VDD.n3704 GND 0.05737f
C12524 VDD.n3705 GND 0.02055f
C12525 VDD.n3706 GND 0.44561f
C12526 VDD.n3707 GND 0.14059f
C12527 VDD.n3708 GND 0.04891f
C12528 VDD.n3709 GND 0.04648f
C12529 VDD.n3710 GND 0.02293f
C12530 VDD.n3711 GND 0.04648f
C12531 VDD.n3712 GND 0.02708f
C12532 VDD.n3713 GND 0.02293f
C12533 VDD.n3714 GND 0.04532f
C12534 VDD.n3715 GND 0.02293f
C12535 VDD.n3716 GND 0.02708f
C12536 VDD.n3717 GND 0.04532f
C12537 VDD.n3718 GND 0.02293f
C12538 VDD.n3719 GND 0.04891f
C12539 VDD.n3720 GND 0.05737f
C12540 VDD.n3721 GND 0.02813f
C12541 VDD.n3722 GND 0.02324f
C12542 VDD.n3723 GND 0.05737f
C12543 VDD.n3724 GND 0.04891f
C12544 VDD.n3725 GND 0.02293f
C12545 VDD.n3726 GND 0.02708f
C12546 VDD.n3727 GND 0.04648f
C12547 VDD.n3728 GND 0.02293f
C12548 VDD.n3729 GND 0.02293f
C12549 VDD.n3730 GND 0.02708f
C12550 VDD.n3731 GND 0.04648f
C12551 VDD.n3732 GND 0.02708f
C12552 VDD.n3733 GND 0.04648f
C12553 VDD.n3734 GND 3.19829f
C12554 VDD.n3735 GND 0.04648f
C12555 VDD.n3736 GND 0.04532f
C12556 VDD.n3737 GND 0.02293f
C12557 VDD.n3738 GND 0.04891f
C12558 VDD.n3739 GND 0.05737f
C12559 VDD.n3740 GND 0.02813f
C12560 VDD.n3741 GND 0.14059f
C12561 VDD.n3742 GND 0.44561f
C12562 VDD.n3743 GND 0.02055f
C12563 VDD.n3744 GND 0.05737f
C12564 VDD.n3745 GND 0.04891f
C12565 VDD.n3746 GND 0.02293f
C12566 VDD.n3747 GND 0.02708f
C12567 VDD.n3748 GND 0.02293f
C12568 VDD.n3749 GND 0.04532f
C12569 VDD.t14 GND 4.12913f
C12570 VDD.n3750 GND 0.04532f
C12571 VDD.n3751 GND 0.04648f
C12572 VDD.n3752 GND 0.05737f
C12573 VDD.n3753 GND 0.01303f
C12574 VDD.n3754 GND 0.95576f
C12575 VDD.n3755 GND 0.08471f
C12576 VDD.n3756 GND 0.01566f
C12577 VDD.n3757 GND 0.08328f
C12578 VDD.n3758 GND 0.04648f
C12579 VDD.n3759 GND 3.47277f
C12580 VDD.n3760 GND 0.04648f
C12581 VDD.n3761 GND 0.05737f
C12582 VDD.n3762 GND 0.0171f
C12583 VDD.n3763 GND 0.064f
C12584 VDD.n3766 GND 0.06555f
C12585 VDD.n3767 GND 0.03083f
C12586 VDD.t113 GND 0.08047f
C12587 VDD.n3768 GND 0.03534f
C12588 VDD.t950 GND 0.15471f
C12589 VDD.n3769 GND 0.03238f
C12590 VDD.n3770 GND 0.02607f
C12591 VDD.n3771 GND 0.09595f
C12592 VDD.t153 GND 0.08047f
C12593 VDD.n3772 GND 0.03534f
C12594 VDD.t937 GND 0.15471f
C12595 VDD.n3773 GND 0.03238f
C12596 VDD.n3774 GND 0.02607f
C12597 VDD.n3776 GND 0.24365f
C12598 VDD.n3777 GND 0.03496f
C12599 VDD.n3778 GND 0.58129f
C12600 VDD.n3779 GND 0.43824f
C12601 VDD.t946 GND 0.15539f
C12602 VDD.n3780 GND 0.06697f
C12603 VDD.t198 GND 0.07226f
C12604 VDD.n3781 GND 0.05627f
C12605 VDD.n3782 GND 0.05442f
C12606 VDD.n3783 GND 0.04255f
C12607 VDD.n3784 GND 0.05152f
C12608 VDD.t272 GND 0.02114f
C12609 VDD.t887 GND 0.02114f
C12610 VDD.n3785 GND 0.14059f
C12611 VDD.n3786 GND 0.04891f
C12612 VDD.n3787 GND 0.04648f
C12613 VDD.n3788 GND 0.04891f
C12614 VDD.n3789 GND 0.04532f
C12615 VDD.n3790 GND 0.04532f
C12616 VDD.t199 GND 4.12913f
C12617 VDD.n3791 GND 0.04648f
C12618 VDD.n3792 GND 0.04648f
C12619 VDD.n3793 GND 0.04648f
C12620 VDD.n3794 GND 0.04648f
C12621 VDD.n3795 GND 0.04648f
C12622 VDD.n3796 GND 0.04648f
C12623 VDD.n3797 GND 3.47277f
C12624 VDD.n3798 GND 0.04648f
C12625 VDD.n3799 GND 0.04648f
C12626 VDD.n3800 GND 0.04648f
C12627 VDD.n3801 GND 0.04648f
C12628 VDD.n3802 GND 0.04532f
C12629 VDD.n3803 GND 0.04532f
C12630 VDD.n3804 GND 0.02497f
C12631 VDD.n3805 GND 0.02497f
C12632 VDD.t890 GND 0.02104f
C12633 VDD.n3806 GND 0.22365f
C12634 VDD.t200 GND 0.02104f
C12635 VDD.t649 GND 0.02104f
C12636 VDD.n3807 GND 0.04891f
C12637 VDD.n3808 GND 0.04891f
C12638 VDD.n3809 GND 0.04532f
C12639 VDD.n3810 GND 0.04648f
C12640 VDD.n3811 GND 0.02293f
C12641 VDD.n3812 GND 0.02708f
C12642 VDD.n3813 GND 0.02293f
C12643 VDD.n3814 GND 0.04532f
C12644 VDD.n3815 GND 0.04532f
C12645 VDD.n3816 GND 0.04532f
C12646 VDD.n3817 GND 0.04532f
C12647 VDD.n3818 GND 0.04532f
C12648 VDD.n3819 GND 0.04532f
C12649 VDD.n3820 GND 0.04532f
C12650 VDD.n3821 GND 0.04532f
C12651 VDD.n3822 GND 0.04532f
C12652 VDD.n3823 GND 0.04532f
C12653 VDD.n3824 GND 0.04532f
C12654 VDD.n3825 GND 0.04532f
C12655 VDD.n3826 GND 0.04532f
C12656 VDD.n3827 GND 0.04532f
C12657 VDD.n3828 GND 0.04532f
C12658 VDD.n3829 GND 0.04532f
C12659 VDD.n3830 GND 0.04532f
C12660 VDD.n3831 GND 0.04532f
C12661 VDD.n3832 GND 0.04532f
C12662 VDD.n3833 GND 0.04532f
C12663 VDD.n3834 GND 0.02293f
C12664 VDD.n3835 GND 0.02293f
C12665 VDD.n3836 GND 0.02708f
C12666 VDD.n3837 GND 0.04648f
C12667 VDD.n3838 GND 3.19829f
C12668 VDD.n3839 GND 0.04532f
C12669 VDD.n3840 GND 0.04648f
C12670 VDD.n3841 GND 0.04648f
C12671 VDD.n3842 GND 0.04891f
C12672 VDD.n3843 GND 0.02293f
C12673 VDD.t271 GND 0.02114f
C12674 VDD.t865 GND 0.02114f
C12675 VDD.t834 GND 0.02114f
C12676 VDD.t609 GND 0.02114f
C12677 VDD.n3844 GND 0.02324f
C12678 VDD.n3845 GND 0.04891f
C12679 VDD.n3846 GND 0.04648f
C12680 VDD.n3847 GND 0.02293f
C12681 VDD.n3848 GND 0.04648f
C12682 VDD.n3849 GND 0.02708f
C12683 VDD.n3850 GND 0.02293f
C12684 VDD.n3851 GND 0.02708f
C12685 VDD.n3852 GND 0.02293f
C12686 VDD.n3853 GND 0.04532f
C12687 VDD.n3854 GND 0.04532f
C12688 VDD.n3855 GND 0.04532f
C12689 VDD.n3856 GND 0.02293f
C12690 VDD.n3857 GND 0.02293f
C12691 VDD.n3858 GND 0.02708f
C12692 VDD.n3859 GND 0.04648f
C12693 VDD.n3860 GND 0.04648f
C12694 VDD.n3861 GND 0.04648f
C12695 VDD.n3862 GND 0.04648f
C12696 VDD.n3863 GND 0.04532f
C12697 VDD.n3864 GND 0.04532f
C12698 VDD.n3865 GND 0.02293f
C12699 VDD.n3866 GND 0.02293f
C12700 VDD.n3867 GND 0.04648f
C12701 VDD.n3868 GND 0.02708f
C12702 VDD.n3869 GND 0.02293f
C12703 VDD.n3870 GND 0.04891f
C12704 VDD.n3871 GND 0.04648f
C12705 VDD.n3872 GND 0.05737f
C12706 VDD.n3873 GND 0.04891f
C12707 VDD.n3874 GND 0.02293f
C12708 VDD.n3875 GND 0.02708f
C12709 VDD.n3876 GND 0.04648f
C12710 VDD.n3877 GND 0.04532f
C12711 VDD.n3878 GND 0.04532f
C12712 VDD.n3879 GND 0.02293f
C12713 VDD.n3880 GND 0.02708f
C12714 VDD.n3881 GND 0.04648f
C12715 VDD.n3882 GND 0.04648f
C12716 VDD.n3883 GND 0.04648f
C12717 VDD.n3884 GND 0.04532f
C12718 VDD.n3885 GND 0.04532f
C12719 VDD.n3886 GND 0.02293f
C12720 VDD.n3887 GND 0.02293f
C12721 VDD.n3888 GND 0.04648f
C12722 VDD.n3889 GND 0.02708f
C12723 VDD.n3890 GND 0.02293f
C12724 VDD.n3891 GND 0.04891f
C12725 VDD.n3892 GND 0.04648f
C12726 VDD.t117 GND 0.02104f
C12727 VDD.t695 GND 0.02104f
C12728 VDD.t816 GND 0.02114f
C12729 VDD.t833 GND 0.02114f
C12730 VDD.n3893 GND 0.44561f
C12731 VDD.n3894 GND 0.04891f
C12732 VDD.n3895 GND 0.04648f
C12733 VDD.n3896 GND 0.02293f
C12734 VDD.n3897 GND 0.04648f
C12735 VDD.n3898 GND 0.02708f
C12736 VDD.n3899 GND 0.02293f
C12737 VDD.n3900 GND 0.04532f
C12738 VDD.n3901 GND 0.02293f
C12739 VDD.n3902 GND 0.02708f
C12740 VDD.n3903 GND 0.04532f
C12741 VDD.n3904 GND 0.02293f
C12742 VDD.n3905 GND 0.04891f
C12743 VDD.n3906 GND 0.05737f
C12744 VDD.n3907 GND 0.02055f
C12745 VDD.n3908 GND 0.08471f
C12746 VDD.n3909 GND 0.95576f
C12747 VDD.t730 GND 0.02114f
C12748 VDD.t777 GND 0.02114f
C12749 VDD.t814 GND 0.02114f
C12750 VDD.t778 GND 0.02114f
C12751 VDD.t249 GND 0.02104f
C12752 VDD.t779 GND 0.02114f
C12753 VDD.t825 GND 0.02114f
C12754 VDD.t518 GND 0.02114f
C12755 VDD.t517 GND 0.02114f
C12756 VDD.t204 GND 0.02104f
C12757 VDD.t688 GND 0.02104f
C12758 VDD.n3910 GND 0.95576f
C12759 VDD.n3911 GND 0.08471f
C12760 VDD.n3912 GND 0.04891f
C12761 VDD.n3913 GND 0.04648f
C12762 VDD.n3914 GND 0.02293f
C12763 VDD.n3915 GND 0.04648f
C12764 VDD.n3916 GND 0.02708f
C12765 VDD.n3917 GND 0.02293f
C12766 VDD.n3918 GND 0.04532f
C12767 VDD.n3919 GND 0.02293f
C12768 VDD.n3920 GND 0.02708f
C12769 VDD.n3921 GND 0.04532f
C12770 VDD.n3922 GND 0.02293f
C12771 VDD.n3923 GND 0.04891f
C12772 VDD.n3924 GND 0.05737f
C12773 VDD.n3925 GND 0.02055f
C12774 VDD.n3926 GND 0.44561f
C12775 VDD.n3927 GND 0.14059f
C12776 VDD.n3928 GND 0.04891f
C12777 VDD.n3929 GND 0.04648f
C12778 VDD.n3930 GND 0.02293f
C12779 VDD.n3931 GND 0.04648f
C12780 VDD.n3932 GND 0.02708f
C12781 VDD.n3933 GND 0.02293f
C12782 VDD.n3934 GND 0.04532f
C12783 VDD.n3935 GND 0.02293f
C12784 VDD.n3936 GND 0.02708f
C12785 VDD.n3937 GND 0.04532f
C12786 VDD.n3938 GND 0.02293f
C12787 VDD.n3939 GND 0.04891f
C12788 VDD.n3940 GND 0.05737f
C12789 VDD.n3941 GND 0.02055f
C12790 VDD.n3942 GND 0.02497f
C12791 VDD.n3943 GND 0.04648f
C12792 VDD.n3944 GND 0.04648f
C12793 VDD.n3945 GND 0.02708f
C12794 VDD.n3946 GND 0.02497f
C12795 VDD.n3947 GND 0.08328f
C12796 VDD.n3948 GND 0.01566f
C12797 VDD.n3949 GND 0.18236f
C12798 VDD.n3950 GND 0.03549f
C12799 VDD.n3951 GND 0.04891f
C12800 VDD.n3952 GND 0.04648f
C12801 VDD.n3953 GND 0.02293f
C12802 VDD.n3954 GND 0.04648f
C12803 VDD.n3955 GND 0.02708f
C12804 VDD.n3956 GND 0.02293f
C12805 VDD.n3957 GND 0.04532f
C12806 VDD.n3958 GND 0.02293f
C12807 VDD.n3959 GND 0.02708f
C12808 VDD.n3960 GND 0.04532f
C12809 VDD.n3961 GND 0.02293f
C12810 VDD.n3962 GND 0.04891f
C12811 VDD.n3963 GND 0.05737f
C12812 VDD.n3964 GND 0.02055f
C12813 VDD.n3965 GND 0.44561f
C12814 VDD.n3966 GND 0.14059f
C12815 VDD.n3967 GND 0.04891f
C12816 VDD.n3968 GND 0.04648f
C12817 VDD.n3969 GND 0.02293f
C12818 VDD.n3970 GND 0.04648f
C12819 VDD.n3971 GND 0.02708f
C12820 VDD.n3972 GND 0.02293f
C12821 VDD.n3973 GND 0.04532f
C12822 VDD.n3974 GND 0.02293f
C12823 VDD.n3975 GND 0.02708f
C12824 VDD.n3976 GND 0.04532f
C12825 VDD.n3977 GND 0.02293f
C12826 VDD.n3978 GND 0.04891f
C12827 VDD.n3979 GND 0.05737f
C12828 VDD.n3980 GND 0.02813f
C12829 VDD.n3981 GND 0.02324f
C12830 VDD.n3982 GND 0.05737f
C12831 VDD.n3983 GND 0.04891f
C12832 VDD.n3984 GND 0.02293f
C12833 VDD.n3985 GND 0.02708f
C12834 VDD.n3986 GND 0.04648f
C12835 VDD.n3987 GND 0.02293f
C12836 VDD.n3988 GND 0.02293f
C12837 VDD.n3989 GND 0.02708f
C12838 VDD.n3990 GND 0.04648f
C12839 VDD.n3991 GND 0.02708f
C12840 VDD.n3992 GND 0.04648f
C12841 VDD.n3993 GND 3.19829f
C12842 VDD.n3994 GND 0.04648f
C12843 VDD.n3995 GND 0.04532f
C12844 VDD.n3996 GND 0.02293f
C12845 VDD.n3997 GND 0.04891f
C12846 VDD.n3998 GND 0.05737f
C12847 VDD.n3999 GND 0.02813f
C12848 VDD.n4000 GND 0.14059f
C12849 VDD.n4001 GND 0.44561f
C12850 VDD.n4002 GND 0.02055f
C12851 VDD.n4003 GND 0.05737f
C12852 VDD.n4004 GND 0.04891f
C12853 VDD.n4005 GND 0.02293f
C12854 VDD.n4006 GND 0.02708f
C12855 VDD.n4007 GND 0.02293f
C12856 VDD.n4008 GND 0.04532f
C12857 VDD.t116 GND 4.12913f
C12858 VDD.n4009 GND 0.04532f
C12859 VDD.n4010 GND 0.04648f
C12860 VDD.n4011 GND 0.05737f
C12861 VDD.n4012 GND 0.01303f
C12862 VDD.n4013 GND 0.95576f
C12863 VDD.n4014 GND 0.08471f
C12864 VDD.n4015 GND 0.01566f
C12865 VDD.n4016 GND 0.08328f
C12866 VDD.n4017 GND 0.04648f
C12867 VDD.n4018 GND 3.47277f
C12868 VDD.n4019 GND 0.04648f
C12869 VDD.n4020 GND 0.05737f
C12870 VDD.n4021 GND 0.0171f
C12871 VDD.n4022 GND 0.064f
C12872 VDD.n4025 GND 0.06555f
C12873 VDD.n4026 GND 0.03083f
C12874 VDD.t203 GND 0.08047f
C12875 VDD.n4027 GND 0.03534f
C12876 VDD.t960 GND 0.15471f
C12877 VDD.n4028 GND 0.03238f
C12878 VDD.n4029 GND 0.02607f
C12879 VDD.n4030 GND 0.09595f
C12880 VDD.t115 GND 0.08047f
C12881 VDD.n4031 GND 0.03534f
C12882 VDD.t957 GND 0.15471f
C12883 VDD.n4032 GND 0.03238f
C12884 VDD.n4033 GND 0.02607f
C12885 VDD.n4035 GND 0.24365f
C12886 VDD.n4036 GND 0.03496f
C12887 VDD.n4037 GND 0.4211f
C12888 VDD.n4038 GND 0.29261f
C12889 VDD.t958 GND 0.15539f
C12890 VDD.n4039 GND 0.06697f
C12891 VDD.t187 GND 0.07226f
C12892 VDD.n4040 GND 0.05627f
C12893 VDD.n4041 GND 0.05442f
C12894 VDD.n4042 GND 0.04255f
C12895 VDD.n4043 GND 0.05152f
C12896 VDD.t319 GND 0.02114f
C12897 VDD.t912 GND 0.02114f
C12898 VDD.n4044 GND 0.14059f
C12899 VDD.n4045 GND 0.04891f
C12900 VDD.n4046 GND 0.04648f
C12901 VDD.n4047 GND 0.04891f
C12902 VDD.n4048 GND 0.04532f
C12903 VDD.n4049 GND 0.04532f
C12904 VDD.t8 GND 4.12913f
C12905 VDD.n4050 GND 0.04648f
C12906 VDD.n4051 GND 0.04648f
C12907 VDD.n4052 GND 0.04648f
C12908 VDD.n4053 GND 0.04648f
C12909 VDD.n4054 GND 0.04648f
C12910 VDD.n4055 GND 0.04648f
C12911 VDD.n4056 GND 3.47277f
C12912 VDD.n4057 GND 0.04648f
C12913 VDD.n4058 GND 0.04648f
C12914 VDD.n4059 GND 0.04648f
C12915 VDD.n4060 GND 0.04648f
C12916 VDD.n4061 GND 0.04532f
C12917 VDD.n4062 GND 0.04532f
C12918 VDD.n4063 GND 0.02497f
C12919 VDD.n4064 GND 0.02497f
C12920 VDD.t407 GND 0.02104f
C12921 VDD.n4065 GND 0.22365f
C12922 VDD.t188 GND 0.02104f
C12923 VDD.t686 GND 0.02104f
C12924 VDD.n4066 GND 0.04891f
C12925 VDD.n4067 GND 0.04891f
C12926 VDD.n4068 GND 0.04532f
C12927 VDD.n4069 GND 0.04648f
C12928 VDD.n4070 GND 0.02293f
C12929 VDD.n4071 GND 0.02708f
C12930 VDD.n4072 GND 0.02293f
C12931 VDD.n4073 GND 0.04532f
C12932 VDD.n4074 GND 0.04532f
C12933 VDD.n4075 GND 0.04532f
C12934 VDD.n4076 GND 0.04532f
C12935 VDD.n4077 GND 0.04532f
C12936 VDD.n4078 GND 0.04532f
C12937 VDD.n4079 GND 0.04532f
C12938 VDD.n4080 GND 0.04532f
C12939 VDD.n4081 GND 0.04532f
C12940 VDD.n4082 GND 0.04532f
C12941 VDD.n4083 GND 0.04532f
C12942 VDD.n4084 GND 0.04532f
C12943 VDD.n4085 GND 0.04532f
C12944 VDD.n4086 GND 0.04532f
C12945 VDD.n4087 GND 0.04532f
C12946 VDD.n4088 GND 0.04532f
C12947 VDD.n4089 GND 0.04532f
C12948 VDD.n4090 GND 0.04532f
C12949 VDD.n4091 GND 0.04532f
C12950 VDD.n4092 GND 0.04532f
C12951 VDD.n4093 GND 0.02293f
C12952 VDD.n4094 GND 0.02293f
C12953 VDD.n4095 GND 0.02708f
C12954 VDD.n4096 GND 0.04648f
C12955 VDD.n4097 GND 3.19829f
C12956 VDD.n4098 GND 0.04532f
C12957 VDD.n4099 GND 0.04648f
C12958 VDD.n4100 GND 0.04648f
C12959 VDD.n4101 GND 0.04891f
C12960 VDD.n4102 GND 0.02293f
C12961 VDD.t471 GND 0.02114f
C12962 VDD.t601 GND 0.02114f
C12963 VDD.t481 GND 0.02114f
C12964 VDD.t799 GND 0.02114f
C12965 VDD.n4103 GND 0.02324f
C12966 VDD.n4104 GND 0.04891f
C12967 VDD.n4105 GND 0.04648f
C12968 VDD.n4106 GND 0.02293f
C12969 VDD.n4107 GND 0.04648f
C12970 VDD.n4108 GND 0.02708f
C12971 VDD.n4109 GND 0.02293f
C12972 VDD.n4110 GND 0.02708f
C12973 VDD.n4111 GND 0.02293f
C12974 VDD.n4112 GND 0.04532f
C12975 VDD.n4113 GND 0.04532f
C12976 VDD.n4114 GND 0.04532f
C12977 VDD.n4115 GND 0.02293f
C12978 VDD.n4116 GND 0.02293f
C12979 VDD.n4117 GND 0.02708f
C12980 VDD.n4118 GND 0.04648f
C12981 VDD.n4119 GND 0.04648f
C12982 VDD.n4120 GND 0.04648f
C12983 VDD.n4121 GND 0.04648f
C12984 VDD.n4122 GND 0.04532f
C12985 VDD.n4123 GND 0.04532f
C12986 VDD.n4124 GND 0.02293f
C12987 VDD.n4125 GND 0.02293f
C12988 VDD.n4126 GND 0.04648f
C12989 VDD.n4127 GND 0.02708f
C12990 VDD.n4128 GND 0.02293f
C12991 VDD.n4129 GND 0.04891f
C12992 VDD.n4130 GND 0.04648f
C12993 VDD.n4131 GND 0.05737f
C12994 VDD.n4132 GND 0.04891f
C12995 VDD.n4133 GND 0.02293f
C12996 VDD.n4134 GND 0.02708f
C12997 VDD.n4135 GND 0.04648f
C12998 VDD.n4136 GND 0.04532f
C12999 VDD.n4137 GND 0.04532f
C13000 VDD.n4138 GND 0.02293f
C13001 VDD.n4139 GND 0.02708f
C13002 VDD.n4140 GND 0.04648f
C13003 VDD.n4141 GND 0.04648f
C13004 VDD.n4142 GND 0.04648f
C13005 VDD.n4143 GND 0.04532f
C13006 VDD.n4144 GND 0.04532f
C13007 VDD.n4145 GND 0.02293f
C13008 VDD.n4146 GND 0.02293f
C13009 VDD.n4147 GND 0.04648f
C13010 VDD.n4148 GND 0.02708f
C13011 VDD.n4149 GND 0.02293f
C13012 VDD.n4150 GND 0.04891f
C13013 VDD.n4151 GND 0.04648f
C13014 VDD.t195 GND 0.02104f
C13015 VDD.t687 GND 0.02104f
C13016 VDD.t239 GND 0.02114f
C13017 VDD.t242 GND 0.02114f
C13018 VDD.n4152 GND 0.44561f
C13019 VDD.n4153 GND 0.04891f
C13020 VDD.n4154 GND 0.04648f
C13021 VDD.n4155 GND 0.02293f
C13022 VDD.n4156 GND 0.04648f
C13023 VDD.n4157 GND 0.02708f
C13024 VDD.n4158 GND 0.02293f
C13025 VDD.n4159 GND 0.04532f
C13026 VDD.n4160 GND 0.02293f
C13027 VDD.n4161 GND 0.02708f
C13028 VDD.n4162 GND 0.04532f
C13029 VDD.n4163 GND 0.02293f
C13030 VDD.n4164 GND 0.04891f
C13031 VDD.n4165 GND 0.05737f
C13032 VDD.n4166 GND 0.02055f
C13033 VDD.n4167 GND 0.08471f
C13034 VDD.n4168 GND 0.95576f
C13035 VDD.t378 GND 0.02114f
C13036 VDD.t580 GND 0.02114f
C13037 VDD.t221 GND 0.02114f
C13038 VDD.t415 GND 0.02114f
C13039 VDD.t811 GND 0.02104f
C13040 VDD.t416 GND 0.02114f
C13041 VDD.t783 GND 0.02114f
C13042 VDD.t7 GND 0.02114f
C13043 VDD.t9 GND 0.02114f
C13044 VDD.t182 GND 0.02104f
C13045 VDD.t682 GND 0.02104f
C13046 VDD.n4169 GND 0.95576f
C13047 VDD.n4170 GND 0.08471f
C13048 VDD.n4171 GND 0.04891f
C13049 VDD.n4172 GND 0.04648f
C13050 VDD.n4173 GND 0.02293f
C13051 VDD.n4174 GND 0.04648f
C13052 VDD.n4175 GND 0.02708f
C13053 VDD.n4176 GND 0.02293f
C13054 VDD.n4177 GND 0.04532f
C13055 VDD.n4178 GND 0.02293f
C13056 VDD.n4179 GND 0.02708f
C13057 VDD.n4180 GND 0.04532f
C13058 VDD.n4181 GND 0.02293f
C13059 VDD.n4182 GND 0.04891f
C13060 VDD.n4183 GND 0.05737f
C13061 VDD.n4184 GND 0.02055f
C13062 VDD.n4185 GND 0.44561f
C13063 VDD.n4186 GND 0.14059f
C13064 VDD.n4187 GND 0.04891f
C13065 VDD.n4188 GND 0.04648f
C13066 VDD.n4189 GND 0.02293f
C13067 VDD.n4190 GND 0.04648f
C13068 VDD.n4191 GND 0.02708f
C13069 VDD.n4192 GND 0.02293f
C13070 VDD.n4193 GND 0.04532f
C13071 VDD.n4194 GND 0.02293f
C13072 VDD.n4195 GND 0.02708f
C13073 VDD.n4196 GND 0.04532f
C13074 VDD.n4197 GND 0.02293f
C13075 VDD.n4198 GND 0.04891f
C13076 VDD.n4199 GND 0.05737f
C13077 VDD.n4200 GND 0.02055f
C13078 VDD.n4201 GND 0.02497f
C13079 VDD.n4202 GND 0.04648f
C13080 VDD.n4203 GND 0.04648f
C13081 VDD.n4204 GND 0.02708f
C13082 VDD.n4205 GND 0.02497f
C13083 VDD.n4206 GND 0.08328f
C13084 VDD.n4207 GND 0.01566f
C13085 VDD.n4208 GND 0.18236f
C13086 VDD.n4209 GND 0.03549f
C13087 VDD.n4210 GND 0.04891f
C13088 VDD.n4211 GND 0.04648f
C13089 VDD.n4212 GND 0.02293f
C13090 VDD.n4213 GND 0.04648f
C13091 VDD.n4214 GND 0.02708f
C13092 VDD.n4215 GND 0.02293f
C13093 VDD.n4216 GND 0.04532f
C13094 VDD.n4217 GND 0.02293f
C13095 VDD.n4218 GND 0.02708f
C13096 VDD.n4219 GND 0.04532f
C13097 VDD.n4220 GND 0.02293f
C13098 VDD.n4221 GND 0.04891f
C13099 VDD.n4222 GND 0.05737f
C13100 VDD.n4223 GND 0.02055f
C13101 VDD.n4224 GND 0.44561f
C13102 VDD.n4225 GND 0.14059f
C13103 VDD.n4226 GND 0.04891f
C13104 VDD.n4227 GND 0.04648f
C13105 VDD.n4228 GND 0.02293f
C13106 VDD.n4229 GND 0.04648f
C13107 VDD.n4230 GND 0.02708f
C13108 VDD.n4231 GND 0.02293f
C13109 VDD.n4232 GND 0.04532f
C13110 VDD.n4233 GND 0.02293f
C13111 VDD.n4234 GND 0.02708f
C13112 VDD.n4235 GND 0.04532f
C13113 VDD.n4236 GND 0.02293f
C13114 VDD.n4237 GND 0.04891f
C13115 VDD.n4238 GND 0.05737f
C13116 VDD.n4239 GND 0.02813f
C13117 VDD.n4240 GND 0.02324f
C13118 VDD.n4241 GND 0.05737f
C13119 VDD.n4242 GND 0.04891f
C13120 VDD.n4243 GND 0.02293f
C13121 VDD.n4244 GND 0.02708f
C13122 VDD.n4245 GND 0.04648f
C13123 VDD.n4246 GND 0.02293f
C13124 VDD.n4247 GND 0.02293f
C13125 VDD.n4248 GND 0.02708f
C13126 VDD.n4249 GND 0.04648f
C13127 VDD.n4250 GND 0.02708f
C13128 VDD.n4251 GND 0.04648f
C13129 VDD.n4252 GND 3.19829f
C13130 VDD.n4253 GND 0.04648f
C13131 VDD.n4254 GND 0.04532f
C13132 VDD.n4255 GND 0.02293f
C13133 VDD.n4256 GND 0.04891f
C13134 VDD.n4257 GND 0.05737f
C13135 VDD.n4258 GND 0.02813f
C13136 VDD.n4259 GND 0.14059f
C13137 VDD.n4260 GND 0.44561f
C13138 VDD.n4261 GND 0.02055f
C13139 VDD.n4262 GND 0.05737f
C13140 VDD.n4263 GND 0.04891f
C13141 VDD.n4264 GND 0.02293f
C13142 VDD.n4265 GND 0.02708f
C13143 VDD.n4266 GND 0.02293f
C13144 VDD.n4267 GND 0.04532f
C13145 VDD.t6 GND 4.12913f
C13146 VDD.n4268 GND 0.04532f
C13147 VDD.n4269 GND 0.04648f
C13148 VDD.n4270 GND 0.05737f
C13149 VDD.n4271 GND 0.01303f
C13150 VDD.n4272 GND 0.95576f
C13151 VDD.n4273 GND 0.08471f
C13152 VDD.n4274 GND 0.01566f
C13153 VDD.n4275 GND 0.08328f
C13154 VDD.n4276 GND 0.04648f
C13155 VDD.n4277 GND 3.47277f
C13156 VDD.n4278 GND 0.04648f
C13157 VDD.n4279 GND 0.05737f
C13158 VDD.n4280 GND 0.0171f
C13159 VDD.n4281 GND 0.064f
C13160 VDD.n4284 GND 0.06555f
C13161 VDD.n4285 GND 0.03083f
C13162 VDD.t181 GND 0.08047f
C13163 VDD.n4286 GND 0.03534f
C13164 VDD.t956 GND 0.15471f
C13165 VDD.n4287 GND 0.03238f
C13166 VDD.n4288 GND 0.02607f
C13167 VDD.n4289 GND 0.09595f
C13168 VDD.t194 GND 0.08047f
C13169 VDD.n4290 GND 0.03534f
C13170 VDD.t951 GND 0.15471f
C13171 VDD.n4291 GND 0.03238f
C13172 VDD.n4292 GND 0.02607f
C13173 VDD.n4294 GND 0.24365f
C13174 VDD.n4295 GND 0.03496f
C13175 VDD.n4296 GND 0.26091f
C13176 VDD.n4297 GND 0.14699f
C13177 VDD.t962 GND 0.15539f
C13178 VDD.n4298 GND 0.06697f
C13179 VDD.t192 GND 0.07226f
C13180 VDD.n4299 GND 0.05627f
C13181 VDD.n4300 GND 0.05442f
C13182 VDD.n4301 GND 0.04255f
C13183 VDD.n4302 GND 0.05152f
C13184 VDD.t437 GND 0.02114f
C13185 VDD.t467 GND 0.02114f
C13186 VDD.n4303 GND 0.14059f
C13187 VDD.n4304 GND 0.04891f
C13188 VDD.n4305 GND 0.04648f
C13189 VDD.n4306 GND 0.04891f
C13190 VDD.n4307 GND 0.04532f
C13191 VDD.n4308 GND 0.04532f
C13192 VDD.t76 GND 4.12913f
C13193 VDD.n4309 GND 0.04648f
C13194 VDD.n4310 GND 0.04648f
C13195 VDD.n4311 GND 0.04648f
C13196 VDD.n4312 GND 0.04648f
C13197 VDD.n4313 GND 0.04648f
C13198 VDD.n4314 GND 0.04648f
C13199 VDD.n4315 GND 3.47277f
C13200 VDD.n4316 GND 0.04648f
C13201 VDD.n4317 GND 0.04648f
C13202 VDD.n4318 GND 0.04648f
C13203 VDD.n4319 GND 0.04648f
C13204 VDD.n4320 GND 0.04532f
C13205 VDD.n4321 GND 0.04532f
C13206 VDD.n4322 GND 0.02497f
C13207 VDD.n4323 GND 0.02497f
C13208 VDD.t470 GND 0.02104f
C13209 VDD.n4324 GND 0.22365f
C13210 VDD.t193 GND 0.02104f
C13211 VDD.t683 GND 0.02104f
C13212 VDD.n4325 GND 0.04891f
C13213 VDD.n4326 GND 0.04891f
C13214 VDD.n4327 GND 0.04532f
C13215 VDD.n4328 GND 0.04648f
C13216 VDD.n4329 GND 0.02293f
C13217 VDD.n4330 GND 0.02708f
C13218 VDD.n4331 GND 0.02293f
C13219 VDD.n4332 GND 0.04532f
C13220 VDD.n4333 GND 0.04532f
C13221 VDD.n4334 GND 0.04532f
C13222 VDD.n4335 GND 0.04532f
C13223 VDD.n4336 GND 0.04532f
C13224 VDD.n4337 GND 0.04532f
C13225 VDD.n4338 GND 0.04532f
C13226 VDD.n4339 GND 0.04532f
C13227 VDD.n4340 GND 0.04532f
C13228 VDD.n4341 GND 0.04532f
C13229 VDD.n4342 GND 0.04532f
C13230 VDD.n4343 GND 0.04532f
C13231 VDD.n4344 GND 0.04532f
C13232 VDD.n4345 GND 0.04532f
C13233 VDD.n4346 GND 0.04532f
C13234 VDD.n4347 GND 0.04532f
C13235 VDD.n4348 GND 0.04532f
C13236 VDD.n4349 GND 0.04532f
C13237 VDD.n4350 GND 0.04532f
C13238 VDD.n4351 GND 0.04532f
C13239 VDD.n4352 GND 0.02293f
C13240 VDD.n4353 GND 0.02293f
C13241 VDD.n4354 GND 0.02708f
C13242 VDD.n4355 GND 0.04648f
C13243 VDD.n4356 GND 3.19829f
C13244 VDD.n4357 GND 0.04532f
C13245 VDD.n4358 GND 0.04648f
C13246 VDD.n4359 GND 0.04648f
C13247 VDD.n4360 GND 0.04891f
C13248 VDD.n4361 GND 0.02293f
C13249 VDD.t808 GND 0.02114f
C13250 VDD.t871 GND 0.02114f
C13251 VDD.t846 GND 0.02114f
C13252 VDD.t413 GND 0.02114f
C13253 VDD.n4362 GND 0.02324f
C13254 VDD.n4363 GND 0.04891f
C13255 VDD.n4364 GND 0.04648f
C13256 VDD.n4365 GND 0.02293f
C13257 VDD.n4366 GND 0.04648f
C13258 VDD.n4367 GND 0.02708f
C13259 VDD.n4368 GND 0.02293f
C13260 VDD.n4369 GND 0.02708f
C13261 VDD.n4370 GND 0.02293f
C13262 VDD.n4371 GND 0.04532f
C13263 VDD.n4372 GND 0.04532f
C13264 VDD.n4373 GND 0.04532f
C13265 VDD.n4374 GND 0.02293f
C13266 VDD.n4375 GND 0.02293f
C13267 VDD.n4376 GND 0.02708f
C13268 VDD.n4377 GND 0.04648f
C13269 VDD.n4378 GND 0.04648f
C13270 VDD.n4379 GND 0.04648f
C13271 VDD.n4380 GND 0.04648f
C13272 VDD.n4381 GND 0.04532f
C13273 VDD.n4382 GND 0.04532f
C13274 VDD.n4383 GND 0.02293f
C13275 VDD.n4384 GND 0.02293f
C13276 VDD.n4385 GND 0.04648f
C13277 VDD.n4386 GND 0.02708f
C13278 VDD.n4387 GND 0.02293f
C13279 VDD.n4388 GND 0.04891f
C13280 VDD.n4389 GND 0.04648f
C13281 VDD.n4390 GND 0.05737f
C13282 VDD.n4391 GND 0.04891f
C13283 VDD.n4392 GND 0.02293f
C13284 VDD.n4393 GND 0.02708f
C13285 VDD.n4394 GND 0.04648f
C13286 VDD.n4395 GND 0.04532f
C13287 VDD.n4396 GND 0.04532f
C13288 VDD.n4397 GND 0.02293f
C13289 VDD.n4398 GND 0.02708f
C13290 VDD.n4399 GND 0.04648f
C13291 VDD.n4400 GND 0.04648f
C13292 VDD.n4401 GND 0.04648f
C13293 VDD.n4402 GND 0.04532f
C13294 VDD.n4403 GND 0.04532f
C13295 VDD.n4404 GND 0.02293f
C13296 VDD.n4405 GND 0.02293f
C13297 VDD.n4406 GND 0.04648f
C13298 VDD.n4407 GND 0.02708f
C13299 VDD.n4408 GND 0.02293f
C13300 VDD.n4409 GND 0.04891f
C13301 VDD.n4410 GND 0.04648f
C13302 VDD.t184 GND 0.02104f
C13303 VDD.t691 GND 0.02104f
C13304 VDD.t236 GND 0.02114f
C13305 VDD.t254 GND 0.02114f
C13306 VDD.n4411 GND 0.44561f
C13307 VDD.n4412 GND 0.04891f
C13308 VDD.n4413 GND 0.04648f
C13309 VDD.n4414 GND 0.02293f
C13310 VDD.n4415 GND 0.04648f
C13311 VDD.n4416 GND 0.02708f
C13312 VDD.n4417 GND 0.02293f
C13313 VDD.n4418 GND 0.04532f
C13314 VDD.n4419 GND 0.02293f
C13315 VDD.n4420 GND 0.02708f
C13316 VDD.n4421 GND 0.04532f
C13317 VDD.n4422 GND 0.02293f
C13318 VDD.n4423 GND 0.04891f
C13319 VDD.n4424 GND 0.05737f
C13320 VDD.n4425 GND 0.02055f
C13321 VDD.n4426 GND 0.08471f
C13322 VDD.n4427 GND 0.95576f
C13323 VDD.t346 GND 0.02114f
C13324 VDD.t77 GND 0.02114f
C13325 VDD.t259 GND 0.02114f
C13326 VDD.t742 GND 0.02114f
C13327 VDD.t830 GND 0.02104f
C13328 VDD.t761 GND 0.02114f
C13329 VDD.t260 GND 0.02114f
C13330 VDD.t579 GND 0.02114f
C13331 VDD.t379 GND 0.02114f
C13332 VDD.t176 GND 0.02104f
C13333 VDD.t685 GND 0.02104f
C13334 VDD.n4428 GND 0.95576f
C13335 VDD.n4429 GND 0.08471f
C13336 VDD.n4430 GND 0.04891f
C13337 VDD.n4431 GND 0.04648f
C13338 VDD.n4432 GND 0.02293f
C13339 VDD.n4433 GND 0.04648f
C13340 VDD.n4434 GND 0.02708f
C13341 VDD.n4435 GND 0.02293f
C13342 VDD.n4436 GND 0.04532f
C13343 VDD.n4437 GND 0.02293f
C13344 VDD.n4438 GND 0.02708f
C13345 VDD.n4439 GND 0.04532f
C13346 VDD.n4440 GND 0.02293f
C13347 VDD.n4441 GND 0.04891f
C13348 VDD.n4442 GND 0.05737f
C13349 VDD.n4443 GND 0.02055f
C13350 VDD.n4444 GND 0.44561f
C13351 VDD.n4445 GND 0.14059f
C13352 VDD.n4446 GND 0.04891f
C13353 VDD.n4447 GND 0.04648f
C13354 VDD.n4448 GND 0.02293f
C13355 VDD.n4449 GND 0.04648f
C13356 VDD.n4450 GND 0.02708f
C13357 VDD.n4451 GND 0.02293f
C13358 VDD.n4452 GND 0.04532f
C13359 VDD.n4453 GND 0.02293f
C13360 VDD.n4454 GND 0.02708f
C13361 VDD.n4455 GND 0.04532f
C13362 VDD.n4456 GND 0.02293f
C13363 VDD.n4457 GND 0.04891f
C13364 VDD.n4458 GND 0.05737f
C13365 VDD.n4459 GND 0.02055f
C13366 VDD.n4460 GND 0.02497f
C13367 VDD.n4461 GND 0.04648f
C13368 VDD.n4462 GND 0.04648f
C13369 VDD.n4463 GND 0.02708f
C13370 VDD.n4464 GND 0.02497f
C13371 VDD.n4465 GND 0.08328f
C13372 VDD.n4466 GND 0.01566f
C13373 VDD.n4467 GND 0.18236f
C13374 VDD.n4468 GND 0.03549f
C13375 VDD.n4469 GND 0.04891f
C13376 VDD.n4470 GND 0.04648f
C13377 VDD.n4471 GND 0.02293f
C13378 VDD.n4472 GND 0.04648f
C13379 VDD.n4473 GND 0.02708f
C13380 VDD.n4474 GND 0.02293f
C13381 VDD.n4475 GND 0.04532f
C13382 VDD.n4476 GND 0.02293f
C13383 VDD.n4477 GND 0.02708f
C13384 VDD.n4478 GND 0.04532f
C13385 VDD.n4479 GND 0.02293f
C13386 VDD.n4480 GND 0.04891f
C13387 VDD.n4481 GND 0.05737f
C13388 VDD.n4482 GND 0.02055f
C13389 VDD.n4483 GND 0.44561f
C13390 VDD.n4484 GND 0.14059f
C13391 VDD.n4485 GND 0.04891f
C13392 VDD.n4486 GND 0.04648f
C13393 VDD.n4487 GND 0.02293f
C13394 VDD.n4488 GND 0.04648f
C13395 VDD.n4489 GND 0.02708f
C13396 VDD.n4490 GND 0.02293f
C13397 VDD.n4491 GND 0.04532f
C13398 VDD.n4492 GND 0.02293f
C13399 VDD.n4493 GND 0.02708f
C13400 VDD.n4494 GND 0.04532f
C13401 VDD.n4495 GND 0.02293f
C13402 VDD.n4496 GND 0.04891f
C13403 VDD.n4497 GND 0.05737f
C13404 VDD.n4498 GND 0.02813f
C13405 VDD.n4499 GND 0.02324f
C13406 VDD.n4500 GND 0.05737f
C13407 VDD.n4501 GND 0.04891f
C13408 VDD.n4502 GND 0.02293f
C13409 VDD.n4503 GND 0.02708f
C13410 VDD.n4504 GND 0.04648f
C13411 VDD.n4505 GND 0.02293f
C13412 VDD.n4506 GND 0.02293f
C13413 VDD.n4507 GND 0.02708f
C13414 VDD.n4508 GND 0.04648f
C13415 VDD.n4509 GND 0.02708f
C13416 VDD.n4510 GND 0.04648f
C13417 VDD.n4511 GND 3.19829f
C13418 VDD.n4512 GND 0.04648f
C13419 VDD.n4513 GND 0.04532f
C13420 VDD.n4514 GND 0.02293f
C13421 VDD.n4515 GND 0.04891f
C13422 VDD.n4516 GND 0.05737f
C13423 VDD.n4517 GND 0.02813f
C13424 VDD.n4518 GND 0.14059f
C13425 VDD.n4519 GND 0.44561f
C13426 VDD.n4520 GND 0.02055f
C13427 VDD.n4521 GND 0.05737f
C13428 VDD.n4522 GND 0.04891f
C13429 VDD.n4523 GND 0.02293f
C13430 VDD.n4524 GND 0.02708f
C13431 VDD.n4525 GND 0.02293f
C13432 VDD.n4526 GND 0.04532f
C13433 VDD.t175 GND 4.12913f
C13434 VDD.n4527 GND 0.04532f
C13435 VDD.n4528 GND 0.04648f
C13436 VDD.n4529 GND 0.05737f
C13437 VDD.n4530 GND 0.01303f
C13438 VDD.n4531 GND 0.95576f
C13439 VDD.n4532 GND 0.08471f
C13440 VDD.n4533 GND 0.01566f
C13441 VDD.n4534 GND 0.08328f
C13442 VDD.n4535 GND 0.04648f
C13443 VDD.n4536 GND 3.47277f
C13444 VDD.n4537 GND 0.04648f
C13445 VDD.n4538 GND 0.05737f
C13446 VDD.n4539 GND 0.0171f
C13447 VDD.n4540 GND 0.064f
C13448 VDD.n4543 GND 0.06555f
C13449 VDD.n4544 GND 0.03083f
C13450 VDD.t174 GND 0.08047f
C13451 VDD.n4545 GND 0.03534f
C13452 VDD.t953 GND 0.15471f
C13453 VDD.n4546 GND 0.03238f
C13454 VDD.n4547 GND 0.02607f
C13455 VDD.n4548 GND 0.09595f
C13456 VDD.t183 GND 0.08047f
C13457 VDD.n4549 GND 0.03534f
C13458 VDD.t945 GND 0.15471f
C13459 VDD.n4550 GND 0.03238f
C13460 VDD.n4551 GND 0.02607f
C13461 VDD.n4553 GND 0.24365f
C13462 VDD.n4554 GND 0.03483f
C13463 VDD.t820 GND 0.02116f
C13464 VDD.t797 GND 0.02116f
C13465 VDD.n4555 GND 0.09893f
C13466 VDD.n4556 GND 0.02854f
C13467 VDD.n4557 GND 0.02503f
C13468 VDD.n4558 GND 0.02503f
C13469 VDD.n4559 GND 0.04556f
C13470 VDD.n4560 GND 0.32569f
C13471 VDD.t819 GND 0.2823f
C13472 VDD.n4561 GND 0.04624f
C13473 VDD.n4562 GND 0.04624f
C13474 VDD.n4563 GND 0.08322f
C13475 VDD.t332 GND 0.3079f
C13476 VDD.n4564 GND 0.04624f
C13477 VDD.n4565 GND 0.04624f
C13478 VDD.t469 GND 0.02116f
C13479 VDD.t270 GND 0.02116f
C13480 VDD.n4566 GND 0.09893f
C13481 VDD.n4567 GND 0.02854f
C13482 VDD.n4568 GND 0.02503f
C13483 VDD.n4569 GND 0.02503f
C13484 VDD.n4570 GND 0.04556f
C13485 VDD.n4571 GND 0.32569f
C13486 VDD.t468 GND 0.3079f
C13487 VDD.n4572 GND 0.04624f
C13488 VDD.n4573 GND 0.04624f
C13489 VDD.t253 GND 0.02116f
C13490 VDD.t584 GND 0.02116f
C13491 VDD.n4574 GND 0.09893f
C13492 VDD.n4575 GND 0.02854f
C13493 VDD.n4576 GND 0.02503f
C13494 VDD.n4577 GND 0.02503f
C13495 VDD.n4578 GND 0.04556f
C13496 VDD.n4579 GND 0.32569f
C13497 VDD.t252 GND 0.2823f
C13498 VDD.n4580 GND 0.04624f
C13499 VDD.n4581 GND 0.04624f
C13500 VDD.n4582 GND 0.08322f
C13501 VDD.t585 GND 0.3079f
C13502 VDD.n4583 GND 0.04624f
C13503 VDD.n4584 GND 0.04624f
C13504 VDD.t889 GND 0.02116f
C13505 VDD.t704 GND 0.02116f
C13506 VDD.n4585 GND 0.09893f
C13507 VDD.n4586 GND 0.02854f
C13508 VDD.n4587 GND 0.02503f
C13509 VDD.n4588 GND 0.02503f
C13510 VDD.n4589 GND 0.04556f
C13511 VDD.n4590 GND 0.32569f
C13512 VDD.t888 GND 0.3079f
C13513 VDD.n4591 GND 0.04624f
C13514 VDD.n4592 GND 0.04624f
C13515 VDD.t293 GND 0.02116f
C13516 VDD.t599 GND 0.02116f
C13517 VDD.n4593 GND 0.09893f
C13518 VDD.n4594 GND 0.02854f
C13519 VDD.n4595 GND 0.02503f
C13520 VDD.n4596 GND 0.02503f
C13521 VDD.n4597 GND 0.04556f
C13522 VDD.n4598 GND 0.32569f
C13523 VDD.t292 GND 0.2823f
C13524 VDD.n4599 GND 0.04624f
C13525 VDD.n4600 GND 0.04624f
C13526 VDD.n4601 GND 0.08322f
C13527 VDD.t549 GND 0.3079f
C13528 VDD.n4602 GND 0.04624f
C13529 VDD.n4603 GND 0.04624f
C13530 VDD.t32 GND 0.02116f
C13531 VDD.t733 GND 0.02116f
C13532 VDD.n4604 GND 0.09893f
C13533 VDD.n4605 GND 0.02854f
C13534 VDD.n4606 GND 0.02503f
C13535 VDD.n4607 GND 0.02503f
C13536 VDD.n4608 GND 0.04556f
C13537 VDD.n4609 GND 0.32569f
C13538 VDD.t31 GND 0.3079f
C13539 VDD.n4610 GND 0.04624f
C13540 VDD.n4611 GND 0.04624f
C13541 VDD.t829 GND 0.02116f
C13542 VDD.t892 GND 0.02116f
C13543 VDD.n4612 GND 0.09893f
C13544 VDD.n4613 GND 0.02854f
C13545 VDD.n4614 GND 0.02503f
C13546 VDD.n4615 GND 0.02503f
C13547 VDD.n4616 GND 0.04556f
C13548 VDD.n4617 GND 0.32569f
C13549 VDD.t828 GND 0.2823f
C13550 VDD.n4618 GND 0.04624f
C13551 VDD.n4619 GND 0.04624f
C13552 VDD.n4620 GND 0.08322f
C13553 VDD.t526 GND 0.3079f
C13554 VDD.n4621 GND 0.04624f
C13555 VDD.n4622 GND 0.04624f
C13556 VDD.t60 GND 0.02116f
C13557 VDD.t455 GND 0.02116f
C13558 VDD.n4623 GND 0.09893f
C13559 VDD.n4624 GND 0.02854f
C13560 VDD.n4625 GND 0.02503f
C13561 VDD.n4626 GND 0.02503f
C13562 VDD.n4627 GND 0.04556f
C13563 VDD.n4628 GND 0.32569f
C13564 VDD.t59 GND 0.3079f
C13565 VDD.n4629 GND 0.04624f
C13566 VDD.n4630 GND 0.04624f
C13567 VDD.t745 GND 0.02116f
C13568 VDD.t595 GND 0.02116f
C13569 VDD.n4631 GND 0.09893f
C13570 VDD.n4632 GND 0.02854f
C13571 VDD.n4633 GND 0.02503f
C13572 VDD.n4634 GND 0.02503f
C13573 VDD.n4635 GND 0.04556f
C13574 VDD.n4636 GND 0.32569f
C13575 VDD.t744 GND 0.2823f
C13576 VDD.n4637 GND 0.04624f
C13577 VDD.n4638 GND 0.04624f
C13578 VDD.n4639 GND 0.08322f
C13579 VDD.t596 GND 0.3079f
C13580 VDD.n4640 GND 0.04624f
C13581 VDD.n4641 GND 0.04624f
C13582 VDD.t554 GND 0.02116f
C13583 VDD.t369 GND 0.02116f
C13584 VDD.n4642 GND 0.09893f
C13585 VDD.n4643 GND 0.02854f
C13586 VDD.n4644 GND 0.02503f
C13587 VDD.n4645 GND 0.02503f
C13588 VDD.n4646 GND 0.04556f
C13589 VDD.n4647 GND 0.32569f
C13590 VDD.t553 GND 0.3079f
C13591 VDD.n4648 GND 0.04624f
C13592 VDD.n4649 GND 0.04624f
C13593 VDD.t823 GND 0.02116f
C13594 VDD.t297 GND 0.02116f
C13595 VDD.n4650 GND 0.09893f
C13596 VDD.n4651 GND 0.02854f
C13597 VDD.n4652 GND 0.02503f
C13598 VDD.n4653 GND 0.02503f
C13599 VDD.n4654 GND 0.04556f
C13600 VDD.n4655 GND 0.32569f
C13601 VDD.t822 GND 0.2823f
C13602 VDD.n4656 GND 0.04624f
C13603 VDD.n4657 GND 0.04624f
C13604 VDD.n4658 GND 0.08322f
C13605 VDD.t645 GND 0.3079f
C13606 VDD.n4659 GND 0.04624f
C13607 VDD.n4660 GND 0.04624f
C13608 VDD.t88 GND 0.02116f
C13609 VDD.t795 GND 0.02116f
C13610 VDD.n4661 GND 0.09893f
C13611 VDD.n4662 GND 0.02854f
C13612 VDD.n4663 GND 0.02503f
C13613 VDD.n4664 GND 0.02503f
C13614 VDD.n4665 GND 0.04556f
C13615 VDD.n4666 GND 0.32569f
C13616 VDD.t87 GND 0.3079f
C13617 VDD.n4667 GND 0.04624f
C13618 VDD.n4668 GND 0.04624f
C13619 VDD.t225 GND 0.02116f
C13620 VDD.t423 GND 0.02116f
C13621 VDD.n4669 GND 0.09893f
C13622 VDD.n4670 GND 0.02854f
C13623 VDD.n4671 GND 0.02503f
C13624 VDD.n4672 GND 0.02503f
C13625 VDD.n4673 GND 0.04556f
C13626 VDD.n4674 GND 0.32569f
C13627 VDD.t224 GND 0.2823f
C13628 VDD.n4675 GND 0.04624f
C13629 VDD.n4676 GND 0.04624f
C13630 VDD.n4677 GND 0.08322f
C13631 VDD.t725 GND 0.3079f
C13632 VDD.n4678 GND 0.04624f
C13633 VDD.n4679 GND 0.04624f
C13634 VDD.t748 GND 0.02116f
C13635 VDD.t879 GND 0.02116f
C13636 VDD.n4680 GND 0.09893f
C13637 VDD.n4681 GND 0.02854f
C13638 VDD.n4682 GND 0.02503f
C13639 VDD.n4683 GND 0.02503f
C13640 VDD.n4684 GND 0.04556f
C13641 VDD.n4685 GND 0.32569f
C13642 VDD.t747 GND 0.3079f
C13643 VDD.n4686 GND 0.04624f
C13644 VDD.n4687 GND 0.04624f
C13645 VDD.t813 GND 0.02116f
C13646 VDD.t843 GND 0.02116f
C13647 VDD.n4688 GND 0.09893f
C13648 VDD.n4689 GND 0.02854f
C13649 VDD.n4690 GND 0.02503f
C13650 VDD.n4691 GND 0.02503f
C13651 VDD.n4692 GND 0.04556f
C13652 VDD.n4693 GND 0.32569f
C13653 VDD.t812 GND 0.2823f
C13654 VDD.n4694 GND 0.04624f
C13655 VDD.n4695 GND 0.04624f
C13656 VDD.n4696 GND 0.08322f
C13657 VDD.t869 GND 0.3079f
C13658 VDD.n4697 GND 0.04624f
C13659 VDD.n4698 GND 0.04624f
C13660 VDD.t341 GND 0.02116f
C13661 VDD.t572 GND 0.02116f
C13662 VDD.n4699 GND 0.09893f
C13663 VDD.n4700 GND 0.16564f
C13664 VDD.n4701 GND 0.02503f
C13665 VDD.n4702 GND 0.02503f
C13666 VDD.n4703 GND 0.04556f
C13667 VDD.n4704 GND 0.32569f
C13668 VDD.t340 GND 0.3079f
C13669 VDD.n4705 GND 0.04624f
C13670 VDD.n4706 GND 0.04624f
C13671 VDD.n4707 GND 0.13241f
C13672 VDD.n4709 GND 0.32569f
C13673 VDD.n4710 GND 0.02503f
C13674 VDD.n4711 GND 0.02704f
C13675 VDD.n4712 GND 0.02503f
C13676 VDD.n4713 GND 0.04556f
C13677 VDD.n4714 GND 0.22764f
C13678 VDD.n4715 GND 0.22764f
C13679 VDD.n4716 GND 0.02704f
C13680 VDD.n4717 GND 0.04624f
C13681 VDD.t571 GND 0.3079f
C13682 VDD.n4719 GND 0.04624f
C13683 VDD.n4720 GND 0.08322f
C13684 VDD.n4721 GND 0.02127f
C13685 VDD.t870 GND 0.02128f
C13686 VDD.n4722 GND 0.02127f
C13687 VDD.n4723 GND 0.06662f
C13688 VDD.n4724 GND 0.09943f
C13689 VDD.n4725 GND 0.08322f
C13690 VDD.n4727 GND 0.32569f
C13691 VDD.n4728 GND 0.02503f
C13692 VDD.n4729 GND 0.02704f
C13693 VDD.n4730 GND 0.02503f
C13694 VDD.n4731 GND 0.04556f
C13695 VDD.n4732 GND 0.30573f
C13696 VDD.n4733 GND 0.30573f
C13697 VDD.n4734 GND 0.04556f
C13698 VDD.n4735 GND 0.02503f
C13699 VDD.n4736 GND 0.02704f
C13700 VDD.n4737 GND 0.02503f
C13701 VDD.n4738 GND 0.04556f
C13702 VDD.n4739 GND 0.22764f
C13703 VDD.n4740 GND 0.22764f
C13704 VDD.n4741 GND 0.02704f
C13705 VDD.n4742 GND 0.04624f
C13706 VDD.t842 GND 0.3079f
C13707 VDD.n4744 GND 0.04624f
C13708 VDD.n4745 GND 0.08322f
C13709 VDD.n4746 GND 0.02127f
C13710 VDD.n4747 GND 0.10432f
C13711 VDD.n4748 GND 0.08322f
C13712 VDD.n4750 GND 0.32569f
C13713 VDD.n4751 GND 0.02503f
C13714 VDD.n4752 GND 0.02704f
C13715 VDD.n4753 GND 0.02503f
C13716 VDD.n4754 GND 0.04556f
C13717 VDD.n4755 GND 0.22764f
C13718 VDD.n4756 GND 0.22764f
C13719 VDD.n4757 GND 0.02704f
C13720 VDD.n4758 GND 0.04624f
C13721 VDD.t878 GND 0.3079f
C13722 VDD.n4760 GND 0.04624f
C13723 VDD.n4761 GND 0.08322f
C13724 VDD.n4762 GND 0.02127f
C13725 VDD.t726 GND 0.02128f
C13726 VDD.n4763 GND 0.02127f
C13727 VDD.n4764 GND 0.06662f
C13728 VDD.n4765 GND 0.09943f
C13729 VDD.n4766 GND 0.08322f
C13730 VDD.n4768 GND 0.32569f
C13731 VDD.n4769 GND 0.02503f
C13732 VDD.n4770 GND 0.02704f
C13733 VDD.n4771 GND 0.02503f
C13734 VDD.n4772 GND 0.04556f
C13735 VDD.n4773 GND 0.30573f
C13736 VDD.n4774 GND 0.30573f
C13737 VDD.n4775 GND 0.04556f
C13738 VDD.n4776 GND 0.02503f
C13739 VDD.n4777 GND 0.02704f
C13740 VDD.n4778 GND 0.02503f
C13741 VDD.n4779 GND 0.04556f
C13742 VDD.n4780 GND 0.22764f
C13743 VDD.n4781 GND 0.22764f
C13744 VDD.n4782 GND 0.02704f
C13745 VDD.n4783 GND 0.04624f
C13746 VDD.t422 GND 0.3079f
C13747 VDD.n4785 GND 0.04624f
C13748 VDD.n4786 GND 0.08322f
C13749 VDD.n4787 GND 0.02127f
C13750 VDD.n4788 GND 0.10432f
C13751 VDD.n4789 GND 0.08322f
C13752 VDD.n4791 GND 0.32569f
C13753 VDD.n4792 GND 0.02503f
C13754 VDD.n4793 GND 0.02704f
C13755 VDD.n4794 GND 0.02503f
C13756 VDD.n4795 GND 0.04556f
C13757 VDD.n4796 GND 0.22764f
C13758 VDD.n4797 GND 0.22764f
C13759 VDD.n4798 GND 0.02704f
C13760 VDD.n4799 GND 0.04624f
C13761 VDD.t794 GND 0.3079f
C13762 VDD.n4801 GND 0.04624f
C13763 VDD.n4802 GND 0.08322f
C13764 VDD.n4803 GND 0.02127f
C13765 VDD.t646 GND 0.02128f
C13766 VDD.n4804 GND 0.02127f
C13767 VDD.n4805 GND 0.06662f
C13768 VDD.n4806 GND 0.09943f
C13769 VDD.n4807 GND 0.08322f
C13770 VDD.n4809 GND 0.32569f
C13771 VDD.n4810 GND 0.02503f
C13772 VDD.n4811 GND 0.02704f
C13773 VDD.n4812 GND 0.02503f
C13774 VDD.n4813 GND 0.04556f
C13775 VDD.n4814 GND 0.30573f
C13776 VDD.n4815 GND 0.30573f
C13777 VDD.n4816 GND 0.04556f
C13778 VDD.n4817 GND 0.02503f
C13779 VDD.n4818 GND 0.02704f
C13780 VDD.n4819 GND 0.02503f
C13781 VDD.n4820 GND 0.04556f
C13782 VDD.n4821 GND 0.22764f
C13783 VDD.n4822 GND 0.22764f
C13784 VDD.n4823 GND 0.02704f
C13785 VDD.n4824 GND 0.04624f
C13786 VDD.t296 GND 0.3079f
C13787 VDD.n4826 GND 0.04624f
C13788 VDD.n4827 GND 0.08322f
C13789 VDD.n4828 GND 0.02127f
C13790 VDD.n4829 GND 0.10432f
C13791 VDD.n4830 GND 0.08322f
C13792 VDD.n4832 GND 0.32569f
C13793 VDD.n4833 GND 0.02503f
C13794 VDD.n4834 GND 0.02704f
C13795 VDD.n4835 GND 0.02503f
C13796 VDD.n4836 GND 0.04556f
C13797 VDD.n4837 GND 0.22764f
C13798 VDD.n4838 GND 0.22764f
C13799 VDD.n4839 GND 0.02704f
C13800 VDD.n4840 GND 0.04624f
C13801 VDD.t368 GND 0.3079f
C13802 VDD.n4842 GND 0.04624f
C13803 VDD.n4843 GND 0.08322f
C13804 VDD.n4844 GND 0.02127f
C13805 VDD.t597 GND 0.02128f
C13806 VDD.n4845 GND 0.02127f
C13807 VDD.n4846 GND 0.06662f
C13808 VDD.n4847 GND 0.09943f
C13809 VDD.n4848 GND 0.08322f
C13810 VDD.n4850 GND 0.32569f
C13811 VDD.n4851 GND 0.02503f
C13812 VDD.n4852 GND 0.02704f
C13813 VDD.n4853 GND 0.02503f
C13814 VDD.n4854 GND 0.04556f
C13815 VDD.n4855 GND 0.30573f
C13816 VDD.n4856 GND 0.30573f
C13817 VDD.n4857 GND 0.04556f
C13818 VDD.n4858 GND 0.02503f
C13819 VDD.n4859 GND 0.02704f
C13820 VDD.n4860 GND 0.02503f
C13821 VDD.n4861 GND 0.04556f
C13822 VDD.n4862 GND 0.22764f
C13823 VDD.n4863 GND 0.22764f
C13824 VDD.n4864 GND 0.02704f
C13825 VDD.n4865 GND 0.04624f
C13826 VDD.t594 GND 0.3079f
C13827 VDD.n4867 GND 0.04624f
C13828 VDD.n4868 GND 0.08322f
C13829 VDD.n4869 GND 0.02127f
C13830 VDD.n4870 GND 0.10432f
C13831 VDD.n4871 GND 0.08322f
C13832 VDD.n4873 GND 0.32569f
C13833 VDD.n4874 GND 0.02503f
C13834 VDD.n4875 GND 0.02704f
C13835 VDD.n4876 GND 0.02503f
C13836 VDD.n4877 GND 0.04556f
C13837 VDD.n4878 GND 0.22764f
C13838 VDD.n4879 GND 0.22764f
C13839 VDD.n4880 GND 0.02704f
C13840 VDD.n4881 GND 0.04624f
C13841 VDD.t454 GND 0.3079f
C13842 VDD.n4883 GND 0.04624f
C13843 VDD.n4884 GND 0.08322f
C13844 VDD.n4885 GND 0.02127f
C13845 VDD.t527 GND 0.02128f
C13846 VDD.n4886 GND 0.02127f
C13847 VDD.n4887 GND 0.06662f
C13848 VDD.n4888 GND 0.09943f
C13849 VDD.n4889 GND 0.08322f
C13850 VDD.n4891 GND 0.32569f
C13851 VDD.n4892 GND 0.02503f
C13852 VDD.n4893 GND 0.02704f
C13853 VDD.n4894 GND 0.02503f
C13854 VDD.n4895 GND 0.04556f
C13855 VDD.n4896 GND 0.30573f
C13856 VDD.n4897 GND 0.30573f
C13857 VDD.n4898 GND 0.04556f
C13858 VDD.n4899 GND 0.02503f
C13859 VDD.n4900 GND 0.02704f
C13860 VDD.n4901 GND 0.02503f
C13861 VDD.n4902 GND 0.04556f
C13862 VDD.n4903 GND 0.22764f
C13863 VDD.n4904 GND 0.22764f
C13864 VDD.n4905 GND 0.02704f
C13865 VDD.n4906 GND 0.04624f
C13866 VDD.t891 GND 0.3079f
C13867 VDD.n4908 GND 0.04624f
C13868 VDD.n4909 GND 0.08322f
C13869 VDD.n4910 GND 0.02127f
C13870 VDD.n4911 GND 0.10432f
C13871 VDD.n4912 GND 0.08322f
C13872 VDD.n4914 GND 0.32569f
C13873 VDD.n4915 GND 0.02503f
C13874 VDD.n4916 GND 0.02704f
C13875 VDD.n4917 GND 0.02503f
C13876 VDD.n4918 GND 0.04556f
C13877 VDD.n4919 GND 0.22764f
C13878 VDD.n4920 GND 0.22764f
C13879 VDD.n4921 GND 0.02704f
C13880 VDD.n4922 GND 0.04624f
C13881 VDD.t732 GND 0.3079f
C13882 VDD.n4924 GND 0.04624f
C13883 VDD.n4925 GND 0.08322f
C13884 VDD.n4926 GND 0.02127f
C13885 VDD.t550 GND 0.02128f
C13886 VDD.n4927 GND 0.02127f
C13887 VDD.n4928 GND 0.06662f
C13888 VDD.n4929 GND 0.09943f
C13889 VDD.n4930 GND 0.08322f
C13890 VDD.n4932 GND 0.32569f
C13891 VDD.n4933 GND 0.02503f
C13892 VDD.n4934 GND 0.02704f
C13893 VDD.n4935 GND 0.02503f
C13894 VDD.n4936 GND 0.04556f
C13895 VDD.n4937 GND 0.30573f
C13896 VDD.n4938 GND 0.30573f
C13897 VDD.n4939 GND 0.04556f
C13898 VDD.n4940 GND 0.02503f
C13899 VDD.n4941 GND 0.02704f
C13900 VDD.n4942 GND 0.02503f
C13901 VDD.n4943 GND 0.04556f
C13902 VDD.n4944 GND 0.22764f
C13903 VDD.n4945 GND 0.22764f
C13904 VDD.n4946 GND 0.02704f
C13905 VDD.n4947 GND 0.04624f
C13906 VDD.t598 GND 0.3079f
C13907 VDD.n4949 GND 0.04624f
C13908 VDD.n4950 GND 0.08322f
C13909 VDD.n4951 GND 0.02127f
C13910 VDD.n4952 GND 0.10432f
C13911 VDD.n4953 GND 0.08322f
C13912 VDD.n4955 GND 0.32569f
C13913 VDD.n4956 GND 0.02503f
C13914 VDD.n4957 GND 0.02704f
C13915 VDD.n4958 GND 0.02503f
C13916 VDD.n4959 GND 0.04556f
C13917 VDD.n4960 GND 0.22764f
C13918 VDD.n4961 GND 0.22764f
C13919 VDD.n4962 GND 0.02704f
C13920 VDD.n4963 GND 0.04624f
C13921 VDD.t703 GND 0.3079f
C13922 VDD.n4965 GND 0.04624f
C13923 VDD.n4966 GND 0.08322f
C13924 VDD.n4967 GND 0.02127f
C13925 VDD.t586 GND 0.02128f
C13926 VDD.n4968 GND 0.02127f
C13927 VDD.n4969 GND 0.06662f
C13928 VDD.n4970 GND 0.09943f
C13929 VDD.n4971 GND 0.08322f
C13930 VDD.n4973 GND 0.32569f
C13931 VDD.n4974 GND 0.02503f
C13932 VDD.n4975 GND 0.02704f
C13933 VDD.n4976 GND 0.02503f
C13934 VDD.n4977 GND 0.04556f
C13935 VDD.n4978 GND 0.30573f
C13936 VDD.n4979 GND 0.30573f
C13937 VDD.n4980 GND 0.04556f
C13938 VDD.n4981 GND 0.02503f
C13939 VDD.n4982 GND 0.02704f
C13940 VDD.n4983 GND 0.02503f
C13941 VDD.n4984 GND 0.04556f
C13942 VDD.n4985 GND 0.22764f
C13943 VDD.n4986 GND 0.22764f
C13944 VDD.n4987 GND 0.02704f
C13945 VDD.n4988 GND 0.04624f
C13946 VDD.t583 GND 0.3079f
C13947 VDD.n4990 GND 0.04624f
C13948 VDD.n4991 GND 0.08322f
C13949 VDD.n4992 GND 0.02127f
C13950 VDD.n4993 GND 0.10432f
C13951 VDD.n4994 GND 0.08322f
C13952 VDD.n4996 GND 0.32569f
C13953 VDD.n4997 GND 0.02503f
C13954 VDD.n4998 GND 0.02704f
C13955 VDD.n4999 GND 0.02503f
C13956 VDD.n5000 GND 0.04556f
C13957 VDD.n5001 GND 0.22764f
C13958 VDD.n5002 GND 0.22764f
C13959 VDD.n5003 GND 0.02704f
C13960 VDD.n5004 GND 0.04624f
C13961 VDD.t269 GND 0.3079f
C13962 VDD.n5006 GND 0.04624f
C13963 VDD.n5007 GND 0.08322f
C13964 VDD.n5008 GND 0.02127f
C13965 VDD.t333 GND 0.02128f
C13966 VDD.n5009 GND 0.02127f
C13967 VDD.n5010 GND 0.06662f
C13968 VDD.n5011 GND 0.09943f
C13969 VDD.n5012 GND 0.08322f
C13970 VDD.n5014 GND 0.32569f
C13971 VDD.n5015 GND 0.02503f
C13972 VDD.n5016 GND 0.02704f
C13973 VDD.n5017 GND 0.02503f
C13974 VDD.n5018 GND 0.04556f
C13975 VDD.n5019 GND 0.30573f
C13976 VDD.n5020 GND 0.30573f
C13977 VDD.n5021 GND 0.04556f
C13978 VDD.n5022 GND 0.02503f
C13979 VDD.n5023 GND 0.02704f
C13980 VDD.n5024 GND 0.02503f
C13981 VDD.n5025 GND 0.04556f
C13982 VDD.n5026 GND 0.22764f
C13983 VDD.n5027 GND 0.22764f
C13984 VDD.n5028 GND 0.02704f
C13985 VDD.n5029 GND 0.04624f
C13986 VDD.t796 GND 0.3079f
C13987 VDD.n5031 GND 0.04624f
C13988 VDD.n5032 GND 0.08322f
C13989 VDD.n5033 GND 0.02127f
C13990 VDD.n5034 GND 0.88136f
C13991 VDD.t756 GND 0.02128f
C13992 VDD.n5035 GND 0.02503f
C13993 VDD.n5036 GND 0.04624f
C13994 VDD.n5037 GND 0.02704f
C13995 VDD.n5038 GND 0.04624f
C13996 VDD.t643 GND 0.57933f
C13997 VDD.n5039 GND 0.04556f
C13998 VDD.n5040 GND 0.04624f
C13999 VDD.n5041 GND 0.04624f
C14000 VDD.n5042 GND 0.02704f
C14001 VDD.n5043 GND 0.02299f
C14002 VDD.n5044 GND 0.04885f
C14003 VDD.t644 GND 0.02128f
C14004 VDD.t913 GND 0.02128f
C14005 VDD.n5045 GND 0.12159f
C14006 VDD.n5046 GND 0.02396f
C14007 VDD.n5047 GND 0.04624f
C14008 VDD.n5048 GND 0.02704f
C14009 VDD.n5049 GND 0.02299f
C14010 VDD.t628 GND 0.57933f
C14011 VDD.n5050 GND 0.04556f
C14012 VDD.n5051 GND 0.04624f
C14013 VDD.n5052 GND 0.04624f
C14014 VDD.n5053 GND 0.02704f
C14015 VDD.n5054 GND 0.02299f
C14016 VDD.n5055 GND 0.04885f
C14017 VDD.n5056 GND 0.02885f
C14018 VDD.n5057 GND 0.04624f
C14019 VDD.n5058 GND 0.02704f
C14020 VDD.n5059 GND 0.02299f
C14021 VDD.t611 GND 0.57933f
C14022 VDD.n5060 GND 0.04556f
C14023 VDD.n5061 GND 0.04624f
C14024 VDD.n5062 GND 0.04624f
C14025 VDD.n5063 GND 0.02704f
C14026 VDD.n5064 GND 0.02299f
C14027 VDD.n5065 GND 0.04885f
C14028 VDD.t612 GND 0.02116f
C14029 VDD.t759 GND 0.02116f
C14030 VDD.n5066 GND 0.09893f
C14031 VDD.t613 GND 0.02116f
C14032 VDD.t629 GND 0.02116f
C14033 VDD.n5067 GND 0.09893f
C14034 VDD.n5068 GND 0.03784f
C14035 VDD.n5069 GND 0.02127f
C14036 VDD.n5070 GND 0.04624f
C14037 VDD.n5071 GND 0.02704f
C14038 VDD.n5072 GND 0.02299f
C14039 VDD.t408 GND 0.57933f
C14040 VDD.n5073 GND 0.04556f
C14041 VDD.n5074 GND 0.04624f
C14042 VDD.n5075 GND 0.04624f
C14043 VDD.n5076 GND 0.02704f
C14044 VDD.n5077 GND 0.02299f
C14045 VDD.n5078 GND 0.04885f
C14046 VDD.t409 GND 0.02128f
C14047 VDD.t476 GND 0.02128f
C14048 VDD.n5079 GND 0.12159f
C14049 VDD.n5080 GND 0.02396f
C14050 VDD.n5081 GND 0.04624f
C14051 VDD.n5082 GND 0.02704f
C14052 VDD.n5083 GND 0.02299f
C14053 VDD.t62 GND 0.57933f
C14054 VDD.n5084 GND 0.04556f
C14055 VDD.n5085 GND 0.04624f
C14056 VDD.n5086 GND 0.04624f
C14057 VDD.n5087 GND 0.02704f
C14058 VDD.n5088 GND 0.02299f
C14059 VDD.n5089 GND 0.04885f
C14060 VDD.n5090 GND 0.02885f
C14061 VDD.n5091 GND 0.04624f
C14062 VDD.n5092 GND 0.02704f
C14063 VDD.n5093 GND 0.02299f
C14064 VDD.t303 GND 0.57933f
C14065 VDD.n5094 GND 0.04556f
C14066 VDD.n5095 GND 0.04624f
C14067 VDD.n5096 GND 0.04624f
C14068 VDD.n5097 GND 0.02704f
C14069 VDD.n5098 GND 0.02299f
C14070 VDD.n5099 GND 0.04885f
C14071 VDD.t617 GND 0.02116f
C14072 VDD.t63 GND 0.02116f
C14073 VDD.n5100 GND 0.09893f
C14074 VDD.t304 GND 0.02116f
C14075 VDD.t558 GND 0.02116f
C14076 VDD.n5101 GND 0.09893f
C14077 VDD.n5102 GND 0.03784f
C14078 VDD.n5103 GND 0.02127f
C14079 VDD.n5104 GND 0.04624f
C14080 VDD.n5105 GND 0.02704f
C14081 VDD.n5106 GND 0.02299f
C14082 VDD.t614 GND 0.57933f
C14083 VDD.n5107 GND 0.04624f
C14084 VDD.n5108 GND 0.04624f
C14085 VDD.n5109 GND 0.08322f
C14086 VDD.t222 GND 0.57933f
C14087 VDD.n5110 GND 0.04556f
C14088 VDD.n5111 GND 0.04624f
C14089 VDD.n5112 GND 0.04624f
C14090 VDD.n5113 GND 0.02704f
C14091 VDD.n5114 GND 0.02299f
C14092 VDD.n5115 GND 0.04885f
C14093 VDD.t615 GND 0.02128f
C14094 VDD.n5116 GND 0.06662f
C14095 VDD.n5117 GND 0.01638f
C14096 VDD.n5118 GND 0.02127f
C14097 VDD.n5119 GND 0.04624f
C14098 VDD.n5120 GND 0.02704f
C14099 VDD.n5121 GND 0.02299f
C14100 VDD.t529 GND 0.57933f
C14101 VDD.n5122 GND 0.04556f
C14102 VDD.n5123 GND 0.04624f
C14103 VDD.n5124 GND 0.04624f
C14104 VDD.n5125 GND 0.02704f
C14105 VDD.n5126 GND 0.02299f
C14106 VDD.n5127 GND 0.04885f
C14107 VDD.t530 GND 0.02116f
C14108 VDD.t330 GND 0.02116f
C14109 VDD.n5128 GND 0.09893f
C14110 VDD.t531 GND 0.02116f
C14111 VDD.t223 GND 0.02116f
C14112 VDD.n5129 GND 0.09893f
C14113 VDD.n5130 GND 0.03784f
C14114 VDD.n5131 GND 0.02127f
C14115 VDD.n5132 GND 0.04624f
C14116 VDD.n5133 GND 0.02704f
C14117 VDD.n5134 GND 0.02299f
C14118 VDD.t763 GND 0.57933f
C14119 VDD.n5135 GND 0.04556f
C14120 VDD.n5136 GND 0.04624f
C14121 VDD.n5137 GND 0.04624f
C14122 VDD.n5138 GND 0.02704f
C14123 VDD.n5139 GND 0.02299f
C14124 VDD.n5140 GND 0.04885f
C14125 VDD.t914 GND 0.02128f
C14126 VDD.t764 GND 0.02128f
C14127 VDD.n5141 GND 0.12159f
C14128 VDD.n5142 GND 0.02396f
C14129 VDD.n5143 GND 0.04624f
C14130 VDD.n5144 GND 0.02704f
C14131 VDD.n5145 GND 0.02299f
C14132 VDD.t506 GND 0.57933f
C14133 VDD.n5146 GND 0.04556f
C14134 VDD.n5147 GND 0.04624f
C14135 VDD.n5148 GND 0.04624f
C14136 VDD.n5149 GND 0.02704f
C14137 VDD.n5150 GND 0.02299f
C14138 VDD.n5151 GND 0.04885f
C14139 VDD.n5152 GND 0.02885f
C14140 VDD.n5153 GND 0.04624f
C14141 VDD.n5154 GND 0.02704f
C14142 VDD.n5155 GND 0.02299f
C14143 VDD.t425 GND 0.57933f
C14144 VDD.n5156 GND 0.04556f
C14145 VDD.n5157 GND 0.04624f
C14146 VDD.n5158 GND 0.04624f
C14147 VDD.n5159 GND 0.02704f
C14148 VDD.n5160 GND 0.02299f
C14149 VDD.n5161 GND 0.04885f
C14150 VDD.t426 GND 0.02116f
C14151 VDD.t507 GND 0.02116f
C14152 VDD.n5162 GND 0.09893f
C14153 VDD.t772 GND 0.02116f
C14154 VDD.t578 GND 0.02116f
C14155 VDD.n5163 GND 0.09893f
C14156 VDD.n5164 GND 0.03784f
C14157 VDD.n5165 GND 0.02127f
C14158 VDD.n5166 GND 0.04624f
C14159 VDD.n5167 GND 0.02704f
C14160 VDD.n5168 GND 0.02299f
C14161 VDD.t452 GND 0.57933f
C14162 VDD.n5169 GND 0.04624f
C14163 VDD.n5170 GND 0.04624f
C14164 VDD.n5171 GND 0.02704f
C14165 VDD.n5172 GND 0.02503f
C14166 VDD.t767 GND 0.02128f
C14167 VDD.t479 GND 0.02128f
C14168 VDD.n5173 GND 0.02885f
C14169 VDD.n5174 GND 0.04885f
C14170 VDD.n5175 GND 0.04624f
C14171 VDD.n5176 GND 0.04885f
C14172 VDD.n5177 GND 0.04556f
C14173 VDD.n5178 GND 0.04556f
C14174 VDD.t487 GND 0.57933f
C14175 VDD.n5179 GND 0.04556f
C14176 VDD.n5180 GND 0.04624f
C14177 VDD.n5181 GND 0.04624f
C14178 VDD.n5182 GND 0.02704f
C14179 VDD.n5183 GND 0.02299f
C14180 VDD.n5184 GND 0.04885f
C14181 VDD.n5185 GND 0.04624f
C14182 VDD.n5186 GND 0.02704f
C14183 VDD.n5187 GND 0.02299f
C14184 VDD.t343 GND 0.57933f
C14185 VDD.n5188 GND 0.04556f
C14186 VDD.n5189 GND 0.04624f
C14187 VDD.n5190 GND 0.04624f
C14188 VDD.n5191 GND 0.02704f
C14189 VDD.n5192 GND 0.02299f
C14190 VDD.n5193 GND 0.04885f
C14191 VDD.t344 GND 0.02116f
C14192 VDD.t722 GND 0.02116f
C14193 VDD.n5194 GND 0.09893f
C14194 VDD.t375 GND 0.02116f
C14195 VDD.t488 GND 0.02116f
C14196 VDD.n5195 GND 0.09893f
C14197 VDD.n5196 GND 0.03784f
C14198 VDD.n5197 GND 0.02127f
C14199 VDD.n5198 GND 0.04624f
C14200 VDD.n5199 GND 0.02704f
C14201 VDD.n5200 GND 0.02299f
C14202 VDD.t566 GND 0.57933f
C14203 VDD.n5201 GND 0.04556f
C14204 VDD.n5202 GND 0.04624f
C14205 VDD.n5203 GND 0.04624f
C14206 VDD.n5204 GND 0.02704f
C14207 VDD.n5205 GND 0.02299f
C14208 VDD.n5206 GND 0.04885f
C14209 VDD.t705 GND 0.02128f
C14210 VDD.t567 GND 0.02128f
C14211 VDD.n5207 GND 0.12159f
C14212 VDD.n5208 GND 0.02396f
C14213 VDD.n5209 GND 0.04624f
C14214 VDD.n5210 GND 0.02704f
C14215 VDD.n5211 GND 0.02299f
C14216 VDD.t335 GND 0.57933f
C14217 VDD.n5212 GND 0.04556f
C14218 VDD.n5213 GND 0.04624f
C14219 VDD.n5214 GND 0.04624f
C14220 VDD.n5215 GND 0.02704f
C14221 VDD.n5216 GND 0.02299f
C14222 VDD.n5217 GND 0.04885f
C14223 VDD.n5218 GND 0.02885f
C14224 VDD.n5219 GND 0.04624f
C14225 VDD.n5220 GND 0.02704f
C14226 VDD.n5221 GND 0.02299f
C14227 VDD.t261 GND 0.57933f
C14228 VDD.n5222 GND 0.04556f
C14229 VDD.n5223 GND 0.04624f
C14230 VDD.n5224 GND 0.04624f
C14231 VDD.n5225 GND 0.02704f
C14232 VDD.n5226 GND 0.02299f
C14233 VDD.n5227 GND 0.04885f
C14234 VDD.t394 GND 0.02116f
C14235 VDD.t336 GND 0.02116f
C14236 VDD.n5228 GND 0.09893f
C14237 VDD.t262 GND 0.02116f
C14238 VDD.t877 GND 0.02116f
C14239 VDD.n5229 GND 0.09893f
C14240 VDD.n5230 GND 0.03784f
C14241 VDD.n5231 GND 0.02127f
C14242 VDD.n5232 GND 0.04624f
C14243 VDD.n5233 GND 0.02704f
C14244 VDD.n5234 GND 0.02299f
C14245 VDD.t376 GND 0.57933f
C14246 VDD.n5235 GND 0.04624f
C14247 VDD.n5236 GND 0.04624f
C14248 VDD.n5237 GND 0.08322f
C14249 VDD.t501 GND 0.57933f
C14250 VDD.n5238 GND 0.04556f
C14251 VDD.n5239 GND 0.04624f
C14252 VDD.n5240 GND 0.04624f
C14253 VDD.n5241 GND 0.02704f
C14254 VDD.n5242 GND 0.02299f
C14255 VDD.n5243 GND 0.04885f
C14256 VDD.t377 GND 0.02128f
C14257 VDD.n5244 GND 0.06662f
C14258 VDD.n5245 GND 0.01638f
C14259 VDD.n5246 GND 0.02127f
C14260 VDD.n5247 GND 0.04624f
C14261 VDD.n5248 GND 0.02704f
C14262 VDD.n5249 GND 0.02299f
C14263 VDD.t442 GND 0.57933f
C14264 VDD.n5250 GND 0.04556f
C14265 VDD.n5251 GND 0.04624f
C14266 VDD.n5252 GND 0.04624f
C14267 VDD.n5253 GND 0.02704f
C14268 VDD.n5254 GND 0.02299f
C14269 VDD.n5255 GND 0.04885f
C14270 VDD.t444 GND 0.02116f
C14271 VDD.t502 GND 0.02116f
C14272 VDD.n5256 GND 0.09893f
C14273 VDD.t443 GND 0.02116f
C14274 VDD.t782 GND 0.02116f
C14275 VDD.n5257 GND 0.09893f
C14276 VDD.n5258 GND 0.03784f
C14277 VDD.n5259 GND 0.02127f
C14278 VDD.n5260 GND 0.04624f
C14279 VDD.n5261 GND 0.02704f
C14280 VDD.n5262 GND 0.02299f
C14281 VDD.t90 GND 0.57933f
C14282 VDD.n5263 GND 0.04556f
C14283 VDD.n5264 GND 0.04624f
C14284 VDD.n5265 GND 0.04624f
C14285 VDD.n5266 GND 0.02704f
C14286 VDD.n5267 GND 0.02299f
C14287 VDD.n5268 GND 0.04885f
C14288 VDD.t91 GND 0.02128f
C14289 VDD.t392 GND 0.02128f
C14290 VDD.n5269 GND 0.12159f
C14291 VDD.n5270 GND 0.02396f
C14292 VDD.n5271 GND 0.04624f
C14293 VDD.n5272 GND 0.02704f
C14294 VDD.n5273 GND 0.02299f
C14295 VDD.t418 GND 0.57933f
C14296 VDD.n5274 GND 0.04556f
C14297 VDD.n5275 GND 0.04624f
C14298 VDD.n5276 GND 0.04624f
C14299 VDD.n5277 GND 0.02704f
C14300 VDD.n5278 GND 0.02299f
C14301 VDD.n5279 GND 0.04885f
C14302 VDD.n5280 GND 0.02885f
C14303 VDD.n5281 GND 0.04624f
C14304 VDD.n5282 GND 0.02704f
C14305 VDD.n5283 GND 0.02299f
C14306 VDD.t308 GND 0.57933f
C14307 VDD.n5284 GND 0.04556f
C14308 VDD.n5285 GND 0.04624f
C14309 VDD.n5286 GND 0.04624f
C14310 VDD.n5287 GND 0.02704f
C14311 VDD.n5288 GND 0.02299f
C14312 VDD.n5289 GND 0.04885f
C14313 VDD.t309 GND 0.02116f
C14314 VDD.t902 GND 0.02116f
C14315 VDD.n5290 GND 0.09893f
C14316 VDD.t449 GND 0.02116f
C14317 VDD.t419 GND 0.02116f
C14318 VDD.n5291 GND 0.09893f
C14319 VDD.n5292 GND 0.03784f
C14320 VDD.n5293 GND 0.02127f
C14321 VDD.n5294 GND 0.04624f
C14322 VDD.n5295 GND 0.02704f
C14323 VDD.n5296 GND 0.02299f
C14324 VDD.t275 GND 0.57933f
C14325 VDD.n5297 GND 0.04624f
C14326 VDD.n5298 GND 0.04624f
C14327 VDD.n5299 GND 0.02704f
C14328 VDD.n5300 GND 0.02503f
C14329 VDD.t565 GND 0.02128f
C14330 VDD.t494 GND 0.02128f
C14331 VDD.n5301 GND 0.02885f
C14332 VDD.n5302 GND 0.04885f
C14333 VDD.n5303 GND 0.04624f
C14334 VDD.n5304 GND 0.04885f
C14335 VDD.n5305 GND 0.04556f
C14336 VDD.n5306 GND 0.04556f
C14337 VDD.t94 GND 0.57933f
C14338 VDD.n5307 GND 0.04556f
C14339 VDD.n5308 GND 0.04624f
C14340 VDD.n5309 GND 0.04624f
C14341 VDD.n5310 GND 0.02704f
C14342 VDD.n5311 GND 0.02299f
C14343 VDD.n5312 GND 0.04885f
C14344 VDD.n5313 GND 0.04624f
C14345 VDD.n5314 GND 0.02704f
C14346 VDD.n5315 GND 0.02299f
C14347 VDD.t482 GND 0.57933f
C14348 VDD.n5316 GND 0.04556f
C14349 VDD.n5317 GND 0.04624f
C14350 VDD.n5318 GND 0.04624f
C14351 VDD.n5319 GND 0.02704f
C14352 VDD.n5320 GND 0.02299f
C14353 VDD.n5321 GND 0.04885f
C14354 VDD.t483 GND 0.02116f
C14355 VDD.t758 GND 0.02116f
C14356 VDD.n5322 GND 0.09893f
C14357 VDD.t484 GND 0.02116f
C14358 VDD.t95 GND 0.02116f
C14359 VDD.n5323 GND 0.09893f
C14360 VDD.n5324 GND 0.03784f
C14361 VDD.n5325 GND 0.02127f
C14362 VDD.n5326 GND 0.04624f
C14363 VDD.n5327 GND 0.02704f
C14364 VDD.n5328 GND 0.02299f
C14365 VDD.t358 GND 0.57933f
C14366 VDD.n5329 GND 0.04556f
C14367 VDD.n5330 GND 0.04624f
C14368 VDD.n5331 GND 0.04624f
C14369 VDD.n5332 GND 0.02704f
C14370 VDD.n5333 GND 0.02299f
C14371 VDD.n5334 GND 0.04885f
C14372 VDD.t590 GND 0.02128f
C14373 VDD.t359 GND 0.02128f
C14374 VDD.n5335 GND 0.12159f
C14375 VDD.n5336 GND 0.02396f
C14376 VDD.n5337 GND 0.04624f
C14377 VDD.n5338 GND 0.02704f
C14378 VDD.n5339 GND 0.02299f
C14379 VDD.t604 GND 0.57933f
C14380 VDD.n5340 GND 0.04556f
C14381 VDD.n5341 GND 0.04624f
C14382 VDD.n5342 GND 0.04624f
C14383 VDD.n5343 GND 0.02704f
C14384 VDD.n5344 GND 0.02299f
C14385 VDD.n5345 GND 0.04885f
C14386 VDD.n5346 GND 0.02885f
C14387 VDD.n5347 GND 0.04624f
C14388 VDD.n5348 GND 0.02704f
C14389 VDD.n5349 GND 0.02299f
C14390 VDD.t74 GND 0.57933f
C14391 VDD.n5350 GND 0.04556f
C14392 VDD.n5351 GND 0.04624f
C14393 VDD.n5352 GND 0.04624f
C14394 VDD.n5353 GND 0.02704f
C14395 VDD.n5354 GND 0.02299f
C14396 VDD.n5355 GND 0.04885f
C14397 VDD.t826 GND 0.02116f
C14398 VDD.t770 GND 0.02116f
C14399 VDD.n5356 GND 0.09893f
C14400 VDD.t75 GND 0.02116f
C14401 VDD.t605 GND 0.02116f
C14402 VDD.n5357 GND 0.09893f
C14403 VDD.n5358 GND 0.03784f
C14404 VDD.n5359 GND 0.02127f
C14405 VDD.n5360 GND 0.04624f
C14406 VDD.n5361 GND 0.02704f
C14407 VDD.n5362 GND 0.02299f
C14408 VDD.t485 GND 0.57933f
C14409 VDD.n5363 GND 0.04624f
C14410 VDD.n5364 GND 0.04624f
C14411 VDD.n5365 GND 0.08322f
C14412 VDD.t215 GND 0.57933f
C14413 VDD.n5366 GND 0.04556f
C14414 VDD.n5367 GND 0.04624f
C14415 VDD.n5368 GND 0.04624f
C14416 VDD.n5369 GND 0.02704f
C14417 VDD.n5370 GND 0.02299f
C14418 VDD.n5371 GND 0.04885f
C14419 VDD.t486 GND 0.02128f
C14420 VDD.n5372 GND 0.06662f
C14421 VDD.n5373 GND 0.01638f
C14422 VDD.n5374 GND 0.02127f
C14423 VDD.n5375 GND 0.04624f
C14424 VDD.n5376 GND 0.02704f
C14425 VDD.n5377 GND 0.02299f
C14426 VDD.t439 GND 0.57933f
C14427 VDD.n5378 GND 0.04556f
C14428 VDD.n5379 GND 0.04624f
C14429 VDD.n5380 GND 0.04624f
C14430 VDD.n5381 GND 0.02704f
C14431 VDD.n5382 GND 0.02299f
C14432 VDD.n5383 GND 0.04885f
C14433 VDD.t441 GND 0.02116f
C14434 VDD.t216 GND 0.02116f
C14435 VDD.n5384 GND 0.09893f
C14436 VDD.t440 GND 0.02116f
C14437 VDD.t827 GND 0.02116f
C14438 VDD.n5385 GND 0.09893f
C14439 VDD.n5386 GND 0.03784f
C14440 VDD.n5387 GND 0.02127f
C14441 VDD.n5388 GND 0.04624f
C14442 VDD.n5389 GND 0.02704f
C14443 VDD.n5390 GND 0.02299f
C14444 VDD.t568 GND 0.57933f
C14445 VDD.n5391 GND 0.04556f
C14446 VDD.n5392 GND 0.04624f
C14447 VDD.n5393 GND 0.04624f
C14448 VDD.n5394 GND 0.02704f
C14449 VDD.n5395 GND 0.02299f
C14450 VDD.n5396 GND 0.04885f
C14451 VDD.t731 GND 0.02128f
C14452 VDD.t569 GND 0.02128f
C14453 VDD.n5397 GND 0.12159f
C14454 VDD.n5398 GND 0.02396f
C14455 VDD.n5399 GND 0.04624f
C14456 VDD.n5400 GND 0.02704f
C14457 VDD.n5401 GND 0.02299f
C14458 VDD.t287 GND 0.57933f
C14459 VDD.n5402 GND 0.04556f
C14460 VDD.n5403 GND 0.04624f
C14461 VDD.n5404 GND 0.04624f
C14462 VDD.n5405 GND 0.02704f
C14463 VDD.n5406 GND 0.02299f
C14464 VDD.n5407 GND 0.04885f
C14465 VDD.n5408 GND 0.02885f
C14466 VDD.n5409 GND 0.04624f
C14467 VDD.n5410 GND 0.02704f
C14468 VDD.n5411 GND 0.02299f
C14469 VDD.t411 GND 0.57933f
C14470 VDD.n5412 GND 0.04556f
C14471 VDD.n5413 GND 0.04624f
C14472 VDD.n5414 GND 0.04624f
C14473 VDD.n5415 GND 0.02704f
C14474 VDD.n5416 GND 0.02299f
C14475 VDD.n5417 GND 0.04885f
C14476 VDD.t412 GND 0.02116f
C14477 VDD.t499 GND 0.02116f
C14478 VDD.n5418 GND 0.09893f
C14479 VDD.t854 GND 0.02116f
C14480 VDD.t288 GND 0.02116f
C14481 VDD.n5419 GND 0.09893f
C14482 VDD.n5420 GND 0.03784f
C14483 VDD.n5421 GND 0.02127f
C14484 VDD.n5422 GND 0.04624f
C14485 VDD.n5423 GND 0.02704f
C14486 VDD.n5424 GND 0.02299f
C14487 VDD.t718 GND 0.57933f
C14488 VDD.n5425 GND 0.04624f
C14489 VDD.n5426 GND 0.04624f
C14490 VDD.n5427 GND 0.02704f
C14491 VDD.n5428 GND 0.02503f
C14492 VDD.t560 GND 0.02128f
C14493 VDD.t365 GND 0.02128f
C14494 VDD.n5429 GND 0.02885f
C14495 VDD.n5430 GND 0.04885f
C14496 VDD.n5431 GND 0.04624f
C14497 VDD.n5432 GND 0.04885f
C14498 VDD.n5433 GND 0.04556f
C14499 VDD.n5434 GND 0.04556f
C14500 VDD.t68 GND 0.57933f
C14501 VDD.n5435 GND 0.04556f
C14502 VDD.n5436 GND 0.04624f
C14503 VDD.n5437 GND 0.04624f
C14504 VDD.n5438 GND 0.02704f
C14505 VDD.n5439 GND 0.02299f
C14506 VDD.n5440 GND 0.04885f
C14507 VDD.n5441 GND 0.04624f
C14508 VDD.n5442 GND 0.02704f
C14509 VDD.n5443 GND 0.02299f
C14510 VDD.t37 GND 0.57933f
C14511 VDD.n5444 GND 0.04556f
C14512 VDD.n5445 GND 0.04624f
C14513 VDD.n5446 GND 0.04624f
C14514 VDD.n5447 GND 0.02704f
C14515 VDD.n5448 GND 0.02299f
C14516 VDD.n5449 GND 0.04885f
C14517 VDD.t38 GND 0.02116f
C14518 VDD.t757 GND 0.02116f
C14519 VDD.n5450 GND 0.09893f
C14520 VDD.t39 GND 0.02116f
C14521 VDD.t69 GND 0.02116f
C14522 VDD.n5451 GND 0.09893f
C14523 VDD.n5452 GND 0.03784f
C14524 VDD.n5453 GND 0.02127f
C14525 VDD.n5454 GND 0.04624f
C14526 VDD.n5455 GND 0.02704f
C14527 VDD.n5456 GND 0.02299f
C14528 VDD.t352 GND 0.57933f
C14529 VDD.n5457 GND 0.04556f
C14530 VDD.n5458 GND 0.04624f
C14531 VDD.n5459 GND 0.04624f
C14532 VDD.n5460 GND 0.02704f
C14533 VDD.n5461 GND 0.02299f
C14534 VDD.n5462 GND 0.04885f
C14535 VDD.t353 GND 0.02128f
C14536 VDD.t898 GND 0.02128f
C14537 VDD.n5463 GND 0.12159f
C14538 VDD.n5464 GND 0.02396f
C14539 VDD.n5465 GND 0.04624f
C14540 VDD.n5466 GND 0.02704f
C14541 VDD.n5467 GND 0.02299f
C14542 VDD.t465 GND 0.57933f
C14543 VDD.n5468 GND 0.04556f
C14544 VDD.n5469 GND 0.04624f
C14545 VDD.n5470 GND 0.04624f
C14546 VDD.n5471 GND 0.02704f
C14547 VDD.n5472 GND 0.02299f
C14548 VDD.n5473 GND 0.04885f
C14549 VDD.n5474 GND 0.02885f
C14550 VDD.n5475 GND 0.04624f
C14551 VDD.n5476 GND 0.02704f
C14552 VDD.n5477 GND 0.02299f
C14553 VDD.t420 GND 0.57933f
C14554 VDD.n5478 GND 0.04556f
C14555 VDD.n5479 GND 0.04624f
C14556 VDD.n5480 GND 0.04624f
C14557 VDD.n5481 GND 0.02704f
C14558 VDD.n5482 GND 0.02299f
C14559 VDD.n5483 GND 0.04885f
C14560 VDD.t737 GND 0.02116f
C14561 VDD.t922 GND 0.02116f
C14562 VDD.n5484 GND 0.09893f
C14563 VDD.t421 GND 0.02116f
C14564 VDD.t466 GND 0.02116f
C14565 VDD.n5485 GND 0.09893f
C14566 VDD.n5486 GND 0.03784f
C14567 VDD.n5487 GND 0.02127f
C14568 VDD.n5488 GND 0.04624f
C14569 VDD.n5489 GND 0.02704f
C14570 VDD.n5490 GND 0.02299f
C14571 VDD.t40 GND 0.57933f
C14572 VDD.n5491 GND 0.04624f
C14573 VDD.n5492 GND 0.04624f
C14574 VDD.n5493 GND 0.08322f
C14575 VDD.t306 GND 0.57933f
C14576 VDD.n5494 GND 0.04556f
C14577 VDD.n5495 GND 0.04624f
C14578 VDD.n5496 GND 0.04624f
C14579 VDD.n5497 GND 0.02704f
C14580 VDD.n5498 GND 0.02299f
C14581 VDD.n5499 GND 0.04885f
C14582 VDD.t41 GND 0.02128f
C14583 VDD.n5500 GND 0.06662f
C14584 VDD.n5501 GND 0.01638f
C14585 VDD.n5502 GND 0.02127f
C14586 VDD.n5503 GND 0.04624f
C14587 VDD.n5504 GND 0.02704f
C14588 VDD.n5505 GND 0.02299f
C14589 VDD.t625 GND 0.57933f
C14590 VDD.n5506 GND 0.04556f
C14591 VDD.n5507 GND 0.04624f
C14592 VDD.n5508 GND 0.04624f
C14593 VDD.n5509 GND 0.02704f
C14594 VDD.n5510 GND 0.02299f
C14595 VDD.n5511 GND 0.04885f
C14596 VDD.t627 GND 0.02116f
C14597 VDD.t307 GND 0.02116f
C14598 VDD.n5512 GND 0.09893f
C14599 VDD.t626 GND 0.02116f
C14600 VDD.t738 GND 0.02116f
C14601 VDD.n5513 GND 0.09893f
C14602 VDD.n5514 GND 0.03784f
C14603 VDD.n5515 GND 0.02127f
C14604 VDD.n5516 GND 0.04624f
C14605 VDD.n5517 GND 0.02704f
C14606 VDD.n5518 GND 0.02299f
C14607 VDD.t635 GND 0.57933f
C14608 VDD.n5519 GND 0.04556f
C14609 VDD.n5520 GND 0.04624f
C14610 VDD.n5521 GND 0.04624f
C14611 VDD.n5522 GND 0.02704f
C14612 VDD.n5523 GND 0.02299f
C14613 VDD.n5524 GND 0.04885f
C14614 VDD.t788 GND 0.02128f
C14615 VDD.t636 GND 0.02128f
C14616 VDD.n5525 GND 0.12159f
C14617 VDD.n5526 GND 0.02396f
C14618 VDD.n5527 GND 0.04624f
C14619 VDD.n5528 GND 0.02704f
C14620 VDD.n5529 GND 0.02299f
C14621 VDD.t400 GND 0.57933f
C14622 VDD.n5530 GND 0.04556f
C14623 VDD.n5531 GND 0.04624f
C14624 VDD.n5532 GND 0.04624f
C14625 VDD.n5533 GND 0.02704f
C14626 VDD.n5534 GND 0.02299f
C14627 VDD.n5535 GND 0.04885f
C14628 VDD.n5536 GND 0.02885f
C14629 VDD.n5537 GND 0.04624f
C14630 VDD.n5538 GND 0.02704f
C14631 VDD.n5539 GND 0.02299f
C14632 VDD.t70 GND 0.57933f
C14633 VDD.n5540 GND 0.04556f
C14634 VDD.n5541 GND 0.04624f
C14635 VDD.n5542 GND 0.04624f
C14636 VDD.n5543 GND 0.02704f
C14637 VDD.n5544 GND 0.02299f
C14638 VDD.n5545 GND 0.04885f
C14639 VDD.t71 GND 0.02116f
C14640 VDD.t438 GND 0.02116f
C14641 VDD.n5546 GND 0.09893f
C14642 VDD.t300 GND 0.02116f
C14643 VDD.t401 GND 0.02116f
C14644 VDD.n5547 GND 0.09893f
C14645 VDD.n5548 GND 0.03784f
C14646 VDD.n5549 GND 0.02127f
C14647 VDD.n5550 GND 0.04624f
C14648 VDD.n5551 GND 0.02704f
C14649 VDD.n5552 GND 0.02299f
C14650 VDD.t16 GND 0.57933f
C14651 VDD.n5553 GND 0.04624f
C14652 VDD.n5554 GND 0.04624f
C14653 VDD.n5555 GND 0.02704f
C14654 VDD.n5556 GND 0.02503f
C14655 VDD.t564 GND 0.02128f
C14656 VDD.t754 GND 0.02128f
C14657 VDD.n5557 GND 0.02885f
C14658 VDD.n5558 GND 0.04885f
C14659 VDD.n5559 GND 0.04624f
C14660 VDD.n5560 GND 0.04885f
C14661 VDD.n5561 GND 0.04556f
C14662 VDD.n5562 GND 0.04556f
C14663 VDD.t18 GND 0.57933f
C14664 VDD.n5563 GND 0.04556f
C14665 VDD.n5564 GND 0.04624f
C14666 VDD.n5565 GND 0.04624f
C14667 VDD.n5566 GND 0.02704f
C14668 VDD.n5567 GND 0.02299f
C14669 VDD.n5568 GND 0.04885f
C14670 VDD.n5569 GND 0.04624f
C14671 VDD.n5570 GND 0.02704f
C14672 VDD.n5571 GND 0.02299f
C14673 VDD.t257 GND 0.57933f
C14674 VDD.n5572 GND 0.04556f
C14675 VDD.n5573 GND 0.04624f
C14676 VDD.n5574 GND 0.04624f
C14677 VDD.n5575 GND 0.02704f
C14678 VDD.n5576 GND 0.02299f
C14679 VDD.n5577 GND 0.04885f
C14680 VDD.t901 GND 0.02116f
C14681 VDD.t19 GND 0.02116f
C14682 VDD.n5578 GND 0.09893f
C14683 VDD.t258 GND 0.02116f
C14684 VDD.t576 GND 0.02116f
C14685 VDD.n5579 GND 0.09893f
C14686 VDD.n5580 GND 0.03784f
C14687 VDD.n5581 GND 0.02127f
C14688 VDD.n5582 GND 0.04624f
C14689 VDD.n5583 GND 0.02704f
C14690 VDD.n5584 GND 0.02299f
C14691 VDD.t637 GND 0.57933f
C14692 VDD.n5585 GND 0.04556f
C14693 VDD.n5586 GND 0.04624f
C14694 VDD.n5587 GND 0.04624f
C14695 VDD.n5588 GND 0.02704f
C14696 VDD.n5589 GND 0.02299f
C14697 VDD.n5590 GND 0.04885f
C14698 VDD.t752 GND 0.02128f
C14699 VDD.t638 GND 0.02128f
C14700 VDD.n5591 GND 0.12159f
C14701 VDD.n5592 GND 0.02396f
C14702 VDD.n5593 GND 0.04624f
C14703 VDD.n5594 GND 0.02704f
C14704 VDD.n5595 GND 0.02299f
C14705 VDD.t78 GND 0.57933f
C14706 VDD.n5596 GND 0.04556f
C14707 VDD.n5597 GND 0.04624f
C14708 VDD.n5598 GND 0.04624f
C14709 VDD.n5599 GND 0.02704f
C14710 VDD.n5600 GND 0.02299f
C14711 VDD.n5601 GND 0.04885f
C14712 VDD.n5602 GND 0.02885f
C14713 VDD.n5603 GND 0.04624f
C14714 VDD.n5604 GND 0.02704f
C14715 VDD.n5605 GND 0.02299f
C14716 VDD.t428 GND 0.57933f
C14717 VDD.n5606 GND 0.04556f
C14718 VDD.n5607 GND 0.04624f
C14719 VDD.n5608 GND 0.04624f
C14720 VDD.n5609 GND 0.02704f
C14721 VDD.n5610 GND 0.02299f
C14722 VDD.n5611 GND 0.04885f
C14723 VDD.t429 GND 0.02116f
C14724 VDD.t79 GND 0.02116f
C14725 VDD.n5612 GND 0.09893f
C14726 VDD.t432 GND 0.02116f
C14727 VDD.t528 GND 0.02116f
C14728 VDD.n5613 GND 0.09893f
C14729 VDD.n5614 GND 0.03784f
C14730 VDD.n5615 GND 0.02127f
C14731 VDD.n5616 GND 0.04624f
C14732 VDD.n5617 GND 0.02704f
C14733 VDD.n5618 GND 0.02299f
C14734 VDD.t899 GND 0.57933f
C14735 VDD.n5619 GND 0.04624f
C14736 VDD.n5620 GND 0.04624f
C14737 VDD.n5621 GND 0.08322f
C14738 VDD.t430 GND 0.57933f
C14739 VDD.n5622 GND 0.04556f
C14740 VDD.n5623 GND 0.04624f
C14741 VDD.n5624 GND 0.04624f
C14742 VDD.n5625 GND 0.02704f
C14743 VDD.n5626 GND 0.02299f
C14744 VDD.n5627 GND 0.04885f
C14745 VDD.t900 GND 0.02128f
C14746 VDD.n5628 GND 0.06662f
C14747 VDD.n5629 GND 0.01638f
C14748 VDD.n5630 GND 0.02127f
C14749 VDD.n5631 GND 0.04624f
C14750 VDD.n5632 GND 0.02704f
C14751 VDD.n5633 GND 0.02299f
C14752 VDD.t503 GND 0.57933f
C14753 VDD.n5634 GND 0.04556f
C14754 VDD.n5635 GND 0.04624f
C14755 VDD.n5636 GND 0.04624f
C14756 VDD.n5637 GND 0.02704f
C14757 VDD.n5638 GND 0.02299f
C14758 VDD.n5639 GND 0.04885f
C14759 VDD.t505 GND 0.02116f
C14760 VDD.t610 GND 0.02116f
C14761 VDD.n5640 GND 0.09893f
C14762 VDD.t504 GND 0.02116f
C14763 VDD.t431 GND 0.02116f
C14764 VDD.n5641 GND 0.09893f
C14765 VDD.n5642 GND 0.03784f
C14766 VDD.n5643 GND 0.02127f
C14767 VDD.n5644 GND 0.04624f
C14768 VDD.n5645 GND 0.02704f
C14769 VDD.n5646 GND 0.02299f
C14770 VDD.t639 GND 0.57933f
C14771 VDD.n5647 GND 0.04556f
C14772 VDD.n5648 GND 0.04624f
C14773 VDD.n5649 GND 0.04624f
C14774 VDD.n5650 GND 0.02704f
C14775 VDD.n5651 GND 0.02299f
C14776 VDD.n5652 GND 0.04885f
C14777 VDD.t753 GND 0.02128f
C14778 VDD.t640 GND 0.02128f
C14779 VDD.n5653 GND 0.12159f
C14780 VDD.n5654 GND 0.02396f
C14781 VDD.n5655 GND 0.04624f
C14782 VDD.n5656 GND 0.02704f
C14783 VDD.n5657 GND 0.02299f
C14784 VDD.t347 GND 0.57933f
C14785 VDD.n5658 GND 0.04556f
C14786 VDD.n5659 GND 0.04624f
C14787 VDD.n5660 GND 0.04624f
C14788 VDD.n5661 GND 0.02704f
C14789 VDD.n5662 GND 0.02299f
C14790 VDD.n5663 GND 0.04885f
C14791 VDD.n5664 GND 0.02885f
C14792 VDD.n5665 GND 0.04624f
C14793 VDD.n5666 GND 0.02704f
C14794 VDD.n5667 GND 0.02299f
C14795 VDD.t495 GND 0.57933f
C14796 VDD.n5668 GND 0.04556f
C14797 VDD.n5669 GND 0.04624f
C14798 VDD.n5670 GND 0.04624f
C14799 VDD.n5671 GND 0.02704f
C14800 VDD.n5672 GND 0.02299f
C14801 VDD.n5673 GND 0.04885f
C14802 VDD.t496 GND 0.02116f
C14803 VDD.t348 GND 0.02116f
C14804 VDD.n5674 GND 0.09893f
C14805 VDD.t712 GND 0.02116f
C14806 VDD.t577 GND 0.02116f
C14807 VDD.n5675 GND 0.09893f
C14808 VDD.n5676 GND 0.03784f
C14809 VDD.n5677 GND 0.02127f
C14810 VDD.n5678 GND 0.04624f
C14811 VDD.n5679 GND 0.02704f
C14812 VDD.n5680 GND 0.02299f
C14813 VDD.t450 GND 0.57933f
C14814 VDD.n5681 GND 0.04624f
C14815 VDD.n5682 GND 0.04624f
C14816 VDD.n5683 GND 0.02704f
C14817 VDD.n5684 GND 0.02503f
C14818 VDD.t765 GND 0.02128f
C14819 VDD.t286 GND 0.02128f
C14820 VDD.n5685 GND 0.02885f
C14821 VDD.n5686 GND 0.04885f
C14822 VDD.n5687 GND 0.04624f
C14823 VDD.n5688 GND 0.04885f
C14824 VDD.n5689 GND 0.04556f
C14825 VDD.n5690 GND 0.04556f
C14826 VDD.t277 GND 0.57933f
C14827 VDD.n5691 GND 0.04556f
C14828 VDD.n5692 GND 0.04624f
C14829 VDD.n5693 GND 0.04624f
C14830 VDD.n5694 GND 0.02704f
C14831 VDD.n5695 GND 0.02299f
C14832 VDD.n5696 GND 0.04885f
C14833 VDD.n5697 GND 0.04624f
C14834 VDD.n5698 GND 0.02704f
C14835 VDD.n5699 GND 0.02299f
C14836 VDD.t862 GND 0.57933f
C14837 VDD.n5700 GND 0.04556f
C14838 VDD.n5701 GND 0.04624f
C14839 VDD.n5702 GND 0.04624f
C14840 VDD.n5703 GND 0.02704f
C14841 VDD.n5704 GND 0.02299f
C14842 VDD.n5705 GND 0.04885f
C14843 VDD.t863 GND 0.02116f
C14844 VDD.t278 GND 0.02116f
C14845 VDD.n5706 GND 0.09893f
C14846 VDD.t864 GND 0.02116f
C14847 VDD.t424 GND 0.02116f
C14848 VDD.n5707 GND 0.09893f
C14849 VDD.n5708 GND 0.03784f
C14850 VDD.n5709 GND 0.02127f
C14851 VDD.n5710 GND 0.04624f
C14852 VDD.n5711 GND 0.02704f
C14853 VDD.n5712 GND 0.02299f
C14854 VDD.t561 GND 0.57933f
C14855 VDD.n5713 GND 0.04556f
C14856 VDD.n5714 GND 0.04624f
C14857 VDD.n5715 GND 0.04624f
C14858 VDD.n5716 GND 0.02704f
C14859 VDD.n5717 GND 0.02299f
C14860 VDD.n5718 GND 0.04885f
C14861 VDD.t792 GND 0.02128f
C14862 VDD.t562 GND 0.02128f
C14863 VDD.n5719 GND 0.12159f
C14864 VDD.n5720 GND 0.02396f
C14865 VDD.n5721 GND 0.04624f
C14866 VDD.n5722 GND 0.02704f
C14867 VDD.n5723 GND 0.02299f
C14868 VDD.t349 GND 0.57933f
C14869 VDD.n5724 GND 0.04556f
C14870 VDD.n5725 GND 0.04624f
C14871 VDD.n5726 GND 0.04624f
C14872 VDD.n5727 GND 0.02704f
C14873 VDD.n5728 GND 0.02299f
C14874 VDD.n5729 GND 0.04885f
C14875 VDD.n5730 GND 0.02885f
C14876 VDD.n5731 GND 0.04624f
C14877 VDD.n5732 GND 0.02704f
C14878 VDD.n5733 GND 0.02299f
C14879 VDD.t2 GND 0.57933f
C14880 VDD.n5734 GND 0.04556f
C14881 VDD.n5735 GND 0.04624f
C14882 VDD.n5736 GND 0.04624f
C14883 VDD.n5737 GND 0.02704f
C14884 VDD.n5738 GND 0.02299f
C14885 VDD.n5739 GND 0.04885f
C14886 VDD.t535 GND 0.02116f
C14887 VDD.t350 GND 0.02116f
C14888 VDD.n5740 GND 0.09893f
C14889 VDD.t3 GND 0.02116f
C14890 VDD.t701 GND 0.02116f
C14891 VDD.n5741 GND 0.09893f
C14892 VDD.n5742 GND 0.03784f
C14893 VDD.n5743 GND 0.02127f
C14894 VDD.n5744 GND 0.04624f
C14895 VDD.n5745 GND 0.02704f
C14896 VDD.n5746 GND 0.02299f
C14897 VDD.t735 GND 0.57933f
C14898 VDD.n5747 GND 0.04624f
C14899 VDD.n5748 GND 0.04624f
C14900 VDD.n5749 GND 0.08322f
C14901 VDD.t0 GND 0.57933f
C14902 VDD.n5750 GND 0.04556f
C14903 VDD.n5751 GND 0.04624f
C14904 VDD.n5752 GND 0.04624f
C14905 VDD.n5753 GND 0.02704f
C14906 VDD.n5754 GND 0.02299f
C14907 VDD.n5755 GND 0.04885f
C14908 VDD.t736 GND 0.02128f
C14909 VDD.n5756 GND 0.06662f
C14910 VDD.n5757 GND 0.01638f
C14911 VDD.n5758 GND 0.02127f
C14912 VDD.n5759 GND 0.04624f
C14913 VDD.n5760 GND 0.02704f
C14914 VDD.n5761 GND 0.02299f
C14915 VDD.t64 GND 0.57933f
C14916 VDD.n5762 GND 0.04556f
C14917 VDD.n5763 GND 0.04624f
C14918 VDD.n5764 GND 0.04624f
C14919 VDD.n5765 GND 0.02704f
C14920 VDD.n5766 GND 0.02299f
C14921 VDD.n5767 GND 0.04885f
C14922 VDD.t66 GND 0.02116f
C14923 VDD.t1 GND 0.02116f
C14924 VDD.n5768 GND 0.09893f
C14925 VDD.t65 GND 0.02116f
C14926 VDD.t534 GND 0.02116f
C14927 VDD.n5769 GND 0.09893f
C14928 VDD.n5770 GND 0.03784f
C14929 VDD.n5771 GND 0.02127f
C14930 VDD.n5772 GND 0.04624f
C14931 VDD.n5773 GND 0.02704f
C14932 VDD.n5774 GND 0.02299f
C14933 VDD.t390 GND 0.57933f
C14934 VDD.n5775 GND 0.04556f
C14935 VDD.n5776 GND 0.04624f
C14936 VDD.n5777 GND 0.04624f
C14937 VDD.n5778 GND 0.02704f
C14938 VDD.n5779 GND 0.02299f
C14939 VDD.n5780 GND 0.04885f
C14940 VDD.t739 GND 0.02128f
C14941 VDD.t391 GND 0.02128f
C14942 VDD.n5781 GND 0.12159f
C14943 VDD.n5782 GND 0.02396f
C14944 VDD.n5783 GND 0.04624f
C14945 VDD.n5784 GND 0.02704f
C14946 VDD.n5785 GND 0.02299f
C14947 VDD.t804 GND 0.57933f
C14948 VDD.n5786 GND 0.04556f
C14949 VDD.n5787 GND 0.04624f
C14950 VDD.n5788 GND 0.04624f
C14951 VDD.n5789 GND 0.02704f
C14952 VDD.n5790 GND 0.02299f
C14953 VDD.n5791 GND 0.04885f
C14954 VDD.n5792 GND 0.02885f
C14955 VDD.n5793 GND 0.04624f
C14956 VDD.n5794 GND 0.02704f
C14957 VDD.n5795 GND 0.02299f
C14958 VDD.t385 GND 0.57933f
C14959 VDD.n5796 GND 0.04556f
C14960 VDD.n5797 GND 0.04624f
C14961 VDD.n5798 GND 0.04624f
C14962 VDD.n5799 GND 0.02704f
C14963 VDD.n5800 GND 0.02299f
C14964 VDD.n5801 GND 0.04885f
C14965 VDD.t847 GND 0.02116f
C14966 VDD.t805 GND 0.02116f
C14967 VDD.n5802 GND 0.09893f
C14968 VDD.t386 GND 0.02116f
C14969 VDD.t875 GND 0.02116f
C14970 VDD.n5803 GND 0.09893f
C14971 VDD.n5804 GND 0.03784f
C14972 VDD.n5805 GND 0.02127f
C14973 VDD.n5806 GND 0.04624f
C14974 VDD.n5807 GND 0.02704f
C14975 VDD.n5808 GND 0.02299f
C14976 VDD.t720 GND 0.57933f
C14977 VDD.n5809 GND 0.04624f
C14978 VDD.n5810 GND 0.04624f
C14979 VDD.n5811 GND 0.02704f
C14980 VDD.n5812 GND 0.02503f
C14981 VDD.t570 GND 0.02128f
C14982 VDD.t537 GND 0.02128f
C14983 VDD.n5813 GND 0.02885f
C14984 VDD.n5814 GND 0.04885f
C14985 VDD.n5815 GND 0.04624f
C14986 VDD.n5816 GND 0.04885f
C14987 VDD.n5817 GND 0.04556f
C14988 VDD.n5818 GND 0.04556f
C14989 VDD.t542 GND 0.57933f
C14990 VDD.n5819 GND 0.04556f
C14991 VDD.n5820 GND 0.04624f
C14992 VDD.n5821 GND 0.04624f
C14993 VDD.n5822 GND 0.02704f
C14994 VDD.n5823 GND 0.02299f
C14995 VDD.n5824 GND 0.04885f
C14996 VDD.n5825 GND 0.04624f
C14997 VDD.n5826 GND 0.02704f
C14998 VDD.n5827 GND 0.02299f
C14999 VDD.t836 GND 0.57933f
C15000 VDD.n5828 GND 0.04556f
C15001 VDD.n5829 GND 0.04624f
C15002 VDD.n5830 GND 0.04624f
C15003 VDD.n5831 GND 0.02704f
C15004 VDD.n5832 GND 0.02299f
C15005 VDD.n5833 GND 0.04885f
C15006 VDD.t837 GND 0.02116f
C15007 VDD.t760 GND 0.02116f
C15008 VDD.n5834 GND 0.09893f
C15009 VDD.t838 GND 0.02116f
C15010 VDD.t543 GND 0.02116f
C15011 VDD.n5835 GND 0.09893f
C15012 VDD.n5836 GND 0.03784f
C15013 VDD.n5837 GND 0.02127f
C15014 VDD.n5838 GND 0.04624f
C15015 VDD.n5839 GND 0.02704f
C15016 VDD.n5840 GND 0.02299f
C15017 VDD.t538 GND 0.57933f
C15018 VDD.n5841 GND 0.04556f
C15019 VDD.n5842 GND 0.04624f
C15020 VDD.n5843 GND 0.04624f
C15021 VDD.n5844 GND 0.02704f
C15022 VDD.n5845 GND 0.02299f
C15023 VDD.n5846 GND 0.04885f
C15024 VDD.t539 GND 0.02128f
C15025 VDD.t766 GND 0.02128f
C15026 VDD.n5847 GND 0.12159f
C15027 VDD.n5848 GND 0.02396f
C15028 VDD.n5849 GND 0.04624f
C15029 VDD.n5850 GND 0.02704f
C15030 VDD.n5851 GND 0.02299f
C15031 VDD.t547 GND 0.57933f
C15032 VDD.n5852 GND 0.04556f
C15033 VDD.n5853 GND 0.04624f
C15034 VDD.n5854 GND 0.04624f
C15035 VDD.n5855 GND 0.02704f
C15036 VDD.n5856 GND 0.02299f
C15037 VDD.n5857 GND 0.04885f
C15038 VDD.n5858 GND 0.02885f
C15039 VDD.n5859 GND 0.04624f
C15040 VDD.n5860 GND 0.02704f
C15041 VDD.n5861 GND 0.02299f
C15042 VDD.t280 GND 0.57933f
C15043 VDD.n5862 GND 0.04556f
C15044 VDD.n5863 GND 0.04624f
C15045 VDD.n5864 GND 0.04624f
C15046 VDD.n5865 GND 0.02704f
C15047 VDD.n5866 GND 0.02299f
C15048 VDD.n5867 GND 0.04885f
C15049 VDD.t281 GND 0.02116f
C15050 VDD.t548 GND 0.02116f
C15051 VDD.n5868 GND 0.09893f
C15052 VDD.t457 GND 0.02116f
C15053 VDD.t573 GND 0.02116f
C15054 VDD.n5869 GND 0.09893f
C15055 VDD.n5870 GND 0.03784f
C15056 VDD.n5871 GND 0.02127f
C15057 VDD.n5872 GND 0.04624f
C15058 VDD.n5873 GND 0.02704f
C15059 VDD.n5874 GND 0.02299f
C15060 VDD.t839 GND 0.57933f
C15061 VDD.n5875 GND 0.04624f
C15062 VDD.n5876 GND 0.04624f
C15063 VDD.n5877 GND 0.08322f
C15064 VDD.t282 GND 0.57933f
C15065 VDD.n5878 GND 0.04556f
C15066 VDD.n5879 GND 0.04624f
C15067 VDD.n5880 GND 0.04624f
C15068 VDD.n5881 GND 0.02704f
C15069 VDD.n5882 GND 0.02299f
C15070 VDD.n5883 GND 0.04885f
C15071 VDD.t840 GND 0.02128f
C15072 VDD.n5884 GND 0.06662f
C15073 VDD.n5885 GND 0.01638f
C15074 VDD.n5886 GND 0.02127f
C15075 VDD.n5887 GND 0.04624f
C15076 VDD.n5888 GND 0.02704f
C15077 VDD.n5889 GND 0.02299f
C15078 VDD.t395 GND 0.57933f
C15079 VDD.n5890 GND 0.04556f
C15080 VDD.n5891 GND 0.04624f
C15081 VDD.n5892 GND 0.04624f
C15082 VDD.n5893 GND 0.02704f
C15083 VDD.n5894 GND 0.02299f
C15084 VDD.n5895 GND 0.04885f
C15085 VDD.t397 GND 0.02116f
C15086 VDD.t574 GND 0.02116f
C15087 VDD.n5896 GND 0.09893f
C15088 VDD.t396 GND 0.02116f
C15089 VDD.t283 GND 0.02116f
C15090 VDD.n5897 GND 0.09893f
C15091 VDD.n5898 GND 0.03784f
C15092 VDD.n5899 GND 0.02127f
C15093 VDD.n5900 GND 0.04624f
C15094 VDD.n5901 GND 0.02704f
C15095 VDD.n5902 GND 0.02299f
C15096 VDD.t540 GND 0.57933f
C15097 VDD.n5903 GND 0.04556f
C15098 VDD.n5904 GND 0.04624f
C15099 VDD.n5905 GND 0.04624f
C15100 VDD.n5906 GND 0.02704f
C15101 VDD.n5907 GND 0.02299f
C15102 VDD.n5908 GND 0.04885f
C15103 VDD.t541 GND 0.02128f
C15104 VDD.t559 GND 0.02128f
C15105 VDD.n5909 GND 0.12159f
C15106 VDD.n5910 GND 0.02396f
C15107 VDD.n5911 GND 0.04624f
C15108 VDD.n5912 GND 0.02704f
C15109 VDD.n5913 GND 0.02299f
C15110 VDD.t81 GND 0.57933f
C15111 VDD.n5914 GND 0.04556f
C15112 VDD.n5915 GND 0.04624f
C15113 VDD.n5916 GND 0.04624f
C15114 VDD.n5917 GND 0.02704f
C15115 VDD.n5918 GND 0.02299f
C15116 VDD.n5919 GND 0.04885f
C15117 VDD.n5920 GND 0.02885f
C15118 VDD.n5921 GND 0.04624f
C15119 VDD.n5922 GND 0.02704f
C15120 VDD.n5923 GND 0.02299f
C15121 VDD.t27 GND 0.57933f
C15122 VDD.n5924 GND 0.04556f
C15123 VDD.n5925 GND 0.04624f
C15124 VDD.n5926 GND 0.04624f
C15125 VDD.n5927 GND 0.02704f
C15126 VDD.n5928 GND 0.02299f
C15127 VDD.n5929 GND 0.04885f
C15128 VDD.t477 GND 0.02116f
C15129 VDD.t532 GND 0.02116f
C15130 VDD.n5930 GND 0.09893f
C15131 VDD.t28 GND 0.02116f
C15132 VDD.t82 GND 0.02116f
C15133 VDD.n5931 GND 0.09893f
C15134 VDD.n5932 GND 0.03784f
C15135 VDD.n5933 GND 0.02127f
C15136 VDD.n5934 GND 0.04624f
C15137 VDD.n5935 GND 0.02704f
C15138 VDD.n5936 GND 0.02299f
C15139 VDD.t716 GND 0.57933f
C15140 VDD.n5937 GND 0.04624f
C15141 VDD.n5938 GND 0.04624f
C15142 VDD.n5939 GND 0.02704f
C15143 VDD.n5940 GND 0.02503f
C15144 VDD.t656 GND 0.02128f
C15145 VDD.t475 GND 0.02128f
C15146 VDD.n5941 GND 0.02885f
C15147 VDD.n5942 GND 0.04885f
C15148 VDD.n5943 GND 0.04624f
C15149 VDD.n5944 GND 0.04885f
C15150 VDD.n5945 GND 0.04556f
C15151 VDD.n5946 GND 0.04556f
C15152 VDD.t20 GND 0.57933f
C15153 VDD.n5947 GND 0.04556f
C15154 VDD.n5948 GND 0.04624f
C15155 VDD.n5949 GND 0.04624f
C15156 VDD.n5950 GND 0.02704f
C15157 VDD.n5951 GND 0.02299f
C15158 VDD.n5952 GND 0.04885f
C15159 VDD.n5953 GND 0.04624f
C15160 VDD.n5954 GND 0.02704f
C15161 VDD.n5955 GND 0.02299f
C15162 VDD.t458 GND 0.57933f
C15163 VDD.n5956 GND 0.04556f
C15164 VDD.n5957 GND 0.04624f
C15165 VDD.n5958 GND 0.04624f
C15166 VDD.n5959 GND 0.02704f
C15167 VDD.n5960 GND 0.02299f
C15168 VDD.n5961 GND 0.04885f
C15169 VDD.t784 GND 0.02116f
C15170 VDD.t21 GND 0.02116f
C15171 VDD.n5962 GND 0.09893f
C15172 VDD.t459 GND 0.02116f
C15173 VDD.t289 GND 0.02116f
C15174 VDD.n5963 GND 0.09893f
C15175 VDD.n5964 GND 0.03784f
C15176 VDD.n5965 GND 0.02127f
C15177 VDD.n5966 GND 0.04624f
C15178 VDD.n5967 GND 0.02704f
C15179 VDD.n5968 GND 0.02299f
C15180 VDD.t388 GND 0.57933f
C15181 VDD.n5969 GND 0.04556f
C15182 VDD.n5970 GND 0.04624f
C15183 VDD.n5971 GND 0.04624f
C15184 VDD.n5972 GND 0.02704f
C15185 VDD.n5973 GND 0.02299f
C15186 VDD.n5974 GND 0.04885f
C15187 VDD.t389 GND 0.02128f
C15188 VDD.t697 GND 0.02128f
C15189 VDD.n5975 GND 0.12159f
C15190 VDD.n5976 GND 0.02396f
C15191 VDD.n5977 GND 0.04624f
C15192 VDD.n5978 GND 0.02704f
C15193 VDD.n5979 GND 0.02299f
C15194 VDD.t618 GND 0.57933f
C15195 VDD.n5980 GND 0.04556f
C15196 VDD.n5981 GND 0.04624f
C15197 VDD.n5982 GND 0.04624f
C15198 VDD.n5983 GND 0.02704f
C15199 VDD.n5984 GND 0.02299f
C15200 VDD.n5985 GND 0.04885f
C15201 VDD.n5986 GND 0.02885f
C15202 VDD.n5987 GND 0.04624f
C15203 VDD.n5988 GND 0.02704f
C15204 VDD.n5989 GND 0.02299f
C15205 VDD.t4 GND 0.57933f
C15206 VDD.n5990 GND 0.04556f
C15207 VDD.n5991 GND 0.04624f
C15208 VDD.n5992 GND 0.04624f
C15209 VDD.n5993 GND 0.02704f
C15210 VDD.n5994 GND 0.02299f
C15211 VDD.n5995 GND 0.04885f
C15212 VDD.t325 GND 0.02116f
C15213 VDD.t885 GND 0.02116f
C15214 VDD.n5996 GND 0.09893f
C15215 VDD.t5 GND 0.02116f
C15216 VDD.t619 GND 0.02116f
C15217 VDD.n5997 GND 0.09893f
C15218 VDD.n5998 GND 0.03784f
C15219 VDD.n5999 GND 0.02127f
C15220 VDD.n6000 GND 0.04624f
C15221 VDD.n6001 GND 0.02704f
C15222 VDD.n6002 GND 0.02299f
C15223 VDD.t460 GND 0.57933f
C15224 VDD.n6003 GND 0.04624f
C15225 VDD.n6004 GND 0.04624f
C15226 VDD.n6005 GND 0.08322f
C15227 VDD.t326 GND 0.57933f
C15228 VDD.n6006 GND 0.04556f
C15229 VDD.n6007 GND 0.04624f
C15230 VDD.n6008 GND 0.04624f
C15231 VDD.n6009 GND 0.02704f
C15232 VDD.n6010 GND 0.02299f
C15233 VDD.n6011 GND 0.04885f
C15234 VDD.t461 GND 0.02128f
C15235 VDD.n6012 GND 0.06662f
C15236 VDD.n6013 GND 0.01638f
C15237 VDD.n6014 GND 0.02127f
C15238 VDD.n6015 GND 0.04624f
C15239 VDD.n6016 GND 0.02704f
C15240 VDD.n6017 GND 0.02299f
C15241 VDD.t316 GND 0.57933f
C15242 VDD.n6018 GND 0.04556f
C15243 VDD.n6019 GND 0.04624f
C15244 VDD.n6020 GND 0.04624f
C15245 VDD.n6021 GND 0.02704f
C15246 VDD.n6022 GND 0.02299f
C15247 VDD.n6023 GND 0.04885f
C15248 VDD.t318 GND 0.02116f
C15249 VDD.t546 GND 0.02116f
C15250 VDD.n6024 GND 0.09893f
C15251 VDD.t317 GND 0.02116f
C15252 VDD.t327 GND 0.02116f
C15253 VDD.n6025 GND 0.09893f
C15254 VDD.n6026 GND 0.03784f
C15255 VDD.n6027 GND 0.02127f
C15256 VDD.n6028 GND 0.04624f
C15257 VDD.n6029 GND 0.02704f
C15258 VDD.n6030 GND 0.02299f
C15259 VDD.t356 GND 0.57933f
C15260 VDD.n6031 GND 0.04556f
C15261 VDD.n6032 GND 0.04624f
C15262 VDD.n6033 GND 0.04624f
C15263 VDD.n6034 GND 0.02704f
C15264 VDD.n6035 GND 0.02299f
C15265 VDD.n6036 GND 0.04885f
C15266 VDD.t357 GND 0.02128f
C15267 VDD.t692 GND 0.02128f
C15268 VDD.n6037 GND 0.12159f
C15269 VDD.n6038 GND 0.02396f
C15270 VDD.n6039 GND 0.04624f
C15271 VDD.n6040 GND 0.02704f
C15272 VDD.n6041 GND 0.02299f
C15273 VDD.t371 GND 0.57933f
C15274 VDD.n6042 GND 0.04556f
C15275 VDD.n6043 GND 0.04624f
C15276 VDD.n6044 GND 0.04624f
C15277 VDD.n6045 GND 0.02704f
C15278 VDD.n6046 GND 0.02299f
C15279 VDD.n6047 GND 0.04885f
C15280 VDD.n6048 GND 0.02885f
C15281 VDD.n6049 GND 0.04624f
C15282 VDD.n6050 GND 0.02704f
C15283 VDD.n6051 GND 0.02299f
C15284 VDD.t523 GND 0.57933f
C15285 VDD.n6052 GND 0.04556f
C15286 VDD.n6053 GND 0.04624f
C15287 VDD.n6054 GND 0.04624f
C15288 VDD.n6055 GND 0.02704f
C15289 VDD.n6056 GND 0.02299f
C15290 VDD.n6057 GND 0.04885f
C15291 VDD.n6058 GND 0.04624f
C15292 VDD.n6059 GND 0.02704f
C15293 VDD.n6060 GND 0.02299f
C15294 VDD.n6061 GND 0.02299f
C15295 VDD.n6062 GND 0.04556f
C15296 VDD.n6063 GND 0.6274f
C15297 VDD.n6064 GND 0.04556f
C15298 VDD.n6065 GND 0.04624f
C15299 VDD.t524 GND 0.02116f
C15300 VDD.t873 GND 0.02116f
C15301 VDD.n6066 GND 0.09893f
C15302 VDD.t910 GND 0.02116f
C15303 VDD.t372 GND 0.02116f
C15304 VDD.n6067 GND 0.09893f
C15305 VDD.n6068 GND 0.07074f
C15306 VDD.n6069 GND 0.06917f
C15307 VDD.n6070 GND 0.04885f
C15308 VDD.n6071 GND 0.02299f
C15309 VDD.n6072 GND 0.04556f
C15310 VDD.n6073 GND 0.46716f
C15311 VDD.n6074 GND 0.02299f
C15312 VDD.n6075 GND 0.04556f
C15313 VDD.n6076 GND 0.46716f
C15314 VDD.n6077 GND 0.04556f
C15315 VDD.n6078 GND 0.04624f
C15316 VDD.n6079 GND 0.05737f
C15317 VDD.n6080 GND 0.04885f
C15318 VDD.n6081 GND 0.02299f
C15319 VDD.n6082 GND 0.04556f
C15320 VDD.n6083 GND 0.46716f
C15321 VDD.n6084 GND 0.02299f
C15322 VDD.n6085 GND 0.04556f
C15323 VDD.n6086 GND 0.46716f
C15324 VDD.n6087 GND 0.04556f
C15325 VDD.n6088 GND 0.04624f
C15326 VDD.n6089 GND 0.05737f
C15327 VDD.n6090 GND 0.04885f
C15328 VDD.n6091 GND 0.02299f
C15329 VDD.n6092 GND 0.04556f
C15330 VDD.n6093 GND 0.6274f
C15331 VDD.n6094 GND 0.02299f
C15332 VDD.n6095 GND 0.04556f
C15333 VDD.n6096 GND 0.6274f
C15334 VDD.n6097 GND 0.04556f
C15335 VDD.n6098 GND 0.04624f
C15336 VDD.n6099 GND 0.05737f
C15337 VDD.n6100 GND 0.04885f
C15338 VDD.n6101 GND 0.02299f
C15339 VDD.n6102 GND 0.04556f
C15340 VDD.n6103 GND 0.46716f
C15341 VDD.n6104 GND 0.02299f
C15342 VDD.n6105 GND 0.04556f
C15343 VDD.n6106 GND 0.46716f
C15344 VDD.n6107 GND 0.04556f
C15345 VDD.n6108 GND 0.04624f
C15346 VDD.n6109 GND 0.05737f
C15347 VDD.n6110 GND 0.04885f
C15348 VDD.n6111 GND 0.02299f
C15349 VDD.n6112 GND 0.04556f
C15350 VDD.n6113 GND 0.6274f
C15351 VDD.n6114 GND 0.6274f
C15352 VDD.n6115 GND 0.04556f
C15353 VDD.n6116 GND 0.02503f
C15354 VDD.n6117 GND 0.02704f
C15355 VDD.n6118 GND 0.02503f
C15356 VDD.n6119 GND 0.04556f
C15357 VDD.n6120 GND 0.6274f
C15358 VDD.n6121 GND 0.02299f
C15359 VDD.n6122 GND 0.04556f
C15360 VDD.n6123 GND 0.6274f
C15361 VDD.n6124 GND 0.04556f
C15362 VDD.n6125 GND 0.04624f
C15363 VDD.n6126 GND 0.05737f
C15364 VDD.n6127 GND 0.04885f
C15365 VDD.n6128 GND 0.02299f
C15366 VDD.n6129 GND 0.04556f
C15367 VDD.n6130 GND 0.46716f
C15368 VDD.n6131 GND 0.02299f
C15369 VDD.n6132 GND 0.04556f
C15370 VDD.n6133 GND 0.46716f
C15371 VDD.n6134 GND 0.04556f
C15372 VDD.n6135 GND 0.04624f
C15373 VDD.n6136 GND 0.05737f
C15374 VDD.n6137 GND 0.04885f
C15375 VDD.n6138 GND 0.02299f
C15376 VDD.n6139 GND 0.04556f
C15377 VDD.n6140 GND 0.46716f
C15378 VDD.n6141 GND 0.02299f
C15379 VDD.n6142 GND 0.04556f
C15380 VDD.n6143 GND 0.46716f
C15381 VDD.n6144 GND 0.04556f
C15382 VDD.n6145 GND 0.04624f
C15383 VDD.n6146 GND 0.05737f
C15384 VDD.n6147 GND 0.04885f
C15385 VDD.n6148 GND 0.02299f
C15386 VDD.n6149 GND 0.04556f
C15387 VDD.n6150 GND 0.6274f
C15388 VDD.n6151 GND 0.02299f
C15389 VDD.n6152 GND 0.04556f
C15390 VDD.n6153 GND 0.6274f
C15391 VDD.n6154 GND 0.04556f
C15392 VDD.n6155 GND 0.04624f
C15393 VDD.n6156 GND 0.05737f
C15394 VDD.n6157 GND 0.04885f
C15395 VDD.n6158 GND 0.02299f
C15396 VDD.n6159 GND 0.04556f
C15397 VDD.n6160 GND 0.46716f
C15398 VDD.n6161 GND 0.02299f
C15399 VDD.n6162 GND 0.04556f
C15400 VDD.n6163 GND 0.46716f
C15401 VDD.n6164 GND 0.04556f
C15402 VDD.n6165 GND 0.04624f
C15403 VDD.n6166 GND 0.05737f
C15404 VDD.n6167 GND 0.04885f
C15405 VDD.n6168 GND 0.02299f
C15406 VDD.n6169 GND 0.04556f
C15407 VDD.n6170 GND 0.46716f
C15408 VDD.n6171 GND 0.46716f
C15409 VDD.n6172 GND 0.02299f
C15410 VDD.n6173 GND 0.02299f
C15411 VDD.n6174 GND 0.02704f
C15412 VDD.n6175 GND 0.04624f
C15413 VDD.n6176 GND 0.04556f
C15414 VDD.n6177 GND 0.6274f
C15415 VDD.n6178 GND 0.6274f
C15416 VDD.n6179 GND 0.04556f
C15417 VDD.n6180 GND 0.04556f
C15418 VDD.n6181 GND 0.02299f
C15419 VDD.n6182 GND 0.02299f
C15420 VDD.n6183 GND 0.02704f
C15421 VDD.n6184 GND 0.04624f
C15422 VDD.t474 GND 0.57933f
C15423 VDD.n6185 GND 0.04624f
C15424 VDD.n6186 GND 0.05737f
C15425 VDD.n6187 GND 0.02396f
C15426 VDD.n6188 GND 0.12159f
C15427 VDD.t717 GND 0.02128f
C15428 VDD.n6189 GND 0.06662f
C15429 VDD.n6190 GND 0.01638f
C15430 VDD.n6191 GND 0.08322f
C15431 VDD.n6192 GND 0.02503f
C15432 VDD.n6193 GND 0.04556f
C15433 VDD.n6194 GND 0.6274f
C15434 VDD.n6195 GND 0.02299f
C15435 VDD.n6196 GND 0.04556f
C15436 VDD.n6197 GND 0.6274f
C15437 VDD.n6198 GND 0.04556f
C15438 VDD.n6199 GND 0.04624f
C15439 VDD.n6200 GND 0.05737f
C15440 VDD.n6201 GND 0.04885f
C15441 VDD.n6202 GND 0.02299f
C15442 VDD.n6203 GND 0.04556f
C15443 VDD.n6204 GND 0.46716f
C15444 VDD.n6205 GND 0.02299f
C15445 VDD.n6206 GND 0.04556f
C15446 VDD.n6207 GND 0.46716f
C15447 VDD.n6208 GND 0.04556f
C15448 VDD.n6209 GND 0.04624f
C15449 VDD.n6210 GND 0.05737f
C15450 VDD.n6211 GND 0.04885f
C15451 VDD.n6212 GND 0.02299f
C15452 VDD.n6213 GND 0.04556f
C15453 VDD.n6214 GND 0.46716f
C15454 VDD.n6215 GND 0.02299f
C15455 VDD.n6216 GND 0.04556f
C15456 VDD.n6217 GND 0.46716f
C15457 VDD.n6218 GND 0.04556f
C15458 VDD.n6219 GND 0.04624f
C15459 VDD.n6220 GND 0.05737f
C15460 VDD.n6221 GND 0.04885f
C15461 VDD.n6222 GND 0.02299f
C15462 VDD.n6223 GND 0.04556f
C15463 VDD.n6224 GND 0.6274f
C15464 VDD.n6225 GND 0.02299f
C15465 VDD.n6226 GND 0.04556f
C15466 VDD.n6227 GND 0.6274f
C15467 VDD.n6228 GND 0.04556f
C15468 VDD.n6229 GND 0.04624f
C15469 VDD.n6230 GND 0.05737f
C15470 VDD.n6231 GND 0.04885f
C15471 VDD.n6232 GND 0.02299f
C15472 VDD.n6233 GND 0.04556f
C15473 VDD.n6234 GND 0.46716f
C15474 VDD.n6235 GND 0.02299f
C15475 VDD.n6236 GND 0.04556f
C15476 VDD.n6237 GND 0.46716f
C15477 VDD.n6238 GND 0.04556f
C15478 VDD.n6239 GND 0.04624f
C15479 VDD.n6240 GND 0.05737f
C15480 VDD.n6241 GND 0.04885f
C15481 VDD.n6242 GND 0.02299f
C15482 VDD.n6243 GND 0.04556f
C15483 VDD.n6244 GND 0.6274f
C15484 VDD.n6245 GND 0.6274f
C15485 VDD.n6246 GND 0.04556f
C15486 VDD.n6247 GND 0.02503f
C15487 VDD.n6248 GND 0.02704f
C15488 VDD.n6249 GND 0.02503f
C15489 VDD.n6250 GND 0.04556f
C15490 VDD.n6251 GND 0.6274f
C15491 VDD.n6252 GND 0.02299f
C15492 VDD.n6253 GND 0.04556f
C15493 VDD.n6254 GND 0.6274f
C15494 VDD.n6255 GND 0.04556f
C15495 VDD.n6256 GND 0.04624f
C15496 VDD.n6257 GND 0.05737f
C15497 VDD.n6258 GND 0.04885f
C15498 VDD.n6259 GND 0.02299f
C15499 VDD.n6260 GND 0.04556f
C15500 VDD.n6261 GND 0.46716f
C15501 VDD.n6262 GND 0.02299f
C15502 VDD.n6263 GND 0.04556f
C15503 VDD.n6264 GND 0.46716f
C15504 VDD.n6265 GND 0.04556f
C15505 VDD.n6266 GND 0.04624f
C15506 VDD.n6267 GND 0.05737f
C15507 VDD.n6268 GND 0.04885f
C15508 VDD.n6269 GND 0.02299f
C15509 VDD.n6270 GND 0.04556f
C15510 VDD.n6271 GND 0.46716f
C15511 VDD.n6272 GND 0.02299f
C15512 VDD.n6273 GND 0.04556f
C15513 VDD.n6274 GND 0.46716f
C15514 VDD.n6275 GND 0.04556f
C15515 VDD.n6276 GND 0.04624f
C15516 VDD.n6277 GND 0.05737f
C15517 VDD.n6278 GND 0.04885f
C15518 VDD.n6279 GND 0.02299f
C15519 VDD.n6280 GND 0.04556f
C15520 VDD.n6281 GND 0.6274f
C15521 VDD.n6282 GND 0.02299f
C15522 VDD.n6283 GND 0.04556f
C15523 VDD.n6284 GND 0.6274f
C15524 VDD.n6285 GND 0.04556f
C15525 VDD.n6286 GND 0.04624f
C15526 VDD.n6287 GND 0.05737f
C15527 VDD.n6288 GND 0.04885f
C15528 VDD.n6289 GND 0.02299f
C15529 VDD.n6290 GND 0.04556f
C15530 VDD.n6291 GND 0.46716f
C15531 VDD.n6292 GND 0.02299f
C15532 VDD.n6293 GND 0.04556f
C15533 VDD.n6294 GND 0.46716f
C15534 VDD.n6295 GND 0.04556f
C15535 VDD.n6296 GND 0.04624f
C15536 VDD.n6297 GND 0.05737f
C15537 VDD.n6298 GND 0.04885f
C15538 VDD.n6299 GND 0.02299f
C15539 VDD.n6300 GND 0.04556f
C15540 VDD.n6301 GND 0.46716f
C15541 VDD.n6302 GND 0.46716f
C15542 VDD.n6303 GND 0.02299f
C15543 VDD.n6304 GND 0.02299f
C15544 VDD.n6305 GND 0.02704f
C15545 VDD.n6306 GND 0.04624f
C15546 VDD.n6307 GND 0.04556f
C15547 VDD.n6308 GND 0.6274f
C15548 VDD.n6309 GND 0.6274f
C15549 VDD.n6310 GND 0.04556f
C15550 VDD.n6311 GND 0.04556f
C15551 VDD.n6312 GND 0.02299f
C15552 VDD.n6313 GND 0.02299f
C15553 VDD.n6314 GND 0.02704f
C15554 VDD.n6315 GND 0.04624f
C15555 VDD.t536 GND 0.57933f
C15556 VDD.n6316 GND 0.04624f
C15557 VDD.n6317 GND 0.05737f
C15558 VDD.n6318 GND 0.02396f
C15559 VDD.n6319 GND 0.12159f
C15560 VDD.t721 GND 0.02128f
C15561 VDD.n6320 GND 0.06662f
C15562 VDD.n6321 GND 0.01638f
C15563 VDD.n6322 GND 0.08322f
C15564 VDD.n6323 GND 0.02503f
C15565 VDD.n6324 GND 0.04556f
C15566 VDD.n6325 GND 0.6274f
C15567 VDD.n6326 GND 0.02299f
C15568 VDD.n6327 GND 0.04556f
C15569 VDD.n6328 GND 0.6274f
C15570 VDD.n6329 GND 0.04556f
C15571 VDD.n6330 GND 0.04624f
C15572 VDD.n6331 GND 0.05737f
C15573 VDD.n6332 GND 0.04885f
C15574 VDD.n6333 GND 0.02299f
C15575 VDD.n6334 GND 0.04556f
C15576 VDD.n6335 GND 0.46716f
C15577 VDD.n6336 GND 0.02299f
C15578 VDD.n6337 GND 0.04556f
C15579 VDD.n6338 GND 0.46716f
C15580 VDD.n6339 GND 0.04556f
C15581 VDD.n6340 GND 0.04624f
C15582 VDD.n6341 GND 0.05737f
C15583 VDD.n6342 GND 0.04885f
C15584 VDD.n6343 GND 0.02299f
C15585 VDD.n6344 GND 0.04556f
C15586 VDD.n6345 GND 0.46716f
C15587 VDD.n6346 GND 0.02299f
C15588 VDD.n6347 GND 0.04556f
C15589 VDD.n6348 GND 0.46716f
C15590 VDD.n6349 GND 0.04556f
C15591 VDD.n6350 GND 0.04624f
C15592 VDD.n6351 GND 0.05737f
C15593 VDD.n6352 GND 0.04885f
C15594 VDD.n6353 GND 0.02299f
C15595 VDD.n6354 GND 0.04556f
C15596 VDD.n6355 GND 0.6274f
C15597 VDD.n6356 GND 0.02299f
C15598 VDD.n6357 GND 0.04556f
C15599 VDD.n6358 GND 0.6274f
C15600 VDD.n6359 GND 0.04556f
C15601 VDD.n6360 GND 0.04624f
C15602 VDD.n6361 GND 0.05737f
C15603 VDD.n6362 GND 0.04885f
C15604 VDD.n6363 GND 0.02299f
C15605 VDD.n6364 GND 0.04556f
C15606 VDD.n6365 GND 0.46716f
C15607 VDD.n6366 GND 0.02299f
C15608 VDD.n6367 GND 0.04556f
C15609 VDD.n6368 GND 0.46716f
C15610 VDD.n6369 GND 0.04556f
C15611 VDD.n6370 GND 0.04624f
C15612 VDD.n6371 GND 0.05737f
C15613 VDD.n6372 GND 0.04885f
C15614 VDD.n6373 GND 0.02299f
C15615 VDD.n6374 GND 0.04556f
C15616 VDD.n6375 GND 0.6274f
C15617 VDD.n6376 GND 0.6274f
C15618 VDD.n6377 GND 0.04556f
C15619 VDD.n6378 GND 0.02503f
C15620 VDD.n6379 GND 0.02704f
C15621 VDD.n6380 GND 0.02503f
C15622 VDD.n6381 GND 0.04556f
C15623 VDD.n6382 GND 0.6274f
C15624 VDD.n6383 GND 0.02299f
C15625 VDD.n6384 GND 0.04556f
C15626 VDD.n6385 GND 0.6274f
C15627 VDD.n6386 GND 0.04556f
C15628 VDD.n6387 GND 0.04624f
C15629 VDD.n6388 GND 0.05737f
C15630 VDD.n6389 GND 0.04885f
C15631 VDD.n6390 GND 0.02299f
C15632 VDD.n6391 GND 0.04556f
C15633 VDD.n6392 GND 0.46716f
C15634 VDD.n6393 GND 0.02299f
C15635 VDD.n6394 GND 0.04556f
C15636 VDD.n6395 GND 0.46716f
C15637 VDD.n6396 GND 0.04556f
C15638 VDD.n6397 GND 0.04624f
C15639 VDD.n6398 GND 0.05737f
C15640 VDD.n6399 GND 0.04885f
C15641 VDD.n6400 GND 0.02299f
C15642 VDD.n6401 GND 0.04556f
C15643 VDD.n6402 GND 0.46716f
C15644 VDD.n6403 GND 0.02299f
C15645 VDD.n6404 GND 0.04556f
C15646 VDD.n6405 GND 0.46716f
C15647 VDD.n6406 GND 0.04556f
C15648 VDD.n6407 GND 0.04624f
C15649 VDD.n6408 GND 0.05737f
C15650 VDD.n6409 GND 0.04885f
C15651 VDD.n6410 GND 0.02299f
C15652 VDD.n6411 GND 0.04556f
C15653 VDD.n6412 GND 0.6274f
C15654 VDD.n6413 GND 0.02299f
C15655 VDD.n6414 GND 0.04556f
C15656 VDD.n6415 GND 0.6274f
C15657 VDD.n6416 GND 0.04556f
C15658 VDD.n6417 GND 0.04624f
C15659 VDD.n6418 GND 0.05737f
C15660 VDD.n6419 GND 0.04885f
C15661 VDD.n6420 GND 0.02299f
C15662 VDD.n6421 GND 0.04556f
C15663 VDD.n6422 GND 0.46716f
C15664 VDD.n6423 GND 0.02299f
C15665 VDD.n6424 GND 0.04556f
C15666 VDD.n6425 GND 0.46716f
C15667 VDD.n6426 GND 0.04556f
C15668 VDD.n6427 GND 0.04624f
C15669 VDD.n6428 GND 0.05737f
C15670 VDD.n6429 GND 0.04885f
C15671 VDD.n6430 GND 0.02299f
C15672 VDD.n6431 GND 0.04556f
C15673 VDD.n6432 GND 0.46716f
C15674 VDD.n6433 GND 0.46716f
C15675 VDD.n6434 GND 0.02299f
C15676 VDD.n6435 GND 0.02299f
C15677 VDD.n6436 GND 0.02704f
C15678 VDD.n6437 GND 0.04624f
C15679 VDD.n6438 GND 0.04556f
C15680 VDD.n6439 GND 0.6274f
C15681 VDD.n6440 GND 0.6274f
C15682 VDD.n6441 GND 0.04556f
C15683 VDD.n6442 GND 0.04556f
C15684 VDD.n6443 GND 0.02299f
C15685 VDD.n6444 GND 0.02299f
C15686 VDD.n6445 GND 0.02704f
C15687 VDD.n6446 GND 0.04624f
C15688 VDD.t285 GND 0.57933f
C15689 VDD.n6447 GND 0.04624f
C15690 VDD.n6448 GND 0.05737f
C15691 VDD.n6449 GND 0.02396f
C15692 VDD.n6450 GND 0.12159f
C15693 VDD.t451 GND 0.02128f
C15694 VDD.n6451 GND 0.06662f
C15695 VDD.n6452 GND 0.01638f
C15696 VDD.n6453 GND 0.08322f
C15697 VDD.n6454 GND 0.02503f
C15698 VDD.n6455 GND 0.04556f
C15699 VDD.n6456 GND 0.6274f
C15700 VDD.n6457 GND 0.02299f
C15701 VDD.n6458 GND 0.04556f
C15702 VDD.n6459 GND 0.6274f
C15703 VDD.n6460 GND 0.04556f
C15704 VDD.n6461 GND 0.04624f
C15705 VDD.n6462 GND 0.05737f
C15706 VDD.n6463 GND 0.04885f
C15707 VDD.n6464 GND 0.02299f
C15708 VDD.n6465 GND 0.04556f
C15709 VDD.n6466 GND 0.46716f
C15710 VDD.n6467 GND 0.02299f
C15711 VDD.n6468 GND 0.04556f
C15712 VDD.n6469 GND 0.46716f
C15713 VDD.n6470 GND 0.04556f
C15714 VDD.n6471 GND 0.04624f
C15715 VDD.n6472 GND 0.05737f
C15716 VDD.n6473 GND 0.04885f
C15717 VDD.n6474 GND 0.02299f
C15718 VDD.n6475 GND 0.04556f
C15719 VDD.n6476 GND 0.46716f
C15720 VDD.n6477 GND 0.02299f
C15721 VDD.n6478 GND 0.04556f
C15722 VDD.n6479 GND 0.46716f
C15723 VDD.n6480 GND 0.04556f
C15724 VDD.n6481 GND 0.04624f
C15725 VDD.n6482 GND 0.05737f
C15726 VDD.n6483 GND 0.04885f
C15727 VDD.n6484 GND 0.02299f
C15728 VDD.n6485 GND 0.04556f
C15729 VDD.n6486 GND 0.6274f
C15730 VDD.n6487 GND 0.02299f
C15731 VDD.n6488 GND 0.04556f
C15732 VDD.n6489 GND 0.6274f
C15733 VDD.n6490 GND 0.04556f
C15734 VDD.n6491 GND 0.04624f
C15735 VDD.n6492 GND 0.05737f
C15736 VDD.n6493 GND 0.04885f
C15737 VDD.n6494 GND 0.02299f
C15738 VDD.n6495 GND 0.04556f
C15739 VDD.n6496 GND 0.46716f
C15740 VDD.n6497 GND 0.02299f
C15741 VDD.n6498 GND 0.04556f
C15742 VDD.n6499 GND 0.46716f
C15743 VDD.n6500 GND 0.04556f
C15744 VDD.n6501 GND 0.04624f
C15745 VDD.n6502 GND 0.05737f
C15746 VDD.n6503 GND 0.04885f
C15747 VDD.n6504 GND 0.02299f
C15748 VDD.n6505 GND 0.04556f
C15749 VDD.n6506 GND 0.6274f
C15750 VDD.n6507 GND 0.6274f
C15751 VDD.n6508 GND 0.04556f
C15752 VDD.n6509 GND 0.02503f
C15753 VDD.n6510 GND 0.02704f
C15754 VDD.n6511 GND 0.02503f
C15755 VDD.n6512 GND 0.04556f
C15756 VDD.n6513 GND 0.6274f
C15757 VDD.n6514 GND 0.02299f
C15758 VDD.n6515 GND 0.04556f
C15759 VDD.n6516 GND 0.6274f
C15760 VDD.n6517 GND 0.04556f
C15761 VDD.n6518 GND 0.04624f
C15762 VDD.n6519 GND 0.05737f
C15763 VDD.n6520 GND 0.04885f
C15764 VDD.n6521 GND 0.02299f
C15765 VDD.n6522 GND 0.04556f
C15766 VDD.n6523 GND 0.46716f
C15767 VDD.n6524 GND 0.02299f
C15768 VDD.n6525 GND 0.04556f
C15769 VDD.n6526 GND 0.46716f
C15770 VDD.n6527 GND 0.04556f
C15771 VDD.n6528 GND 0.04624f
C15772 VDD.n6529 GND 0.05737f
C15773 VDD.n6530 GND 0.04885f
C15774 VDD.n6531 GND 0.02299f
C15775 VDD.n6532 GND 0.04556f
C15776 VDD.n6533 GND 0.46716f
C15777 VDD.n6534 GND 0.02299f
C15778 VDD.n6535 GND 0.04556f
C15779 VDD.n6536 GND 0.46716f
C15780 VDD.n6537 GND 0.04556f
C15781 VDD.n6538 GND 0.04624f
C15782 VDD.n6539 GND 0.05737f
C15783 VDD.n6540 GND 0.04885f
C15784 VDD.n6541 GND 0.02299f
C15785 VDD.n6542 GND 0.04556f
C15786 VDD.n6543 GND 0.6274f
C15787 VDD.n6544 GND 0.02299f
C15788 VDD.n6545 GND 0.04556f
C15789 VDD.n6546 GND 0.6274f
C15790 VDD.n6547 GND 0.04556f
C15791 VDD.n6548 GND 0.04624f
C15792 VDD.n6549 GND 0.05737f
C15793 VDD.n6550 GND 0.04885f
C15794 VDD.n6551 GND 0.02299f
C15795 VDD.n6552 GND 0.04556f
C15796 VDD.n6553 GND 0.46716f
C15797 VDD.n6554 GND 0.02299f
C15798 VDD.n6555 GND 0.04556f
C15799 VDD.n6556 GND 0.46716f
C15800 VDD.n6557 GND 0.04556f
C15801 VDD.n6558 GND 0.04624f
C15802 VDD.n6559 GND 0.05737f
C15803 VDD.n6560 GND 0.04885f
C15804 VDD.n6561 GND 0.02299f
C15805 VDD.n6562 GND 0.04556f
C15806 VDD.n6563 GND 0.46716f
C15807 VDD.n6564 GND 0.46716f
C15808 VDD.n6565 GND 0.02299f
C15809 VDD.n6566 GND 0.02299f
C15810 VDD.n6567 GND 0.02704f
C15811 VDD.n6568 GND 0.04624f
C15812 VDD.n6569 GND 0.04556f
C15813 VDD.n6570 GND 0.6274f
C15814 VDD.n6571 GND 0.6274f
C15815 VDD.n6572 GND 0.04556f
C15816 VDD.n6573 GND 0.04556f
C15817 VDD.n6574 GND 0.02299f
C15818 VDD.n6575 GND 0.02299f
C15819 VDD.n6576 GND 0.02704f
C15820 VDD.n6577 GND 0.04624f
C15821 VDD.t563 GND 0.57933f
C15822 VDD.n6578 GND 0.04624f
C15823 VDD.n6579 GND 0.05737f
C15824 VDD.n6580 GND 0.02396f
C15825 VDD.n6581 GND 0.12159f
C15826 VDD.t17 GND 0.02128f
C15827 VDD.n6582 GND 0.06662f
C15828 VDD.n6583 GND 0.01638f
C15829 VDD.n6584 GND 0.08322f
C15830 VDD.n6585 GND 0.02503f
C15831 VDD.n6586 GND 0.04556f
C15832 VDD.n6587 GND 0.6274f
C15833 VDD.n6588 GND 0.02299f
C15834 VDD.n6589 GND 0.04556f
C15835 VDD.n6590 GND 0.6274f
C15836 VDD.n6591 GND 0.04556f
C15837 VDD.n6592 GND 0.04624f
C15838 VDD.n6593 GND 0.05737f
C15839 VDD.n6594 GND 0.04885f
C15840 VDD.n6595 GND 0.02299f
C15841 VDD.n6596 GND 0.04556f
C15842 VDD.n6597 GND 0.46716f
C15843 VDD.n6598 GND 0.02299f
C15844 VDD.n6599 GND 0.04556f
C15845 VDD.n6600 GND 0.46716f
C15846 VDD.n6601 GND 0.04556f
C15847 VDD.n6602 GND 0.04624f
C15848 VDD.n6603 GND 0.05737f
C15849 VDD.n6604 GND 0.04885f
C15850 VDD.n6605 GND 0.02299f
C15851 VDD.n6606 GND 0.04556f
C15852 VDD.n6607 GND 0.46716f
C15853 VDD.n6608 GND 0.02299f
C15854 VDD.n6609 GND 0.04556f
C15855 VDD.n6610 GND 0.46716f
C15856 VDD.n6611 GND 0.04556f
C15857 VDD.n6612 GND 0.04624f
C15858 VDD.n6613 GND 0.05737f
C15859 VDD.n6614 GND 0.04885f
C15860 VDD.n6615 GND 0.02299f
C15861 VDD.n6616 GND 0.04556f
C15862 VDD.n6617 GND 0.6274f
C15863 VDD.n6618 GND 0.02299f
C15864 VDD.n6619 GND 0.04556f
C15865 VDD.n6620 GND 0.6274f
C15866 VDD.n6621 GND 0.04556f
C15867 VDD.n6622 GND 0.04624f
C15868 VDD.n6623 GND 0.05737f
C15869 VDD.n6624 GND 0.04885f
C15870 VDD.n6625 GND 0.02299f
C15871 VDD.n6626 GND 0.04556f
C15872 VDD.n6627 GND 0.46716f
C15873 VDD.n6628 GND 0.02299f
C15874 VDD.n6629 GND 0.04556f
C15875 VDD.n6630 GND 0.46716f
C15876 VDD.n6631 GND 0.04556f
C15877 VDD.n6632 GND 0.04624f
C15878 VDD.n6633 GND 0.05737f
C15879 VDD.n6634 GND 0.04885f
C15880 VDD.n6635 GND 0.02299f
C15881 VDD.n6636 GND 0.04556f
C15882 VDD.n6637 GND 0.6274f
C15883 VDD.n6638 GND 0.6274f
C15884 VDD.n6639 GND 0.04556f
C15885 VDD.n6640 GND 0.02503f
C15886 VDD.n6641 GND 0.02704f
C15887 VDD.n6642 GND 0.02503f
C15888 VDD.n6643 GND 0.04556f
C15889 VDD.n6644 GND 0.6274f
C15890 VDD.n6645 GND 0.02299f
C15891 VDD.n6646 GND 0.04556f
C15892 VDD.n6647 GND 0.6274f
C15893 VDD.n6648 GND 0.04556f
C15894 VDD.n6649 GND 0.04624f
C15895 VDD.n6650 GND 0.05737f
C15896 VDD.n6651 GND 0.04885f
C15897 VDD.n6652 GND 0.02299f
C15898 VDD.n6653 GND 0.04556f
C15899 VDD.n6654 GND 0.46716f
C15900 VDD.n6655 GND 0.02299f
C15901 VDD.n6656 GND 0.04556f
C15902 VDD.n6657 GND 0.46716f
C15903 VDD.n6658 GND 0.04556f
C15904 VDD.n6659 GND 0.04624f
C15905 VDD.n6660 GND 0.05737f
C15906 VDD.n6661 GND 0.04885f
C15907 VDD.n6662 GND 0.02299f
C15908 VDD.n6663 GND 0.04556f
C15909 VDD.n6664 GND 0.46716f
C15910 VDD.n6665 GND 0.02299f
C15911 VDD.n6666 GND 0.04556f
C15912 VDD.n6667 GND 0.46716f
C15913 VDD.n6668 GND 0.04556f
C15914 VDD.n6669 GND 0.04624f
C15915 VDD.n6670 GND 0.05737f
C15916 VDD.n6671 GND 0.04885f
C15917 VDD.n6672 GND 0.02299f
C15918 VDD.n6673 GND 0.04556f
C15919 VDD.n6674 GND 0.6274f
C15920 VDD.n6675 GND 0.02299f
C15921 VDD.n6676 GND 0.04556f
C15922 VDD.n6677 GND 0.6274f
C15923 VDD.n6678 GND 0.04556f
C15924 VDD.n6679 GND 0.04624f
C15925 VDD.n6680 GND 0.05737f
C15926 VDD.n6681 GND 0.04885f
C15927 VDD.n6682 GND 0.02299f
C15928 VDD.n6683 GND 0.04556f
C15929 VDD.n6684 GND 0.46716f
C15930 VDD.n6685 GND 0.02299f
C15931 VDD.n6686 GND 0.04556f
C15932 VDD.n6687 GND 0.46716f
C15933 VDD.n6688 GND 0.04556f
C15934 VDD.n6689 GND 0.04624f
C15935 VDD.n6690 GND 0.05737f
C15936 VDD.n6691 GND 0.04885f
C15937 VDD.n6692 GND 0.02299f
C15938 VDD.n6693 GND 0.04556f
C15939 VDD.n6694 GND 0.46716f
C15940 VDD.n6695 GND 0.46716f
C15941 VDD.n6696 GND 0.02299f
C15942 VDD.n6697 GND 0.02299f
C15943 VDD.n6698 GND 0.02704f
C15944 VDD.n6699 GND 0.04624f
C15945 VDD.n6700 GND 0.04556f
C15946 VDD.n6701 GND 0.6274f
C15947 VDD.n6702 GND 0.6274f
C15948 VDD.n6703 GND 0.04556f
C15949 VDD.n6704 GND 0.04556f
C15950 VDD.n6705 GND 0.02299f
C15951 VDD.n6706 GND 0.02299f
C15952 VDD.n6707 GND 0.02704f
C15953 VDD.n6708 GND 0.04624f
C15954 VDD.t364 GND 0.57933f
C15955 VDD.n6709 GND 0.04624f
C15956 VDD.n6710 GND 0.05737f
C15957 VDD.n6711 GND 0.02396f
C15958 VDD.n6712 GND 0.12159f
C15959 VDD.t719 GND 0.02128f
C15960 VDD.n6713 GND 0.06662f
C15961 VDD.n6714 GND 0.01638f
C15962 VDD.n6715 GND 0.08322f
C15963 VDD.n6716 GND 0.02503f
C15964 VDD.n6717 GND 0.04556f
C15965 VDD.n6718 GND 0.6274f
C15966 VDD.n6719 GND 0.02299f
C15967 VDD.n6720 GND 0.04556f
C15968 VDD.n6721 GND 0.6274f
C15969 VDD.n6722 GND 0.04556f
C15970 VDD.n6723 GND 0.04624f
C15971 VDD.n6724 GND 0.05737f
C15972 VDD.n6725 GND 0.04885f
C15973 VDD.n6726 GND 0.02299f
C15974 VDD.n6727 GND 0.04556f
C15975 VDD.n6728 GND 0.46716f
C15976 VDD.n6729 GND 0.02299f
C15977 VDD.n6730 GND 0.04556f
C15978 VDD.n6731 GND 0.46716f
C15979 VDD.n6732 GND 0.04556f
C15980 VDD.n6733 GND 0.04624f
C15981 VDD.n6734 GND 0.05737f
C15982 VDD.n6735 GND 0.04885f
C15983 VDD.n6736 GND 0.02299f
C15984 VDD.n6737 GND 0.04556f
C15985 VDD.n6738 GND 0.46716f
C15986 VDD.n6739 GND 0.02299f
C15987 VDD.n6740 GND 0.04556f
C15988 VDD.n6741 GND 0.46716f
C15989 VDD.n6742 GND 0.04556f
C15990 VDD.n6743 GND 0.04624f
C15991 VDD.n6744 GND 0.05737f
C15992 VDD.n6745 GND 0.04885f
C15993 VDD.n6746 GND 0.02299f
C15994 VDD.n6747 GND 0.04556f
C15995 VDD.n6748 GND 0.6274f
C15996 VDD.n6749 GND 0.02299f
C15997 VDD.n6750 GND 0.04556f
C15998 VDD.n6751 GND 0.6274f
C15999 VDD.n6752 GND 0.04556f
C16000 VDD.n6753 GND 0.04624f
C16001 VDD.n6754 GND 0.05737f
C16002 VDD.n6755 GND 0.04885f
C16003 VDD.n6756 GND 0.02299f
C16004 VDD.n6757 GND 0.04556f
C16005 VDD.n6758 GND 0.46716f
C16006 VDD.n6759 GND 0.02299f
C16007 VDD.n6760 GND 0.04556f
C16008 VDD.n6761 GND 0.46716f
C16009 VDD.n6762 GND 0.04556f
C16010 VDD.n6763 GND 0.04624f
C16011 VDD.n6764 GND 0.05737f
C16012 VDD.n6765 GND 0.04885f
C16013 VDD.n6766 GND 0.02299f
C16014 VDD.n6767 GND 0.04556f
C16015 VDD.n6768 GND 0.6274f
C16016 VDD.n6769 GND 0.6274f
C16017 VDD.n6770 GND 0.04556f
C16018 VDD.n6771 GND 0.02503f
C16019 VDD.n6772 GND 0.02704f
C16020 VDD.n6773 GND 0.02503f
C16021 VDD.n6774 GND 0.04556f
C16022 VDD.n6775 GND 0.6274f
C16023 VDD.n6776 GND 0.02299f
C16024 VDD.n6777 GND 0.04556f
C16025 VDD.n6778 GND 0.6274f
C16026 VDD.n6779 GND 0.04556f
C16027 VDD.n6780 GND 0.04624f
C16028 VDD.n6781 GND 0.05737f
C16029 VDD.n6782 GND 0.04885f
C16030 VDD.n6783 GND 0.02299f
C16031 VDD.n6784 GND 0.04556f
C16032 VDD.n6785 GND 0.46716f
C16033 VDD.n6786 GND 0.02299f
C16034 VDD.n6787 GND 0.04556f
C16035 VDD.n6788 GND 0.46716f
C16036 VDD.n6789 GND 0.04556f
C16037 VDD.n6790 GND 0.04624f
C16038 VDD.n6791 GND 0.05737f
C16039 VDD.n6792 GND 0.04885f
C16040 VDD.n6793 GND 0.02299f
C16041 VDD.n6794 GND 0.04556f
C16042 VDD.n6795 GND 0.46716f
C16043 VDD.n6796 GND 0.02299f
C16044 VDD.n6797 GND 0.04556f
C16045 VDD.n6798 GND 0.46716f
C16046 VDD.n6799 GND 0.04556f
C16047 VDD.n6800 GND 0.04624f
C16048 VDD.n6801 GND 0.05737f
C16049 VDD.n6802 GND 0.04885f
C16050 VDD.n6803 GND 0.02299f
C16051 VDD.n6804 GND 0.04556f
C16052 VDD.n6805 GND 0.6274f
C16053 VDD.n6806 GND 0.02299f
C16054 VDD.n6807 GND 0.04556f
C16055 VDD.n6808 GND 0.6274f
C16056 VDD.n6809 GND 0.04556f
C16057 VDD.n6810 GND 0.04624f
C16058 VDD.n6811 GND 0.05737f
C16059 VDD.n6812 GND 0.04885f
C16060 VDD.n6813 GND 0.02299f
C16061 VDD.n6814 GND 0.04556f
C16062 VDD.n6815 GND 0.46716f
C16063 VDD.n6816 GND 0.02299f
C16064 VDD.n6817 GND 0.04556f
C16065 VDD.n6818 GND 0.46716f
C16066 VDD.n6819 GND 0.04556f
C16067 VDD.n6820 GND 0.04624f
C16068 VDD.n6821 GND 0.05737f
C16069 VDD.n6822 GND 0.04885f
C16070 VDD.n6823 GND 0.02299f
C16071 VDD.n6824 GND 0.04556f
C16072 VDD.n6825 GND 0.46716f
C16073 VDD.n6826 GND 0.46716f
C16074 VDD.n6827 GND 0.02299f
C16075 VDD.n6828 GND 0.02299f
C16076 VDD.n6829 GND 0.02704f
C16077 VDD.n6830 GND 0.04624f
C16078 VDD.n6831 GND 0.04556f
C16079 VDD.n6832 GND 0.6274f
C16080 VDD.n6833 GND 0.6274f
C16081 VDD.n6834 GND 0.04556f
C16082 VDD.n6835 GND 0.04556f
C16083 VDD.n6836 GND 0.02299f
C16084 VDD.n6837 GND 0.02299f
C16085 VDD.n6838 GND 0.02704f
C16086 VDD.n6839 GND 0.04624f
C16087 VDD.t493 GND 0.57933f
C16088 VDD.n6840 GND 0.04624f
C16089 VDD.n6841 GND 0.05737f
C16090 VDD.n6842 GND 0.02396f
C16091 VDD.n6843 GND 0.12159f
C16092 VDD.t276 GND 0.02128f
C16093 VDD.n6844 GND 0.06662f
C16094 VDD.n6845 GND 0.01638f
C16095 VDD.n6846 GND 0.08322f
C16096 VDD.n6847 GND 0.02503f
C16097 VDD.n6848 GND 0.04556f
C16098 VDD.n6849 GND 0.6274f
C16099 VDD.n6850 GND 0.02299f
C16100 VDD.n6851 GND 0.04556f
C16101 VDD.n6852 GND 0.6274f
C16102 VDD.n6853 GND 0.04556f
C16103 VDD.n6854 GND 0.04624f
C16104 VDD.n6855 GND 0.05737f
C16105 VDD.n6856 GND 0.04885f
C16106 VDD.n6857 GND 0.02299f
C16107 VDD.n6858 GND 0.04556f
C16108 VDD.n6859 GND 0.46716f
C16109 VDD.n6860 GND 0.02299f
C16110 VDD.n6861 GND 0.04556f
C16111 VDD.n6862 GND 0.46716f
C16112 VDD.n6863 GND 0.04556f
C16113 VDD.n6864 GND 0.04624f
C16114 VDD.n6865 GND 0.05737f
C16115 VDD.n6866 GND 0.04885f
C16116 VDD.n6867 GND 0.02299f
C16117 VDD.n6868 GND 0.04556f
C16118 VDD.n6869 GND 0.46716f
C16119 VDD.n6870 GND 0.02299f
C16120 VDD.n6871 GND 0.04556f
C16121 VDD.n6872 GND 0.46716f
C16122 VDD.n6873 GND 0.04556f
C16123 VDD.n6874 GND 0.04624f
C16124 VDD.n6875 GND 0.05737f
C16125 VDD.n6876 GND 0.04885f
C16126 VDD.n6877 GND 0.02299f
C16127 VDD.n6878 GND 0.04556f
C16128 VDD.n6879 GND 0.6274f
C16129 VDD.n6880 GND 0.02299f
C16130 VDD.n6881 GND 0.04556f
C16131 VDD.n6882 GND 0.6274f
C16132 VDD.n6883 GND 0.04556f
C16133 VDD.n6884 GND 0.04624f
C16134 VDD.n6885 GND 0.05737f
C16135 VDD.n6886 GND 0.04885f
C16136 VDD.n6887 GND 0.02299f
C16137 VDD.n6888 GND 0.04556f
C16138 VDD.n6889 GND 0.46716f
C16139 VDD.n6890 GND 0.02299f
C16140 VDD.n6891 GND 0.04556f
C16141 VDD.n6892 GND 0.46716f
C16142 VDD.n6893 GND 0.04556f
C16143 VDD.n6894 GND 0.04624f
C16144 VDD.n6895 GND 0.05737f
C16145 VDD.n6896 GND 0.04885f
C16146 VDD.n6897 GND 0.02299f
C16147 VDD.n6898 GND 0.04556f
C16148 VDD.n6899 GND 0.6274f
C16149 VDD.n6900 GND 0.6274f
C16150 VDD.n6901 GND 0.04556f
C16151 VDD.n6902 GND 0.02503f
C16152 VDD.n6903 GND 0.02704f
C16153 VDD.n6904 GND 0.02503f
C16154 VDD.n6905 GND 0.04556f
C16155 VDD.n6906 GND 0.6274f
C16156 VDD.n6907 GND 0.02299f
C16157 VDD.n6908 GND 0.04556f
C16158 VDD.n6909 GND 0.6274f
C16159 VDD.n6910 GND 0.04556f
C16160 VDD.n6911 GND 0.04624f
C16161 VDD.n6912 GND 0.05737f
C16162 VDD.n6913 GND 0.04885f
C16163 VDD.n6914 GND 0.02299f
C16164 VDD.n6915 GND 0.04556f
C16165 VDD.n6916 GND 0.46716f
C16166 VDD.n6917 GND 0.02299f
C16167 VDD.n6918 GND 0.04556f
C16168 VDD.n6919 GND 0.46716f
C16169 VDD.n6920 GND 0.04556f
C16170 VDD.n6921 GND 0.04624f
C16171 VDD.n6922 GND 0.05737f
C16172 VDD.n6923 GND 0.04885f
C16173 VDD.n6924 GND 0.02299f
C16174 VDD.n6925 GND 0.04556f
C16175 VDD.n6926 GND 0.46716f
C16176 VDD.n6927 GND 0.02299f
C16177 VDD.n6928 GND 0.04556f
C16178 VDD.n6929 GND 0.46716f
C16179 VDD.n6930 GND 0.04556f
C16180 VDD.n6931 GND 0.04624f
C16181 VDD.n6932 GND 0.05737f
C16182 VDD.n6933 GND 0.04885f
C16183 VDD.n6934 GND 0.02299f
C16184 VDD.n6935 GND 0.04556f
C16185 VDD.n6936 GND 0.6274f
C16186 VDD.n6937 GND 0.02299f
C16187 VDD.n6938 GND 0.04556f
C16188 VDD.n6939 GND 0.6274f
C16189 VDD.n6940 GND 0.04556f
C16190 VDD.n6941 GND 0.04624f
C16191 VDD.n6942 GND 0.05737f
C16192 VDD.n6943 GND 0.04885f
C16193 VDD.n6944 GND 0.02299f
C16194 VDD.n6945 GND 0.04556f
C16195 VDD.n6946 GND 0.46716f
C16196 VDD.n6947 GND 0.02299f
C16197 VDD.n6948 GND 0.04556f
C16198 VDD.n6949 GND 0.46716f
C16199 VDD.n6950 GND 0.04556f
C16200 VDD.n6951 GND 0.04624f
C16201 VDD.n6952 GND 0.05737f
C16202 VDD.n6953 GND 0.04885f
C16203 VDD.n6954 GND 0.02299f
C16204 VDD.n6955 GND 0.04556f
C16205 VDD.n6956 GND 0.46716f
C16206 VDD.n6957 GND 0.46716f
C16207 VDD.n6958 GND 0.02299f
C16208 VDD.n6959 GND 0.02299f
C16209 VDD.n6960 GND 0.02704f
C16210 VDD.n6961 GND 0.04624f
C16211 VDD.n6962 GND 0.04556f
C16212 VDD.n6963 GND 0.6274f
C16213 VDD.n6964 GND 0.6274f
C16214 VDD.n6965 GND 0.04556f
C16215 VDD.n6966 GND 0.04556f
C16216 VDD.n6967 GND 0.02299f
C16217 VDD.n6968 GND 0.02299f
C16218 VDD.n6969 GND 0.02704f
C16219 VDD.n6970 GND 0.04624f
C16220 VDD.t478 GND 0.57933f
C16221 VDD.n6971 GND 0.04624f
C16222 VDD.n6972 GND 0.05737f
C16223 VDD.n6973 GND 0.02396f
C16224 VDD.n6974 GND 0.12159f
C16225 VDD.t453 GND 0.02128f
C16226 VDD.n6975 GND 0.06662f
C16227 VDD.n6976 GND 0.01638f
C16228 VDD.n6977 GND 0.08322f
C16229 VDD.n6978 GND 0.02503f
C16230 VDD.n6979 GND 0.04556f
C16231 VDD.n6980 GND 0.6274f
C16232 VDD.n6981 GND 0.02299f
C16233 VDD.n6982 GND 0.04556f
C16234 VDD.n6983 GND 0.6274f
C16235 VDD.n6984 GND 0.04556f
C16236 VDD.n6985 GND 0.04624f
C16237 VDD.n6986 GND 0.05737f
C16238 VDD.n6987 GND 0.04885f
C16239 VDD.n6988 GND 0.02299f
C16240 VDD.n6989 GND 0.04556f
C16241 VDD.n6990 GND 0.46716f
C16242 VDD.n6991 GND 0.02299f
C16243 VDD.n6992 GND 0.04556f
C16244 VDD.n6993 GND 0.46716f
C16245 VDD.n6994 GND 0.04556f
C16246 VDD.n6995 GND 0.04624f
C16247 VDD.n6996 GND 0.05737f
C16248 VDD.n6997 GND 0.04885f
C16249 VDD.n6998 GND 0.02299f
C16250 VDD.n6999 GND 0.04556f
C16251 VDD.n7000 GND 0.46716f
C16252 VDD.n7001 GND 0.02299f
C16253 VDD.n7002 GND 0.04556f
C16254 VDD.n7003 GND 0.46716f
C16255 VDD.n7004 GND 0.04556f
C16256 VDD.n7005 GND 0.04624f
C16257 VDD.n7006 GND 0.05737f
C16258 VDD.n7007 GND 0.04885f
C16259 VDD.n7008 GND 0.02299f
C16260 VDD.n7009 GND 0.04556f
C16261 VDD.n7010 GND 0.6274f
C16262 VDD.n7011 GND 0.02299f
C16263 VDD.n7012 GND 0.04556f
C16264 VDD.n7013 GND 0.6274f
C16265 VDD.n7014 GND 0.04556f
C16266 VDD.n7015 GND 0.04624f
C16267 VDD.n7016 GND 0.05737f
C16268 VDD.n7017 GND 0.04885f
C16269 VDD.n7018 GND 0.02299f
C16270 VDD.n7019 GND 0.04556f
C16271 VDD.n7020 GND 0.46716f
C16272 VDD.n7021 GND 0.02299f
C16273 VDD.n7022 GND 0.04556f
C16274 VDD.n7023 GND 0.46716f
C16275 VDD.n7024 GND 0.04556f
C16276 VDD.n7025 GND 0.04624f
C16277 VDD.n7026 GND 0.05737f
C16278 VDD.n7027 GND 0.04885f
C16279 VDD.n7028 GND 0.02299f
C16280 VDD.n7029 GND 0.04556f
C16281 VDD.n7030 GND 0.6274f
C16282 VDD.n7031 GND 0.6274f
C16283 VDD.n7032 GND 0.04556f
C16284 VDD.n7033 GND 0.02503f
C16285 VDD.n7034 GND 0.02704f
C16286 VDD.n7035 GND 0.02503f
C16287 VDD.n7036 GND 0.04556f
C16288 VDD.n7037 GND 0.6274f
C16289 VDD.n7038 GND 0.02299f
C16290 VDD.n7039 GND 0.04556f
C16291 VDD.n7040 GND 0.6274f
C16292 VDD.n7041 GND 0.04556f
C16293 VDD.n7042 GND 0.04624f
C16294 VDD.n7043 GND 0.05737f
C16295 VDD.n7044 GND 0.04885f
C16296 VDD.n7045 GND 0.02299f
C16297 VDD.n7046 GND 0.04556f
C16298 VDD.n7047 GND 0.46716f
C16299 VDD.n7048 GND 0.02299f
C16300 VDD.n7049 GND 0.04556f
C16301 VDD.n7050 GND 0.46716f
C16302 VDD.n7051 GND 0.04556f
C16303 VDD.n7052 GND 0.04624f
C16304 VDD.n7053 GND 0.05737f
C16305 VDD.n7054 GND 0.04885f
C16306 VDD.n7055 GND 0.02299f
C16307 VDD.n7056 GND 0.04556f
C16308 VDD.n7057 GND 0.46716f
C16309 VDD.n7058 GND 0.02299f
C16310 VDD.n7059 GND 0.04556f
C16311 VDD.n7060 GND 0.46716f
C16312 VDD.n7061 GND 0.04556f
C16313 VDD.n7062 GND 0.04624f
C16314 VDD.n7063 GND 0.05737f
C16315 VDD.n7064 GND 0.04885f
C16316 VDD.n7065 GND 0.02299f
C16317 VDD.n7066 GND 0.04556f
C16318 VDD.n7067 GND 0.6274f
C16319 VDD.n7068 GND 0.02299f
C16320 VDD.n7069 GND 0.04556f
C16321 VDD.n7070 GND 0.6274f
C16322 VDD.n7071 GND 0.04556f
C16323 VDD.n7072 GND 0.04624f
C16324 VDD.n7073 GND 0.05737f
C16325 VDD.n7074 GND 0.04885f
C16326 VDD.n7075 GND 0.02299f
C16327 VDD.n7076 GND 0.04556f
C16328 VDD.n7077 GND 0.46716f
C16329 VDD.n7078 GND 0.02299f
C16330 VDD.n7079 GND 0.04556f
C16331 VDD.n7080 GND 0.46716f
C16332 VDD.n7081 GND 0.04556f
C16333 VDD.n7082 GND 0.04624f
C16334 VDD.n7083 GND 0.05737f
C16335 VDD.n7084 GND 0.04885f
C16336 VDD.n7085 GND 0.02299f
C16337 VDD.n7086 GND 0.04556f
C16338 VDD.n7087 GND 0.46716f
C16339 VDD.n7088 GND 0.02299f
C16340 VDD.n7089 GND 0.04556f
C16341 VDD.n7090 GND 0.46716f
C16342 VDD.n7091 GND 0.04556f
C16343 VDD.n7092 GND 0.04624f
C16344 VDD.n7093 GND 0.05737f
C16345 VDD.n7094 GND 0.04885f
C16346 VDD.n7095 GND 0.02299f
C16347 VDD.n7096 GND 0.04556f
C16348 VDD.n7097 GND 0.6274f
C16349 VDD.n7098 GND 0.04556f
C16350 VDD.n7099 GND 0.6274f
C16351 VDD.t755 GND 0.67839f
C16352 VDD.n7101 GND 0.5739f
C16353 VDD.n7102 GND 0.02503f
C16354 VDD.n7103 GND 0.08322f
C16355 VDD.n7104 GND 0.01638f
C16356 VDD.n7105 GND 0.06662f
C16357 VDD.n7106 GND 0.9404f
C16358 VDD.n7107 GND 0.01573f
C16359 VDD.n7108 GND 0.08322f
C16360 VDD.n7110 GND 0.32569f
C16361 VDD.n7111 GND 0.02503f
C16362 VDD.n7112 GND 0.02704f
C16363 VDD.n7113 GND 0.02503f
C16364 VDD.n7114 GND 0.04556f
C16365 VDD.n7115 GND 0.22764f
C16366 VDD.n7116 GND 0.22764f
C16367 VDD.n7117 GND 0.04556f
C16368 VDD.n7118 GND 0.02503f
C16369 VDD.n7119 GND 0.02704f
C16370 VDD.n7120 GND 0.02503f
C16371 VDD.n7121 GND 0.04556f
C16372 VDD.n7122 GND 0.22764f
C16373 VDD.n7123 GND 0.22764f
C16374 VDD.n7124 GND 0.04556f
C16375 VDD.n7125 GND 0.02503f
C16376 VDD.n7126 GND 0.08322f
C16377 VDD.n7127 GND 0.0781f
C16378 VDD.n7128 GND 0.01573f
C16379 VDD.n7129 GND 0.08322f
C16380 VDD.n7131 GND 0.32569f
C16381 VDD.n7132 GND 0.02503f
C16382 VDD.n7133 GND 0.02704f
C16383 VDD.n7134 GND 0.02503f
C16384 VDD.n7135 GND 0.04556f
C16385 VDD.n7136 GND 0.22764f
C16386 VDD.n7137 GND 0.22764f
C16387 VDD.n7138 GND 0.04556f
C16388 VDD.n7139 GND 0.02503f
C16389 VDD.n7140 GND 0.02704f
C16390 VDD.n7141 GND 0.02503f
C16391 VDD.n7142 GND 0.04556f
C16392 VDD.n7143 GND 0.22764f
C16393 VDD.n7144 GND 0.22764f
C16394 VDD.n7145 GND 0.04556f
C16395 VDD.n7146 GND 0.02503f
C16396 VDD.n7147 GND 0.08322f
C16397 VDD.n7148 GND 0.0781f
C16398 VDD.n7149 GND 0.01573f
C16399 VDD.n7150 GND 0.08322f
C16400 VDD.n7152 GND 0.32569f
C16401 VDD.n7153 GND 0.02503f
C16402 VDD.n7154 GND 0.02704f
C16403 VDD.n7155 GND 0.02503f
C16404 VDD.n7156 GND 0.04556f
C16405 VDD.n7157 GND 0.22764f
C16406 VDD.n7158 GND 0.22764f
C16407 VDD.n7159 GND 0.04556f
C16408 VDD.n7160 GND 0.02503f
C16409 VDD.n7161 GND 0.02704f
C16410 VDD.n7162 GND 0.02503f
C16411 VDD.n7163 GND 0.04556f
C16412 VDD.n7164 GND 0.22764f
C16413 VDD.n7165 GND 0.22764f
C16414 VDD.n7166 GND 0.04556f
C16415 VDD.n7167 GND 0.02503f
C16416 VDD.n7168 GND 0.08322f
C16417 VDD.n7169 GND 0.0781f
C16418 VDD.n7170 GND 0.01573f
C16419 VDD.n7171 GND 0.08322f
C16420 VDD.n7173 GND 0.32569f
C16421 VDD.n7174 GND 0.02503f
C16422 VDD.n7175 GND 0.02704f
C16423 VDD.n7176 GND 0.02503f
C16424 VDD.n7177 GND 0.04556f
C16425 VDD.n7178 GND 0.22764f
C16426 VDD.n7179 GND 0.22764f
C16427 VDD.n7180 GND 0.04556f
C16428 VDD.n7181 GND 0.02503f
C16429 VDD.n7182 GND 0.02704f
C16430 VDD.n7183 GND 0.02503f
C16431 VDD.n7184 GND 0.04556f
C16432 VDD.n7185 GND 0.22764f
C16433 VDD.n7186 GND 0.22764f
C16434 VDD.n7187 GND 0.04556f
C16435 VDD.n7188 GND 0.02503f
C16436 VDD.n7189 GND 0.08322f
C16437 VDD.n7190 GND 0.0781f
C16438 VDD.n7191 GND 0.01573f
C16439 VDD.n7192 GND 0.08322f
C16440 VDD.n7194 GND 0.32569f
C16441 VDD.n7195 GND 0.02503f
C16442 VDD.n7196 GND 0.02704f
C16443 VDD.n7197 GND 0.02503f
C16444 VDD.n7198 GND 0.04556f
C16445 VDD.n7199 GND 0.22764f
C16446 VDD.n7200 GND 0.22764f
C16447 VDD.n7201 GND 0.04556f
C16448 VDD.n7202 GND 0.02503f
C16449 VDD.n7203 GND 0.02704f
C16450 VDD.n7204 GND 0.02503f
C16451 VDD.n7205 GND 0.04556f
C16452 VDD.n7206 GND 0.22764f
C16453 VDD.n7207 GND 0.22764f
C16454 VDD.n7208 GND 0.04556f
C16455 VDD.n7209 GND 0.02503f
C16456 VDD.n7210 GND 0.08322f
C16457 VDD.n7211 GND 0.0781f
C16458 VDD.n7212 GND 0.01573f
C16459 VDD.n7213 GND 0.08322f
C16460 VDD.n7215 GND 0.32569f
C16461 VDD.n7216 GND 0.02503f
C16462 VDD.n7217 GND 0.02704f
C16463 VDD.n7218 GND 0.02503f
C16464 VDD.n7219 GND 0.04556f
C16465 VDD.n7220 GND 0.22764f
C16466 VDD.n7221 GND 0.22764f
C16467 VDD.n7222 GND 0.04556f
C16468 VDD.n7223 GND 0.02503f
C16469 VDD.n7224 GND 0.02704f
C16470 VDD.n7225 GND 0.02503f
C16471 VDD.n7226 GND 0.04556f
C16472 VDD.n7227 GND 0.22764f
C16473 VDD.n7228 GND 0.22764f
C16474 VDD.n7229 GND 0.04556f
C16475 VDD.n7230 GND 0.02503f
C16476 VDD.n7231 GND 0.08322f
C16477 VDD.n7232 GND 0.0781f
C16478 VDD.n7233 GND 0.01573f
C16479 VDD.n7234 GND 0.08322f
C16480 VDD.n7236 GND 0.32569f
C16481 VDD.n7237 GND 0.02503f
C16482 VDD.n7238 GND 0.02704f
C16483 VDD.n7239 GND 0.02503f
C16484 VDD.n7240 GND 0.04556f
C16485 VDD.n7241 GND 0.22764f
C16486 VDD.n7242 GND 0.22764f
C16487 VDD.n7243 GND 0.04556f
C16488 VDD.n7244 GND 0.02503f
C16489 VDD.n7245 GND 0.02704f
C16490 VDD.n7246 GND 0.02503f
C16491 VDD.n7247 GND 0.04556f
C16492 VDD.n7248 GND 0.22764f
C16493 VDD.n7249 GND 0.22764f
C16494 VDD.n7250 GND 0.04556f
C16495 VDD.n7251 GND 0.02503f
C16496 VDD.n7252 GND 0.08322f
C16497 VDD.n7253 GND 0.0781f
C16498 VDD.n7254 GND 0.01573f
C16499 VDD.n7255 GND 0.08322f
C16500 VDD.n7257 GND 0.32569f
C16501 VDD.n7258 GND 0.02503f
C16502 VDD.n7259 GND 0.02704f
C16503 VDD.n7260 GND 0.02503f
C16504 VDD.n7261 GND 0.04556f
C16505 VDD.n7262 GND 0.22764f
C16506 VDD.n7263 GND 0.22764f
C16507 VDD.n7264 GND 0.04556f
C16508 VDD.n7265 GND 0.02503f
C16509 VDD.n7266 GND 0.02704f
C16510 VDD.n7267 GND 0.02503f
C16511 VDD.n7268 GND 0.04556f
C16512 VDD.n7269 GND 0.22764f
C16513 VDD.n7270 GND 0.22764f
C16514 VDD.n7271 GND 0.04556f
C16515 VDD.n7272 GND 0.02503f
C16516 VDD.n7273 GND 0.08322f
C16517 VDD.n7274 GND 0.42619f
C16518 VDD.n7275 GND 0.83549f
C16519 VDD.t43 GND 1.47626f
C16520 VDD.t45 GND 1.47626f
C16521 VDD.n7276 GND 0.83058f
C16522 VDD.t884 GND 1.85633f
C16523 VDD.n7277 GND 0.4649f
C16524 VDD.n7278 GND 0.24011f
C16525 VDD.n7279 GND 0.20697f
C16526 VDD.n7280 GND 0.24788f
C16527 VDD.n7281 GND 0.2251f
C16528 VDD.n7282 GND 0.42965f
C16529 VDD.n7283 GND 3.79486f
C16530 VDD.t883 GND 4.87495f
C16531 VDD.n7284 GND 0.51282f
C16532 VDD.n7285 GND 1.5196f
C16533 VDD.n7286 GND 0.24938f
C16534 VDD.n7287 GND 0.40375f
C16535 VDD.n7289 GND 3.64032f
C16536 VDD.n7290 GND 0.29413f
C16537 VDD.n7291 GND 0.30011f
C16538 VDD.n7292 GND 0.29413f
C16539 VDD.n7293 GND 0.50861f
C16540 VDD.n7294 GND 6.25502f
C16541 VDD.n7295 GND 6.25502f
C16542 VDD.n7296 GND 0.40865f
C16543 VDD.n7297 GND 0.2251f
C16544 VDD.n7298 GND 0.24788f
C16545 VDD.n7299 GND 3.53645f
C16546 VDD.n7300 GND 0.22728f
C16547 VDD.t42 GND 3.95625f
C16548 VDD.n7302 GND 0.22728f
C16549 VDD.n7303 GND 0.13298f
C16550 VDD.n7304 GND 0.13223f
C16551 VDD.n7305 GND 0.13298f
C16552 VDD.n7306 GND 0.22728f
C16553 VDD.t44 GND 3.79486f
C16554 VDD.n7307 GND 0.22728f
C16555 VDD.n7308 GND 0.20697f
C16556 VDD.n7309 GND 0.17665f
C16557 VDD.n7310 GND 0.06416f
C16558 VDD.n7311 GND 0.13559f
C16559 VDD.n7312 GND 0.95867f
C16560 VDD.n7313 GND 1.35274f
C16561 VDD.n7314 GND 0.46498f
C16562 VDD.n7315 GND 1.01318f
C16563 VDD.n7316 GND 5.58872f
C16564 VDD.n7317 GND 6.61419f
C16565 VDD.n7318 GND 7.77316f
C16566 VDD.n7319 GND 1.9565f
C16567 VDD.n7320 GND 1.63616f
C16568 VDD.n7321 GND 0.80951f
C16569 VDD.n7322 GND 0.49254f
C16570 VDD.n7323 GND 1.07656f
C16571 VDD.n7324 GND 4.54112f
C16572 VDD.n7325 GND 4.35649f
C16573 VDD.n7326 GND 3.94958f
C16574 VDD.n7327 GND 0.93302f
C16575 VDD.n7328 GND 0.41396f
C16576 VDD.n7329 GND 1.04097f
C16577 VDD.n7330 GND 0.83835f
C16578 VDD.t728 GND 0.23053f
C16579 VDD.n7331 GND 2.08406f
C16580 VDD.n7332 GND 0.59333f
C16581 VDD.n7333 GND 0.11704f
C16582 CDAC_v3_0.switch_8.Z.t1 GND 0.09736f
C16583 CDAC_v3_0.switch_8.Z.t4 GND 0.09736f
C16584 CDAC_v3_0.switch_8.Z.n0 GND 0.34968f
C16585 CDAC_v3_0.switch_8.Z.n1 GND 1.07811f
C16586 CDAC_v3_0.switch_8.Z.n2 GND 0.10087f
C16587 CDAC_v3_0.switch_8.Z.t2 GND 24.2603f
C16588 CDAC_v3_0.switch_8.Z.n3 GND 10.09f
C16589 CDAC_v3_0.switch_8.Z.n4 GND 0.03204f
C16590 CDAC_v3_0.switch_8.Z.t0 GND 0.0943f
C16591 CDAC_v3_0.switch_8.Z.n5 GND 0.20705f
C16592 CDAC_v3_0.switch_8.Z.t3 GND 0.09411f
C16593 Q0.t7 GND 0.16953f
C16594 Q0.t9 GND 0.32734f
C16595 Q0.n0 GND 0.24301f
C16596 Q0.n1 GND 0.04497f
C16597 Q0.t4 GND 0.16953f
C16598 Q0.t6 GND 0.32734f
C16599 Q0.n2 GND 0.24149f
C16600 Q0.n3 GND 0.04844f
C16601 Q0.n4 GND 0.07131f
C16602 Q0.n5 GND 2.48828f
C16603 Q0.t1 GND 0.0425f
C16604 Q0.n6 GND 0.20844f
C16605 Q0.n7 GND 0.0475f
C16606 Q0.t3 GND 0.04512f
C16607 Q0.t2 GND 0.0442f
C16608 Q0.n8 GND 0.25136f
C16609 Q0.n9 GND 0.08202f
C16610 Q0.t0 GND 0.0442f
C16611 Q0.n10 GND 0.06808f
C16612 Q0.n11 GND 0.12055f
C16613 Q0.n12 GND 0.04755f
C16614 Q0.t5 GND 0.32586f
C16615 Q0.n13 GND 0.09519f
C16616 Q0.n14 GND 0.0413f
C16617 Q0.n15 GND 0.1816f
C16618 Q0.t8 GND 0.15155f
C16619 Q0.n16 GND 0.46052f
C16620 Q0.n17 GND 1.11843f
C16621 EN.t104 GND 0.45234f
C16622 EN.n0 GND 0.14601f
C16623 EN.t17 GND 0.23461f
C16624 EN.n1 GND 0.0505f
C16625 EN.n2 GND 0.03015f
C16626 EN.n3 GND 0.27984f
C16627 EN.t73 GND 0.45234f
C16628 EN.n4 GND 0.14601f
C16629 EN.t99 GND 0.23461f
C16630 EN.n5 GND 0.0505f
C16631 EN.n6 GND 0.03015f
C16632 EN.n8 GND 0.63823f
C16633 EN.t36 GND 0.45321f
C16634 EN.n9 GND 0.19532f
C16635 EN.t28 GND 0.21077f
C16636 EN.n10 GND 0.42365f
C16637 EN.n11 GND 0.12042f
C16638 EN.t47 GND 0.45123f
C16639 EN.n12 GND 0.13182f
C16640 EN.n13 GND 0.04376f
C16641 EN.n14 GND 0.07393f
C16642 EN.t23 GND 0.23462f
C16643 EN.n15 GND 0.21886f
C16644 EN.n16 GND 0.04847f
C16645 EN.t48 GND 0.45123f
C16646 EN.n17 GND 0.13182f
C16647 EN.n18 GND 0.04376f
C16648 EN.n19 GND 0.07393f
C16649 EN.n20 GND 0.27984f
C16650 EN.t42 GND 0.45125f
C16651 EN.n21 GND 0.46786f
C16652 EN.n22 GND 0.05062f
C16653 EN.n23 GND 0.06758f
C16654 EN.t87 GND 0.21077f
C16655 EN.n24 GND 0.42365f
C16656 EN.n25 GND 0.12042f
C16657 EN.n26 GND 0.71089f
C16658 EN.n28 GND 0.04847f
C16659 EN.n29 GND 0.21886f
C16660 EN.t10 GND 1.16452f
C16661 EN.t5 GND 1.16469f
C16662 EN.n30 GND 0.10307f
C16663 EN.t92 GND 0.45123f
C16664 EN.n31 GND 0.09445f
C16665 EN.n32 GND 0.07603f
C16666 EN.n33 GND 0.27984f
C16667 EN.t89 GND 0.23471f
C16668 EN.n34 GND 0.10307f
C16669 EN.t66 GND 0.45123f
C16670 EN.n35 GND 0.09445f
C16671 EN.n36 GND 0.07603f
C16672 EN.n38 GND 0.71062f
C16673 EN.n39 GND 0.49693f
C16674 EN.n40 GND 0.27368f
C16675 EN.n41 GND 0.27064f
C16676 EN.n42 GND 0.12042f
C16677 EN.t37 GND 0.45123f
C16678 EN.n43 GND 0.19654f
C16679 EN.t80 GND 0.21059f
C16680 EN.n44 GND 0.13677f
C16681 EN.n45 GND 7.30175f
C16682 EN.n46 GND 6.37487f
C16683 EN.t20 GND 0.45234f
C16684 EN.n47 GND 0.14601f
C16685 EN.t102 GND 0.23461f
C16686 EN.n48 GND 0.0505f
C16687 EN.n49 GND 0.03015f
C16688 EN.n50 GND 0.27984f
C16689 EN.t1 GND 0.45234f
C16690 EN.n51 GND 0.14601f
C16691 EN.t72 GND 0.23461f
C16692 EN.n52 GND 0.0505f
C16693 EN.n53 GND 0.03015f
C16694 EN.n55 GND 0.72631f
C16695 EN.n56 GND 0.11416f
C16696 EN.n57 GND 0.25524f
C16697 EN.n58 GND 0.12042f
C16698 EN.t22 GND 0.45123f
C16699 EN.n59 GND 0.19654f
C16700 EN.t93 GND 0.21059f
C16701 EN.n60 GND 0.13677f
C16702 EN.n61 GND 6.83455f
C16703 EN.n62 GND 5.95015f
C16704 EN.t38 GND 0.45234f
C16705 EN.n63 GND 0.14601f
C16706 EN.t30 GND 0.23461f
C16707 EN.n64 GND 0.0505f
C16708 EN.n65 GND 0.03015f
C16709 EN.n66 GND 0.27984f
C16710 EN.t21 GND 0.45234f
C16711 EN.n67 GND 0.14601f
C16712 EN.t7 GND 0.23461f
C16713 EN.n68 GND 0.0505f
C16714 EN.n69 GND 0.03015f
C16715 EN.n71 GND 0.72631f
C16716 EN.n72 GND 0.11416f
C16717 EN.n73 GND 0.25524f
C16718 EN.n74 GND 0.12042f
C16719 EN.t100 GND 0.45123f
C16720 EN.n75 GND 0.19654f
C16721 EN.t43 GND 0.21059f
C16722 EN.n76 GND 0.13677f
C16723 EN.n77 GND 6.36735f
C16724 EN.n78 GND 5.52542f
C16725 EN.t16 GND 0.45234f
C16726 EN.n79 GND 0.14601f
C16727 EN.t3 GND 0.23461f
C16728 EN.n80 GND 0.0505f
C16729 EN.n81 GND 0.03015f
C16730 EN.n82 GND 0.27984f
C16731 EN.t98 GND 0.45234f
C16732 EN.n83 GND 0.14601f
C16733 EN.t83 GND 0.23461f
C16734 EN.n84 GND 0.0505f
C16735 EN.n85 GND 0.03015f
C16736 EN.n87 GND 0.72631f
C16737 EN.n88 GND 0.11416f
C16738 EN.n89 GND 0.25524f
C16739 EN.n90 GND 0.12042f
C16740 EN.t18 GND 0.45123f
C16741 EN.n91 GND 0.19654f
C16742 EN.t86 GND 0.21059f
C16743 EN.n92 GND 0.13677f
C16744 EN.n93 GND 5.90015f
C16745 EN.n94 GND 5.10069f
C16746 EN.t101 GND 0.45234f
C16747 EN.n95 GND 0.14601f
C16748 EN.t85 GND 0.23461f
C16749 EN.n96 GND 0.0505f
C16750 EN.n97 GND 0.03015f
C16751 EN.n98 GND 0.27984f
C16752 EN.t71 GND 0.45234f
C16753 EN.n99 GND 0.14601f
C16754 EN.t59 GND 0.23461f
C16755 EN.n100 GND 0.0505f
C16756 EN.n101 GND 0.03015f
C16757 EN.n103 GND 0.72631f
C16758 EN.n104 GND 0.11416f
C16759 EN.n105 GND 0.25524f
C16760 EN.n106 GND 0.12042f
C16761 EN.t8 GND 0.45123f
C16762 EN.n107 GND 0.19654f
C16763 EN.t78 GND 0.21059f
C16764 EN.n108 GND 0.13677f
C16765 EN.n109 GND 5.43295f
C16766 EN.n110 GND 4.67596f
C16767 EN.t29 GND 0.45234f
C16768 EN.n111 GND 0.14601f
C16769 EN.t106 GND 0.23461f
C16770 EN.n112 GND 0.0505f
C16771 EN.n113 GND 0.03015f
C16772 EN.n114 GND 0.27984f
C16773 EN.t6 GND 0.45234f
C16774 EN.n115 GND 0.14601f
C16775 EN.t75 GND 0.23461f
C16776 EN.n116 GND 0.0505f
C16777 EN.n117 GND 0.03015f
C16778 EN.n119 GND 0.72631f
C16779 EN.n120 GND 0.11416f
C16780 EN.n121 GND 0.25524f
C16781 EN.n122 GND 0.12042f
C16782 EN.t9 GND 0.45123f
C16783 EN.n123 GND 0.19654f
C16784 EN.t57 GND 0.21059f
C16785 EN.n124 GND 0.13677f
C16786 EN.n125 GND 4.96575f
C16787 EN.n126 GND 4.25124f
C16788 EN.t91 GND 0.45234f
C16789 EN.n127 GND 0.14601f
C16790 EN.t77 GND 0.23461f
C16791 EN.n128 GND 0.0505f
C16792 EN.n129 GND 0.03015f
C16793 EN.n130 GND 0.27984f
C16794 EN.t65 GND 0.45234f
C16795 EN.n131 GND 0.14601f
C16796 EN.t54 GND 0.23461f
C16797 EN.n132 GND 0.0505f
C16798 EN.n133 GND 0.03015f
C16799 EN.n135 GND 0.72631f
C16800 EN.n136 GND 0.11416f
C16801 EN.n137 GND 0.25524f
C16802 EN.n138 GND 0.12042f
C16803 EN.t4 GND 0.45123f
C16804 EN.n139 GND 0.19654f
C16805 EN.t69 GND 0.21059f
C16806 EN.n140 GND 0.13677f
C16807 EN.n141 GND 4.49855f
C16808 EN.n142 GND 3.82651f
C16809 EN.t84 GND 0.45234f
C16810 EN.n143 GND 0.14601f
C16811 EN.t12 GND 0.23461f
C16812 EN.n144 GND 0.0505f
C16813 EN.n145 GND 0.03015f
C16814 EN.n146 GND 0.27984f
C16815 EN.t58 GND 0.45234f
C16816 EN.n147 GND 0.14601f
C16817 EN.t95 GND 0.23461f
C16818 EN.n148 GND 0.0505f
C16819 EN.n149 GND 0.03015f
C16820 EN.n151 GND 0.72631f
C16821 EN.n152 GND 0.11416f
C16822 EN.n153 GND 0.25524f
C16823 EN.n154 GND 0.12042f
C16824 EN.t27 GND 0.45123f
C16825 EN.n155 GND 0.19654f
C16826 EN.t62 GND 0.21059f
C16827 EN.n156 GND 0.13677f
C16828 EN.n157 GND 4.03135f
C16829 EN.n158 GND 3.40178f
C16830 EN.t32 GND 0.45234f
C16831 EN.n159 GND 0.14601f
C16832 EN.t68 GND 0.23461f
C16833 EN.n160 GND 0.0505f
C16834 EN.n161 GND 0.03015f
C16835 EN.n162 GND 0.27984f
C16836 EN.t14 GND 0.45234f
C16837 EN.n163 GND 0.14601f
C16838 EN.t51 GND 0.23461f
C16839 EN.n164 GND 0.0505f
C16840 EN.n165 GND 0.03015f
C16841 EN.n167 GND 0.72631f
C16842 EN.n168 GND 0.11416f
C16843 EN.n169 GND 0.25524f
C16844 EN.n170 GND 0.12042f
C16845 EN.t107 GND 0.45123f
C16846 EN.n171 GND 0.19654f
C16847 EN.t61 GND 0.21059f
C16848 EN.n172 GND 0.13677f
C16849 EN.n173 GND 3.56415f
C16850 EN.n174 GND 2.97706f
C16851 EN.t76 GND 0.45234f
C16852 EN.n175 GND 0.14601f
C16853 EN.t60 GND 0.23461f
C16854 EN.n176 GND 0.0505f
C16855 EN.n177 GND 0.03015f
C16856 EN.n178 GND 0.27984f
C16857 EN.t53 GND 0.45234f
C16858 EN.n179 GND 0.14601f
C16859 EN.t49 GND 0.23461f
C16860 EN.n180 GND 0.0505f
C16861 EN.n181 GND 0.03015f
C16862 EN.n183 GND 0.72631f
C16863 EN.n184 GND 0.11416f
C16864 EN.n185 GND 0.25524f
C16865 EN.n186 GND 0.12042f
C16866 EN.t96 GND 0.45123f
C16867 EN.n187 GND 0.19654f
C16868 EN.t55 GND 0.21059f
C16869 EN.n188 GND 0.13677f
C16870 EN.n189 GND 3.09696f
C16871 EN.n190 GND 2.55233f
C16872 EN.t11 GND 0.45234f
C16873 EN.n191 GND 0.14601f
C16874 EN.t19 GND 0.23461f
C16875 EN.n192 GND 0.0505f
C16876 EN.n193 GND 0.03015f
C16877 EN.n194 GND 0.27984f
C16878 EN.t94 GND 0.45234f
C16879 EN.n195 GND 0.14601f
C16880 EN.t105 GND 0.23461f
C16881 EN.n196 GND 0.0505f
C16882 EN.n197 GND 0.03015f
C16883 EN.n199 GND 0.72631f
C16884 EN.n200 GND 0.11416f
C16885 EN.n201 GND 0.25524f
C16886 EN.n202 GND 0.12042f
C16887 EN.t2 GND 0.45123f
C16888 EN.n203 GND 0.19654f
C16889 EN.t46 GND 0.21059f
C16890 EN.n204 GND 0.13677f
C16891 EN.n205 GND 2.62976f
C16892 EN.n206 GND 2.1276f
C16893 EN.t0 GND 0.45234f
C16894 EN.n207 GND 0.14601f
C16895 EN.t88 GND 0.23461f
C16896 EN.n208 GND 0.0505f
C16897 EN.n209 GND 0.03015f
C16898 EN.n210 GND 0.27984f
C16899 EN.t79 GND 0.45234f
C16900 EN.n211 GND 0.14601f
C16901 EN.t63 GND 0.23461f
C16902 EN.n212 GND 0.0505f
C16903 EN.n213 GND 0.03015f
C16904 EN.n215 GND 0.72631f
C16905 EN.n216 GND 0.11416f
C16906 EN.n217 GND 0.25524f
C16907 EN.n218 GND 0.12042f
C16908 EN.t15 GND 0.45123f
C16909 EN.n219 GND 0.19654f
C16910 EN.t82 GND 0.21059f
C16911 EN.n220 GND 0.13677f
C16912 EN.n221 GND 2.16256f
C16913 EN.n222 GND 1.70288f
C16914 EN.t97 GND 0.45234f
C16915 EN.n223 GND 0.14601f
C16916 EN.t81 GND 0.23461f
C16917 EN.n224 GND 0.0505f
C16918 EN.n225 GND 0.03015f
C16919 EN.n226 GND 0.27984f
C16920 EN.t70 GND 0.45234f
C16921 EN.n227 GND 0.14601f
C16922 EN.t56 GND 0.23461f
C16923 EN.n228 GND 0.0505f
C16924 EN.n229 GND 0.03015f
C16925 EN.n231 GND 0.72631f
C16926 EN.n232 GND 0.11416f
C16927 EN.n233 GND 0.25524f
C16928 EN.n234 GND 0.12042f
C16929 EN.t25 GND 0.45123f
C16930 EN.n235 GND 0.19654f
C16931 EN.t74 GND 0.21059f
C16932 EN.n236 GND 0.13677f
C16933 EN.n237 GND 1.69536f
C16934 EN.n238 GND 1.27815f
C16935 EN.t39 GND 0.45234f
C16936 EN.n239 GND 0.14601f
C16937 EN.t31 GND 0.23461f
C16938 EN.n240 GND 0.0505f
C16939 EN.n241 GND 0.03015f
C16940 EN.n242 GND 0.27984f
C16941 EN.t24 GND 0.45234f
C16942 EN.n243 GND 0.14601f
C16943 EN.t13 GND 0.23461f
C16944 EN.n244 GND 0.0505f
C16945 EN.n245 GND 0.03015f
C16946 EN.n247 GND 0.72631f
C16947 EN.n248 GND 0.11416f
C16948 EN.n249 GND 0.25524f
C16949 EN.n250 GND 0.12042f
C16950 EN.t52 GND 0.45123f
C16951 EN.n251 GND 0.19654f
C16952 EN.t103 GND 0.21059f
C16953 EN.n252 GND 0.13677f
C16954 EN.n253 GND 1.22816f
C16955 EN.n254 GND 0.85342f
C16956 EN.t67 GND 0.45234f
C16957 EN.n255 GND 0.14601f
C16958 EN.t45 GND 0.23461f
C16959 EN.n256 GND 0.0505f
C16960 EN.n257 GND 0.03015f
C16961 EN.n258 GND 0.27984f
C16962 EN.t50 GND 0.45234f
C16963 EN.n259 GND 0.14601f
C16964 EN.t33 GND 0.23461f
C16965 EN.n260 GND 0.0505f
C16966 EN.n261 GND 0.03015f
C16967 EN.n263 GND 0.72631f
C16968 EN.n264 GND 0.11416f
C16969 EN.n265 GND 0.25524f
C16970 EN.n266 GND 0.12042f
C16971 EN.t41 GND 0.45123f
C16972 EN.n267 GND 0.19654f
C16973 EN.t34 GND 0.21059f
C16974 EN.n268 GND 0.13677f
C16975 EN.n269 GND 0.76096f
C16976 EN.n270 GND 0.42869f
C16977 EN.t90 GND 0.45234f
C16978 EN.n271 GND 0.14601f
C16979 EN.t40 GND 0.23461f
C16980 EN.n272 GND 0.0505f
C16981 EN.n273 GND 0.03015f
C16982 EN.n274 GND 0.27984f
C16983 EN.t64 GND 0.45234f
C16984 EN.n275 GND 0.14601f
C16985 EN.t26 GND 0.23461f
C16986 EN.n276 GND 0.0505f
C16987 EN.n277 GND 0.03015f
C16988 EN.n279 GND 0.72631f
C16989 EN.n280 GND 0.11416f
C16990 EN.n281 GND 0.25524f
C16991 EN.n282 GND 0.12042f
C16992 EN.t35 GND 0.45123f
C16993 EN.n283 GND 0.19654f
C16994 EN.t44 GND 0.21059f
C16995 EN.n284 GND 0.13638f
C16996 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t2 GND 0.04916f
C16997 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n0 GND 0.12652f
C16998 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n1 GND 0.10289f
C16999 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t4 GND 0.19589f
C17000 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t7 GND 0.37676f
C17001 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n2 GND 0.08939f
C17002 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n3 GND 0.08866f
C17003 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n4 GND 0.15046f
C17004 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n5 GND 0.112f
C17005 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t6 GND 0.37841f
C17006 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n6 GND 0.16309f
C17007 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t5 GND 0.18751f
C17008 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t1 GND 0.0511f
C17009 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n7 GND 0.32233f
C17010 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t0 GND 0.05217f
C17011 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.t3 GND 0.0511f
C17012 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n8 GND 0.29063f
C17013 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n9 GND 0.10073f
C17014 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.C.n10 GND 0.06269f
C17015 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t4 GND 0.48439f
C17016 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n0 GND 0.21098f
C17017 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t5 GND 0.24285f
C17018 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t3 GND 0.0657f
C17019 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n1 GND 0.41359f
C17020 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t2 GND 0.06708f
C17021 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t1 GND 0.0657f
C17022 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n2 GND 0.37365f
C17023 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n3 GND 0.12192f
C17024 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n4 GND 0.01546f
C17025 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n5 GND 0.0204f
C17026 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t6 GND 0.48632f
C17027 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t7 GND 0.25185f
C17028 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n6 GND 0.36445f
C17029 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n7 GND 0.14399f
C17030 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.t0 GND 0.06705f
C17031 Ring_Counter_0.D_FlipFlop_0.3-input-nand_2.Vout.n8 GND 0.23153f
.ends

