** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-12_21-01-12/parameters/DNL/run_1/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.494117647 8.5u 0.494117647 8.500001u 0.495882352875 17.0u 0.495882352875 17.000001u 0.49764705875 25.5u
+ 0.49764705875 25.500001u 0.499411764625 34.0u 0.499411764625 34.000001u 0.5011764705 42.5u 0.5011764705 42.500001u 0.502941176375 51.0u
+ 0.502941176375 51.000001u 0.50470588225 59.5u 0.50470588225 59.500001u 0.506470588125 68.0u 0.506470588125 68.000001u 0.508235294 76.5u
+ 0.508235294 76.500001u 0.51 85.0u 0.51 85.000001u 0.511764705875 93.5u 0.511764705875 93.500001u 0.51352941175 102.0u 0.51352941175
+ 102.000001u 0.515294117625 110.5u 0.515294117625 110.500001u 0.5170588235 119.0u 0.5170588235 119.000001u 0.518823529375 127.5u
+ 0.518823529375 127.500001u 0.52058823525 136.0u 0.52058823525 136.000001u 0.522352941125 144.5u 0.522352941125 144.500001u 0.524117647 153.0u
+ 0.524117647 153.000001u 0.525882352875 161.5u 0.525882352875 161.500001u 0.52764705875 170.0u 0.52764705875 170.000001u 0.529411764625 178.5u
+ 0.529411764625)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_1
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ss

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 178.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-12_21-01-12/parameters/DNL/run_1/sar_output_dnl_1.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
