magic
tech sky130A
magscale 1 2
timestamp 1757220954
<< metal3 >>
rect 274 -435 334 -399
rect -54 -763 1378 -435
rect -54 -823 1414 -763
rect -54 -1479 1378 -823
rect -90 -1539 1378 -1479
rect -54 -1867 1378 -1539
rect 990 -1903 1050 -1867
<< mimcap >>
rect -26 -503 1350 -463
rect -26 -1799 14 -503
rect 1310 -1799 1350 -503
rect -26 -1839 1350 -1799
<< mimcapcontact >>
rect 14 -1799 1310 -503
<< metal4 >>
rect 632 -502 692 -398
rect 13 -503 1311 -502
rect 13 -1121 14 -503
rect -90 -1181 14 -1121
rect 13 -1799 14 -1181
rect 1310 -1121 1311 -503
rect 1310 -1181 1414 -1121
rect 1310 -1799 1311 -1181
rect 13 -1800 1311 -1799
rect 632 -1904 692 -1800
<< end >>
