magic
tech sky130A
magscale 1 2
timestamp 1761392116
<< nwell >>
rect 0 -882 8762 928
<< pwell >>
rect 0 978 8762 1782
rect 0 -1736 8762 -932
<< metal1 >>
rect 0 1831 8762 1845
rect 0 1779 33 1831
rect 85 1779 8762 1831
rect 0 1765 8762 1779
rect 349 985 395 1204
rect 340 979 404 985
rect 340 927 346 979
rect 398 927 404 979
rect 340 921 404 927
rect 1698 979 1762 985
rect 1698 927 1704 979
rect 1756 927 1762 979
rect 1698 921 1762 927
rect 2578 979 2658 993
rect 2578 927 2592 979
rect 2644 927 2658 979
rect 349 672 395 921
rect 2578 913 2658 927
rect 3670 979 3734 985
rect 3670 927 3676 979
rect 3728 927 3734 979
rect 3670 921 3734 927
rect 6652 979 6732 993
rect 6652 927 6666 979
rect 6718 927 6732 979
rect 6652 913 6732 927
rect 7744 979 7808 985
rect 7744 927 7750 979
rect 7802 927 7808 979
rect 7744 921 7808 927
rect 3056 859 3120 865
rect 3056 807 3062 859
rect 3114 807 3120 859
rect 3056 801 3120 807
rect 7130 859 7194 865
rect 7130 807 7136 859
rect 7188 807 7194 859
rect 7130 801 7194 807
rect 4550 738 4630 752
rect 4550 686 4564 738
rect 4616 686 4630 738
rect 4550 672 4630 686
rect 5764 738 5844 752
rect 5764 686 5778 738
rect 5830 686 5844 738
rect 5764 672 5844 686
rect 450 409 530 423
rect 450 357 464 409
rect 516 357 530 409
rect 450 343 530 357
rect 4394 409 4474 423
rect 4394 357 4408 409
rect 4460 357 4474 409
rect 4394 343 4474 357
rect 8468 409 8548 423
rect 8468 357 8482 409
rect 8534 357 8548 409
rect 8468 343 8548 357
rect 1108 288 1188 302
rect 1108 236 1122 288
rect 1174 236 1188 288
rect 1108 222 1188 236
rect 2304 288 2384 302
rect 2304 236 2318 288
rect 2370 236 2384 288
rect 2304 222 2384 236
rect 4244 288 4324 302
rect 4244 236 4258 288
rect 4310 236 4324 288
rect 4244 222 4324 236
rect 6378 288 6458 302
rect 6378 236 6392 288
rect 6444 236 6458 288
rect 6378 222 6458 236
rect 8318 288 8398 302
rect 8318 236 8332 288
rect 8384 236 8398 288
rect 8318 222 8398 236
rect 0 -17 8762 63
rect 1108 -190 1188 -176
rect 1108 -242 1122 -190
rect 1174 -242 1188 -190
rect 1108 -256 1188 -242
rect 2304 -190 2384 -176
rect 2304 -242 2318 -190
rect 2370 -242 2384 -190
rect 2304 -256 2384 -242
rect 4244 -190 4324 -176
rect 4244 -242 4258 -190
rect 4310 -242 4324 -190
rect 4244 -256 4324 -242
rect 6378 -190 6458 -176
rect 6378 -242 6392 -190
rect 6444 -242 6458 -190
rect 6378 -256 6458 -242
rect 8318 -190 8398 -176
rect 8318 -242 8332 -190
rect 8384 -242 8398 -190
rect 8318 -256 8398 -242
rect 4394 -311 4474 -297
rect 4394 -363 4408 -311
rect 4460 -363 4474 -311
rect 4394 -377 4474 -363
rect 8468 -311 8548 -297
rect 8468 -363 8482 -311
rect 8534 -363 8548 -311
rect 8468 -377 8548 -363
rect 4550 -640 4630 -626
rect 4550 -692 4564 -640
rect 4616 -692 4630 -640
rect 4550 -706 4630 -692
rect 5764 -640 5844 -626
rect 5764 -692 5778 -640
rect 5830 -692 5844 -640
rect 5764 -706 5844 -692
rect 3056 -761 3120 -755
rect 3056 -813 3062 -761
rect 3114 -813 3120 -761
rect 3056 -819 3120 -813
rect 7130 -761 7194 -755
rect 7130 -813 7136 -761
rect 7188 -813 7194 -761
rect 7130 -819 7194 -813
rect 1698 -881 1762 -875
rect 1698 -933 1704 -881
rect 1756 -933 1762 -881
rect 1698 -939 1762 -933
rect 2578 -881 2658 -867
rect 2578 -933 2592 -881
rect 2644 -933 2658 -881
rect 2578 -947 2658 -933
rect 3670 -881 3734 -875
rect 3670 -933 3676 -881
rect 3728 -933 3734 -881
rect 3670 -939 3734 -933
rect 5294 -881 5374 -867
rect 5294 -933 5308 -881
rect 5360 -933 5374 -881
rect 5294 -947 5374 -933
rect 6386 -881 6450 -875
rect 6386 -933 6392 -881
rect 6444 -933 6450 -881
rect 6386 -939 6450 -933
rect 6652 -881 6732 -867
rect 6652 -933 6666 -881
rect 6718 -933 6732 -881
rect 6652 -947 6732 -933
rect 7744 -881 7808 -875
rect 7744 -933 7750 -881
rect 7802 -933 7808 -881
rect 7744 -939 7808 -933
rect 2304 -1092 2384 -1078
rect 2304 -1144 2318 -1092
rect 2370 -1144 2384 -1092
rect 2304 -1158 2384 -1144
rect 5020 -1092 5100 -1078
rect 5020 -1144 5034 -1092
rect 5086 -1144 5100 -1092
rect 5020 -1158 5100 -1144
rect 0 -1733 8762 -1719
rect 0 -1785 33 -1733
rect 85 -1785 8762 -1733
rect 0 -1799 8762 -1785
<< via1 >>
rect 33 1779 85 1831
rect 346 927 398 979
rect 1704 927 1756 979
rect 2592 927 2644 979
rect 3676 927 3728 979
rect 6666 927 6718 979
rect 7750 927 7802 979
rect 3062 807 3114 859
rect 7136 807 7188 859
rect 4564 686 4616 738
rect 5778 686 5830 738
rect 464 357 516 409
rect 4408 357 4460 409
rect 8482 357 8534 409
rect 1122 236 1174 288
rect 2318 236 2370 288
rect 4258 236 4310 288
rect 6392 236 6444 288
rect 8332 236 8384 288
rect 1122 -242 1174 -190
rect 2318 -242 2370 -190
rect 4258 -242 4310 -190
rect 6392 -242 6444 -190
rect 8332 -242 8384 -190
rect 4408 -363 4460 -311
rect 8482 -363 8534 -311
rect 4564 -692 4616 -640
rect 5778 -692 5830 -640
rect 3062 -813 3114 -761
rect 7136 -813 7188 -761
rect 1704 -933 1756 -881
rect 2592 -933 2644 -881
rect 3676 -933 3728 -881
rect 5308 -933 5360 -881
rect 6392 -933 6444 -881
rect 6666 -933 6718 -881
rect 7750 -933 7802 -881
rect 2318 -1144 2370 -1092
rect 5034 -1144 5086 -1092
rect 33 -1785 85 -1733
<< metal2 >>
rect 19 1833 99 1845
rect 19 1777 31 1833
rect 87 1777 99 1833
rect 19 1765 99 1777
rect 332 979 1770 993
rect 332 927 346 979
rect 398 927 1704 979
rect 1756 927 1770 979
rect 332 913 1770 927
rect 2578 979 3742 993
rect 2578 927 2592 979
rect 2644 927 3676 979
rect 3728 927 3742 979
rect 2578 913 3742 927
rect 6652 979 7816 993
rect 6652 927 6666 979
rect 6718 927 7750 979
rect 7802 927 7816 979
rect 6652 913 7816 927
rect 1247 861 7202 873
rect 1247 805 1259 861
rect 1315 859 7202 861
rect 1315 807 3062 859
rect 3114 807 7136 859
rect 7188 807 7202 859
rect 1315 805 7202 807
rect 1247 793 7202 805
rect 4550 738 5844 752
rect 4550 686 4564 738
rect 4616 686 5778 738
rect 5830 686 5844 738
rect 4550 672 5844 686
rect 450 411 642 423
rect 450 409 574 411
rect 450 357 464 409
rect 516 357 574 409
rect 450 355 574 357
rect 630 355 642 411
rect 450 343 642 355
rect 4394 411 4474 423
rect 4394 355 4406 411
rect 4462 355 4474 411
rect 4394 343 4474 355
rect 8468 411 8548 423
rect 8468 355 8480 411
rect 8536 355 8548 411
rect 8468 343 8548 355
rect 1108 290 1476 302
rect 1108 288 1408 290
rect 1108 236 1122 288
rect 1174 236 1408 288
rect 1108 234 1408 236
rect 1464 234 1476 290
rect 1108 222 1476 234
rect 2304 290 2384 302
rect 2304 234 2316 290
rect 2372 234 2384 290
rect 2304 222 2384 234
rect 4244 290 4324 302
rect 4244 234 4256 290
rect 4312 234 4324 290
rect 4244 222 4324 234
rect 6378 290 6458 302
rect 6378 234 6390 290
rect 6446 234 6458 290
rect 6378 222 6458 234
rect 8318 290 8398 302
rect 8318 234 8330 290
rect 8386 234 8398 290
rect 8318 222 8398 234
rect 1108 -188 1327 -176
rect 1108 -190 1259 -188
rect 1108 -242 1122 -190
rect 1174 -242 1259 -190
rect 1108 -244 1259 -242
rect 1315 -244 1327 -188
rect 1108 -256 1327 -244
rect 2304 -188 2384 -176
rect 2304 -244 2316 -188
rect 2372 -244 2384 -188
rect 2304 -256 2384 -244
rect 4244 -188 4474 -176
rect 4244 -190 4406 -188
rect 4244 -242 4258 -190
rect 4310 -242 4406 -190
rect 4244 -244 4406 -242
rect 4462 -244 4474 -188
rect 4244 -256 4474 -244
rect 6378 -188 6458 -176
rect 6378 -244 6390 -188
rect 6446 -244 6458 -188
rect 6378 -256 6458 -244
rect 8318 -188 8548 -176
rect 8318 -190 8480 -188
rect 8318 -242 8332 -190
rect 8384 -242 8480 -190
rect 8318 -244 8480 -242
rect 8536 -244 8548 -188
rect 8318 -256 8548 -244
rect 4244 -309 4474 -297
rect 4244 -365 4256 -309
rect 4312 -311 4474 -309
rect 4312 -363 4408 -311
rect 4460 -363 4474 -311
rect 4312 -365 4474 -363
rect 4244 -377 4474 -365
rect 8318 -309 8548 -297
rect 8318 -365 8330 -309
rect 8386 -311 8548 -309
rect 8386 -363 8482 -311
rect 8534 -363 8548 -311
rect 8386 -365 8548 -363
rect 8318 -377 8548 -365
rect 4550 -640 5844 -626
rect 4550 -692 4564 -640
rect 4616 -692 5778 -640
rect 5830 -692 5844 -640
rect 4550 -706 5844 -692
rect 1396 -759 7202 -747
rect 1396 -815 1408 -759
rect 1464 -761 7202 -759
rect 1464 -813 3062 -761
rect 3114 -813 7136 -761
rect 7188 -813 7202 -761
rect 1464 -815 7202 -813
rect 1396 -827 7202 -815
rect 562 -879 1770 -867
rect 562 -935 574 -879
rect 630 -881 1770 -879
rect 630 -933 1704 -881
rect 1756 -933 1770 -881
rect 630 -935 1770 -933
rect 562 -947 1770 -935
rect 2578 -881 3742 -867
rect 2578 -933 2592 -881
rect 2644 -933 3676 -881
rect 3728 -933 3742 -881
rect 2578 -947 3742 -933
rect 5294 -881 6458 -867
rect 5294 -933 5308 -881
rect 5360 -933 6392 -881
rect 6444 -933 6458 -881
rect 5294 -947 6458 -933
rect 6652 -881 7816 -867
rect 6652 -933 6666 -881
rect 6718 -933 7750 -881
rect 7802 -933 7816 -881
rect 6652 -947 7816 -933
rect 2304 -1092 5100 -1078
rect 2304 -1144 2318 -1092
rect 2370 -1144 5034 -1092
rect 5086 -1144 5100 -1092
rect 2304 -1158 5100 -1144
rect 19 -1731 99 -1719
rect 19 -1787 31 -1731
rect 87 -1787 99 -1731
rect 19 -1799 99 -1787
<< via2 >>
rect 31 1831 87 1833
rect 31 1779 33 1831
rect 33 1779 85 1831
rect 85 1779 87 1831
rect 31 1777 87 1779
rect 1259 805 1315 861
rect 574 355 630 411
rect 4406 409 4462 411
rect 4406 357 4408 409
rect 4408 357 4460 409
rect 4460 357 4462 409
rect 4406 355 4462 357
rect 8480 409 8536 411
rect 8480 357 8482 409
rect 8482 357 8534 409
rect 8534 357 8536 409
rect 8480 355 8536 357
rect 1408 234 1464 290
rect 2316 288 2372 290
rect 2316 236 2318 288
rect 2318 236 2370 288
rect 2370 236 2372 288
rect 2316 234 2372 236
rect 4256 288 4312 290
rect 4256 236 4258 288
rect 4258 236 4310 288
rect 4310 236 4312 288
rect 4256 234 4312 236
rect 6390 288 6446 290
rect 6390 236 6392 288
rect 6392 236 6444 288
rect 6444 236 6446 288
rect 6390 234 6446 236
rect 8330 288 8386 290
rect 8330 236 8332 288
rect 8332 236 8384 288
rect 8384 236 8386 288
rect 8330 234 8386 236
rect 1259 -244 1315 -188
rect 2316 -190 2372 -188
rect 2316 -242 2318 -190
rect 2318 -242 2370 -190
rect 2370 -242 2372 -190
rect 2316 -244 2372 -242
rect 4406 -244 4462 -188
rect 6390 -190 6446 -188
rect 6390 -242 6392 -190
rect 6392 -242 6444 -190
rect 6444 -242 6446 -190
rect 6390 -244 6446 -242
rect 8480 -244 8536 -188
rect 4256 -365 4312 -309
rect 8330 -365 8386 -309
rect 1408 -815 1464 -759
rect 574 -935 630 -879
rect 31 -1733 87 -1731
rect 31 -1785 33 -1733
rect 33 -1785 85 -1733
rect 85 -1785 87 -1733
rect 31 -1787 87 -1785
<< metal3 >>
rect 26 1833 92 1838
rect 26 1777 31 1833
rect 87 1777 92 1833
rect 26 1772 92 1777
rect 29 -1726 89 1772
rect 1254 861 1320 866
rect 1254 805 1259 861
rect 1315 805 1320 861
rect 1254 800 1320 805
rect 569 411 635 416
rect 569 355 574 411
rect 630 355 635 411
rect 569 350 635 355
rect 572 -874 632 350
rect 1257 -183 1317 800
rect 4401 411 4467 416
rect 4401 355 4406 411
rect 4462 355 4467 411
rect 4401 350 4467 355
rect 8475 411 8541 416
rect 8475 355 8480 411
rect 8536 355 8541 411
rect 8475 350 8541 355
rect 1403 290 1469 295
rect 1403 234 1408 290
rect 1464 234 1469 290
rect 1403 229 1469 234
rect 2311 290 2377 295
rect 2311 234 2316 290
rect 2372 234 2377 290
rect 2311 229 2377 234
rect 4251 290 4317 295
rect 4251 234 4256 290
rect 4312 234 4317 290
rect 4251 229 4317 234
rect 1254 -188 1320 -183
rect 1254 -244 1259 -188
rect 1315 -244 1320 -188
rect 1254 -249 1320 -244
rect 1406 -754 1466 229
rect 2314 -183 2374 229
rect 2311 -188 2377 -183
rect 2311 -244 2316 -188
rect 2372 -244 2377 -188
rect 2311 -249 2377 -244
rect 4254 -304 4314 229
rect 4404 -183 4464 350
rect 6385 290 6451 295
rect 6385 234 6390 290
rect 6446 234 6451 290
rect 6385 229 6451 234
rect 8325 290 8391 295
rect 8325 234 8330 290
rect 8386 234 8391 290
rect 8325 229 8391 234
rect 6388 -183 6448 229
rect 4401 -188 4467 -183
rect 4401 -244 4406 -188
rect 4462 -244 4467 -188
rect 4401 -249 4467 -244
rect 6385 -188 6451 -183
rect 6385 -244 6390 -188
rect 6446 -244 6451 -188
rect 6385 -249 6451 -244
rect 8328 -304 8388 229
rect 8478 -183 8538 350
rect 8475 -188 8541 -183
rect 8475 -244 8480 -188
rect 8536 -244 8541 -188
rect 8475 -249 8541 -244
rect 4251 -309 4317 -304
rect 4251 -365 4256 -309
rect 4312 -365 4317 -309
rect 4251 -370 4317 -365
rect 8325 -309 8391 -304
rect 8325 -365 8330 -309
rect 8386 -365 8391 -309
rect 8325 -370 8391 -365
rect 1403 -759 1469 -754
rect 1403 -815 1408 -759
rect 1464 -815 1469 -759
rect 1403 -820 1469 -815
rect 569 -879 635 -874
rect 569 -935 574 -879
rect 630 -935 635 -879
rect 569 -940 635 -935
rect 26 -1731 92 -1726
rect 26 -1787 31 -1731
rect 87 -1787 92 -1731
rect 26 -1792 92 -1787
use 3-input-nand  3-input-nand_0
timestamp 1761375837
transform 1 0 -1279 0 -1 400
box 2023 -1445 3995 417
use 3-input-nand  3-input-nand_1
timestamp 1761375837
transform 1 0 -1279 0 1 -354
box 2023 -1445 3995 417
use 3-input-nand  3-input-nand_2
timestamp 1761375837
transform 1 0 693 0 -1 400
box 2023 -1445 3995 417
use 3-input-nand  3-input-nand_3
timestamp 1761375837
transform 1 0 693 0 1 -354
box 2023 -1445 3995 417
use 3-input-nand  3-input-nand_4
timestamp 1761375837
transform 1 0 4767 0 -1 400
box 2023 -1445 3995 417
use 3-input-nand  3-input-nand_5
timestamp 1761375837
transform 1 0 4767 0 1 -354
box 2023 -1445 3995 417
use Inverter  Inverter_0
timestamp 1761294637
transform 1 0 -1366 0 -1 942
box 1366 -903 2110 959
use Inverter  Inverter_1
timestamp 1761294637
transform 1 0 3322 0 1 -896
box 1366 -903 2110 959
use Nand_Gate  Nand_Gate_0
timestamp 1761392116
transform 1 0 3526 0 -1 1298
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_1
timestamp 1761392116
transform 1 0 3526 0 1 -1252
box 1906 -547 3264 1315
<< labels >>
flabel metal1 349 672 395 1204 0 FreeSans 160 0 0 0 D
port 1 nsew
flabel metal3 1406 -759 1466 239 0 FreeSans 160 90 0 0 nCLR
port 3 nsew
flabel metal1 0 0 8762 46 0 FreeSans 160 0 0 0 VDD
port 7 nsew
flabel metal1 0 1782 8762 1828 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal3 1257 -193 1317 805 0 FreeSans 160 90 0 0 nPRE
port 4 nsew
flabel metal3 2314 -205 2374 239 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 8478 -188 8538 355 0 FreeSans 160 0 0 0 Q
port 6 nsew
flabel metal3 8328 -309 8388 234 0 FreeSans 160 0 0 0 Qbar
port 5 nsew
<< end >>
