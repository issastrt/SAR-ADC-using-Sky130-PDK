magic
tech sky130A
magscale 1 2
timestamp 1761294637
<< nwell >>
rect 1366 892 2110 896
rect 1366 14 1408 892
rect 2068 14 2110 892
<< mvpsubdiff >>
rect 1414 -118 1474 -84
rect 2002 -118 2062 -84
rect 1414 -144 1448 -118
rect 1414 -758 1448 -732
rect 2028 -144 2062 -118
rect 2028 -758 2062 -732
rect 1414 -792 1474 -758
rect 2002 -792 2062 -758
<< mvpsubdiffcont >>
rect 1474 -118 2002 -84
rect 1414 -732 1448 -144
rect 2028 -732 2062 -144
rect 1474 -792 2002 -758
<< locali >>
rect 1582 936 1894 942
rect 1582 902 1588 936
rect 1888 902 1894 936
rect 1582 784 1894 902
rect 1414 -118 1474 -84
rect 2002 -118 2062 -84
rect 1414 -144 1448 -118
rect 1414 -758 1448 -732
rect 2028 -144 2062 -118
rect 2028 -758 2062 -732
rect 1414 -792 1474 -758
rect 2002 -792 2062 -758
rect 1510 -846 1966 -792
rect 1510 -880 1516 -846
rect 1960 -880 1966 -846
rect 1510 -886 1966 -880
<< viali >>
rect 1588 902 1888 936
rect 1516 -880 1960 -846
<< metal1 >>
rect 1366 936 2110 959
rect 1366 902 1588 936
rect 1888 902 2110 936
rect 1366 879 2110 902
rect 1496 599 1576 879
rect 1666 640 1810 720
rect 1496 519 1660 599
rect 1580 311 1660 519
rect 1816 391 1896 599
rect 1816 311 2052 391
rect 1666 190 1810 270
rect 1698 -182 1778 190
rect 1594 -262 1882 -182
rect 1972 -294 2052 311
rect 1508 -502 1588 -294
rect 1424 -582 1588 -502
rect 1888 -374 2052 -294
rect 1888 -582 1968 -374
rect 1424 -823 1504 -582
rect 1594 -694 1882 -614
rect 1366 -846 2110 -823
rect 1366 -880 1516 -846
rect 1960 -880 2110 -846
rect 1366 -903 2110 -880
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1757220954
transform 1 0 1738 0 1 455
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM2
timestamp 1757220954
transform 1 0 1738 0 1 -438
box -372 -402 372 402
<< labels >>
flabel metal1 1366 -886 2110 -840 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 1972 -374 2052 391 0 FreeSans 160 0 0 0 Vout
port 3 nsew
flabel metal1 1366 879 2110 959 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 1698 -262 1778 270 0 FreeSans 160 0 0 0 Vin
port 2 nsew
<< end >>
