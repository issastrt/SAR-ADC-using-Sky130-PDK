** sch_path: /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-03_11-29-22/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0 8.5u 0 8.500001u 0.001764705875 17u 0.001764705875 17.000001u 0.00352941175 25.5u 0.00352941175 25.500001u
+ 0.005294117625 34u 0.005294117625 34.000001u 0.0070588235 42.5u 0.0070588235 42.500001u 0.008823529375 51u 0.008823529375 51.000001u
+ 0.01058823525 59.5u 0.01058823525 59.500001u 0.012352941125 68u 0.012352941125 68.000001u 0.014117647 76.5u 0.014117647 76.500001u
+ 0.015882352875 85u 0.015882352875 85.000001u 0.01764705875 93.5u 0.01764705875 93.500001u 0.019411764625 102u 0.019411764625 102.000001u
+ 0.0211764705 110.5u 0.0211764705 110.500001u 0.022941176375 119u 0.022941176375 119.000001u 0.02470588225 127.5u 0.02470588225 127.500001u
+ 0.026470588125 136u 0.026470588125 136.000001u 0.028235294 144.5u 0.028235294 144.500001u 0.03 153u 0.03 153.000001u 0.031764705875 161.5u
+ 0.031764705875 161.500001u 0.03352941175 170u 0.03352941175 170.000001u 0.035294117625 178.5u 0.035294117625 178.500001u 0.0370588235 187u
+ 0.0370588235 187.000001u 0.038823529375 195.5u 0.038823529375 195.500001u 0.04058823525 204u 0.04058823525 204.000001u 0.042352941125 212.5u
+ 0.042352941125 212.500001u 0.044117647 221u 0.044117647 221.000001u 0.045882352875 229.5u 0.045882352875 229.500001u 0.04764705875 238u
+ 0.04764705875 238.000001u 0.049411764625 246.5u 0.049411764625 246.500001u 0.0511764705 255u 0.0511764705 255.000001u 0.052941176375 263.5u
+ 0.052941176375 263.500001u 0.05470588225 272u 0.05470588225 272.000001u 0.056470588125 280.5u 0.056470588125 280.500001u 0.058235294 289u
+ 0.058235294 289.000001u 0.06 297.5u 0.06 297.500001u 0.061764705875 306u 0.061764705875 306.000001u 0.06352941175 314.5u 0.06352941175
+ 314.500001u 0.065294117625 323u 0.065294117625 323.000001u 0.0670588235 331.5u 0.0670588235 331.500001u 0.068823529375 340u 0.068823529375)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/madra/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 340u uic
  wrdata /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-03_11-29-22/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
