magic
tech sky130A
magscale 1 2
timestamp 1761401821
<< nwell >>
rect -2503 49987 -2429 50061
rect 6259 49987 6333 50061
rect 15021 49987 15095 50061
rect 23783 49987 23857 50061
rect 32545 49987 32619 50061
rect 12794 46139 12868 46213
rect 16738 46139 16812 46213
rect 20682 46139 20756 46213
rect 24626 46139 24700 46213
rect 28570 46139 28644 46213
rect 32514 46139 32588 46213
rect 36458 46139 36532 46213
<< mvnsubdiff >>
rect -2436 49995 -2429 50061
rect 6326 49995 6333 50061
rect 15088 49995 15095 50061
rect 23850 49995 23857 50061
rect 32612 49995 32619 50061
<< metal1 >>
rect 50621 55861 50685 55867
rect 50621 55809 50627 55861
rect 50679 55809 50685 55861
rect 50621 55803 50685 55809
rect -12812 53576 57722 53590
rect -12812 53524 -12798 53576
rect -12746 53524 57656 53576
rect 57708 53524 57722 53576
rect -12812 53510 57722 53524
rect -7188 53337 -7108 53351
rect -7188 53285 -7174 53337
rect -7122 53285 -7108 53337
rect -7188 53271 -7108 53285
rect -6574 53337 -6494 53351
rect -6574 53285 -6560 53337
rect -6508 53285 -6494 53337
rect -6574 53271 -6494 53285
rect 1574 53337 1654 53351
rect 1574 53285 1588 53337
rect 1640 53285 1654 53337
rect 1574 53271 1654 53285
rect 2188 53337 2268 53351
rect 2188 53285 2202 53337
rect 2254 53285 2268 53337
rect 2188 53271 2268 53285
rect 10336 53337 10416 53351
rect 10336 53285 10350 53337
rect 10402 53285 10416 53337
rect 10336 53271 10416 53285
rect 10950 53337 11030 53351
rect 10950 53285 10964 53337
rect 11016 53285 11030 53337
rect 10950 53271 11030 53285
rect 19098 53337 19178 53351
rect 19098 53285 19112 53337
rect 19164 53285 19178 53337
rect 19098 53271 19178 53285
rect 19712 53337 19792 53351
rect 19712 53285 19726 53337
rect 19778 53285 19792 53337
rect 19712 53271 19792 53285
rect 27860 53337 27940 53351
rect 27860 53285 27874 53337
rect 27926 53285 27940 53337
rect 27860 53271 27940 53285
rect 28474 53337 28554 53351
rect 28474 53285 28488 53337
rect 28540 53285 28554 53337
rect 28474 53271 28554 53285
rect 36622 53337 36702 53351
rect 36622 53285 36636 53337
rect 36688 53285 36702 53337
rect 36622 53271 36702 53285
rect 37236 53337 37316 53351
rect 37236 53285 37250 53337
rect 37302 53285 37316 53337
rect 37236 53271 37316 53285
rect 45384 53337 45464 53351
rect 45384 53285 45398 53337
rect 45450 53285 45464 53337
rect 45384 53271 45464 53285
rect 45998 53337 46078 53351
rect 45998 53285 46012 53337
rect 46064 53285 46078 53337
rect 45998 53271 46078 53285
rect 54146 53337 54226 53351
rect 54146 53285 54160 53337
rect 54212 53285 54226 53337
rect 54146 53271 54226 53285
rect 54760 53336 54840 53350
rect 54760 53284 54774 53336
rect 54826 53284 54840 53336
rect 54760 53270 54840 53284
rect -11327 52887 -11247 52901
rect -11327 52835 -11313 52887
rect -11261 52835 -11247 52887
rect -11327 52821 -11247 52835
rect -2565 52887 -2485 52901
rect -2565 52835 -2551 52887
rect -2499 52835 -2485 52887
rect -2565 52821 -2485 52835
rect 6197 52887 6277 52901
rect 6197 52835 6211 52887
rect 6263 52835 6277 52887
rect 6197 52821 6277 52835
rect 14959 52887 15039 52901
rect 14959 52835 14973 52887
rect 15025 52835 15039 52887
rect 14959 52821 15039 52835
rect 23721 52887 23801 52901
rect 23721 52835 23735 52887
rect 23787 52835 23801 52887
rect 23721 52821 23801 52835
rect 32483 52887 32563 52901
rect 32483 52835 32497 52887
rect 32549 52835 32563 52887
rect 32483 52821 32563 52835
rect 41245 52887 41325 52901
rect 41245 52835 41259 52887
rect 41311 52835 41325 52887
rect 41245 52821 41325 52835
rect 50007 52887 50087 52901
rect 50007 52835 50021 52887
rect 50073 52835 50087 52887
rect 50007 52821 50087 52835
rect -11933 52646 -11869 52652
rect -11933 52594 -11927 52646
rect -11875 52594 -11869 52646
rect -11933 52588 -11869 52594
rect -7462 52646 -7382 52660
rect -7462 52594 -7448 52646
rect -7396 52594 -7382 52646
rect -7462 52580 -7382 52594
rect -3171 52646 -3107 52652
rect -3171 52594 -3165 52646
rect -3113 52594 -3107 52646
rect -3171 52588 -3107 52594
rect 1300 52646 1380 52660
rect 1300 52594 1314 52646
rect 1366 52594 1380 52646
rect 1300 52580 1380 52594
rect 5591 52646 5655 52652
rect 5591 52594 5597 52646
rect 5649 52594 5655 52646
rect 5591 52588 5655 52594
rect 10062 52646 10142 52660
rect 10062 52594 10076 52646
rect 10128 52594 10142 52646
rect 10062 52580 10142 52594
rect 14353 52646 14417 52652
rect 14353 52594 14359 52646
rect 14411 52594 14417 52646
rect 14353 52588 14417 52594
rect 18824 52646 18904 52660
rect 18824 52594 18838 52646
rect 18890 52594 18904 52646
rect 18824 52580 18904 52594
rect 23115 52646 23179 52652
rect 23115 52594 23121 52646
rect 23173 52594 23179 52646
rect 23115 52588 23179 52594
rect 27586 52646 27666 52660
rect 27586 52594 27600 52646
rect 27652 52594 27666 52646
rect 27586 52580 27666 52594
rect 31877 52646 31941 52652
rect 31877 52594 31883 52646
rect 31935 52594 31941 52646
rect 31877 52588 31941 52594
rect 36348 52646 36428 52660
rect 36348 52594 36362 52646
rect 36414 52594 36428 52646
rect 36348 52580 36428 52594
rect 40639 52646 40703 52652
rect 40639 52594 40645 52646
rect 40697 52594 40703 52646
rect 40639 52588 40703 52594
rect 45110 52646 45190 52660
rect 45110 52594 45124 52646
rect 45176 52594 45190 52646
rect 45110 52580 45190 52594
rect 49401 52646 49465 52652
rect 49401 52594 49407 52646
rect 49459 52594 49465 52646
rect 49401 52588 49465 52594
rect 53872 52646 53952 52660
rect 53872 52594 53886 52646
rect 53938 52594 53952 52646
rect 53872 52580 53952 52594
rect -10360 52340 -10280 52354
rect -10360 52288 -10346 52340
rect -10294 52288 -10280 52340
rect -10360 52274 -10280 52288
rect -1598 52340 -1518 52354
rect -1598 52288 -1584 52340
rect -1532 52288 -1518 52340
rect -1598 52274 -1518 52288
rect 7164 52340 7244 52354
rect 7164 52288 7178 52340
rect 7230 52288 7244 52340
rect 7164 52274 7244 52288
rect 15926 52340 16006 52354
rect 15926 52288 15940 52340
rect 15992 52288 16006 52340
rect 15926 52274 16006 52288
rect 24688 52340 24768 52354
rect 24688 52288 24702 52340
rect 24754 52288 24768 52340
rect 24688 52274 24768 52288
rect 33450 52340 33530 52354
rect 33450 52288 33464 52340
rect 33516 52288 33530 52340
rect 33450 52274 33530 52288
rect 42212 52340 42292 52354
rect 42212 52288 42226 52340
rect 42278 52288 42292 52340
rect 42212 52274 42292 52288
rect 50974 52340 51054 52354
rect 50974 52288 50988 52340
rect 51040 52288 51054 52340
rect 50974 52274 51054 52288
rect -12957 51754 57585 51791
rect -12957 51702 -12940 51754
rect -12888 51702 57516 51754
rect 57568 51702 57585 51754
rect -12957 51648 57585 51702
rect -10360 51505 -10280 51519
rect -10360 51453 -10346 51505
rect -10294 51453 -10280 51505
rect -10360 51439 -10280 51453
rect -1598 51505 -1518 51519
rect -1598 51453 -1584 51505
rect -1532 51453 -1518 51505
rect -1598 51439 -1518 51453
rect 7164 51505 7244 51519
rect 7164 51453 7178 51505
rect 7230 51453 7244 51505
rect 7164 51439 7244 51453
rect 15926 51505 16006 51519
rect 15926 51453 15940 51505
rect 15992 51453 16006 51505
rect 15926 51439 16006 51453
rect 24688 51505 24768 51519
rect 24688 51453 24702 51505
rect 24754 51453 24768 51505
rect 24688 51439 24768 51453
rect 33450 51505 33530 51519
rect 33450 51453 33464 51505
rect 33516 51453 33530 51505
rect 33450 51439 33530 51453
rect 42212 51505 42292 51519
rect 42212 51453 42226 51505
rect 42278 51453 42292 51505
rect 42212 51439 42292 51453
rect 50974 51505 51054 51519
rect 50974 51453 50988 51505
rect 51040 51453 51054 51505
rect 50974 51439 51054 51453
rect -12332 50971 -12252 50985
rect -12332 50919 -12318 50971
rect -12266 50919 -12252 50971
rect -12332 50905 -12252 50919
rect -3570 50971 -3490 50985
rect -3570 50919 -3556 50971
rect -3504 50919 -3490 50971
rect -3570 50905 -3490 50919
rect 5192 50971 5272 50985
rect 5192 50919 5206 50971
rect 5258 50919 5272 50971
rect 5192 50905 5272 50919
rect 13954 50971 14034 50985
rect 13954 50919 13968 50971
rect 14020 50919 14034 50971
rect 13954 50905 14034 50919
rect 22716 50971 22796 50985
rect 22716 50919 22730 50971
rect 22782 50919 22796 50971
rect 22716 50905 22796 50919
rect 31478 50971 31558 50985
rect 31478 50919 31492 50971
rect 31544 50919 31558 50971
rect 31478 50905 31558 50919
rect 40240 50971 40320 50985
rect 40240 50919 40254 50971
rect 40306 50919 40320 50971
rect 40240 50905 40320 50919
rect 49002 50971 49082 50985
rect 49002 50919 49016 50971
rect 49068 50919 49082 50971
rect 49002 50905 49082 50919
rect 49002 50171 49082 50185
rect 49002 50119 49016 50171
rect 49068 50119 49082 50171
rect 49002 50105 49082 50119
rect -12812 49932 -12664 49946
rect -12812 49880 -12798 49932
rect -12746 49880 -12664 49932
rect -12812 49866 -12664 49880
rect 57431 49932 57722 49946
rect 57431 49880 57656 49932
rect 57708 49880 57722 49932
rect 57431 49866 57722 49880
rect 51721 49693 51795 49704
rect 51721 49641 51732 49693
rect 51784 49641 51795 49693
rect 51721 49630 51795 49641
rect 57432 48150 57582 48164
rect 57432 48098 57516 48150
rect 57568 48098 57582 48150
rect 57432 48084 57582 48098
rect -12812 47012 57722 47026
rect -12812 46960 -12798 47012
rect -12746 46960 50241 47012
rect 50293 46960 55673 47012
rect 55725 46960 57656 47012
rect 57708 46960 57722 47012
rect -12812 46946 57722 46960
rect 8855 46202 8919 46208
rect 8855 46150 8861 46202
rect 8913 46150 8919 46202
rect 12799 46202 12863 46208
rect 12799 46199 12805 46202
rect 12794 46153 12805 46199
rect 8855 46144 8919 46150
rect 12799 46150 12805 46153
rect 12857 46199 12863 46202
rect 16743 46202 16807 46208
rect 16743 46199 16749 46202
rect 12857 46153 12868 46199
rect 16738 46153 16749 46199
rect 12857 46150 12863 46153
rect 12799 46144 12863 46150
rect 16743 46150 16749 46153
rect 16801 46199 16807 46202
rect 20687 46202 20751 46208
rect 20687 46199 20693 46202
rect 16801 46153 16812 46199
rect 20682 46153 20693 46199
rect 16801 46150 16807 46153
rect 16743 46144 16807 46150
rect 20687 46150 20693 46153
rect 20745 46199 20751 46202
rect 24631 46202 24695 46208
rect 24631 46199 24637 46202
rect 20745 46153 20756 46199
rect 24626 46153 24637 46199
rect 20745 46150 20751 46153
rect 20687 46144 20751 46150
rect 24631 46150 24637 46153
rect 24689 46199 24695 46202
rect 28575 46202 28639 46208
rect 28575 46199 28581 46202
rect 24689 46153 24700 46199
rect 28570 46153 28581 46199
rect 24689 46150 24695 46153
rect 24631 46144 24695 46150
rect 28575 46150 28581 46153
rect 28633 46199 28639 46202
rect 32519 46202 32583 46208
rect 32519 46199 32525 46202
rect 28633 46153 28644 46199
rect 32514 46153 32525 46199
rect 28633 46150 28639 46153
rect 28575 46144 28639 46150
rect 32519 46150 32525 46153
rect 32577 46199 32583 46202
rect 36463 46202 36527 46208
rect 36463 46199 36469 46202
rect 32577 46153 32588 46199
rect 36458 46153 36469 46199
rect 32577 46150 32583 46153
rect 32519 46144 32583 46150
rect 36463 46150 36469 46153
rect 36521 46199 36527 46202
rect 36521 46153 36532 46199
rect 36521 46150 36527 46153
rect 36463 46144 36527 46150
rect -12954 45230 57582 45244
rect -12954 45178 -12940 45230
rect -12888 45178 57516 45230
rect 57568 45178 57582 45230
rect -12954 45164 57582 45178
rect 50227 42090 50307 42104
rect 50227 42038 50241 42090
rect 50293 42038 50307 42090
rect 50227 42024 50307 42038
rect 55659 42090 55739 42104
rect 55659 42038 55673 42090
rect 55725 42038 55739 42090
rect 55659 42024 55739 42038
rect 50226 10356 55345 10402
<< via1 >>
rect 50627 55809 50679 55861
rect -12798 53524 -12746 53576
rect 57656 53524 57708 53576
rect -7174 53285 -7122 53337
rect -6560 53285 -6508 53337
rect 1588 53285 1640 53337
rect 2202 53285 2254 53337
rect 10350 53285 10402 53337
rect 10964 53285 11016 53337
rect 19112 53285 19164 53337
rect 19726 53285 19778 53337
rect 27874 53285 27926 53337
rect 28488 53285 28540 53337
rect 36636 53285 36688 53337
rect 37250 53285 37302 53337
rect 45398 53285 45450 53337
rect 46012 53285 46064 53337
rect 54160 53285 54212 53337
rect 54774 53284 54826 53336
rect -11313 52835 -11261 52887
rect -2551 52835 -2499 52887
rect 6211 52835 6263 52887
rect 14973 52835 15025 52887
rect 23735 52835 23787 52887
rect 32497 52835 32549 52887
rect 41259 52835 41311 52887
rect 50021 52835 50073 52887
rect -11927 52594 -11875 52646
rect -7448 52594 -7396 52646
rect -3165 52594 -3113 52646
rect 1314 52594 1366 52646
rect 5597 52594 5649 52646
rect 10076 52594 10128 52646
rect 14359 52594 14411 52646
rect 18838 52594 18890 52646
rect 23121 52594 23173 52646
rect 27600 52594 27652 52646
rect 31883 52594 31935 52646
rect 36362 52594 36414 52646
rect 40645 52594 40697 52646
rect 45124 52594 45176 52646
rect 49407 52594 49459 52646
rect 53886 52594 53938 52646
rect -10346 52288 -10294 52340
rect -1584 52288 -1532 52340
rect 7178 52288 7230 52340
rect 15940 52288 15992 52340
rect 24702 52288 24754 52340
rect 33464 52288 33516 52340
rect 42226 52288 42278 52340
rect 50988 52288 51040 52340
rect -12940 51702 -12888 51754
rect 57516 51702 57568 51754
rect -10346 51453 -10294 51505
rect -1584 51453 -1532 51505
rect 7178 51453 7230 51505
rect 15940 51453 15992 51505
rect 24702 51453 24754 51505
rect 33464 51453 33516 51505
rect 42226 51453 42278 51505
rect 50988 51453 51040 51505
rect -12318 50919 -12266 50971
rect -3556 50919 -3504 50971
rect 5206 50919 5258 50971
rect 13968 50919 14020 50971
rect 22730 50919 22782 50971
rect 31492 50919 31544 50971
rect 40254 50919 40306 50971
rect 49016 50919 49068 50971
rect 49016 50119 49068 50171
rect -12798 49880 -12746 49932
rect 57656 49880 57708 49932
rect 51732 49641 51784 49693
rect 57516 48098 57568 48150
rect -12798 46960 -12746 47012
rect 50241 46960 50293 47012
rect 55673 46960 55725 47012
rect 57656 46960 57708 47012
rect 8861 46150 8913 46202
rect 12805 46150 12857 46202
rect 16749 46150 16801 46202
rect 20693 46150 20745 46202
rect 24637 46150 24689 46202
rect 28581 46150 28633 46202
rect 32525 46150 32577 46202
rect 36469 46150 36521 46202
rect -12940 45178 -12888 45230
rect 57516 45178 57568 45230
rect 50241 42038 50293 42090
rect 55673 42038 55725 42090
<< metal2 >>
rect -12954 62966 -7874 62978
rect -12954 62910 -12942 62966
rect -12886 62910 -7874 62966
rect -12954 62898 -7874 62910
rect 51941 61738 57722 61750
rect 51941 61682 51953 61738
rect 52009 61682 57654 61738
rect 57710 61682 57722 61738
rect 51941 61670 57722 61682
rect -12812 61589 -7214 61601
rect -12812 61533 -12800 61589
rect -12744 61533 -7282 61589
rect -7226 61533 -7214 61589
rect -12812 61521 -7214 61533
rect 50613 55863 50693 55875
rect 50613 55807 50625 55863
rect 50681 55807 50693 55863
rect 50613 55795 50693 55807
rect -12812 53578 -12732 53590
rect -12812 53522 -12800 53578
rect -12744 53522 -12732 53578
rect -12812 53510 -12732 53522
rect 57642 53576 57722 53590
rect 57642 53524 57656 53576
rect 57708 53524 57722 53576
rect 57642 53510 57722 53524
rect -7188 53339 -7108 53351
rect -7188 53283 -7176 53339
rect -7120 53283 -7108 53339
rect -7188 53271 -7108 53283
rect -6574 53339 -6494 53351
rect -6574 53283 -6562 53339
rect -6506 53283 -6494 53339
rect -6574 53271 -6494 53283
rect 1574 53339 1654 53351
rect 1574 53283 1586 53339
rect 1642 53283 1654 53339
rect 1574 53271 1654 53283
rect 2188 53339 2268 53351
rect 2188 53283 2200 53339
rect 2256 53283 2268 53339
rect 2188 53271 2268 53283
rect 10336 53339 10416 53351
rect 10336 53283 10348 53339
rect 10404 53283 10416 53339
rect 10336 53271 10416 53283
rect 10950 53339 11030 53351
rect 10950 53283 10962 53339
rect 11018 53283 11030 53339
rect 10950 53271 11030 53283
rect 19098 53339 19178 53351
rect 19098 53283 19110 53339
rect 19166 53283 19178 53339
rect 19098 53271 19178 53283
rect 19712 53339 19792 53351
rect 19712 53283 19724 53339
rect 19780 53283 19792 53339
rect 19712 53271 19792 53283
rect 27860 53339 27940 53351
rect 27860 53283 27872 53339
rect 27928 53283 27940 53339
rect 27860 53271 27940 53283
rect 28474 53339 28554 53351
rect 28474 53283 28486 53339
rect 28542 53283 28554 53339
rect 28474 53271 28554 53283
rect 36622 53339 36702 53351
rect 36622 53283 36634 53339
rect 36690 53283 36702 53339
rect 36622 53271 36702 53283
rect 37236 53339 37316 53351
rect 37236 53283 37248 53339
rect 37304 53283 37316 53339
rect 37236 53271 37316 53283
rect 45384 53339 45464 53351
rect 45384 53283 45396 53339
rect 45452 53283 45464 53339
rect 45384 53271 45464 53283
rect 45998 53339 46078 53351
rect 45998 53283 46010 53339
rect 46066 53283 46078 53339
rect 45998 53271 46078 53283
rect 54146 53339 54226 53351
rect 54146 53283 54158 53339
rect 54214 53283 54226 53339
rect 54146 53271 54226 53283
rect 54760 53338 54840 53350
rect 54760 53282 54772 53338
rect 54828 53282 54840 53338
rect 54760 53270 54840 53282
rect -11327 52889 50119 52901
rect -11327 52887 19352 52889
rect -11327 52835 -11313 52887
rect -11261 52835 -2551 52887
rect -2499 52835 6211 52887
rect 6263 52835 14973 52887
rect 15025 52835 19352 52887
rect -11327 52833 19352 52835
rect 19408 52887 50119 52889
rect 19408 52835 23735 52887
rect 23787 52835 32497 52887
rect 32549 52835 41259 52887
rect 41311 52835 50021 52887
rect 50073 52835 50119 52887
rect 19408 52833 50119 52835
rect -11327 52821 50119 52833
rect -11941 52646 -7382 52660
rect -11941 52594 -11927 52646
rect -11875 52594 -7448 52646
rect -7396 52594 -7382 52646
rect -11941 52580 -7382 52594
rect -3179 52646 1380 52660
rect -3179 52594 -3165 52646
rect -3113 52594 1314 52646
rect 1366 52594 1380 52646
rect -3179 52580 1380 52594
rect 5583 52646 10142 52660
rect 5583 52594 5597 52646
rect 5649 52594 10076 52646
rect 10128 52594 10142 52646
rect 5583 52580 10142 52594
rect 14345 52646 18904 52660
rect 14345 52594 14359 52646
rect 14411 52594 18838 52646
rect 18890 52594 18904 52646
rect 14345 52580 18904 52594
rect 23107 52646 27666 52660
rect 23107 52594 23121 52646
rect 23173 52594 27600 52646
rect 27652 52594 27666 52646
rect 23107 52580 27666 52594
rect 31869 52646 36428 52660
rect 31869 52594 31883 52646
rect 31935 52594 36362 52646
rect 36414 52594 36428 52646
rect 31869 52580 36428 52594
rect 40631 52646 45190 52660
rect 40631 52594 40645 52646
rect 40697 52594 45124 52646
rect 45176 52594 45190 52646
rect 40631 52580 45190 52594
rect 49393 52646 53952 52660
rect 49393 52594 49407 52646
rect 49459 52594 53886 52646
rect 53938 52594 53952 52646
rect 49393 52580 53952 52594
rect -10360 52342 -10280 52354
rect -10360 52286 -10348 52342
rect -10292 52286 -10280 52342
rect -10360 52274 -10280 52286
rect -1598 52342 -1518 52354
rect -1598 52286 -1586 52342
rect -1530 52286 -1518 52342
rect -1598 52274 -1518 52286
rect 7164 52342 7244 52354
rect 7164 52286 7176 52342
rect 7232 52286 7244 52342
rect 7164 52274 7244 52286
rect 15926 52342 16006 52354
rect 15926 52286 15938 52342
rect 15994 52286 16006 52342
rect 15926 52274 16006 52286
rect 24688 52342 24768 52354
rect 24688 52286 24700 52342
rect 24756 52286 24768 52342
rect 24688 52274 24768 52286
rect 33450 52342 33530 52354
rect 33450 52286 33462 52342
rect 33518 52286 33530 52342
rect 33450 52274 33530 52286
rect 42212 52342 42292 52354
rect 42212 52286 42224 52342
rect 42280 52286 42292 52342
rect 42212 52274 42292 52286
rect 50974 52342 51054 52354
rect 50974 52286 50986 52342
rect 51042 52286 51054 52342
rect 50974 52274 51054 52286
rect -12954 51756 -12874 51768
rect -12954 51700 -12942 51756
rect -12886 51700 -12874 51756
rect -12954 51688 -12874 51700
rect 57502 51756 57582 51768
rect 57502 51700 57514 51756
rect 57570 51700 57582 51756
rect 57502 51688 57582 51700
rect -10360 51507 -10280 51519
rect -10360 51451 -10348 51507
rect -10292 51451 -10280 51507
rect -10360 51439 -10280 51451
rect -1598 51507 -1518 51519
rect -1598 51451 -1586 51507
rect -1530 51451 -1518 51507
rect -1598 51439 -1518 51451
rect 7164 51507 7244 51519
rect 7164 51451 7176 51507
rect 7232 51451 7244 51507
rect 7164 51439 7244 51451
rect 15926 51507 16006 51519
rect 15926 51451 15938 51507
rect 15994 51451 16006 51507
rect 15926 51439 16006 51451
rect 24688 51507 24768 51519
rect 24688 51451 24700 51507
rect 24756 51451 24768 51507
rect 24688 51439 24768 51451
rect 33450 51507 33530 51519
rect 33450 51451 33462 51507
rect 33518 51451 33530 51507
rect 33450 51439 33530 51451
rect 42212 51507 42292 51519
rect 42212 51451 42224 51507
rect 42280 51451 42292 51507
rect 42212 51439 42292 51451
rect 50974 51507 51054 51519
rect 50974 51451 50986 51507
rect 51042 51451 51054 51507
rect 50974 51439 51054 51451
rect -12332 50971 49082 50985
rect -12332 50919 -12318 50971
rect -12266 50919 -3556 50971
rect -3504 50919 5206 50971
rect 5258 50919 13968 50971
rect 14020 50919 22730 50971
rect 22782 50919 31492 50971
rect 31544 50919 40254 50971
rect 40306 50919 49016 50971
rect 49068 50919 49082 50971
rect -12332 50905 49082 50919
rect 49002 50173 49082 50185
rect 49002 50117 49014 50173
rect 49070 50117 49082 50173
rect 49002 50105 49082 50117
rect -11268 50052 49997 50064
rect -11268 49996 -11256 50052
rect -11200 49996 -2494 50052
rect -2438 49996 6268 50052
rect 6324 49996 15030 50052
rect 15086 49996 23792 50052
rect 23848 49996 32554 50052
rect 32610 49996 41316 50052
rect 41372 49996 49929 50052
rect 49985 49996 49997 50052
rect -11268 49984 49997 49996
rect -12812 49934 -12732 49946
rect -12812 49878 -12800 49934
rect -12744 49878 -12732 49934
rect -12812 49866 -12732 49878
rect 57642 49932 57722 49946
rect 57642 49880 57656 49932
rect 57708 49880 57722 49932
rect 57642 49866 57722 49880
rect 51718 49695 51798 49707
rect 51718 49639 51730 49695
rect 51786 49639 51798 49695
rect 51718 49627 51798 49639
rect 57502 48152 57582 48164
rect 57502 48096 57514 48152
rect 57570 48096 57582 48152
rect 57502 48084 57582 48096
rect -12812 47014 -12732 47026
rect -12812 46958 -12800 47014
rect -12744 46958 -12732 47014
rect -12812 46946 -12732 46958
rect 50227 47014 50307 47026
rect 50227 46958 50239 47014
rect 50295 46958 50307 47014
rect 50227 46946 50307 46958
rect 55659 47014 55739 47026
rect 55659 46958 55671 47014
rect 55727 46958 55739 47014
rect 55659 46946 55739 46958
rect 57642 47014 57722 47026
rect 57642 46958 57654 47014
rect 57710 46958 57722 47014
rect 57642 46946 57722 46958
rect 8847 46204 8927 46216
rect 8847 46148 8859 46204
rect 8915 46148 8927 46204
rect 8847 46136 8927 46148
rect 12791 46204 12871 46216
rect 12791 46148 12803 46204
rect 12859 46148 12871 46204
rect 12791 46136 12871 46148
rect 16735 46204 16815 46216
rect 16735 46148 16747 46204
rect 16803 46148 16815 46204
rect 16735 46136 16815 46148
rect 20679 46204 20759 46216
rect 20679 46148 20691 46204
rect 20747 46148 20759 46204
rect 20679 46136 20759 46148
rect 24623 46204 24703 46216
rect 24623 46148 24635 46204
rect 24691 46148 24703 46204
rect 24623 46136 24703 46148
rect 28567 46204 28647 46216
rect 28567 46148 28579 46204
rect 28635 46148 28647 46204
rect 28567 46136 28647 46148
rect 32511 46204 32591 46216
rect 32511 46148 32523 46204
rect 32579 46148 32591 46204
rect 32511 46136 32591 46148
rect 36455 46204 36535 46216
rect 36455 46148 36467 46204
rect 36523 46148 36535 46204
rect 36455 46136 36535 46148
rect -12954 45232 -12874 45244
rect -12954 45176 -12942 45232
rect -12886 45176 -12874 45232
rect -12954 45164 -12874 45176
rect 57502 45232 57582 45244
rect 57502 45176 57514 45232
rect 57570 45176 57582 45232
rect 57502 45164 57582 45176
rect 50227 42092 50307 42104
rect 50227 42036 50239 42092
rect 50295 42036 50307 42092
rect 50227 42024 50307 42036
rect 55659 42092 55739 42104
rect 55659 42036 55671 42092
rect 55727 42036 55739 42092
rect 55659 42024 55739 42036
rect 49002 29812 50027 29824
rect 49002 29756 49014 29812
rect 49070 29756 50027 29812
rect 49002 29744 50027 29756
<< via2 >>
rect -12942 62910 -12886 62966
rect 51953 61682 52009 61738
rect 57654 61682 57710 61738
rect -12800 61533 -12744 61589
rect -7282 61533 -7226 61589
rect 50625 55861 50681 55863
rect 50625 55809 50627 55861
rect 50627 55809 50679 55861
rect 50679 55809 50681 55861
rect 50625 55807 50681 55809
rect -12800 53576 -12744 53578
rect -12800 53524 -12798 53576
rect -12798 53524 -12746 53576
rect -12746 53524 -12744 53576
rect -12800 53522 -12744 53524
rect -7176 53337 -7120 53339
rect -7176 53285 -7174 53337
rect -7174 53285 -7122 53337
rect -7122 53285 -7120 53337
rect -7176 53283 -7120 53285
rect -6562 53337 -6506 53339
rect -6562 53285 -6560 53337
rect -6560 53285 -6508 53337
rect -6508 53285 -6506 53337
rect -6562 53283 -6506 53285
rect 1586 53337 1642 53339
rect 1586 53285 1588 53337
rect 1588 53285 1640 53337
rect 1640 53285 1642 53337
rect 1586 53283 1642 53285
rect 2200 53337 2256 53339
rect 2200 53285 2202 53337
rect 2202 53285 2254 53337
rect 2254 53285 2256 53337
rect 2200 53283 2256 53285
rect 10348 53337 10404 53339
rect 10348 53285 10350 53337
rect 10350 53285 10402 53337
rect 10402 53285 10404 53337
rect 10348 53283 10404 53285
rect 10962 53337 11018 53339
rect 10962 53285 10964 53337
rect 10964 53285 11016 53337
rect 11016 53285 11018 53337
rect 10962 53283 11018 53285
rect 19110 53337 19166 53339
rect 19110 53285 19112 53337
rect 19112 53285 19164 53337
rect 19164 53285 19166 53337
rect 19110 53283 19166 53285
rect 19724 53337 19780 53339
rect 19724 53285 19726 53337
rect 19726 53285 19778 53337
rect 19778 53285 19780 53337
rect 19724 53283 19780 53285
rect 27872 53337 27928 53339
rect 27872 53285 27874 53337
rect 27874 53285 27926 53337
rect 27926 53285 27928 53337
rect 27872 53283 27928 53285
rect 28486 53337 28542 53339
rect 28486 53285 28488 53337
rect 28488 53285 28540 53337
rect 28540 53285 28542 53337
rect 28486 53283 28542 53285
rect 36634 53337 36690 53339
rect 36634 53285 36636 53337
rect 36636 53285 36688 53337
rect 36688 53285 36690 53337
rect 36634 53283 36690 53285
rect 37248 53337 37304 53339
rect 37248 53285 37250 53337
rect 37250 53285 37302 53337
rect 37302 53285 37304 53337
rect 37248 53283 37304 53285
rect 45396 53337 45452 53339
rect 45396 53285 45398 53337
rect 45398 53285 45450 53337
rect 45450 53285 45452 53337
rect 45396 53283 45452 53285
rect 46010 53337 46066 53339
rect 46010 53285 46012 53337
rect 46012 53285 46064 53337
rect 46064 53285 46066 53337
rect 46010 53283 46066 53285
rect 54158 53337 54214 53339
rect 54158 53285 54160 53337
rect 54160 53285 54212 53337
rect 54212 53285 54214 53337
rect 54158 53283 54214 53285
rect 54772 53336 54828 53338
rect 54772 53284 54774 53336
rect 54774 53284 54826 53336
rect 54826 53284 54828 53336
rect 54772 53282 54828 53284
rect 19352 52833 19408 52889
rect -10348 52340 -10292 52342
rect -10348 52288 -10346 52340
rect -10346 52288 -10294 52340
rect -10294 52288 -10292 52340
rect -10348 52286 -10292 52288
rect -1586 52340 -1530 52342
rect -1586 52288 -1584 52340
rect -1584 52288 -1532 52340
rect -1532 52288 -1530 52340
rect -1586 52286 -1530 52288
rect 7176 52340 7232 52342
rect 7176 52288 7178 52340
rect 7178 52288 7230 52340
rect 7230 52288 7232 52340
rect 7176 52286 7232 52288
rect 15938 52340 15994 52342
rect 15938 52288 15940 52340
rect 15940 52288 15992 52340
rect 15992 52288 15994 52340
rect 15938 52286 15994 52288
rect 24700 52340 24756 52342
rect 24700 52288 24702 52340
rect 24702 52288 24754 52340
rect 24754 52288 24756 52340
rect 24700 52286 24756 52288
rect 33462 52340 33518 52342
rect 33462 52288 33464 52340
rect 33464 52288 33516 52340
rect 33516 52288 33518 52340
rect 33462 52286 33518 52288
rect 42224 52340 42280 52342
rect 42224 52288 42226 52340
rect 42226 52288 42278 52340
rect 42278 52288 42280 52340
rect 42224 52286 42280 52288
rect 50986 52340 51042 52342
rect 50986 52288 50988 52340
rect 50988 52288 51040 52340
rect 51040 52288 51042 52340
rect 50986 52286 51042 52288
rect -12942 51754 -12886 51756
rect -12942 51702 -12940 51754
rect -12940 51702 -12888 51754
rect -12888 51702 -12886 51754
rect -12942 51700 -12886 51702
rect 57514 51754 57570 51756
rect 57514 51702 57516 51754
rect 57516 51702 57568 51754
rect 57568 51702 57570 51754
rect 57514 51700 57570 51702
rect -10348 51505 -10292 51507
rect -10348 51453 -10346 51505
rect -10346 51453 -10294 51505
rect -10294 51453 -10292 51505
rect -10348 51451 -10292 51453
rect -1586 51505 -1530 51507
rect -1586 51453 -1584 51505
rect -1584 51453 -1532 51505
rect -1532 51453 -1530 51505
rect -1586 51451 -1530 51453
rect 7176 51505 7232 51507
rect 7176 51453 7178 51505
rect 7178 51453 7230 51505
rect 7230 51453 7232 51505
rect 7176 51451 7232 51453
rect 15938 51505 15994 51507
rect 15938 51453 15940 51505
rect 15940 51453 15992 51505
rect 15992 51453 15994 51505
rect 15938 51451 15994 51453
rect 24700 51505 24756 51507
rect 24700 51453 24702 51505
rect 24702 51453 24754 51505
rect 24754 51453 24756 51505
rect 24700 51451 24756 51453
rect 33462 51505 33518 51507
rect 33462 51453 33464 51505
rect 33464 51453 33516 51505
rect 33516 51453 33518 51505
rect 33462 51451 33518 51453
rect 42224 51505 42280 51507
rect 42224 51453 42226 51505
rect 42226 51453 42278 51505
rect 42278 51453 42280 51505
rect 42224 51451 42280 51453
rect 50986 51505 51042 51507
rect 50986 51453 50988 51505
rect 50988 51453 51040 51505
rect 51040 51453 51042 51505
rect 50986 51451 51042 51453
rect 49014 50171 49070 50173
rect 49014 50119 49016 50171
rect 49016 50119 49068 50171
rect 49068 50119 49070 50171
rect 49014 50117 49070 50119
rect -11256 49996 -11200 50052
rect -2494 49996 -2438 50052
rect 6268 49996 6324 50052
rect 15030 49996 15086 50052
rect 23792 49996 23848 50052
rect 32554 49996 32610 50052
rect 41316 49996 41372 50052
rect 49929 49996 49985 50052
rect -12800 49932 -12744 49934
rect -12800 49880 -12798 49932
rect -12798 49880 -12746 49932
rect -12746 49880 -12744 49932
rect -12800 49878 -12744 49880
rect 51730 49693 51786 49695
rect 51730 49641 51732 49693
rect 51732 49641 51784 49693
rect 51784 49641 51786 49693
rect 51730 49639 51786 49641
rect 57514 48150 57570 48152
rect 57514 48098 57516 48150
rect 57516 48098 57568 48150
rect 57568 48098 57570 48150
rect 57514 48096 57570 48098
rect -12800 47012 -12744 47014
rect -12800 46960 -12798 47012
rect -12798 46960 -12746 47012
rect -12746 46960 -12744 47012
rect -12800 46958 -12744 46960
rect 50239 47012 50295 47014
rect 50239 46960 50241 47012
rect 50241 46960 50293 47012
rect 50293 46960 50295 47012
rect 50239 46958 50295 46960
rect 55671 47012 55727 47014
rect 55671 46960 55673 47012
rect 55673 46960 55725 47012
rect 55725 46960 55727 47012
rect 55671 46958 55727 46960
rect 57654 47012 57710 47014
rect 57654 46960 57656 47012
rect 57656 46960 57708 47012
rect 57708 46960 57710 47012
rect 57654 46958 57710 46960
rect 8859 46202 8915 46204
rect 8859 46150 8861 46202
rect 8861 46150 8913 46202
rect 8913 46150 8915 46202
rect 8859 46148 8915 46150
rect 12803 46202 12859 46204
rect 12803 46150 12805 46202
rect 12805 46150 12857 46202
rect 12857 46150 12859 46202
rect 12803 46148 12859 46150
rect 16747 46202 16803 46204
rect 16747 46150 16749 46202
rect 16749 46150 16801 46202
rect 16801 46150 16803 46202
rect 16747 46148 16803 46150
rect 20691 46202 20747 46204
rect 20691 46150 20693 46202
rect 20693 46150 20745 46202
rect 20745 46150 20747 46202
rect 20691 46148 20747 46150
rect 24635 46202 24691 46204
rect 24635 46150 24637 46202
rect 24637 46150 24689 46202
rect 24689 46150 24691 46202
rect 24635 46148 24691 46150
rect 28579 46202 28635 46204
rect 28579 46150 28581 46202
rect 28581 46150 28633 46202
rect 28633 46150 28635 46202
rect 28579 46148 28635 46150
rect 32523 46202 32579 46204
rect 32523 46150 32525 46202
rect 32525 46150 32577 46202
rect 32577 46150 32579 46202
rect 32523 46148 32579 46150
rect 36467 46202 36523 46204
rect 36467 46150 36469 46202
rect 36469 46150 36521 46202
rect 36521 46150 36523 46202
rect 36467 46148 36523 46150
rect -12942 45230 -12886 45232
rect -12942 45178 -12940 45230
rect -12940 45178 -12888 45230
rect -12888 45178 -12886 45230
rect -12942 45176 -12886 45178
rect 57514 45230 57570 45232
rect 57514 45178 57516 45230
rect 57516 45178 57568 45230
rect 57568 45178 57570 45230
rect 57514 45176 57570 45178
rect 50239 42090 50295 42092
rect 50239 42038 50241 42090
rect 50241 42038 50293 42090
rect 50293 42038 50295 42090
rect 50239 42036 50295 42038
rect 55671 42090 55727 42092
rect 55671 42038 55673 42090
rect 55673 42038 55725 42090
rect 55725 42038 55727 42090
rect 55671 42036 55727 42038
rect 49014 29756 49070 29812
<< metal3 >>
rect -12947 62966 -12881 62971
rect -12947 62910 -12942 62966
rect -12886 62910 -12881 62966
rect -12947 62905 -12881 62910
rect -6944 62908 -1886 62968
rect 52642 62908 57572 62968
rect -12944 51761 -12884 62905
rect 51948 61740 52014 61743
rect -6421 61680 47040 61740
rect 47100 61680 48171 61740
rect 51669 61738 52014 61740
rect 51669 61682 51953 61738
rect 52009 61682 52014 61738
rect 51669 61680 52014 61682
rect 51948 61677 52014 61680
rect -12805 61589 -12739 61594
rect -12805 61533 -12800 61589
rect -12744 61533 -12739 61589
rect -12805 61528 -12739 61533
rect -7287 61591 -7221 61594
rect -7287 61589 -6974 61591
rect -7287 61533 -7282 61589
rect -7226 61533 -6974 61589
rect -7287 61531 -6974 61533
rect -7287 61528 -7221 61531
rect -12802 53583 -12742 61528
rect -6421 60623 47040 60683
rect 47100 60623 51181 60683
rect -4548 54459 -2183 54519
rect -984 54459 1381 54519
rect 2580 54459 4945 54519
rect 6144 54459 8509 54519
rect 9708 54459 12073 54519
rect 13272 54459 15637 54519
rect 16836 54459 19201 54519
rect -3396 53837 -3336 54459
rect -6572 53831 -6496 53837
rect -6572 53767 -6566 53831
rect -6502 53767 -6496 53831
rect -6572 53761 -6496 53767
rect -3404 53831 -3328 53837
rect -3404 53767 -3398 53831
rect -3334 53767 -3328 53831
rect -3404 53761 -3328 53767
rect -2653 53831 -2577 53837
rect -2653 53767 -2647 53831
rect -2583 53767 -2577 53831
rect -2653 53761 -2577 53767
rect -11415 53703 -11339 53709
rect -11415 53639 -11409 53703
rect -11345 53639 -11339 53703
rect -11415 53633 -11339 53639
rect -7186 53703 -7110 53709
rect -7186 53639 -7180 53703
rect -7116 53639 -7110 53703
rect -7186 53633 -7110 53639
rect -12805 53578 -12739 53583
rect -12805 53522 -12800 53578
rect -12744 53522 -12739 53578
rect -12805 53517 -12739 53522
rect -12947 51756 -12881 51761
rect -12947 51700 -12942 51756
rect -12886 51700 -12881 51756
rect -12947 51695 -12881 51700
rect -12944 45237 -12884 51695
rect -12802 49939 -12742 53517
rect -11407 50688 -11347 53633
rect -7178 53344 -7118 53633
rect -6564 53344 -6504 53761
rect -7181 53339 -7115 53344
rect -7181 53283 -7176 53339
rect -7120 53283 -7115 53339
rect -7181 53278 -7115 53283
rect -6567 53339 -6501 53344
rect -6567 53283 -6562 53339
rect -6506 53283 -6501 53339
rect -6567 53278 -6501 53283
rect -10353 52342 -10287 52347
rect -10353 52286 -10348 52342
rect -10292 52286 -10287 52342
rect -10353 52281 -10287 52286
rect -10350 51512 -10290 52281
rect -10353 51507 -10287 51512
rect -10353 51451 -10348 51507
rect -10292 51451 -10287 51507
rect -10353 51446 -10287 51451
rect -2645 50687 -2585 53761
rect 168 53709 228 54459
rect 1584 53837 1644 53846
rect 1576 53831 1652 53837
rect 1576 53767 1582 53831
rect 1646 53767 1652 53831
rect 1576 53761 1652 53767
rect 160 53703 236 53709
rect 160 53639 166 53703
rect 230 53639 236 53703
rect 160 53633 236 53639
rect 1584 53344 1644 53761
rect 3732 53709 3792 54459
rect 7296 53837 7356 54459
rect 7288 53831 7364 53837
rect 7288 53767 7294 53831
rect 7358 53767 7364 53831
rect 7288 53761 7364 53767
rect 2190 53703 2266 53709
rect 2190 53639 2196 53703
rect 2260 53639 2266 53703
rect 2190 53633 2266 53639
rect 3724 53703 3800 53709
rect 3724 53639 3730 53703
rect 3794 53639 3800 53703
rect 3724 53633 3800 53639
rect 6109 53703 6185 53709
rect 6109 53639 6115 53703
rect 6179 53639 6185 53703
rect 6109 53633 6185 53639
rect 10338 53703 10414 53709
rect 10338 53639 10344 53703
rect 10408 53639 10414 53703
rect 10338 53633 10414 53639
rect 2198 53344 2258 53633
rect 1581 53339 1647 53344
rect 1581 53283 1586 53339
rect 1642 53283 1647 53339
rect 1581 53278 1647 53283
rect 2195 53339 2261 53344
rect 2195 53283 2200 53339
rect 2256 53283 2261 53339
rect 2195 53278 2261 53283
rect -1591 52342 -1525 52347
rect -1591 52286 -1586 52342
rect -1530 52286 -1525 52342
rect -1591 52281 -1525 52286
rect -1588 51512 -1528 52281
rect -1591 51507 -1525 51512
rect -1591 51451 -1586 51507
rect -1530 51451 -1525 51507
rect -1591 51446 -1525 51451
rect 6117 50688 6177 53633
rect 10346 53344 10406 53633
rect 10960 53344 11020 54459
rect 14424 53709 14484 54459
rect 17988 53837 18048 54459
rect 17980 53831 18056 53837
rect 17980 53767 17986 53831
rect 18050 53767 18056 53831
rect 17980 53761 18056 53767
rect 14416 53703 14492 53709
rect 14416 53639 14422 53703
rect 14486 53639 14492 53703
rect 14416 53633 14492 53639
rect 14871 53703 14947 53709
rect 14871 53639 14877 53703
rect 14941 53639 14947 53703
rect 14871 53633 14947 53639
rect 19100 53703 19176 53709
rect 19100 53639 19106 53703
rect 19170 53639 19176 53703
rect 19100 53633 19176 53639
rect 10343 53339 10409 53344
rect 10343 53283 10348 53339
rect 10404 53283 10409 53339
rect 10343 53278 10409 53283
rect 10957 53339 11023 53344
rect 10957 53283 10962 53339
rect 11018 53283 11023 53339
rect 10957 53278 11023 53283
rect 7171 52342 7237 52347
rect 7171 52286 7176 52342
rect 7232 52286 7237 52342
rect 7171 52281 7237 52286
rect 7174 51512 7234 52281
rect 7171 51507 7237 51512
rect 7171 51451 7176 51507
rect 7232 51451 7237 51507
rect 7171 51446 7237 51451
rect 14879 50688 14939 53633
rect 19108 53344 19168 53633
rect 19105 53339 19171 53344
rect 19105 53283 19110 53339
rect 19166 53283 19171 53339
rect 19105 53278 19171 53283
rect 19350 52894 19410 60623
rect 50620 55865 50686 55868
rect 50620 55863 51788 55865
rect 50620 55807 50625 55863
rect 50681 55807 51788 55863
rect 50620 55805 51788 55807
rect 50620 55802 50686 55805
rect 20400 54459 22765 54519
rect 23964 54459 26329 54519
rect 27528 54459 29893 54519
rect 31092 54459 33457 54519
rect 34656 54459 37021 54519
rect 38220 54459 40585 54519
rect 41784 54459 44149 54519
rect 45348 54459 47713 54519
rect 48912 54459 51277 54519
rect 19714 53831 19790 53837
rect 19714 53767 19720 53831
rect 19784 53767 19790 53831
rect 19714 53761 19790 53767
rect 19722 53344 19782 53761
rect 21552 53709 21612 54459
rect 25116 53837 25176 54459
rect 25108 53831 25184 53837
rect 25108 53767 25114 53831
rect 25178 53767 25184 53831
rect 25108 53761 25184 53767
rect 28476 53831 28552 53837
rect 28476 53767 28482 53831
rect 28546 53767 28552 53831
rect 28476 53761 28552 53767
rect 27870 53709 27930 53720
rect 21544 53703 21620 53709
rect 21544 53639 21550 53703
rect 21614 53639 21620 53703
rect 21544 53633 21620 53639
rect 23633 53703 23709 53709
rect 23633 53639 23639 53703
rect 23703 53639 23709 53703
rect 23633 53633 23709 53639
rect 27862 53703 27938 53709
rect 27862 53639 27868 53703
rect 27932 53639 27938 53703
rect 27862 53633 27938 53639
rect 19719 53339 19785 53344
rect 19719 53283 19724 53339
rect 19780 53283 19785 53339
rect 19719 53278 19785 53283
rect 19347 52889 19413 52894
rect 19347 52833 19352 52889
rect 19408 52833 19413 52889
rect 19347 52828 19413 52833
rect 15933 52342 15999 52347
rect 15933 52286 15938 52342
rect 15994 52286 15999 52342
rect 15933 52281 15999 52286
rect 15936 51512 15996 52281
rect 15933 51507 15999 51512
rect 15933 51451 15938 51507
rect 15994 51451 15999 51507
rect 15933 51446 15999 51451
rect 23641 50688 23701 53633
rect 27870 53344 27930 53633
rect 28484 53344 28544 53761
rect 28680 53709 28740 54459
rect 32244 53837 32304 54459
rect 32236 53831 32312 53837
rect 32236 53767 32242 53831
rect 32306 53767 32312 53831
rect 32236 53761 32312 53767
rect 35808 53709 35868 54459
rect 39372 53837 39432 54459
rect 37238 53831 37314 53837
rect 37238 53767 37244 53831
rect 37308 53767 37314 53831
rect 37238 53761 37314 53767
rect 39364 53831 39440 53837
rect 39364 53767 39370 53831
rect 39434 53767 39440 53831
rect 39364 53761 39440 53767
rect 28672 53703 28748 53709
rect 28672 53639 28678 53703
rect 28742 53639 28748 53703
rect 28672 53633 28748 53639
rect 32395 53703 32471 53709
rect 32395 53639 32401 53703
rect 32465 53639 32471 53703
rect 32395 53633 32471 53639
rect 35800 53703 35876 53709
rect 35800 53639 35806 53703
rect 35870 53639 35876 53703
rect 35800 53633 35876 53639
rect 36624 53703 36700 53709
rect 36624 53639 36630 53703
rect 36694 53639 36700 53703
rect 36624 53633 36700 53639
rect 27867 53339 27933 53344
rect 27867 53283 27872 53339
rect 27928 53283 27933 53339
rect 27867 53278 27933 53283
rect 28481 53339 28547 53344
rect 28481 53283 28486 53339
rect 28542 53283 28547 53339
rect 28481 53278 28547 53283
rect 24695 52342 24761 52347
rect 24695 52286 24700 52342
rect 24756 52286 24761 52342
rect 24695 52281 24761 52286
rect 24698 51512 24758 52281
rect 24695 51507 24761 51512
rect 24695 51451 24700 51507
rect 24756 51451 24761 51507
rect 24695 51446 24761 51451
rect 32403 50688 32463 53633
rect 36632 53344 36692 53633
rect 37246 53344 37306 53761
rect 42936 53709 42996 54459
rect 46500 53837 46560 54459
rect 46000 53831 46076 53837
rect 46000 53767 46006 53831
rect 46070 53767 46076 53831
rect 46000 53761 46076 53767
rect 46492 53831 46568 53837
rect 46492 53767 46498 53831
rect 46562 53767 46568 53831
rect 46492 53761 46568 53767
rect 41157 53703 41233 53709
rect 41157 53639 41163 53703
rect 41227 53639 41233 53703
rect 41157 53633 41233 53639
rect 42928 53703 43004 53709
rect 42928 53639 42934 53703
rect 42998 53639 43004 53703
rect 42928 53633 43004 53639
rect 45386 53703 45462 53709
rect 45386 53639 45392 53703
rect 45456 53639 45462 53703
rect 45386 53633 45462 53639
rect 36629 53339 36695 53344
rect 36629 53283 36634 53339
rect 36690 53283 36695 53339
rect 36629 53278 36695 53283
rect 37243 53339 37309 53344
rect 37243 53283 37248 53339
rect 37304 53283 37309 53339
rect 37243 53278 37309 53283
rect 33457 52342 33523 52347
rect 33457 52286 33462 52342
rect 33518 52286 33523 52342
rect 33457 52281 33523 52286
rect 33460 51512 33520 52281
rect 33457 51507 33523 51512
rect 33457 51451 33462 51507
rect 33518 51451 33523 51507
rect 33457 51446 33523 51451
rect 41165 50688 41225 53633
rect 45394 53344 45454 53633
rect 46008 53344 46068 53761
rect 50064 53709 50124 54459
rect 49919 53703 49995 53709
rect 49919 53639 49925 53703
rect 49989 53639 49995 53703
rect 49919 53633 49995 53639
rect 50056 53703 50132 53709
rect 50056 53639 50062 53703
rect 50126 53639 50132 53703
rect 50056 53633 50132 53639
rect 45391 53339 45457 53344
rect 45391 53283 45396 53339
rect 45452 53283 45457 53339
rect 45391 53278 45457 53283
rect 46005 53339 46071 53344
rect 46005 53283 46010 53339
rect 46066 53283 46071 53339
rect 46005 53278 46071 53283
rect 42219 52342 42285 52347
rect 42219 52286 42224 52342
rect 42280 52286 42285 52342
rect 42219 52281 42285 52286
rect 42222 51512 42282 52281
rect 42219 51507 42285 51512
rect 42219 51451 42224 51507
rect 42280 51451 42285 51507
rect 42219 51446 42285 51451
rect 49927 50688 49987 53633
rect 50981 52342 51047 52347
rect 50981 52286 50986 52342
rect 51042 52286 51047 52342
rect 50981 52281 51047 52286
rect 50984 51512 51044 52281
rect 50981 51507 51047 51512
rect 50981 51451 50986 51507
rect 51042 51451 51047 51507
rect 50981 51446 51047 51451
rect 49009 50173 49075 50178
rect 49009 50117 49014 50173
rect 49070 50117 49075 50173
rect -11261 50052 -11195 50112
rect -11261 49996 -11256 50052
rect -11200 49996 -11195 50052
rect -11261 49991 -11195 49996
rect -2499 50052 -2433 50117
rect -2499 49996 -2494 50052
rect -2438 49996 -2433 50052
rect -2499 49991 -2433 49996
rect 6263 50052 6329 50117
rect 6263 49996 6268 50052
rect 6324 49996 6329 50052
rect 6263 49991 6329 49996
rect 15025 50052 15091 50117
rect 15025 49996 15030 50052
rect 15086 49996 15091 50052
rect 15025 49991 15091 49996
rect 23787 50052 23853 50117
rect 23787 49996 23792 50052
rect 23848 49996 23853 50052
rect 23787 49991 23853 49996
rect 32549 50052 32615 50117
rect 32549 49996 32554 50052
rect 32610 49996 32615 50052
rect 32549 49991 32615 49996
rect 41311 50052 41377 50117
rect 49009 50112 49075 50117
rect 41311 49996 41316 50052
rect 41372 49996 41377 50052
rect 41311 49991 41377 49996
rect 6266 49987 6326 49991
rect 15028 49987 15088 49991
rect 23790 49987 23850 49991
rect 32552 49987 32612 49991
rect 41314 49987 41374 49991
rect -12805 49934 -12739 49939
rect -12805 49878 -12800 49934
rect -12744 49878 -12739 49934
rect -12805 49873 -12739 49878
rect -12802 47019 -12742 49873
rect -4186 47145 -4126 49684
rect 4576 47273 4636 49684
rect 13338 47401 13398 49685
rect 22100 47529 22160 49684
rect 28569 47779 28645 47785
rect 28569 47715 28575 47779
rect 28639 47715 28645 47779
rect 28569 47709 28645 47715
rect 24625 47651 24701 47657
rect 24625 47587 24631 47651
rect 24695 47587 24701 47651
rect 24625 47581 24701 47587
rect 20681 47523 20757 47529
rect 20681 47459 20687 47523
rect 20751 47459 20757 47523
rect 20681 47453 20757 47459
rect 22092 47523 22168 47529
rect 22092 47459 22098 47523
rect 22162 47459 22168 47523
rect 22092 47453 22168 47459
rect 13330 47395 13406 47401
rect 13330 47331 13336 47395
rect 13400 47331 13406 47395
rect 13330 47325 13406 47331
rect 16737 47395 16813 47401
rect 16737 47331 16743 47395
rect 16807 47331 16813 47395
rect 16737 47325 16813 47331
rect 4568 47267 4644 47273
rect 4568 47203 4574 47267
rect 4638 47203 4644 47267
rect 4568 47197 4644 47203
rect 12793 47267 12869 47273
rect 12793 47203 12799 47267
rect 12863 47203 12869 47267
rect 12793 47197 12869 47203
rect -4194 47139 -4118 47145
rect -4194 47075 -4188 47139
rect -4124 47075 -4118 47139
rect -4194 47069 -4118 47075
rect 8849 47139 8925 47145
rect 8849 47075 8855 47139
rect 8919 47075 8925 47139
rect 8849 47069 8925 47075
rect -12805 47014 -12739 47019
rect -12805 46958 -12800 47014
rect -12744 46958 -12739 47014
rect -12805 46953 -12739 46958
rect 8857 46209 8917 47069
rect 12801 46209 12861 47197
rect 16745 46209 16805 47325
rect 20689 46209 20749 47453
rect 24633 46209 24693 47581
rect 28577 46209 28637 47709
rect 30862 47657 30922 49685
rect 36457 48035 36533 48041
rect 36457 47971 36463 48035
rect 36527 47971 36533 48035
rect 36457 47965 36533 47971
rect 32513 47907 32589 47913
rect 32513 47843 32519 47907
rect 32583 47843 32589 47907
rect 32513 47837 32589 47843
rect 30854 47651 30930 47657
rect 30854 47587 30860 47651
rect 30924 47587 30930 47651
rect 30854 47581 30930 47587
rect 32521 46209 32581 47837
rect 36465 46209 36525 47965
rect 39624 47785 39684 49683
rect 48386 47913 48446 49684
rect 48378 47907 48454 47913
rect 48378 47843 48384 47907
rect 48448 47843 48454 47907
rect 48378 47837 48454 47843
rect 39616 47779 39692 47785
rect 39616 47715 39622 47779
rect 39686 47715 39692 47779
rect 39616 47709 39692 47715
rect 8854 46204 8920 46209
rect 8854 46148 8859 46204
rect 8915 46148 8920 46204
rect 8854 46143 8920 46148
rect 12798 46204 12864 46209
rect 12798 46148 12803 46204
rect 12859 46148 12864 46204
rect 12798 46143 12864 46148
rect 16742 46204 16808 46209
rect 16742 46148 16747 46204
rect 16803 46148 16808 46204
rect 16742 46143 16808 46148
rect 20686 46204 20752 46209
rect 20686 46148 20691 46204
rect 20747 46148 20752 46204
rect 20686 46143 20752 46148
rect 24630 46204 24696 46209
rect 24630 46148 24635 46204
rect 24691 46148 24696 46204
rect 24630 46143 24696 46148
rect 28574 46204 28640 46209
rect 28574 46148 28579 46204
rect 28635 46148 28640 46204
rect 28574 46143 28640 46148
rect 32518 46204 32584 46209
rect 32518 46148 32523 46204
rect 32579 46148 32584 46204
rect 32518 46143 32584 46148
rect 36462 46204 36528 46209
rect 36462 46148 36467 46204
rect 36523 46148 36528 46204
rect 36462 46143 36528 46148
rect -12947 45232 -12881 45237
rect -12947 45176 -12942 45232
rect -12886 45176 -12881 45232
rect -12947 45171 -12881 45176
rect 49012 29817 49072 50112
rect 49924 50052 49990 50057
rect 49924 49996 49929 50052
rect 49985 49996 49990 50052
rect 49924 49991 49990 49996
rect 51728 49700 51788 55805
rect 54762 53831 54838 53837
rect 54762 53767 54768 53831
rect 54832 53767 54838 53831
rect 54762 53761 54838 53767
rect 54148 53703 54224 53709
rect 54148 53639 54154 53703
rect 54218 53639 54224 53703
rect 54148 53633 54224 53639
rect 54156 53344 54216 53633
rect 54153 53339 54219 53344
rect 54770 53343 54830 53761
rect 54153 53283 54158 53339
rect 54214 53283 54219 53339
rect 54153 53278 54219 53283
rect 54767 53338 54833 53343
rect 54767 53282 54772 53338
rect 54828 53282 54833 53338
rect 54767 53277 54833 53282
rect 57512 51761 57572 62908
rect 57649 61738 57715 61743
rect 57649 61682 57654 61738
rect 57710 61682 57715 61738
rect 57649 61677 57715 61682
rect 57652 53583 57712 61677
rect 57649 53517 57715 53583
rect 57509 51756 57575 51761
rect 57509 51700 57514 51756
rect 57570 51700 57575 51756
rect 57509 51695 57575 51700
rect 51725 49695 51791 49700
rect 51725 49639 51730 49695
rect 51786 49639 51791 49695
rect 51725 49634 51791 49639
rect 57148 48041 57208 49678
rect 57512 48157 57572 51695
rect 57652 49939 57712 53517
rect 57649 49873 57715 49939
rect 57509 48152 57575 48157
rect 57509 48096 57514 48152
rect 57570 48096 57575 48152
rect 57509 48091 57575 48096
rect 57140 48035 57216 48041
rect 57140 47971 57146 48035
rect 57210 47971 57216 48035
rect 57140 47965 57216 47971
rect 50234 47014 50300 47019
rect 50234 46958 50239 47014
rect 50295 46958 50300 47014
rect 50234 46953 50300 46958
rect 55666 47014 55732 47019
rect 55666 46958 55671 47014
rect 55727 46958 55732 47014
rect 55666 46953 55732 46958
rect 50237 42097 50297 46953
rect 55669 42097 55729 46953
rect 57512 45237 57572 48091
rect 57652 47019 57712 49873
rect 57649 47014 57715 47019
rect 57649 46958 57654 47014
rect 57710 46958 57715 47014
rect 57649 46953 57715 46958
rect 57509 45232 57575 45237
rect 57509 45176 57514 45232
rect 57570 45176 57575 45232
rect 57509 45171 57575 45176
rect 50234 42092 50300 42097
rect 50234 42036 50239 42092
rect 50295 42036 50300 42092
rect 50234 42031 50300 42036
rect 55666 42092 55732 42097
rect 55666 42036 55671 42092
rect 55727 42036 55732 42092
rect 55666 42031 55732 42036
rect 49009 29812 49075 29817
rect 49009 29756 49014 29812
rect 49070 29756 49075 29812
rect 49009 29751 49075 29756
rect 41580 26826 41656 26832
rect 41580 26762 41586 26826
rect 41650 26824 41656 26826
rect 48674 26826 48750 26832
rect 48674 26824 48680 26826
rect 41650 26764 48680 26824
rect 41650 26762 41656 26764
rect 41580 26756 41656 26762
rect 48674 26762 48680 26764
rect 48744 26762 48750 26826
rect 48674 26756 48750 26762
rect 52220 26826 52296 26832
rect 52220 26762 52226 26826
rect 52290 26762 52296 26826
rect 52220 26756 52296 26762
rect 52228 24771 52288 26756
<< via3 >>
rect -6566 53767 -6502 53831
rect -3398 53767 -3334 53831
rect -2647 53767 -2583 53831
rect -11409 53639 -11345 53703
rect -7180 53639 -7116 53703
rect 1582 53767 1646 53831
rect 166 53639 230 53703
rect 7294 53767 7358 53831
rect 2196 53639 2260 53703
rect 3730 53639 3794 53703
rect 6115 53639 6179 53703
rect 10344 53639 10408 53703
rect 17986 53767 18050 53831
rect 14422 53639 14486 53703
rect 14877 53639 14941 53703
rect 19106 53639 19170 53703
rect 19720 53767 19784 53831
rect 25114 53767 25178 53831
rect 28482 53767 28546 53831
rect 21550 53639 21614 53703
rect 23639 53639 23703 53703
rect 27868 53639 27932 53703
rect 32242 53767 32306 53831
rect 37244 53767 37308 53831
rect 39370 53767 39434 53831
rect 28678 53639 28742 53703
rect 32401 53639 32465 53703
rect 35806 53639 35870 53703
rect 36630 53639 36694 53703
rect 46006 53767 46070 53831
rect 46498 53767 46562 53831
rect 41163 53639 41227 53703
rect 42934 53639 42998 53703
rect 45392 53639 45456 53703
rect 49925 53639 49989 53703
rect 50062 53639 50126 53703
rect 28575 47715 28639 47779
rect 24631 47587 24695 47651
rect 20687 47459 20751 47523
rect 22098 47459 22162 47523
rect 13336 47331 13400 47395
rect 16743 47331 16807 47395
rect 4574 47203 4638 47267
rect 12799 47203 12863 47267
rect -4188 47075 -4124 47139
rect 8855 47075 8919 47139
rect 36463 47971 36527 48035
rect 32519 47843 32583 47907
rect 30860 47587 30924 47651
rect 48384 47843 48448 47907
rect 39622 47715 39686 47779
rect 54768 53767 54832 53831
rect 54154 53639 54218 53703
rect 57146 47971 57210 48035
rect 41586 26762 41650 26826
rect 48680 26762 48744 26826
rect 52226 26762 52290 26826
<< metal4 >>
rect -6567 53831 -6501 53832
rect -6567 53767 -6566 53831
rect -6502 53829 -6501 53831
rect -3399 53831 -3333 53832
rect -3399 53829 -3398 53831
rect -6502 53769 -3398 53829
rect -6502 53767 -6501 53769
rect -6567 53766 -6501 53767
rect -3399 53767 -3398 53769
rect -3334 53767 -3333 53831
rect -3399 53766 -3333 53767
rect -2648 53831 -2582 53832
rect -2648 53767 -2647 53831
rect -2583 53829 -2582 53831
rect 1581 53831 1647 53832
rect 1581 53829 1582 53831
rect -2583 53769 1582 53829
rect -2583 53767 -2582 53769
rect -2648 53766 -2582 53767
rect 1581 53767 1582 53769
rect 1646 53829 1647 53831
rect 7293 53831 7359 53832
rect 7293 53829 7294 53831
rect 1646 53769 7294 53829
rect 1646 53767 1647 53769
rect 1581 53766 1647 53767
rect 7293 53767 7294 53769
rect 7358 53767 7359 53831
rect 7293 53766 7359 53767
rect 17985 53831 18051 53832
rect 17985 53767 17986 53831
rect 18050 53829 18051 53831
rect 19719 53831 19785 53832
rect 19719 53829 19720 53831
rect 18050 53769 19720 53829
rect 18050 53767 18051 53769
rect 17985 53766 18051 53767
rect 19719 53767 19720 53769
rect 19784 53767 19785 53831
rect 19719 53766 19785 53767
rect 25113 53831 25179 53832
rect 25113 53767 25114 53831
rect 25178 53829 25179 53831
rect 28481 53831 28547 53832
rect 28481 53829 28482 53831
rect 25178 53769 28482 53829
rect 25178 53767 25179 53769
rect 25113 53766 25179 53767
rect 28481 53767 28482 53769
rect 28546 53767 28547 53831
rect 28481 53766 28547 53767
rect 32241 53831 32307 53832
rect 32241 53767 32242 53831
rect 32306 53829 32307 53831
rect 37243 53831 37309 53832
rect 37243 53829 37244 53831
rect 32306 53769 37244 53829
rect 32306 53767 32307 53769
rect 32241 53766 32307 53767
rect 37243 53767 37244 53769
rect 37308 53767 37309 53831
rect 37243 53766 37309 53767
rect 39369 53831 39435 53832
rect 39369 53767 39370 53831
rect 39434 53829 39435 53831
rect 46005 53831 46071 53832
rect 46005 53829 46006 53831
rect 39434 53769 46006 53829
rect 39434 53767 39435 53769
rect 39369 53766 39435 53767
rect 46005 53767 46006 53769
rect 46070 53767 46071 53831
rect 46005 53766 46071 53767
rect 46497 53831 46563 53832
rect 46497 53767 46498 53831
rect 46562 53829 46563 53831
rect 54767 53831 54833 53832
rect 54767 53829 54768 53831
rect 46562 53769 54768 53829
rect 46562 53767 46563 53769
rect 46497 53766 46563 53767
rect 54767 53767 54768 53769
rect 54832 53767 54833 53831
rect 54767 53766 54833 53767
rect -11410 53703 -11344 53704
rect -11410 53639 -11409 53703
rect -11345 53701 -11344 53703
rect -7181 53703 -7115 53704
rect -7181 53701 -7180 53703
rect -11345 53641 -7180 53701
rect -11345 53639 -11344 53641
rect -11410 53638 -11344 53639
rect -7181 53639 -7180 53641
rect -7116 53701 -7115 53703
rect 165 53703 231 53704
rect 165 53701 166 53703
rect -7116 53641 166 53701
rect -7116 53639 -7115 53641
rect -7181 53638 -7115 53639
rect 165 53639 166 53641
rect 230 53639 231 53703
rect 165 53638 231 53639
rect 2195 53703 2261 53704
rect 2195 53639 2196 53703
rect 2260 53701 2261 53703
rect 3729 53703 3795 53704
rect 3729 53701 3730 53703
rect 2260 53641 3730 53701
rect 2260 53639 2261 53641
rect 2195 53638 2261 53639
rect 3729 53639 3730 53641
rect 3794 53639 3795 53703
rect 3729 53638 3795 53639
rect 6114 53703 6180 53704
rect 6114 53639 6115 53703
rect 6179 53701 6180 53703
rect 10343 53703 10409 53704
rect 10343 53701 10344 53703
rect 6179 53641 10344 53701
rect 6179 53639 6180 53641
rect 6114 53638 6180 53639
rect 10343 53639 10344 53641
rect 10408 53701 10409 53703
rect 14421 53703 14487 53704
rect 14421 53701 14422 53703
rect 10408 53641 14422 53701
rect 10408 53639 10409 53641
rect 10343 53638 10409 53639
rect 14421 53639 14422 53641
rect 14486 53639 14487 53703
rect 14421 53638 14487 53639
rect 14876 53703 14942 53704
rect 14876 53639 14877 53703
rect 14941 53701 14942 53703
rect 19105 53703 19171 53704
rect 19105 53701 19106 53703
rect 14941 53641 19106 53701
rect 14941 53639 14942 53641
rect 14876 53638 14942 53639
rect 19105 53639 19106 53641
rect 19170 53701 19171 53703
rect 21549 53703 21615 53704
rect 21549 53701 21550 53703
rect 19170 53641 21550 53701
rect 19170 53639 19171 53641
rect 19105 53638 19171 53639
rect 21549 53639 21550 53641
rect 21614 53639 21615 53703
rect 21549 53638 21615 53639
rect 23638 53703 23704 53704
rect 23638 53639 23639 53703
rect 23703 53701 23704 53703
rect 27867 53703 27933 53704
rect 27867 53701 27868 53703
rect 23703 53641 27868 53701
rect 23703 53639 23704 53641
rect 23638 53638 23704 53639
rect 27867 53639 27868 53641
rect 27932 53701 27933 53703
rect 28677 53703 28743 53704
rect 28677 53701 28678 53703
rect 27932 53641 28678 53701
rect 27932 53639 27933 53641
rect 27867 53638 27933 53639
rect 28677 53639 28678 53641
rect 28742 53639 28743 53703
rect 28677 53638 28743 53639
rect 32400 53703 32466 53704
rect 32400 53639 32401 53703
rect 32465 53701 32466 53703
rect 35805 53703 35871 53704
rect 35805 53701 35806 53703
rect 32465 53641 35806 53701
rect 32465 53639 32466 53641
rect 32400 53638 32466 53639
rect 35805 53639 35806 53641
rect 35870 53701 35871 53703
rect 36629 53703 36695 53704
rect 36629 53701 36630 53703
rect 35870 53641 36630 53701
rect 35870 53639 35871 53641
rect 35805 53638 35871 53639
rect 36629 53639 36630 53641
rect 36694 53639 36695 53703
rect 36629 53638 36695 53639
rect 41162 53703 41228 53704
rect 41162 53639 41163 53703
rect 41227 53701 41228 53703
rect 42933 53703 42999 53704
rect 42933 53701 42934 53703
rect 41227 53641 42934 53701
rect 41227 53639 41228 53641
rect 41162 53638 41228 53639
rect 42933 53639 42934 53641
rect 42998 53701 42999 53703
rect 45391 53703 45457 53704
rect 45391 53701 45392 53703
rect 42998 53641 45392 53701
rect 42998 53639 42999 53641
rect 42933 53638 42999 53639
rect 45391 53639 45392 53641
rect 45456 53639 45457 53703
rect 45391 53638 45457 53639
rect 49924 53703 49990 53704
rect 49924 53639 49925 53703
rect 49989 53701 49990 53703
rect 50061 53703 50127 53704
rect 50061 53701 50062 53703
rect 49989 53641 50062 53701
rect 49989 53639 49990 53641
rect 49924 53638 49990 53639
rect 50061 53639 50062 53641
rect 50126 53701 50127 53703
rect 54153 53703 54219 53704
rect 54153 53701 54154 53703
rect 50126 53641 54154 53701
rect 50126 53639 50127 53641
rect 50061 53638 50127 53639
rect 54153 53639 54154 53641
rect 54218 53639 54219 53703
rect 54153 53638 54219 53639
rect 36462 48035 36528 48036
rect 36462 47971 36463 48035
rect 36527 48033 36528 48035
rect 57145 48035 57211 48036
rect 57145 48033 57146 48035
rect 36527 47973 57146 48033
rect 36527 47971 36528 47973
rect 36462 47970 36528 47971
rect 57145 47971 57146 47973
rect 57210 47971 57211 48035
rect 57145 47970 57211 47971
rect 32518 47907 32584 47908
rect 32518 47843 32519 47907
rect 32583 47905 32584 47907
rect 48383 47907 48449 47908
rect 48383 47905 48384 47907
rect 32583 47845 48384 47905
rect 32583 47843 32584 47845
rect 32518 47842 32584 47843
rect 48383 47843 48384 47845
rect 48448 47843 48449 47907
rect 48383 47842 48449 47843
rect 28574 47779 28640 47780
rect 28574 47715 28575 47779
rect 28639 47777 28640 47779
rect 39621 47779 39687 47780
rect 39621 47777 39622 47779
rect 28639 47717 39622 47777
rect 28639 47715 28640 47717
rect 28574 47714 28640 47715
rect 39621 47715 39622 47717
rect 39686 47715 39687 47779
rect 39621 47714 39687 47715
rect 24630 47651 24696 47652
rect 24630 47587 24631 47651
rect 24695 47649 24696 47651
rect 30859 47651 30925 47652
rect 30859 47649 30860 47651
rect 24695 47589 30860 47649
rect 24695 47587 24696 47589
rect 24630 47586 24696 47587
rect 30859 47587 30860 47589
rect 30924 47587 30925 47651
rect 30859 47586 30925 47587
rect 20686 47523 20752 47524
rect 20686 47459 20687 47523
rect 20751 47521 20752 47523
rect 22097 47523 22163 47524
rect 22097 47521 22098 47523
rect 20751 47461 22098 47521
rect 20751 47459 20752 47461
rect 20686 47458 20752 47459
rect 22097 47459 22098 47461
rect 22162 47459 22163 47523
rect 22097 47458 22163 47459
rect 13335 47395 13401 47396
rect 13335 47331 13336 47395
rect 13400 47393 13401 47395
rect 16742 47395 16808 47396
rect 16742 47393 16743 47395
rect 13400 47333 16743 47393
rect 13400 47331 13401 47333
rect 13335 47330 13401 47331
rect 16742 47331 16743 47333
rect 16807 47331 16808 47395
rect 16742 47330 16808 47331
rect 4573 47267 4639 47268
rect 4573 47203 4574 47267
rect 4638 47265 4639 47267
rect 12798 47267 12864 47268
rect 12798 47265 12799 47267
rect 4638 47205 12799 47265
rect 4638 47203 4639 47205
rect 4573 47202 4639 47203
rect 12798 47203 12799 47205
rect 12863 47203 12864 47267
rect 12798 47202 12864 47203
rect -4189 47139 -4123 47140
rect -4189 47075 -4188 47139
rect -4124 47137 -4123 47139
rect 8854 47139 8920 47140
rect 8854 47137 8855 47139
rect -4124 47077 8855 47137
rect -4124 47075 -4123 47077
rect -4189 47074 -4123 47075
rect 8854 47075 8855 47077
rect 8919 47075 8920 47139
rect 8854 47074 8920 47075
rect 688 42540 44080 42600
rect 41585 26826 41651 26827
rect 41585 26762 41586 26826
rect 41650 26762 41651 26826
rect 41585 26761 41651 26762
rect 48679 26826 48745 26827
rect 48679 26762 48680 26826
rect 48744 26824 48745 26826
rect 52225 26826 52291 26827
rect 52225 26824 52226 26826
rect 48744 26764 52226 26824
rect 48744 26762 48745 26764
rect 48679 26761 48745 26762
rect 52225 26762 52226 26764
rect 52290 26762 52291 26826
rect 52225 26761 52291 26762
rect 41588 25576 41648 26761
rect 41272 25516 41648 25576
<< metal5 >>
rect 51500 20625 51820 20945
use And_Gate  And_Gate_0
timestamp 1761392116
transform 1 0 -10715 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_1
timestamp 1761392116
transform 1 0 -1953 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_2
timestamp 1761392116
transform 1 0 6809 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_3
timestamp 1761392116
transform 1 0 15571 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_4
timestamp 1761392116
transform 1 0 24333 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_5
timestamp 1761392116
transform 1 0 33095 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_6
timestamp 1761392116
transform 1 0 41857 0 1 51955
box -1558 -227 544 1635
use And_Gate  And_Gate_7
timestamp 1761392116
transform 1 0 50619 0 1 51955
box -1558 -227 544 1635
use CDAC_v3  CDAC_v3_0
timestamp 1761401821
transform 1 0 960 0 1 288
box -1004 -280 43852 46738
use Comparator  Comparator_0
timestamp 1761291873
transform -1 0 80195 0 1 12366
box 24473 -2307 30902 29738
use D_FlipFlop  D_FlipFlop_0
timestamp 1761392116
transform 1 0 48670 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_1
timestamp 1761392116
transform 1 0 39908 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_2
timestamp 1761392116
transform 1 0 31146 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_3
timestamp 1761392116
transform 1 0 22384 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_4
timestamp 1761392116
transform 1 0 4860 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_5
timestamp 1761392116
transform 1 0 13622 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_6
timestamp 1761392116
transform 1 0 -3902 0 1 49883
box 0 -1799 8762 1845
use D_FlipFlop  D_FlipFlop_7
timestamp 1761392116
transform 1 0 -12664 0 1 49883
box 0 -1799 8762 1845
use Nand_Gate  Nand_Gate_0
timestamp 1761392116
transform -1 0 4506 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_1
timestamp 1761392116
transform -1 0 -4256 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_2
timestamp 1761392116
transform -1 0 13268 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_3
timestamp 1761392116
transform -1 0 30792 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_4
timestamp 1761392116
transform -1 0 39554 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_5
timestamp 1761392116
transform -1 0 48316 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_6
timestamp 1761392116
transform -1 0 22030 0 1 52275
box 1906 -547 3264 1315
use Nand_Gate  Nand_Gate_7
timestamp 1761392116
transform -1 0 57078 0 1 52275
box 1906 -547 3264 1315
use Ring_Counter  Ring_Counter_0
timestamp 1761401228
transform 0 1 60854 -1 0 63603
box 606 -68808 9368 -8140
<< labels >>
flabel metal4 -4141 47077 8855 47137 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal4 4621 47205 12799 47265 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal4 13383 47333 16743 47393 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal4 20751 47461 22081 47521 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal4 24695 47589 30843 47649 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal4 28639 47717 39599 47777 0 FreeSans 160 0 0 0 Q5
port 8 nsew
flabel metal4 32583 47845 48367 47905 0 FreeSans 160 0 0 0 Q6
port 9 nsew
flabel metal4 36527 47973 57129 48033 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal4 688 42540 44080 42600 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal5 51500 20625 51820 20945 0 FreeSans 1120 0 0 0 Vin
port 13 nsew
flabel metal1 50226 10356 55345 10402 0 FreeSans 160 0 0 0 Vbias
port 11 nsew
flabel metal3 -6421 61680 47040 61740 0 FreeSans 160 0 0 0 EN
port 1 nsew
flabel metal3 57652 47014 57712 61677 0 FreeSans 160 90 0 0 VDD
port 12 nsew
flabel metal3 48912 54459 51277 54519 0 FreeSans 160 0 0 0 FFCLR
flabel metal3 19350 52906 19410 60683 0 FreeSans 160 90 0 0 CLK
port 0 nsew
<< properties >>
string SAR-ADC-using-Sky130-PDK gencell
<< end >>
