** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-11_19-22-56/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 1.27058823525 8.5u 1.27058823525 8.500001u 1.272352941125 17.0u 1.272352941125 17.000001u 1.274117647 25.5u
+ 1.274117647 25.500001u 1.275882352875 34.0u 1.275882352875 34.000001u 1.27764705875 42.5u 1.27764705875 42.500001u 1.279411764625 51.0u
+ 1.279411764625 51.000001u 1.2811764705 59.5u 1.2811764705 59.500001u 1.282941176375 68.0u 1.282941176375 68.000001u 1.28470588225 76.5u
+ 1.28470588225 76.500001u 1.286470588125 85.0u 1.286470588125 85.000001u 1.288235294 93.5u 1.288235294 93.500001u 1.29 102.0u 1.29 102.000001u
+ 1.291764705875 110.5u 1.291764705875 110.500001u 1.29352941175 119.0u 1.29352941175 119.000001u 1.295294117625 127.5u 1.295294117625 127.500001u
+ 1.2970588235 136.0u 1.2970588235 136.000001u 1.298823529375 144.5u 1.298823529375 144.500001u 1.30058823525 153.0u 1.30058823525 153.000001u
+ 1.302352941125 161.5u 1.302352941125 161.500001u 1.304117647 170.0u 1.304117647 170.000001u 1.305882352875 178.5u 1.305882352875)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ff

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 178.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-11_19-22-56/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
