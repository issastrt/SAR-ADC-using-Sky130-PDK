* NGSPICE file created from SAR-ADC-using-Sky130-PDK.ext - technology: sky130A

.subckt SAR-ADC-using-Sky130-PDK CLK Q0 Q1 Q2 Q3 Q4 Q6 Q5 Q7 VDD Vin EN GND Vbias
X0 Comparator_0.Vinm CDAC8_0.switch_7.Z.t131 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1 a_64511_52572# EN.t0 Vbias.t123 Vbias.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X2 a_45761_13083# CLK.t0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 Vbias.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X3 Vbias.t117 EN.t1 a_29289_15797# Vbias.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X4 VDD.t698 Nand_Gate_4.A.t4 RingCounter_0.D_FlipFlop_8.Q' VDD.t689 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X5 D_FlipFlop_6.3-input-nand_2.C.t2 D_FlipFlop_6.3-input-nand_1.Vout VDD.t713 VDD.t712 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X6 a_51499_49858# EN.t2 Vbias.t115 Vbias.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X7 Vbias.t121 EN.t3 a_46375_13083# Vbias.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 VDD.t814 VDD.t815 VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X9 a_100961_13083# CLK.t1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 Vbias.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X10 Comparator_0.Vinm CDAC8_0.switch_7.Z.t130 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X11 Comparator_0.Vinm CDAC8_0.switch_8.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X12 D_FlipFlop_7.Q' D_FlipFlop_7.Nand_Gate_1.Vout VDD.t489 VDD.t472 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X13 a_124399_52572# RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_123785_52572# Vbias.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X14 a_68585_52572# EN.t4 Vbias.t119 Vbias.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X15 a_51369_13083# RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 a_50755_13083# Vbias.t753 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X16 Comparator_0.Vinm CDAC8_0.switch_6.Z.t67 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X17 VDD.t239 D_FlipFlop_1.3-input-nand_2.Vout.t4 D_FlipFlop_1.3-input-nand_2.C.t3 VDD.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X18 Vbias.t113 EN.t5 a_101575_13083# Vbias.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X19 a_65125_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_64511_52572# Vbias.t579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X20 Comparator_0.Vinm CDAC8_0.switch_6.Z.t66 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X21 Comparator_0.Vinm CDAC8_0.switch_6.Z.t65 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X22 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_0.D.t3 VDD.t631 VDD.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X23 VDD.t1100 CLK.t2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 VDD.t1048 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X24 Nand_Gate_0.A.t2 RingCounter_0.D_FlipFlop_2.Q' a_69199_52572# Vbias.t361 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X25 Comparator_0.Vinm CDAC8_0.switch_6.Z.t64 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X26 VDD.t130 EN.t6 D_FlipFlop_1.3-input-nand_2.C.t0 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X27 a_52113_49858# RingCounter_0.D_FlipFlop_1.Inverter_0.Vout a_51499_49858# Vbias.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X28 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 a_56187_49858# Vbias.t556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X29 VDD.t366 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 VDD.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X30 VDD.t610 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_2.A.t3 VDD.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X31 a_48565_16975# CLK.t3 Vbias.t329 Vbias.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X32 a_134283_17072# And_Gate_1.Vout.t2 D_FlipFlop_7.3-input-nand_1.Vout Vbias.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X33 VDD.t861 Nand_Gate_2.B.t4 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X34 VDD.t818 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 VDD.t817 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X35 a_123785_52572# EN.t7 Vbias.t111 Vbias.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X36 VDD.t613 And_Gate_4.Vout.t2 D_FlipFlop_2.3-input-nand_1.Vout VDD.t612 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X37 And_Gate_7.Vout.t1 And_Gate_7.Inverter_0.Vin Vbias.t740 Vbias.t739 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X38 a_134283_27764# And_Gate_3.Vout.t2 D_FlipFlop_4.3-input-nand_1.Vout Vbias.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X39 a_71017_47663# Nand_Gate_0.A.t4 Vbias.t724 Vbias.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X40 a_74807_15797# RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout Vbias.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X41 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_2.3-input-nand_2.C.t4 VDD.t137 VDD.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X42 Comparator_0.Vinm CDAC8_0.switch_9.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X43 Nand_Gate_5.B.t3 RingCounter_0.D_FlipFlop_6.Q' a_124399_52572# Vbias.t536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X44 Vbias.t232 VDD.t1108 a_51369_13083# Vbias.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X45 Comparator_0.Vinm CDAC8_0.switch_7.Z.t129 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X46 a_79495_15797# Nand_Gate_6.A.t4 a_78881_15797# Vbias.t712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X47 Nand_Gate_6.A.t3 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t626 VDD.t625 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X48 Vbias.t433 FFCLR.t4 a_132925_37007# Vbias.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X49 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 a_111387_49858# Vbias.t892 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X50 a_107927_13083# RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 Vbias.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X51 a_56187_49858# RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 Vbias.t543 Vbias.t542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X52 Comparator_0.Vinm CDAC8_0.switch_7.Z.t128 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X53 Comparator_0.Vinm CDAC8_0.switch_9.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X54 Vbias.t234 VDD.t1109 a_57415_15797# Vbias.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X55 a_134897_43285# D_FlipFlop_0.D.t4 a_134283_43285# Vbias.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X56 Nand_Gate_2.A.t1 RingCounter_0.D_FlipFlop_4.Q' VDD.t488 VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X57 a_108671_52572# EN.t8 Vbias.t109 Vbias.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X58 VDD.t970 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t969 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X59 Comparator_0.Vinm CDAC8_0.switch_8.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X60 VDD.t128 EN.t9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 VDD.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X61 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 a_109285_52572# Vbias.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X62 Comparator_0.Vinm CDAC8_0.switch_7.Z.t127 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X63 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 VDD.t812 VDD.t813 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X64 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 EN.t10 VDD.t126 VDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X65 D_FlipFlop_1.3-input-nand_2.Vout.t2 D_FlipFlop_1.3-input-nand_0.Vout VDD.t682 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X66 VDD.t487 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 VDD.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X67 a_76909_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 Vbias.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X68 Comparator_0.Vinm CDAC8_0.switch_6.Z.t63 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X69 VDD.t124 EN.t11 Nand_Gate_6.A.t0 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X70 Vbias.t236 VDD.t1110 a_112615_15797# Vbias.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X71 D_FlipFlop_0.3-input-nand_2.Vout.t2 D_FlipFlop_0.3-input-nand_0.Vout VDD.t606 VDD.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X72 a_110029_13083# RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 Vbias.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X73 VDD.t955 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 VDD.t954 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X74 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 CLK.t4 Vbias.t331 Vbias.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X75 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 VDD.t841 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X76 Vbias.t434 D_FlipFlop_5.3-input-nand_2.C.t4 a_130209_24200# Vbias.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X77 a_75898_39392# Q6.t4 Vbias.t759 Vbias.t758 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X78 Comparator_0.Vinm CDAC8_0.switch_7.Z.t126 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X79 CDAC8_0.switch_2.Z.t2 a_75898_21528# VDD.t557 VDD.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X80 Comparator_0.Vinm CDAC8_0.switch_8.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X81 VDD.t402 Q3.t4 CDAC8_0.switch_5.Z.t2 Vbias.t436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X82 Nand_Gate_5.Vout.t2 Nand_Gate_5.B.t4 a_115177_47663# Vbias.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X83 a_109285_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_108671_52572# Vbias.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X84 Vbias.t617 Nand_Gate_6.B.t4 a_134897_24200# Vbias.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X85 VDD.t389 FFCLR.t5 D_FlipFlop_5.3-input-nand_0.Vout VDD.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X86 VDD.t1099 CLK.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 VDD.t1045 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X87 Vbias.t333 CLK.t6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 Vbias.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X88 VDD.t459 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_5.Q' VDD.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X89 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout Nand_Gate_2.A.t4 Vbias.t708 Vbias.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X90 RingCounter_0.D_FlipFlop_17.Q' EN.t12 VDD.t122 VDD.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X91 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t810 VDD.t811 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X92 VDD.t404 Q3.t5 D_FlipFlop_4.Q' VDD.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X93 VDD.t899 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 VDD.t219 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X94 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 CLK.t7 Vbias.t335 Vbias.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X95 VDD.t551 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 VDD.t550 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X96 a_86591_49858# VDD.t1111 Vbias.t238 Vbias.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X97 RingCounter_0.D_FlipFlop_17.Q' FFCLR.t6 VDD.t391 VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X98 VDD.t1098 CLK.t8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 VDD.t1042 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X99 CDAC8_0.switch_5.Z.t1 a_75898_28676# Vbias.t764 Vbias.t763 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X100 a_115177_47663# Nand_Gate_5.A.t4 Vbias.t830 Vbias.t829 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X101 a_118967_15797# RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout Vbias.t858 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X102 RingCounter_0.D_FlipFlop_5.Q' VDD.t808 VDD.t809 VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X103 Nand_Gate_4.B.t0 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X104 Comparator_0.Vinm CDAC8_0.switch_9.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X105 a_132311_40571# D_FlipFlop_3.3-input-nand_2.Vout.t4 D_FlipFlop_3.3-input-nand_2.C.t2 Vbias.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X106 Comparator_0.Vinm CDAC8_0.switch_7.Z.t125 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X107 Vbias.t652 D_FlipFlop_0.D.t5 D_FlipFlop_5.Inverter_0.Vout Vbias.t651 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X108 VDD.t177 D_FlipFlop_3.3-input-nand_2.C.t4 D_FlipFlop_3.3-input-nand_2.Vout.t0 VDD.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X109 Vbias.t856 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 a_85847_13083# Vbias.t855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X110 VDD.t393 FFCLR.t7 D_FlipFlop_2.3-input-nand_0.Vout VDD.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X111 RingCounter_0.D_FlipFlop_5.Q' Nand_Gate_2.B.t5 VDD.t863 VDD.t862 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X112 Comparator_0.Vinm CDAC8_0.switch_7.Z.t124 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X113 a_128237_39721# D_FlipFlop_2.Q' Q6.t3 Vbias.t775 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X114 D_FlipFlop_4.Q' D_FlipFlop_4.Nand_Gate_1.Vout VDD.t888 VDD.t887 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X115 VDD.t708 Nand_Gate_2.A.t5 D_FlipFlop_3.3-input-nand_2.Vout.t2 VDD.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X116 VDD.t383 D_FlipFlop_0.3-input-nand_2.Vout.t4 D_FlipFlop_0.3-input-nand_2.C.t1 VDD.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X117 VDD.t951 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout VDD.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X118 VDD.t892 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout VDD.t890 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X119 a_87205_49858# RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 a_86591_49858# Vbias.t449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X120 a_139496_37417.t1 a_139496_37417.t0 VDD.t700 VDD.t699 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X121 Vbias.t709 Nand_Gate_2.A.t6 a_128851_43285# Vbias.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X122 Vbias.t584 D_FlipFlop_6.3-input-nand_2.C.t4 a_130209_20636# Vbias.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X123 VDD.t395 FFCLR.t8 D_FlipFlop_0.3-input-nand_2.C.t3 VDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X124 VDD.t120 EN.t13 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 VDD.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X125 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 CLK.t9 a_41073_52572# Vbias.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X126 VDD.t118 EN.t14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X127 Comparator_0.Vinm CDAC8_0.switch_8.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X128 a_43789_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 Vbias.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X129 Vbias.t551 Nand_Gate_7.B.t4 a_134897_20636# Vbias.t550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X130 VDD.t397 FFCLR.t9 D_FlipFlop_6.3-input-nand_0.Vout VDD.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X131 a_128237_23350# D_FlipFlop_6.Q' Q1.t3 Vbias.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X132 CDAC8_0.switch_6.Z.t0 a_75898_39392# VDD.t619 VDD.t618 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X133 VDD.t116 EN.t15 Nand_Gate_4.B.t1 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X134 a_139696_27690# Vin.t0 a_138366_35417.t1 Vbias.t548 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X135 Comparator_0.Vinm CDAC8_0.switch_7.Z.t123 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X136 Comparator_0.Vinm CDAC8_0.switch_6.Z.t62 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X137 a_132925_40571# D_FlipFlop_3.3-input-nand_1.Vout a_132311_40571# Vbias.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X138 VDD.t526 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 VDD.t525 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X139 Comparator_0.Vinm CDAC8_0.switch_7.Z.t122 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X140 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 VDD.t952 VDD.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X141 CDAC8_0.switch_1.Z.t0 a_75898_18814# VDD.t283 VDD.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X142 a_75898_28676# Q3.t6 VDD.t406 VDD.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X143 a_134897_19786# D_FlipFlop_0.D.t6 a_134283_19786# Vbias.t653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X144 VDD.t446 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 VDD.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X145 a_103765_47663# Nand_Gate_2.Vout.t3 Vbias.t720 Vbias.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X146 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout Nand_Gate_3.B.t4 Vbias.t421 Vbias.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X147 Vbias.t338 CLK.t10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 Vbias.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X148 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t806 VDD.t807 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X149 VDD.t449 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X150 And_Gate_3.Vout.t0 And_Gate_3.Inverter_0.Vin VDD.t590 VDD.t589 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X151 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 CLK.t11 VDD.t1090 VDD.t1089 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X152 Comparator_0.Vinm CDAC8_0.switch_6.Z.t61 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X153 VDD.t114 EN.t16 Nand_Gate_1.B.t0 VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X154 VDD.t18 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X155 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 CLK.t12 a_96273_49858# Vbias.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X156 Vbias.t284 Q7.t4 CDAC8_0.switch_7.Z.t0 VDD.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X157 VDD.t243 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X158 Vbias.t345 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 a_52727_13083# Vbias.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X159 VDD.t458 And_Gate_5.Vout.t2 D_FlipFlop_1.3-input-nand_1.Vout VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X160 Comparator_0.Vinm CDAC8_0.switch_7.Z.t121 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X161 VDD.t378 Nand_Gate_3.B.t5 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD.t377 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X162 Comparator_0.Vinm CDAC8_0.switch_7.Z.t120 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X163 D_FlipFlop_1.Nand_Gate_1.Vout D_FlipFlop_1.3-input-nand_2.C.t4 VDD.t231 VDD.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X164 a_57545_49858# VDD.t1112 Vbias.t240 Vbias.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X165 Comparator_0.Vinm CDAC8_0.switch_7.Z.t119 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X166 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 VDD.t856 VDD.t855 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X167 Comparator_0.Vinm CDAC8_0.switch_9.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X168 a_138366_35417.t2 D_FlipFlop_0.D.t0 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X169 a_75898_42964# Q5.t4 VDD.t385 VDD.t384 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X170 a_130209_33443# D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout Vbias.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X171 VDD.t444 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout VDD.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X172 VDD.t562 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 VDD.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X173 VDD.t630 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_0.Vout VDD.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X174 a_112745_49858# VDD.t1113 Vbias.t242 Vbias.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X175 VDD.t874 D_FlipFlop_7.3-input-nand_2.C.t4 D_FlipFlop_7.3-input-nand_2.Vout.t3 VDD.t873 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X176 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 VDD.t656 VDD.t655 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X177 Vbias.t129 D_FlipFlop_2.3-input-nand_2.C.t5 a_130209_37007# Vbias.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X178 Nand_Gate_1.Vout.t1 Nand_Gate_1.B.t4 VDD.t368 VDD.t367 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X179 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 VDD.t661 VDD.t660 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X180 Vbias.t725 Nand_Gate_0.A.t5 a_134897_37007# Vbias.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X181 Comparator_0.Vinm CDAC8_0.switch_7.Z.t118 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X182 a_69199_52572# RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_68585_52572# Vbias.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X183 Comparator_0.Vinm CDAC8_0.switch_7.Z.t117 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X184 Vbias.t367 Nand_Gate_7.A.t4 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout Vbias.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X185 VDD.t1101 Nand_Gate_4.B.t4 D_FlipFlop_7.3-input-nand_2.Vout.t1 VDD.t985 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X186 Comparator_0.Vinm CDAC8_0.switch_7.Z.t116 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X187 a_138318_16817# a_138318_16817# Vbias.t473 Vbias.t472 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X188 Comparator_0.Vinm CDAC8_0.switch_9.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X189 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout Nand_Gate_2.B.t6 Vbias.t602 Vbias.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X190 Vbias.t887 Nand_Gate_4.B.t5 a_128851_19786# Vbias.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X191 a_132311_26914# D_FlipFlop_5.3-input-nand_2.C.t5 D_FlipFlop_5.3-input-nand_2.Vout.t1 Vbias.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X192 a_72835_13083# Nand_Gate_7.B.t5 RingCounter_0.D_FlipFlop_13.Q' Vbias.t552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X193 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD.t804 VDD.t805 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X194 a_77523_13083# RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 a_76909_13083# Vbias.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X195 Comparator_0.Vinm CDAC8_0.switch_6.Z.t60 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X196 a_73579_52572# VDD.t1114 Vbias.t244 Vbias.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X197 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK.t13 VDD.t1097 VDD.t1030 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X198 Vbias.t416 Nand_Gate_1.B.t5 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout Vbias.t415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X199 VDD.t195 FFCLR.t10 D_FlipFlop_6.Q' VDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X200 Vbias.t465 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 a_63767_15797# Vbias.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X201 Vbias.t810 And_Gate_2.Vout.t2 D_FlipFlop_5.Inverter_1.Vout Vbias.t809 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X202 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 CLK.t14 a_63153_49858# Vbias.t340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X203 Comparator_0.Vinm CDAC8_0.switch_6.Z.t59 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X204 VDD.t1091 CLK.t15 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 VDD.t1050 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X205 VDD.t16 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X206 Comparator_0.Vinm CDAC8_0.switch_7.Z.t115 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X207 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 CLK.t16 VDD.t1096 VDD.t1060 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X208 Comparator_0.Vinm CDAC8_0.switch_6.Z.t58 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X209 a_132925_26914# D_FlipFlop_5.3-input-nand_0.Vout a_132311_26914# Vbias.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X210 VDD.t8 And_Gate_4.A.t3 And_Gate_4.Inverter_0.Vin VDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X211 Comparator_0.Vinm CDAC8_0.switch_6.Z.t57 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X212 VDD.t1103 Nand_Gate_4.B.t6 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout VDD.t1102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X213 Vbias.t246 VDD.t1115 a_77523_13083# Vbias.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X214 Comparator_0.Vinm CDAC8_0.switch_7.Z.t114 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X215 Comparator_0.Vinm CDAC8_0.switch_7.Z.t113 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X216 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 EN.t17 VDD.t112 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X217 a_84489_15797# RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_83875_15797# Vbias.t648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X218 Comparator_0.Vinm CDAC8_0.switch_9.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X219 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 a_78267_52572# Vbias.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X220 a_75898_25104# Q2.t4 VDD.t641 VDD.t640 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X221 VDD.t709 Nand_Gate_2.A.t7 D_FlipFlop_3.3-input-nand_1.Vout VDD.t648 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X222 a_128237_36157# D_FlipFlop_1.Q' Q7.t0 Vbias.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X223 a_117609_13083# RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 a_116995_13083# Vbias.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X224 RingCounter_0.D_FlipFlop_11.Q' RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 VDD.t461 VDD.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X225 VDD.t110 EN.t18 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X226 VDD.t921 Nand_Gate_1.A.t4 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout VDD.t920 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X227 VDD.t988 Q6.t5 CDAC8_0.switch_6.Z.t2 Vbias.t883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X228 a_128237_46849# D_FlipFlop_0.Q' Q4.t1 Vbias.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X229 Comparator_0.Vinm CDAC8_0.switch_7.Z.t112 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X230 Vbias.t727 Nand_Gate_0.A.t6 a_132925_39721# Vbias.t726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X231 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 VDD.t528 VDD.t527 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X232 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_0.D.t7 VDD.t844 VDD.t843 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X233 a_83875_15797# RingCounter_0.D_FlipFlop_12.Q' Nand_Gate_6.A.t1 Vbias.t494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X234 VDD.t515 And_Gate_6.Vout.t2 D_FlipFlop_3.3-input-nand_0.Vout VDD.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X235 a_88563_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 a_87949_15797# Vbias.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X236 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.3-input-nand_2.Vout.t5 VDD.t287 VDD.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X237 Comparator_0.Vinm CDAC8_0.switch_7.Z.t111 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X238 VDD.t1095 CLK.t17 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 VDD.t1094 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X239 Comparator_0.Vinm CDAC8_0.switch_7.Z.t110 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X240 Vbias.t107 EN.t19 a_84489_15797# Vbias.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X241 VDD.t579 Nand_Gate_6.B.t5 RingCounter_0.D_FlipFlop_11.Q' VDD.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X242 Vbias.t388 And_Gate_0.Vout.t2 D_FlipFlop_6.Inverter_1.Vout Vbias.t387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X243 VDD.t412 And_Gate_7.Vout.t2 D_FlipFlop_0.3-input-nand_1.Vout VDD.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X244 VDD.t889 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Q' VDD.t706 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X245 a_128237_30478# D_FlipFlop_4.Q' Q3.t1 Vbias.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X246 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_0.3-input-nand_2.C.t4 VDD.t479 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X247 a_44403_13083# RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 a_43789_13083# Vbias.t476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X248 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 VDD.t513 VDD.t512 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X249 CDAC8_0.switch_6.Z.t1 a_75898_39392# Vbias.t645 Vbias.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X250 Vbias.t553 Nand_Gate_7.B.t6 a_132925_23350# Vbias.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X251 And_Gate_7.Inverter_0.Vin CLK.t18 VDD.t1093 VDD.t1092 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X252 And_Gate_5.A.t1 Nand_Gate_3.B.t6 VDD.t380 VDD.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X253 a_40459_52572# EN.t20 Vbias.t105 Vbias.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X254 Vbias.t248 VDD.t1116 a_117609_13083# Vbias.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X255 VDD.t803 VDD.t802 RingCounter_0.D_FlipFlop_11.Q' VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X256 a_134283_24200# And_Gate_2.Vout.t3 D_FlipFlop_5.3-input-nand_1.Vout Vbias.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X257 VDD.t801 VDD.t800 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X258 a_130209_44135# D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout Vbias.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X259 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 Nand_Gate_7.A.t5 VDD.t319 VDD.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X260 a_132311_17072# D_FlipFlop_7.3-input-nand_2.Vout.t4 D_FlipFlop_7.3-input-nand_2.C.t1 Vbias.t798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X261 VDD.t196 FFCLR.t11 Q7.t3 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X262 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 EN.t21 VDD.t108 VDD.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X263 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_0.D.t8 VDD.t845 VDD.t585 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X264 a_134897_40571# D_FlipFlop_3.Inverter_0.Vout a_134283_40571# Vbias.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X265 Vbias.t103 EN.t22 a_88563_15797# Vbias.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X266 Comparator_0.Vinm CDAC8_0.switch_8.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X267 a_132311_27764# D_FlipFlop_4.3-input-nand_2.Vout.t4 D_FlipFlop_4.3-input-nand_2.C.t0 Vbias.t435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X268 VDD.t864 D_FlipFlop_4.3-input-nand_2.C.t4 D_FlipFlop_4.3-input-nand_2.Vout.t2 VDD.t687 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X269 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 VDD.t930 VDD.t543 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X270 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 CLK.t19 VDD.t1088 VDD.t1056 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X271 a_29289_13083# RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 a_28675_13083# Vbias.t705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X272 Comparator_0.Vinm CDAC8_0.switch_7.Z.t109 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X273 VDD.t936 Nand_Gate_5.A.t5 Q4.t3 VDD.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X274 Comparator_0.Vinm CDAC8_0.switch_7.Z.t108 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X275 Comparator_0.Vinm CDAC8_0.switch_0.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X276 VDD.t519 RingCounter_0.D_FlipFlop_13.Q' Nand_Gate_7.B.t3 VDD.t355 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X277 a_128851_43285# D_FlipFlop_3.Nand_Gate_0.Vout a_128237_43285# Vbias.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X278 Comparator_0.Vinm CDAC8_0.switch_6.Z.t56 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X279 Vbias.t250 VDD.t1117 a_44403_13083# Vbias.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X280 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 Nand_Gate_1.B.t6 VDD.t880 VDD.t646 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X281 VDD.t882 Nand_Gate_1.B.t7 D_FlipFlop_4.3-input-nand_2.Vout.t0 VDD.t881 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X282 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 VDD.t894 VDD.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X283 Comparator_0.Vinm CDAC8_0.switch_6.Z.t55 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X284 a_41073_52572# RingCounter_0.D_FlipFlop_16.Q.t4 a_40459_52572# Vbias.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X285 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_0.D.t9 VDD.t847 VDD.t846 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X286 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 a_76165_49858# Vbias.t317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X287 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 a_45147_52572# Vbias.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X288 VDD.t10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X289 a_132925_17072# D_FlipFlop_7.3-input-nand_1.Vout a_132311_17072# Vbias.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X290 VDD.t611 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 VDD.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X291 VDD.t106 EN.t23 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X292 a_28675_13083# RingCounter_0.D_FlipFlop_16.Q.t5 RingCounter_0.D_FlipFlop_16.Q' Vbias.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X293 a_122427_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 Vbias.t301 Vbias.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X294 Vbias.t437 Q3.t7 CDAC8_0.switch_5.Z.t3 VDD.t407 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X295 a_95659_49858# EN.t24 Vbias.t101 Vbias.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X296 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 VDD.t530 VDD.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X297 a_132925_27764# D_FlipFlop_4.3-input-nand_1.Vout a_132311_27764# Vbias.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X298 Vbias.t252 VDD.t1118 a_29289_13083# Vbias.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X299 a_82057_16975# Nand_Gate_6.A.t5 Vbias.t714 Vbias.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X300 Comparator_0.Vinm CDAC8_0.switch_7.Z.t107 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X301 a_50755_15797# RingCounter_0.D_FlipFlop_15.Q' Nand_Gate_4.B.t2 Vbias.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X302 a_134283_20636# And_Gate_0.Vout.t3 D_FlipFlop_6.3-input-nand_1.Vout Vbias.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X303 Comparator_0.Vinm CDAC8_0.switch_7.Z.t106 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X304 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 a_100347_52572# Vbias.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X305 Nand_Gate_0.A.t0 EN.t25 VDD.t104 VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X306 a_55443_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 a_54829_15797# Vbias.t847 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X307 VDD.t549 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 VDD.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X308 VDD.t321 Nand_Gate_7.A.t6 RingCounter_0.D_FlipFlop_14.Q' VDD.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X309 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 VDD.t508 VDD.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X310 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 VDD.t477 VDD.t476 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X311 VDD.t1104 Nand_Gate_4.B.t7 D_FlipFlop_7.3-input-nand_1.Vout VDD.t650 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X312 a_107313_52572# Nand_Gate_2.B.t7 a_106699_52572# Vbias.t603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X313 Comparator_0.Vinm CDAC8_0.switch_6.Z.t54 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X314 VDD.t799 VDD.t798 RingCounter_0.D_FlipFlop_14.Q' VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X315 Comparator_0.Vinm CDAC8_0.switch_7.Z.t105 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X316 a_96273_49858# RingCounter_0.D_FlipFlop_5.Inverter_0.Vout a_95659_49858# Vbias.t894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X317 Comparator_0.Vinm CDAC8_0.switch_9.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X318 VDD.t408 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 VDD.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X319 Nand_Gate_5.B.t0 EN.t26 VDD.t102 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X320 a_110643_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 a_110029_15797# Vbias.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X321 CDAC8_0.switch_7.Z.t2 a_75898_35820# VDD.t382 VDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X322 Vbias.t638 And_Gate_4.Vout.t3 D_FlipFlop_2.Inverter_1.Vout Vbias.t637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X323 Comparator_0.Vinm CDAC8_0.switch_9.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X324 VDD.t270 And_Gate_1.Vout.t3 D_FlipFlop_7.3-input-nand_0.Vout VDD.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X325 a_90665_52572# EN.t27 Vbias.t99 Vbias.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X326 Comparator_0.Vinm CDAC8_0.switch_6.Z.t53 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X327 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 VDD.t261 VDD.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X328 Vbias.t97 EN.t28 a_55443_15797# Vbias.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X329 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.3-input-nand_2.Vout.t5 VDD.t922 VDD.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X330 Vbias.t166 FFCLR.t12 a_128851_40571# Vbias.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X331 Nand_Gate_2.A.t2 RingCounter_0.D_FlipFlop_4.Q' a_91279_52572# Vbias.t532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X332 VDD.t481 RingCounter_0.D_FlipFlop_10.Q' Nand_Gate_1.B.t2 VDD.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X333 Comparator_0.Vinm CDAC8_0.switch_7.Z.t104 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X334 Vbias.t426 Q5.t5 CDAC8_0.switch_9.Z.t2 VDD.t386 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X335 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK.t20 a_107313_52572# Vbias.t480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X336 And_Gate_1.Vout.t1 And_Gate_1.Inverter_0.Vin Vbias.t369 Vbias.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X337 a_74807_13083# RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 Vbias.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X338 a_70645_16975# CLK.t21 Vbias.t482 Vbias.t481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X339 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 EN.t29 VDD.t100 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X340 Comparator_0.Vinm CDAC8_0.switch_8.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X341 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 a_43045_49858# Vbias.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X342 a_79495_13083# RingCounter_0.D_FlipFlop_13.Inverter_0.Vout a_78881_13083# Vbias.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X343 Vbias.t91 EN.t30 a_110643_15797# Vbias.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X344 a_120325_49858# RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 a_119711_49858# Vbias.t716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X345 a_75551_52572# EN.t31 Vbias.t95 Vbias.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X346 VDD.t158 Q1.t4 D_FlipFlop_6.Q' VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X347 RingCounter_0.D_FlipFlop_9.Q' RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 VDD.t999 VDD.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X348 VDD.t871 Nand_Gate_1.A.t5 Nand_Gate_1.Vout.t2 VDD.t870 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X349 VDD.t338 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X350 a_62539_49858# EN.t32 Vbias.t93 Vbias.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X351 Vbias.t89 EN.t33 a_57415_13083# Vbias.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X352 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 VDD.t796 VDD.t797 VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X353 a_128851_19786# D_FlipFlop_7.Nand_Gate_0.Vout a_128237_19786# Vbias.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X354 D_FlipFlop_5.3-input-nand_2.C.t2 D_FlipFlop_5.3-input-nand_1.Vout VDD.t594 VDD.t593 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X355 a_134897_26914# D_FlipFlop_0.D.t10 a_134283_26914# Vbias.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X356 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 VDD.t678 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X357 a_76909_13083# RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 Vbias.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X358 Comparator_0.Vinm CDAC8_0.switch_7.Z.t103 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X359 Vbias.t168 FFCLR.t13 a_132925_36157# Vbias.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X360 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 VDD.t165 VDD.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X361 a_89307_49858# RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 Vbias.t12 Vbias.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X362 Vbias.t87 EN.t34 a_112615_13083# Vbias.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X363 VDD.t98 EN.t35 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X364 a_134283_37007# And_Gate_4.Vout.t4 D_FlipFlop_2.3-input-nand_1.Vout Vbias.t502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X365 a_76165_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_75551_52572# Vbias.t852 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X366 D_FlipFlop_6.Q' D_FlipFlop_6.Nand_Gate_1.Vout VDD.t893 VDD.t662 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X367 VDD.t795 VDD.t794 RingCounter_0.D_FlipFlop_9.Q' VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X368 VDD.t537 RingCounter_0.D_FlipFlop_16.Q' RingCounter_0.D_FlipFlop_16.Q.t2 VDD.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X369 Vbias.t832 Nand_Gate_5.A.t6 a_132925_46849# Vbias.t831 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X370 Comparator_0.Vinm CDAC8_0.switch_6.Z.t52 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X371 a_63153_49858# RingCounter_0.D_FlipFlop_2.Inverter_0.Vout a_62539_49858# Vbias.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X372 And_Gate_3.Inverter_0.Vin Nand_Gate_1.Vout.t3 a_114805_16975# Vbias.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X373 And_Gate_1.B.t1 Nand_Gate_4.B.t8 a_37897_16975# Vbias.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X374 VDD.t935 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 VDD.t615 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X375 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 a_67227_49858# Vbias.t756 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X376 Comparator_0.Vinm CDAC8_0.switch_7.Z.t102 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X377 Vbias.t519 D_FlipFlop_2.3-input-nand_2.Vout.t4 a_130209_39721# Vbias.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X378 Comparator_0.Vinm CDAC8_0.switch_9.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X379 VDD.t496 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 VDD.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X380 Vbias.t169 FFCLR.t14 a_134897_39721# Vbias.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X381 Comparator_0.Vinm CDAC8_0.switch_6.Z.t51 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X382 a_85847_15797# RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout Vbias.t401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X383 VDD.t849 D_FlipFlop_0.D.t11 D_FlipFlop_3.Inverter_0.Vout VDD.t848 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X384 Vbias.t771 Nand_Gate_1.B.t8 a_132925_30478# Vbias.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X385 Comparator_0.Vinm CDAC8_0.switch_7.Z.t101 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X386 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 a_122427_49858# Vbias.t679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X387 a_118967_13083# RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 Vbias.t859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X388 Vbias.t661 Q2.t5 CDAC8_0.switch_0.Z.t1 VDD.t642 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X389 Vbias.t149 D_FlipFlop_6.3-input-nand_2.Vout.t4 a_130209_23350# Vbias.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X390 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_3.Inverter_0.Vout VDD.t317 VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X391 Comparator_0.Vinm CDAC8_0.switch_8.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X392 Vbias.t171 FFCLR.t15 a_134897_23350# Vbias.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X393 Vbias.t254 VDD.t1119 a_68455_15797# Vbias.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X394 a_42431_52572# VDD.t1120 Vbias.t256 Vbias.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X395 VDD.t883 Nand_Gate_1.B.t9 D_FlipFlop_4.3-input-nand_1.Vout VDD.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X396 Comparator_0.Vinm CDAC8_0.switch_9.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X397 VDD.t296 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD.t295 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X398 VDD.t189 D_FlipFlop_1.Q' Q7.t1 VDD.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X399 VDD.t96 EN.t36 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 VDD.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X400 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 VDD.t792 VDD.t793 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X401 a_87949_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 Vbias.t857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X402 VDD.t218 D_FlipFlop_0.Q' Q4.t2 VDD.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X403 VDD.t417 And_Gate_3.Vout.t3 D_FlipFlop_4.3-input-nand_0.Vout VDD.t416 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X404 Vbias.t258 VDD.t1121 a_123655_15797# Vbias.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X405 a_43789_13083# RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 Vbias.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X406 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.3-input-nand_2.Vout.t5 VDD.t680 VDD.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X407 VDD.t222 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 VDD.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X408 Comparator_0.Vinm CDAC8_0.switch_7.Z.t100 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X409 Vbias.t618 Nand_Gate_6.B.t6 a_128851_26914# Vbias.t524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X410 VDD.t198 FFCLR.t16 And_Gate_5.A.t2 VDD.t197 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X411 a_102319_52572# RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_101705_52572# Vbias.t347 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X412 Comparator_0.Vinm CDAC8_0.switch_0.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X413 Comparator_0.Vinm CDAC8_0.switch_7.Z.t99 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X414 a_43045_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 a_42431_52572# Vbias.t874 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X415 VDD.t1087 CLK.t22 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 VDD.t1018 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X416 a_91279_49858# RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 a_90665_49858# Vbias.t479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X417 VDD.t145 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_7.Q' VDD.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X418 FFCLR.t2 RingCounter_0.D_FlipFlop_17.Q' a_47119_52572# Vbias.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X419 Q7.t2 D_FlipFlop_1.Nand_Gate_0.Vout VDD.t362 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X420 a_134897_17072# D_FlipFlop_7.Inverter_0.Vout a_134283_17072# Vbias.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X421 VDD.t791 VDD.t790 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X422 VDD.t300 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 VDD.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X423 a_97631_49858# VDD.t1122 Vbias.t260 Vbias.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X424 RingCounter_0.D_FlipFlop_1.Q' Nand_Gate_3.B.t7 VDD.t208 VDD.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X425 VDD.t167 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 VDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X426 Q4.t0 D_FlipFlop_0.Nand_Gate_0.Vout VDD.t193 VDD.t192 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X427 a_134897_27764# D_FlipFlop_4.Inverter_0.Vout a_134283_27764# Vbias.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X428 And_Gate_6.Vout.t1 And_Gate_6.Inverter_0.Vin Vbias.t656 Vbias.t655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X429 VDD.t1086 CLK.t23 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 VDD.t1016 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X430 a_52727_15797# RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout Vbias.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X431 Comparator_0.Vinm CDAC8_0.switch_7.Z.t98 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X432 Nand_Gate_2.B.t2 RingCounter_0.D_FlipFlop_5.Q' a_102319_52572# Vbias.t765 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X433 a_57415_15797# Nand_Gate_7.A.t7 a_56801_15797# Vbias.t769 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X434 Comparator_0.Vinm CDAC8_0.switch_9.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X435 a_128237_33443# Q7.t5 D_FlipFlop_1.Q' Vbias.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X436 Nand_Gate_7.A.t3 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t482 VDD.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X437 Comparator_0.Vinm CDAC8_0.switch_7.Z.t97 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X438 a_75898_42964# Q5.t6 Vbias.t428 Vbias.t427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X439 RingCounter_0.D_FlipFlop_7.Q' Nand_Gate_5.A.t7 VDD.t938 VDD.t937 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X440 Vbias.t144 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 a_30647_15797# Vbias.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X441 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout VDD.t595 VDD.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X442 a_75898_46095# Q4.t4 Vbias.t794 Vbias.t793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X443 Vbias.t262 VDD.t1123 a_35335_15797# Vbias.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X444 CDAC8_0.switch_5.Z.t0 a_75898_28676# VDD.t868 VDD.t867 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X445 VDD.t500 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 VDD.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X446 And_Gate_2.Inverter_0.Vin Nand_Gate_6.Vout.t3 VDD.t959 VDD.t958 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X447 a_98245_49858# RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 a_97631_49858# Vbias.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X448 a_112615_15797# Nand_Gate_1.B.t10 a_112001_15797# Vbias.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X449 a_67227_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 Vbias.t489 Vbias.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X450 Comparator_0.Vinm CDAC8_0.switch_6.Z.t50 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X451 VDD.t94 EN.t37 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X452 Comparator_0.Vinm CDAC8_0.switch_9.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X453 VDD.t92 EN.t38 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X454 a_54829_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 Vbias.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X455 VDD.t851 D_FlipFlop_0.D.t12 D_FlipFlop_7.Inverter_0.Vout VDD.t850 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X456 Comparator_0.Vinm CDAC8_0.switch_7.Z.t96 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X457 VDD.t672 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout VDD.t670 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X458 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout VDD.t456 VDD.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X459 Comparator_0.Vinm CDAC8_0.switch_7.Z.t95 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X460 Comparator_0.Vinm CDAC8_0.switch_5.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X461 D_FlipFlop_7.3-input-nand_1.Vout D_FlipFlop_7.Inverter_0.Vout VDD.t605 VDD.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X462 a_106699_52572# VDD.t1124 Vbias.t264 Vbias.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X463 Comparator_0.Vinm CDAC8_0.switch_7.Z.t94 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X464 VDD.t439 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 VDD.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X465 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout Nand_Gate_2.B.t8 VDD.t567 VDD.t566 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X466 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 VDD.t502 VDD.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X467 VDD.t90 EN.t39 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 VDD.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X468 D_FlipFlop_2.3-input-nand_2.C.t2 D_FlipFlop_2.3-input-nand_1.Vout VDD.t558 VDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X469 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 EN.t40 VDD.t88 VDD.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X470 Comparator_0.Vinm CDAC8_0.switch_2.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X471 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout Nand_Gate_0.A.t7 Vbias.t729 Vbias.t728 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X472 Vbias.t484 CLK.t24 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 Vbias.t483 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X473 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t788 VDD.t789 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X474 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 VDD.t20 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X475 VDD.t424 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 VDD.t423 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X476 Comparator_0.Vinm CDAC8_0.switch_6.Z.t49 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X477 VDD.t279 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X478 Vbias.t523 FFCLR.t17 a_128851_17072# Vbias.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X479 a_132311_24200# D_FlipFlop_5.3-input-nand_2.Vout.t4 D_FlipFlop_5.3-input-nand_2.C.t0 Vbias.t417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X480 a_64511_49858# VDD.t1125 Vbias.t266 Vbias.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X481 VDD.t400 D_FlipFlop_5.3-input-nand_2.C.t6 D_FlipFlop_5.3-input-nand_2.Vout.t2 VDD.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X482 a_128851_40571# D_FlipFlop_3.Nand_Gate_1.Vout a_128237_40571# Vbias.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X483 Comparator_0.Vinm CDAC8_0.switch_6.Z.t48 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X484 Comparator_0.Vinm CDAC8_0.switch_7.Z.t93 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X485 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 CLK.t25 VDD.t1085 VDD.t1084 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X486 Vbias.t785 Nand_Gate_6.A.t6 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout Vbias.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X487 CDAC8_0.switch_9.Z.t0 a_75898_42964# VDD.t308 VDD.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X488 VDD.t581 Nand_Gate_6.B.t7 D_FlipFlop_5.3-input-nand_2.Vout.t0 VDD.t580 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X489 Vbias.t525 FFCLR.t18 a_128851_27764# Vbias.t524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X490 Comparator_0.Vinm CDAC8_0.switch_7.Z.t92 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X491 Vbias.t295 D_FlipFlop_1.3-input-nand_2.Vout.t5 a_130209_36157# Vbias.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X492 Comparator_0.Vinm CDAC8_0.switch_9.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X493 Vbias.t85 EN.t41 a_134897_36157# Vbias.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X494 Vbias.t734 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 a_63767_13083# Vbias.t733 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X495 Comparator_0.Vinm CDAC8_0.switch_7.Z.t91 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X496 VDD.t517 And_Gate_6.Vout.t3 D_FlipFlop_3.Inverter_1.Vout VDD.t516 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X497 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout VDD.t975 VDD.t692 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X498 a_75898_25104# Q2.t6 Vbias.t663 Vbias.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X499 VDD.t825 Nand_Gate_0.A.t8 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X500 Vbias.t425 D_FlipFlop_0.3-input-nand_2.Vout.t5 a_130209_46849# Vbias.t424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X501 a_124399_49858# RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 a_123785_49858# Vbias.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X502 VDD.t1083 CLK.t26 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 VDD.t1082 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X503 a_68585_49858# VDD.t1126 Vbias.t268 Vbias.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X504 VDD.t703 a_138318_16817# Vbias.t702 sky130_fd_pr__res_xhigh_po_5p73 l=150
X505 Vbias.t527 FFCLR.t19 a_134897_46849# Vbias.t526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X506 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 VDD.t429 VDD.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X507 a_116995_15797# RingCounter_0.D_FlipFlop_10.Q' Nand_Gate_1.B.t1 Vbias.t518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X508 a_132925_24200# D_FlipFlop_5.3-input-nand_1.Vout a_132311_24200# Vbias.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X509 a_65125_49858# RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 a_64511_49858# Vbias.t799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X510 VDD.t139 D_FlipFlop_2.3-input-nand_2.C.t6 D_FlipFlop_2.3-input-nand_2.Vout.t1 VDD.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X511 Comparator_0.Vinm CDAC8_0.switch_7.Z.t90 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X512 RingCounter_0.D_FlipFlop_2.Q' Nand_Gate_0.A.t9 a_69199_49858# Vbias.t731 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X513 a_75898_18814# Q0.t4 Vbias.t558 Vbias.t557 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X514 And_Gate_4.Vout.t0 And_Gate_4.Inverter_0.Vin VDD.t327 VDD.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X515 VDD.t463 a_138366_35417.t3 D_FlipFlop_0.D.t2 VDD.t462 sky130_fd_pr__pfet_g5v0d10v5 ad=17.4 pd=120.58 as=17.4 ps=120.58 w=60 l=1
X516 a_84489_13083# RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 a_83875_13083# Vbias.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X517 VDD.t826 Nand_Gate_0.A.t10 D_FlipFlop_2.3-input-nand_2.Vout.t3 VDD.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X518 Vbias.t698 D_FlipFlop_4.3-input-nand_2.Vout.t6 a_130209_30478# Vbias.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X519 Comparator_0.Vinm CDAC8_0.switch_7.Z.t89 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X520 Comparator_0.Vinm CDAC8_0.switch_7.Z.t88 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X521 a_123785_49858# VDD.t1127 Vbias.t270 Vbias.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X522 Vbias.t529 FFCLR.t20 a_134897_30478# Vbias.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X523 Comparator_0.Vinm CDAC8_0.switch_9.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X524 VDD.t163 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X525 Comparator_0.Vinm CDAC8_0.switch_5.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X526 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 VDD.t224 VDD.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X527 a_132311_20636# D_FlipFlop_6.3-input-nand_2.Vout.t5 D_FlipFlop_6.3-input-nand_2.C.t0 Vbias.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X528 VDD.t554 D_FlipFlop_6.3-input-nand_2.C.t5 D_FlipFlop_6.3-input-nand_2.Vout.t1 VDD.t553 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X529 a_80239_52572# RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_79625_52572# Vbias.t569 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X530 RingCounter_0.D_FlipFlop_6.Q' Nand_Gate_5.B.t5 a_124399_49858# Vbias.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X531 a_128237_44135# Q4.t5 D_FlipFlop_0.Q' Vbias.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X532 VDD.t520 Nand_Gate_7.B.t7 D_FlipFlop_6.3-input-nand_2.Vout.t3 VDD.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X533 a_83875_13083# Nand_Gate_6.A.t7 RingCounter_0.D_FlipFlop_12.Q' Vbias.t786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X534 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 EN.t42 VDD.t86 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X535 a_88563_13083# RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 a_87949_13083# Vbias.t614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X536 a_108671_49858# VDD.t1128 Vbias.t272 Vbias.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X537 Vbias.t274 VDD.t1129 a_84489_13083# Vbias.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X538 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK.t27 VDD.t1081 VDD.t1004 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X539 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 CLK.t28 VDD.t1080 VDD.t1079 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X540 a_89921_15797# CLK.t29 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 Vbias.t585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X541 Comparator_0.Vinm CDAC8_0.switch_7.Z.t87 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X542 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 a_109285_49858# Vbias.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X543 a_132925_20636# D_FlipFlop_6.3-input-nand_1.Vout a_132311_20636# Vbias.t692 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X544 CDAC8_0.switch_0.Z.t2 a_75898_25104# VDD.t967 VDD.t966 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X545 VDD.t853 D_FlipFlop_0.D.t13 D_FlipFlop_4.Inverter_0.Vout VDD.t852 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X546 VDD.t832 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD.t665 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X547 VDD.t483 FFCLR.t21 D_FlipFlop_5.Q' VDD.t293 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X548 a_134283_39721# And_Gate_4.Vout.t5 D_FlipFlop_2.3-input-nand_0.Vout Vbias.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X549 And_Gate_4.A.t2 Nand_Gate_0.B.t4 VDD.t994 VDD.t993 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X550 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 CLK.t30 VDD.t1078 VDD.t1032 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X551 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_4.Inverter_0.Vout VDD.t265 VDD.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X552 VDD.t344 RingCounter_0.D_FlipFlop_16.Q.t6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 VDD.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X553 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 CLK.t31 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X554 VDD.t877 Nand_Gate_7.A.t8 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout VDD.t876 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X555 Vbias.t276 VDD.t1130 a_88563_13083# Vbias.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X556 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 VDD.t387 VDD.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X557 a_109285_49858# RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 a_108671_49858# Vbias.t722 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X558 a_95529_15797# RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_94915_15797# Vbias.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X559 Comparator_0.Vinm CDAC8_0.switch_7.Z.t86 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X560 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 CLK.t32 Vbias.t587 Vbias.t586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X561 a_134283_23350# And_Gate_0.Vout.t4 D_FlipFlop_6.3-input-nand_0.Vout Vbias.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X562 Comparator_0.Vinm CDAC8_0.switch_9.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X563 Vbias.t83 EN.t43 a_132925_33443# Vbias.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X564 And_Gate_7.Vout.t0 And_Gate_7.Inverter_0.Vin VDD.t835 VDD.t834 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X565 Comparator_0.Vinm CDAC8_0.switch_7.Z.t85 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X566 a_130209_43285# D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout Vbias.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X567 VDD.t1075 CLK.t33 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 VDD.t1074 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X568 VDD.t3 Nand_Gate_1.B.t11 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X569 a_128851_26914# D_FlipFlop_5.Nand_Gate_0.Vout a_128237_26914# Vbias.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X570 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 VDD.t711 VDD.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X571 Comparator_0.Vinm CDAC8_0.switch_7.Z.t84 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X572 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 VDD.t441 VDD.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X573 VDD.t272 And_Gate_1.Vout.t4 D_FlipFlop_7.Inverter_1.Vout VDD.t271 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X574 RingCounter_0.D_FlipFlop_3.Q' VDD.t786 VDD.t787 VDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X575 Comparator_0.Vinm CDAC8_0.switch_9.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X576 VDD.t677 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout VDD.t675 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X577 a_47119_52572# RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 a_46505_52572# Vbias.t704 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X578 Comparator_0.Vinm CDAC8_0.switch_6.Z.t47 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X579 a_50755_13083# Nand_Gate_4.B.t9 RingCounter_0.D_FlipFlop_15.Q' Vbias.t373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X580 Comparator_0.Vinm CDAC8_0.switch_8.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X581 Vbias.t81 EN.t44 a_95529_15797# Vbias.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X582 VDD.t352 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_1.Q' VDD.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X583 a_132311_37007# D_FlipFlop_2.3-input-nand_2.Vout.t5 D_FlipFlop_2.3-input-nand_2.C.t1 Vbias.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X584 a_55443_13083# RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 a_54829_13083# Vbias.t800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X585 Comparator_0.Vinm CDAC8_0.switch_7.Z.t83 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X586 And_Gate_5.Inverter_0.Vin CLK.t34 VDD.t1072 VDD.t1071 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X587 Comparator_0.Vinm CDAC8_0.switch_6.Z.t46 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X588 Comparator_0.Vinm CDAC8_0.switch_6.Z.t45 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X589 D_FlipFlop_1.3-input-nand_2.C.t1 D_FlipFlop_1.3-input-nand_1.Vout VDD.t191 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X590 Comparator_0.Vinm CDAC8_0.switch_6.Z.t44 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X591 VDD.t785 VDD.t784 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X592 a_56801_15797# CLK.t35 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 Vbias.t657 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X593 VDD.t858 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 VDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X594 Nand_Gate_2.A.t0 EN.t45 VDD.t84 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X595 VDD.t895 Q5.t7 CDAC8_0.switch_9.Z.t3 Vbias.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X596 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK.t36 a_41073_49858# Vbias.t658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X597 VDD.t1073 CLK.t37 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 VDD.t1022 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X598 a_110643_13083# RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 a_110029_13083# Vbias.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X599 Comparator_0.Vinm CDAC8_0.switch_7.Z.t82 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X600 VDD.t916 Q4.t6 CDAC8_0.switch_8.Z.t3 Vbias.t795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X601 Nand_Gate_5.Vout.t1 Nand_Gate_5.B.t6 VDD.t911 VDD.t910 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X602 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 CLK.t38 VDD.t1070 VDD.t1028 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X603 VDD.t454 RingCounter_0.D_FlipFlop_12.Q' Nand_Gate_6.A.t2 VDD.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X604 VDD.t1069 CLK.t39 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 VDD.t1068 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X605 a_112001_15797# CLK.t40 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 Vbias.t659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X606 a_132925_37007# D_FlipFlop_2.3-input-nand_1.Vout a_132311_37007# Vbias.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X607 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK.t41 a_74193_52572# Vbias.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X608 Vbias.t278 VDD.t1131 a_55443_13083# Vbias.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X609 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 VDD.t875 VDD.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X610 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 EN.t46 VDD.t82 VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X611 a_62409_15797# RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_61795_15797# Vbias.t521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X612 CDAC8_0.switch_9.Z.t1 a_75898_42964# Vbias.t359 Vbias.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X613 VDD.t1067 CLK.t42 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 VDD.t1020 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X614 VDD.t132 And_Gate_2.Vout.t4 D_FlipFlop_5.3-input-nand_0.Vout VDD.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X615 CDAC8_0.switch_8.Z.t2 a_75898_46095# Vbias.t561 Vbias.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X616 And_Gate_5.Inverter_0.Vin CLK.t43 a_59605_47663# Vbias.t407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X617 RingCounter_0.D_FlipFlop_13.Q' RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 VDD.t323 VDD.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X618 VDD.t80 EN.t47 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 VDD.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X619 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.3-input-nand_2.Vout.t5 VDD.t370 VDD.t369 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X620 Comparator_0.Vinm CDAC8_0.switch_9.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X621 Comparator_0.Vinm CDAC8_0.switch_7.Z.t81 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X622 Vbias.t173 VDD.t1132 a_110643_13083# Vbias.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X623 And_Gate_0.Vout.t1 And_Gate_0.Inverter_0.Vin Vbias.t616 Vbias.t615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X624 Comparator_0.Vinm CDAC8_0.switch_7.Z.t80 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X625 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 VDD.t247 VDD.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X626 VDD.t288 D_FlipFlop_3.3-input-nand_2.Vout.t6 D_FlipFlop_3.3-input-nand_2.C.t1 VDD.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X627 a_66483_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 a_65869_15797# Vbias.t755 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X628 VDD.t485 FFCLR.t22 D_FlipFlop_3.3-input-nand_2.C.t3 VDD.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X629 Comparator_0.Vinm CDAC8_0.switch_6.Z.t43 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X630 VDD.t608 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 VDD.t607 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X631 VDD.t965 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 VDD.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X632 Vbias.t79 EN.t48 a_62409_15797# Vbias.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X633 a_128851_17072# D_FlipFlop_7.Nand_Gate_1.Vout a_128237_17072# Vbias.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X634 Comparator_0.Vinm CDAC8_0.switch_5.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X635 a_134897_24200# D_FlipFlop_5.Inverter_0.Vout a_134283_24200# Vbias.t575 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X636 a_118353_52572# Nand_Gate_5.A.t8 a_117739_52572# Vbias.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X637 VDD.t614 And_Gate_4.Vout.t6 D_FlipFlop_2.3-input-nand_0.Vout VDD.t612 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X638 And_Gate_6.Inverter_0.Vin CLK.t44 VDD.t1066 VDD.t1065 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X639 VDD.t783 VDD.t782 RingCounter_0.D_FlipFlop_13.Q' VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X640 VDD.t521 Nand_Gate_7.B.t8 D_FlipFlop_6.3-input-nand_1.Vout VDD.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X641 a_130209_19786# D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout Vbias.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X642 a_128851_27764# D_FlipFlop_4.Nand_Gate_1.Vout a_128237_27764# Vbias.t620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X643 Comparator_0.Vinm CDAC8_0.switch_7.Z.t79 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X644 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t961 VDD.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X645 Comparator_0.Vinm CDAC8_0.switch_6.Z.t42 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X646 Comparator_0.Vinm CDAC8_0.switch_6.Z.t41 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X647 a_121683_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 a_121069_15797# Vbias.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X648 VDD.t702 a_139496_37417.t3 a_138366_35417.t0 VDD.t701 sky130_fd_pr__pfet_g5v0d10v5 ad=14.5 pd=100.58 as=14.5 ps=100.58 w=50 l=1
X649 Comparator_0.Vinm CDAC8_0.switch_6.Z.t40 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X650 Comparator_0.Vinm CDAC8_0.switch_7.Z.t78 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X651 Vbias.t530 FFCLR.t23 a_132925_44135# Vbias.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X652 a_75898_46095# Q4.t7 VDD.t212 VDD.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X653 VDD.t1064 CLK.t45 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 VDD.t1014 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X654 VDD.t4 Q2.t7 CDAC8_0.switch_0.Z.t0 Vbias.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X655 VDD.t147 And_Gate_0.Vout.t5 D_FlipFlop_6.3-input-nand_0.Vout VDD.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X656 Comparator_0.Vinm CDAC8_0.switch_6.Z.t39 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X657 Comparator_0.Vinm CDAC8_0.switch_7.Z.t77 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X658 VDD.t879 Nand_Gate_7.A.t9 And_Gate_0.B.t0 VDD.t878 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X659 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.3-input-nand_2.Vout.t6 VDD.t949 VDD.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X660 VDD.t419 And_Gate_3.Vout.t4 D_FlipFlop_4.Inverter_1.Vout VDD.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X661 VDD.t627 RingCounter_0.D_FlipFlop_15.Q' Nand_Gate_4.B.t3 VDD.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X662 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK.t46 a_118353_52572# Vbias.t408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X663 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 VDD.t953 VDD.t925 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X664 a_69199_49858# RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 a_68585_49858# Vbias.t541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X665 And_Gate_0.B.t1 Nand_Gate_7.B.t9 a_59977_16975# Vbias.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X666 a_85847_13083# RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 Vbias.t848 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X667 VDD.t983 FFCLR.t24 D_FlipFlop_2.Q' VDD.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X668 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 VDD.t780 VDD.t781 VDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X669 a_106569_15797# RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_105955_15797# Vbias.t291 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X670 VDD.t532 Q0.t5 CDAC8_0.switch_1.Z.t2 Vbias.t559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X671 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 EN.t49 VDD.t78 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X672 a_134283_36157# And_Gate_5.Vout.t3 D_FlipFlop_1.3-input-nand_0.Vout Vbias.t502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X673 D_FlipFlop_3.3-input-nand_2.Vout.t3 D_FlipFlop_3.3-input-nand_0.Vout VDD.t982 VDD.t635 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X674 CDAC8_0.switch_0.Z.t3 a_75898_25104# Vbias.t854 Vbias.t853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X675 RingCounter_0.D_FlipFlop_10.Q' RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 VDD.t898 VDD.t897 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X676 RingCounter_0.D_FlipFlop_8.Q' RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 VDD.t840 VDD.t704 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X677 VDD.t76 EN.t50 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X678 a_100347_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 Vbias.t665 Vbias.t664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X679 a_134283_46849# And_Gate_7.Vout.t3 D_FlipFlop_0.3-input-nand_0.Vout Vbias.t445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X680 D_FlipFlop_0.3-input-nand_2.C.t2 D_FlipFlop_0.3-input-nand_1.Vout VDD.t597 VDD.t596 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X681 VDD.t686 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t685 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X682 a_73579_49858# EN.t51 Vbias.t77 Vbias.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X683 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 a_87205_52572# Vbias.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X684 Vbias.t75 EN.t52 a_68455_13083# Vbias.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X685 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 VDD.t257 VDD.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X686 And_Gate_3.Vout.t1 And_Gate_3.Inverter_0.Vin Vbias.t622 Vbias.t621 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X687 a_134897_20636# D_FlipFlop_6.Inverter_0.Vout a_134283_20636# Vbias.t653 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X688 Comparator_0.Vinm CDAC8_0.switch_7.Z.t76 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X689 VDD.t6 Q2.t8 D_FlipFlop_5.Q' VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X690 CDAC8_0.switch_1.Z.t1 a_75898_18814# Vbias.t342 Vbias.t341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X691 VDD.t286 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_2.B.t1 VDD.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X692 Comparator_0.Vinm CDAC8_0.switch_9.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X693 Vbias.t834 D_FlipFlop_0.D.t14 D_FlipFlop_2.Inverter_0.Vout Vbias.t833 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X694 FFCLR.t1 VDD.t778 VDD.t779 VDD.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X695 a_33363_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_32749_15797# Vbias.t619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X696 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 VDD.t644 VDD.t643 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X697 Vbias.t175 VDD.t1133 a_90535_15797# Vbias.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X698 a_87949_13083# RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 Vbias.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X699 VDD.t220 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 VDD.t219 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X700 Vbias.t73 EN.t53 a_106569_15797# Vbias.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X701 a_134283_30478# And_Gate_3.Vout.t5 D_FlipFlop_4.3-input-nand_0.Vout Vbias.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X702 FFCLR.t3 RingCounter_0.D_FlipFlop_17.Q' VDD.t918 VDD.t390 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X703 VDD.t777 VDD.t776 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X704 Vbias.t71 EN.t54 a_123655_13083# Vbias.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X705 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 VDD.t1106 VDD.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X706 VDD.t443 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout VDD.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X707 Nand_Gate_2.Vout.t2 Nand_Gate_2.B.t9 a_93097_47663# Vbias.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X708 Vbias.t152 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 a_96887_15797# Vbias.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X709 VDD.t775 VDD.t774 RingCounter_0.D_FlipFlop_8.Q' VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X710 Vbias.t879 FFCLR.t25 a_128851_24200# Vbias.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X711 Vbias.t290 D_FlipFlop_1.3-input-nand_2.C.t5 a_130209_33443# Vbias.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X712 VDD.t200 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 RingCounter_0.D_FlipFlop_3.Q' VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X713 VDD.t690 RingCounter_0.D_FlipFlop_8.Q' Nand_Gate_4.A.t2 VDD.t689 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X714 Vbias.t836 D_FlipFlop_0.D.t15 D_FlipFlop_6.Inverter_0.Vout Vbias.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X715 Nand_Gate_2.B.t0 EN.t55 VDD.t74 VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X716 Vbias.t880 FFCLR.t26 a_134897_33443# Vbias.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X717 VDD.t72 EN.t56 D_FlipFlop_1.3-input-nand_0.Vout VDD.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X718 VDD.t923 D_FlipFlop_7.3-input-nand_2.Vout.t6 D_FlipFlop_7.3-input-nand_2.C.t2 VDD.t873 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X719 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 a_78267_49858# Vbias.t867 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X720 Comparator_0.Vinm CDAC8_0.switch_7.Z.t75 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X721 D_FlipFlop_5.Q' D_FlipFlop_5.Nand_Gate_1.Vout VDD.t963 VDD.t587 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X722 VDD.t828 Nand_Gate_0.A.t11 And_Gate_4.A.t1 VDD.t827 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X723 Comparator_0.Vinm CDAC8_0.switch_7.Z.t74 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X724 Comparator_0.Vinm CDAC8_0.switch_7.Z.t73 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X725 Nand_Gate_2.B.t3 RingCounter_0.D_FlipFlop_5.Q' VDD.t869 VDD.t862 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X726 Comparator_0.Vinm CDAC8_0.switch_7.Z.t72 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X727 VDD.t984 FFCLR.t27 D_FlipFlop_0.3-input-nand_0.Vout VDD.t933 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X728 Vbias.t69 EN.t57 a_33363_15797# Vbias.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X729 VDD.t986 FFCLR.t28 D_FlipFlop_7.3-input-nand_2.C.t3 VDD.t985 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X730 RingCounter_0.D_FlipFlop_16.Q' RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 VDD.t634 VDD.t633 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X731 a_96887_15797# RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout Vbias.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X732 VDD.t275 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 VDD.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X733 Comparator_0.Vinm CDAC8_0.switch_6.Z.t38 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X734 Nand_Gate_1.Vout.t0 Nand_Gate_1.B.t12 a_104137_16975# Vbias.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X735 a_52727_13083# RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 Vbias.t745 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X736 And_Gate_1.Inverter_0.Vin And_Gate_1.B.t3 VDD.t340 VDD.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X737 RingCounter_0.D_FlipFlop_3.Q' Nand_Gate_0.B.t5 VDD.t995 VDD.t658 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X738 a_57415_13083# RingCounter_0.D_FlipFlop_15.Inverter_0.Vout a_56801_13083# Vbias.t654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X739 Comparator_0.Vinm CDAC8_0.switch_5.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X740 a_53471_52572# EN.t58 Vbias.t67 Vbias.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X741 Vbias.t668 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 a_30647_13083# Vbias.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X742 VDD.t819 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD.t817 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X743 a_40459_49858# VDD.t1134 Vbias.t177 Vbias.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X744 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 a_54085_52572# Vbias.t544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X745 Vbias.t65 EN.t59 a_35335_13083# Vbias.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X746 VDD.t1063 CLK.t47 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 VDD.t1062 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X747 Comparator_0.Vinm CDAC8_0.switch_6.Z.t37 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X748 And_Gate_4.Inverter_0.Vin CLK.t48 a_81685_47663# Vbias.t409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X749 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 VDD.t772 VDD.t773 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X750 VDD.t771 VDD.t770 RingCounter_0.D_FlipFlop_16.Q' VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X751 Comparator_0.Vinm CDAC8_0.switch_6.Z.t36 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X752 a_112615_13083# RingCounter_0.D_FlipFlop_9.Inverter_0.Vout a_112001_13083# Vbias.t673 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X753 Vbias.t882 FFCLR.t29 a_128851_20636# Vbias.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X754 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout VDD.t565 VDD.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X755 Comparator_0.Vinm CDAC8_0.switch_7.Z.t71 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X756 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 VDD.t450 VDD.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X757 a_54829_13083# RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 Vbias.t555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X758 Comparator_0.Vinm CDAC8_0.switch_9.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X759 a_134897_37007# D_FlipFlop_2.Inverter_0.Vout a_134283_37007# Vbias.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X760 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout Nand_Gate_0.A.t12 VDD.t830 VDD.t829 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X761 a_113359_52572# RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_112745_52572# Vbias.t762 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X762 D_FlipFlop_7.3-input-nand_2.Vout.t0 D_FlipFlop_7.3-input-nand_0.Vout VDD.t669 VDD.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X763 a_54085_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_53471_52572# Vbias.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X764 Comparator_0.Vinm CDAC8_0.switch_7.Z.t70 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X765 a_81685_47663# And_Gate_4.A.t4 Vbias.t8 Vbias.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X766 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 EN.t60 VDD.t70 VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X767 Nand_Gate_3.B.t2 RingCounter_0.D_FlipFlop_1.Q' a_58159_52572# Vbias.t885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X768 VDD.t349 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_6.Q' VDD.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X769 a_41073_49858# RingCounter_0.D_FlipFlop_17.Inverter_0.Vout a_40459_49858# Vbias.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X770 VDD.t940 D_FlipFlop_0.D.t16 D_FlipFlop_5.Inverter_0.Vout VDD.t939 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X771 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 VDD.t245 VDD.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X772 Comparator_0.Vinm CDAC8_0.switch_7.Z.t69 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X773 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 VDD.t645 VDD.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X774 VDD.t769 VDD.t768 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 VDD.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X775 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 a_45147_49858# Vbias.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X776 And_Gate_2.Vout.t0 And_Gate_2.Inverter_0.Vin VDD.t601 VDD.t600 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X777 VDD.t202 Nand_Gate_5.A.t9 Nand_Gate_5.Vout.t0 VDD.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X778 RingCounter_0.D_FlipFlop_2.Q' Nand_Gate_0.A.t13 VDD.t831 VDD.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X779 a_122427_49858# RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 Vbias.t453 Vbias.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X780 VDD.t518 And_Gate_6.Vout.t4 D_FlipFlop_3.3-input-nand_1.Vout VDD.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X781 Comparator_0.Vinm CDAC8_0.switch_7.Z.t68 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X782 a_74193_52572# Nand_Gate_0.A.t14 a_73579_52572# Vbias.t732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X783 a_63767_15797# RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout Vbias.t748 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X784 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_3.3-input-nand_2.C.t5 VDD.t217 VDD.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X785 VDD.t968 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 VDD.t954 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X786 Nand_Gate_5.A.t3 RingCounter_0.D_FlipFlop_7.Q' a_113359_52572# Vbias.t851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X787 a_68455_15797# Nand_Gate_7.B.t10 a_67841_15797# Vbias.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X788 a_132311_39721# D_FlipFlop_2.3-input-nand_2.C.t7 D_FlipFlop_2.3-input-nand_2.Vout.t2 Vbias.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X789 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 a_100347_49858# Vbias.t406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X790 a_130209_40571# D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout Vbias.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X791 VDD.t268 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout VDD.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X792 RingCounter_0.D_FlipFlop_6.Q' Nand_Gate_5.B.t7 VDD.t912 VDD.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X793 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout VDD.t592 VDD.t591 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X794 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 VDD.t364 VDD.t363 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X795 VDD.t942 D_FlipFlop_0.D.t17 D_FlipFlop_2.Inverter_0.Vout VDD.t941 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X796 VDD.t629 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout VDD.t628 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X797 a_107313_49858# RingCounter_0.D_FlipFlop_7.Inverter_0.Vout a_106699_49858# Vbias.t627 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X798 VDD.t552 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t550 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X799 a_123655_15797# Nand_Gate_5.B.t8 a_123041_15797# Vbias.t790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X800 VDD.t68 EN.t61 D_FlipFlop_1.Q' VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X801 Vbias.t516 D_FlipFlop_0.3-input-nand_2.C.t5 a_130209_44135# Vbias.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X802 a_78267_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 Vbias.t319 Vbias.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X803 a_132311_23350# D_FlipFlop_6.3-input-nand_2.C.t6 D_FlipFlop_6.3-input-nand_2.Vout.t0 Vbias.t417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X804 And_Gate_7.Inverter_0.Vin CLK.t49 a_125845_47663# Vbias.t410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X805 And_Gate_5.A.t0 Nand_Gate_3.B.t8 a_48937_47663# Vbias.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X806 Vbias.t228 Nand_Gate_5.A.t10 a_134897_44135# Vbias.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X807 a_65869_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 Vbias.t735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X808 a_116995_13083# Nand_Gate_1.B.t13 RingCounter_0.D_FlipFlop_10.Q' Vbias.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X809 VDD.t688 D_FlipFlop_4.3-input-nand_2.Vout.t7 D_FlipFlop_4.3-input-nand_2.C.t1 VDD.t687 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X810 VDD.t944 D_FlipFlop_0.D.t18 D_FlipFlop_6.Inverter_0.Vout VDD.t943 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X811 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 VDD.t667 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X812 a_90665_49858# VDD.t1135 Vbias.t179 Vbias.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X813 a_132925_39721# D_FlipFlop_2.3-input-nand_0.Vout a_132311_39721# Vbias.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X814 VDD.t237 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 VDD.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X815 VDD.t987 FFCLR.t30 D_FlipFlop_4.3-input-nand_2.C.t3 VDD.t881 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X816 a_117739_52572# VDD.t1136 Vbias.t181 Vbias.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X817 Nand_Gate_6.Vout.t1 Nand_Gate_6.B.t8 VDD.t583 VDD.t582 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X818 VDD.t989 Q6.t6 D_FlipFlop_2.Q' VDD.t885 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X819 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout Nand_Gate_5.A.t11 VDD.t204 VDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X820 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_6.Inverter_0.Vout VDD.t866 VDD.t846 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X821 RingCounter_0.D_FlipFlop_4.Q' Nand_Gate_2.A.t8 a_91279_49858# Vbias.t710 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X822 VDD.t767 VDD.t766 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X823 Vbias.t432 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 a_107927_15797# Vbias.t431 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X824 Vbias.t508 FFCLR.t31 a_128851_37007# Vbias.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X825 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 CLK.t50 a_107313_49858# Vbias.t411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X826 a_121069_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 Vbias.t538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X827 Vbias.t838 D_FlipFlop_0.D.t19 D_FlipFlop_1.Inverter_0.Vout Vbias.t837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X828 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout Nand_Gate_0.B.t6 Vbias.t743 Vbias.t742 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X829 Comparator_0.Vinm CDAC8_0.switch_7.Z.t67 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X830 Vbias.t279 Q4.t8 CDAC8_0.switch_8.Z.t0 VDD.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X831 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 VDD.t495 VDD.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X832 VDD.t765 VDD.t764 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X833 a_132925_23350# D_FlipFlop_6.3-input-nand_0.Vout a_132311_23350# Vbias.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X834 Comparator_0.Vinm CDAC8_0.switch_7.Z.t66 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X835 Vbias.t840 D_FlipFlop_0.D.t20 D_FlipFlop_0.Inverter_0.Vout Vbias.t839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X836 VDD.t540 Nand_Gate_5.Vout.t3 And_Gate_7.Inverter_0.Vin VDD.t539 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X837 VDD.t679 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X838 Comparator_0.Vinm CDAC8_0.switch_7.Z.t65 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X839 a_75551_49858# VDD.t1137 Vbias.t183 Vbias.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X840 Comparator_0.Vinm CDAC8_0.switch_7.Z.t64 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X841 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK.t51 VDD.t1061 VDD.t1060 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X842 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 CLK.t52 VDD.t1059 VDD.t1058 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X843 a_30647_15797# RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout Vbias.t580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X844 VDD.t559 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 VDD.t525 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X845 D_FlipFlop_2.Q' D_FlipFlop_2.Nand_Gate_1.Vout VDD.t328 VDD.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X846 a_35335_15797# Nand_Gate_4.A.t5 a_34721_15797# Vbias.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X847 a_89921_13083# CLK.t53 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 Vbias.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X848 Comparator_0.Vinm CDAC8_0.switch_6.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X849 Vbias.t574 D_FlipFlop_0.D.t21 D_FlipFlop_4.Inverter_0.Vout Vbias.t573 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X850 Vbias.t504 And_Gate_5.Vout.t4 D_FlipFlop_1.Inverter_1.Vout Vbias.t503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X851 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout VDD.t547 VDD.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X852 a_128237_43285# D_FlipFlop_3.Q' Q5.t0 Vbias.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X853 Comparator_0.Vinm CDAC8_0.switch_7.Z.t63 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X854 Comparator_0.Vinm CDAC8_0.switch_8.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X855 Comparator_0.Vinm CDAC8_0.switch_9.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X856 D_FlipFlop_4.3-input-nand_2.Vout.t1 D_FlipFlop_4.3-input-nand_0.Vout VDD.t524 VDD.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X857 Comparator_0.Vinm CDAC8_0.switch_6.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X858 And_Gate_0.Inverter_0.Vin And_Gate_0.B.t3 VDD.t621 VDD.t620 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X859 a_76165_49858# RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 a_75551_49858# Vbias.t414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X860 Comparator_0.Vinm CDAC8_0.switch_6.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X861 a_45147_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 Vbias.t316 Vbias.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X862 VDD.t273 And_Gate_1.Vout.t5 D_FlipFlop_7.3-input-nand_1.Vout VDD.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X863 a_32749_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 Vbias.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X864 D_FlipFlop_7.Nand_Gate_1.Vout D_FlipFlop_7.3-input-nand_2.C.t5 VDD.t376 VDD.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X865 a_95529_13083# RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 a_94915_13083# Vbias.t505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X866 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout VDD.t187 VDD.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X867 VDD.t904 Nand_Gate_6.A.t8 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout VDD.t903 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X868 VDD.t707 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 FFCLR.t0 VDD.t706 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X869 Comparator_0.Vinm CDAC8_0.switch_8.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X870 VDD.t542 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 VDD.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X871 VDD.t260 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout VDD.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X872 a_128851_24200# D_FlipFlop_5.Nand_Gate_1.Vout a_128237_24200# Vbias.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X873 Comparator_0.Vinm CDAC8_0.switch_6.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X874 VDD.t763 VDD.t762 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X875 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout FFCLR.t32 Vbias.t510 Vbias.t509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X876 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_0.D.t22 VDD.t545 VDD.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X877 Comparator_0.Vinm CDAC8_0.switch_6.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X878 a_130209_26914# D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout Vbias.t545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X879 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t760 VDD.t761 VDD.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X880 a_139696_27690# a_138318_16817# Vbias.t471 Vbias.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=1
X881 Comparator_0.Vinm CDAC8_0.switch_7.Z.t62 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X882 VDD.t710 Nand_Gate_2.A.t9 Q5.t3 VDD.t652 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X883 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.D.t23 VDD.t546 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X884 a_42431_49858# EN.t62 Vbias.t63 Vbias.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X885 Vbias.t185 VDD.t1138 a_95529_13083# Vbias.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X886 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK.t54 VDD.t1057 VDD.t1056 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X887 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 CLK.t55 VDD.t1055 VDD.t1054 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X888 VDD.t467 FFCLR.t33 D_FlipFlop_0.Q' VDD.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X889 a_39715_15797# RingCounter_0.D_FlipFlop_8.Q' Nand_Gate_4.A.t1 Vbias.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X890 a_134283_33443# And_Gate_5.Vout.t5 D_FlipFlop_1.3-input-nand_1.Vout Vbias.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X891 a_56801_13083# CLK.t56 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 Vbias.t442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X892 VDD.t668 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X893 Comparator_0.Vinm CDAC8_0.switch_6.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X894 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 CLK.t57 VDD.t1053 VDD.t1052 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X895 VDD.t469 FFCLR.t34 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X896 a_102319_49858# RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 a_101705_49858# Vbias.t520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X897 VDD.t572 Nand_Gate_7.B.t11 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout VDD.t571 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X898 Comparator_0.Vinm CDAC8_0.switch_7.Z.t61 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X899 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 VDD.t531 VDD.t529 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X900 Comparator_0.Vinm CDAC8_0.switch_8.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X901 Comparator_0.Vinm CDAC8_0.switch_9.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X902 And_Gate_1.B.t2 Nand_Gate_4.B.t10 VDD.t330 VDD.t329 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X903 a_43045_49858# RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_42431_49858# Vbias.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X904 a_132311_36157# D_FlipFlop_1.3-input-nand_2.C.t6 D_FlipFlop_1.3-input-nand_2.Vout.t0 Vbias.t343 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X905 RingCounter_0.D_FlipFlop_17.Q' FFCLR.t35 a_47119_49858# Vbias.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X906 a_112001_13083# CLK.t58 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 Vbias.t443 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X907 a_128851_20636# D_FlipFlop_6.Nand_Gate_1.Vout a_128237_20636# Vbias.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X908 Comparator_0.Vinm CDAC8_0.switch_7.Z.t60 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X909 VDD.t872 Nand_Gate_1.A.t6 RingCounter_0.D_FlipFlop_9.Q' VDD.t602 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X910 And_Gate_5.Vout.t0 And_Gate_5.Inverter_0.Vin VDD.t860 VDD.t859 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X911 a_62409_13083# RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 a_61795_13083# Vbias.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X912 a_79625_52572# EN.t63 Vbias.t61 Vbias.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X913 a_132311_46849# D_FlipFlop_0.3-input-nand_2.C.t6 D_FlipFlop_0.3-input-nand_2.Vout.t1 Vbias.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X914 VDD.t914 Nand_Gate_5.B.t9 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout VDD.t913 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X915 VDD.t1051 CLK.t59 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 VDD.t1050 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X916 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 VDD.t509 VDD.t507 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X917 Comparator_0.Vinm CDAC8_0.switch_8.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X918 a_128237_19786# D_FlipFlop_7.Q' Q0.t3 Vbias.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X919 a_58159_52572# RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_57545_52572# Vbias.t606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X920 RingCounter_0.D_FlipFlop_5.Q' Nand_Gate_2.B.t10 a_102319_49858# Vbias.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X921 VDD.t149 And_Gate_0.Vout.t6 D_FlipFlop_6.Inverter_1.Vout VDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X922 VDD.t206 Nand_Gate_5.A.t12 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X923 Comparator_0.Vinm CDAC8_0.switch_7.Z.t59 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X924 Comparator_0.Vinm CDAC8_0.switch_6.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X925 a_132311_30478# D_FlipFlop_4.3-input-nand_2.C.t5 D_FlipFlop_4.3-input-nand_2.Vout.t3 Vbias.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X926 a_132925_36157# D_FlipFlop_1.3-input-nand_0.Vout a_132311_36157# Vbias.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X927 Vbias.t447 And_Gate_7.Vout.t4 D_FlipFlop_0.Inverter_1.Vout Vbias.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X928 VDD.t278 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_2.Q' VDD.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X929 Comparator_0.Vinm CDAC8_0.switch_6.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X930 VDD.t973 Q7.t6 D_FlipFlop_1.Q' VDD.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X931 a_66483_13083# RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 a_65869_13083# Vbias.t860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X932 Vbias.t187 VDD.t1139 a_62409_13083# Vbias.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X933 a_132925_46849# D_FlipFlop_0.3-input-nand_0.Vout a_132311_46849# Vbias.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X934 Nand_Gate_6.B.t1 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD.t538 VDD.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X935 a_67841_15797# CLK.t60 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 Vbias.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X936 a_37897_16975# Nand_Gate_4.A.t6 Vbias.t718 Vbias.t717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X937 a_114805_16975# CLK.t61 Vbias.t812 Vbias.t811 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X938 VDD.t420 And_Gate_3.Vout.t6 D_FlipFlop_4.3-input-nand_1.Vout VDD.t416 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X939 a_67227_49858# RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 Vbias.t491 Vbias.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X940 VDD.t1107 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 VDD.t398 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X941 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_4.3-input-nand_2.C.t6 VDD.t361 VDD.t360 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X942 a_130209_17072# D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout Vbias.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X943 a_134897_39721# D_FlipFlop_0.D.t24 a_134283_39721# Vbias.t365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X944 a_119711_52572# EN.t64 Vbias.t59 Vbias.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X945 VDD.t1049 CLK.t62 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 VDD.t1048 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X946 a_121683_13083# RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 a_121069_13083# Vbias.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X947 a_132925_30478# D_FlipFlop_4.3-input-nand_0.Vout a_132311_30478# Vbias.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X948 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 CLK.t63 VDD.t1047 VDD.t1002 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X949 a_130209_27764# D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout Vbias.t545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X950 VDD.t506 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_0.Vout VDD.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X951 a_106699_49858# EN.t65 Vbias.t57 Vbias.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X952 Comparator_0.Vinm CDAC8_0.switch_6.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X953 VDD.t617 RingCounter_0.D_FlipFlop_11.Q' Nand_Gate_6.B.t3 VDD.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X954 VDD.t697 Nand_Gate_4.A.t7 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout VDD.t696 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X955 VDD.t332 Nand_Gate_4.B.t11 Q0.t1 VDD.t331 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X956 D_FlipFlop_1.Q' D_FlipFlop_1.Nand_Gate_1.Vout VDD.t14 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X957 Comparator_0.Vinm CDAC8_0.switch_6.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X958 a_123041_15797# CLK.t64 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 Vbias.t813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X959 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK.t65 a_85233_52572# Vbias.t814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X960 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 VDD.t957 VDD.t512 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X961 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 EN.t66 VDD.t66 VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X962 VDD.t64 EN.t67 Nand_Gate_6.B.t0 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X963 a_73449_15797# RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_72835_15797# Vbias.t537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X964 a_134897_23350# D_FlipFlop_0.D.t25 a_134283_23350# Vbias.t575 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X965 Comparator_0.Vinm CDAC8_0.switch_7.Z.t58 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X966 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 CLK.t66 Vbias.t816 Vbias.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X967 Comparator_0.Vinm CDAC8_0.switch_7.Z.t57 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X968 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 VDD.t22 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X969 a_46505_52572# VDD.t1140 Vbias.t189 Vbias.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X970 a_106569_13083# RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 a_105955_13083# Vbias.t886 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X971 Comparator_0.Vinm CDAC8_0.switch_9.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X972 Comparator_0.Vinm CDAC8_0.switch_7.Z.t56 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X973 RingCounter_0.D_FlipFlop_12.Q' RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 VDD.t823 VDD.t625 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X974 VDD.t906 Nand_Gate_6.A.t9 Nand_Gate_6.Vout.t2 VDD.t905 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X975 Comparator_0.Vinm CDAC8_0.switch_7.Z.t55 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X976 Vbias.t818 CLK.t67 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 Vbias.t817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X977 a_128851_37007# D_FlipFlop_2.Nand_Gate_1.Vout a_128237_37007# Vbias.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X978 Vbias.t134 Nand_Gate_2.A.t10 a_132925_43285# Vbias.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X979 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 VDD.t544 VDD.t543 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X980 RingCounter_0.D_FlipFlop_1.Q' VDD.t758 VDD.t759 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X981 a_134283_44135# And_Gate_7.Vout.t5 D_FlipFlop_0.3-input-nand_1.Vout Vbias.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X982 CDAC8_0.switch_8.Z.t1 a_75898_46095# VDD.t534 VDD.t533 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X983 VDD.t971 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 VDD.t969 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X984 VDD.t616 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 VDD.t615 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X985 a_101705_52572# EN.t68 Vbias.t55 Vbias.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X986 Vbias.t53 EN.t69 a_73449_15797# Vbias.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X987 a_33363_13083# RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 a_32749_13083# Vbias.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X988 Vbias.t51 EN.t70 a_90535_13083# Vbias.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X989 Comparator_0.Vinm CDAC8_0.switch_7.Z.t54 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X990 Vbias.t191 VDD.t1141 a_106569_13083# Vbias.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X991 RingCounter_0.D_FlipFlop_7.Q' VDD.t756 VDD.t757 VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X992 VDD.t755 VDD.t754 RingCounter_0.D_FlipFlop_12.Q' VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X993 Comparator_0.Vinm CDAC8_0.switch_1.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X994 a_34721_15797# CLK.t68 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout Vbias.t819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X995 Vbias.t890 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 a_96887_13083# Vbias.t889 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X996 And_Gate_2.Inverter_0.Vin Nand_Gate_6.Vout.t4 a_92725_16975# Vbias.t850 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X997 VDD.t290 Nand_Gate_6.B.t9 D_FlipFlop_5.3-input-nand_1.Vout VDD.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X998 VDD.t1046 CLK.t69 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 VDD.t1045 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X999 Vbias.t613 Nand_Gate_0.A.t15 a_128851_39721# Vbias.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1000 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK.t70 VDD.t1044 VDD.t1000 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1001 VDD.t457 RingCounter_0.D_FlipFlop_14.Q' Nand_Gate_7.A.t1 VDD.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1002 a_59605_47663# And_Gate_5.A.t3 Vbias.t738 Vbias.t737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1003 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK.t71 a_52113_52572# Vbias.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1004 Vbias.t193 VDD.t1142 a_33363_13083# Vbias.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1005 Comparator_0.Vinm CDAC8_0.switch_6.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1006 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 VDD.t854 VDD.t476 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1007 a_80239_49858# RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 a_79625_49858# Vbias.t730 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1008 a_96887_13083# RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 Vbias.t741 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1009 VDD.t241 D_FlipFlop_3.Q' Q5.t1 VDD.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1010 Comparator_0.Vinm CDAC8_0.switch_7.Z.t53 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1011 Comparator_0.Vinm CDAC8_0.switch_6.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1012 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 EN.t71 VDD.t62 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1013 VDD.t60 EN.t72 Nand_Gate_7.A.t0 VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1014 a_40329_15797# RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_39715_15797# Vbias.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1015 VDD.t1043 CLK.t72 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 VDD.t1042 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1016 Comparator_0.Vinm CDAC8_0.switch_7.Z.t52 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1017 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 CLK.t73 Vbias.t499 Vbias.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1018 VDD.t215 Q4.t9 D_FlipFlop_0.Q' VDD.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1019 Vbias.t610 Nand_Gate_7.B.t12 a_128851_23350# Vbias.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1020 VDD.t1041 CLK.t74 And_Gate_2.Inverter_0.Vin VDD.t1040 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1021 RingCounter_0.D_FlipFlop_15.Q' RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 VDD.t842 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1022 Comparator_0.Vinm CDAC8_0.switch_7.Z.t51 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1023 a_111387_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 Vbias.t691 Vbias.t690 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1024 Comparator_0.Vinm CDAC8_0.switch_9.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1025 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 VDD.t229 VDD.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1026 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 a_98245_52572# Vbias.t685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1027 VDD.t865 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_5.A.t1 VDD.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1028 Q5.t2 D_FlipFlop_3.Nand_Gate_0.Vout VDD.t253 VDD.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1029 VDD.t333 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 VDD.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1030 Vbias.t49 EN.t73 a_40329_15797# Vbias.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1031 Comparator_0.Vinm CDAC8_0.switch_7.Z.t50 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1032 Comparator_0.Vinm CDAC8_0.switch_7.Z.t49 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1033 VDD.t753 VDD.t752 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1034 Comparator_0.Vinm CDAC8_0.switch_6.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1035 Nand_Gate_3.B.t3 RingCounter_0.D_FlipFlop_1.Q' VDD.t997 VDD.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1036 VDD.t535 Nand_Gate_1.B.t14 Q3.t0 VDD.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1037 D_FlipFlop_0.Q' D_FlipFlop_0.Nand_Gate_1.Vout VDD.t964 VDD.t192 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1038 VDD.t751 VDD.t750 RingCounter_0.D_FlipFlop_15.Q' VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1039 Nand_Gate_1.A.t1 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t233 VDD.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1040 Vbias.t47 EN.t74 a_121683_15797# Vbias.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1041 Comparator_0.Vinm CDAC8_0.switch_7.Z.t48 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1042 VDD.t448 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 RingCounter_0.D_FlipFlop_4.Q' VDD.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1043 VDD.t599 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 VDD.t598 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1044 Vbias.t375 Nand_Gate_4.B.t12 a_132925_19786# Vbias.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1045 a_128237_40571# Q5.t8 D_FlipFlop_3.Q' Vbias.t775 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1046 Nand_Gate_5.A.t2 RingCounter_0.D_FlipFlop_7.Q' VDD.t960 VDD.t937 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1047 VDD.t950 D_FlipFlop_6.3-input-nand_2.Vout.t7 D_FlipFlop_6.3-input-nand_2.C.t3 VDD.t553 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1048 D_FlipFlop_5.3-input-nand_2.Vout.t3 D_FlipFlop_5.3-input-nand_0.Vout VDD.t681 VDD.t593 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1049 And_Gate_4.Vout.t1 And_Gate_4.Inverter_0.Vin Vbias.t371 Vbias.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1050 VDD.t491 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1051 Nand_Gate_0.B.t3 RingCounter_0.D_FlipFlop_3.Q' a_80239_52572# Vbias.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1052 VDD.t695 Nand_Gate_4.A.t8 And_Gate_1.B.t0 VDD.t694 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1053 VDD.t471 FFCLR.t36 D_FlipFlop_6.3-input-nand_2.C.t1 VDD.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1054 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t584 VDD.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1055 a_47119_49858# RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_46505_49858# Vbias.t776 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1056 VDD.t749 VDD.t748 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1057 a_63767_13083# RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 Vbias.t749 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1058 a_134897_36157# D_FlipFlop_0.D.t26 a_134283_36157# Vbias.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1059 VDD.t58 EN.t75 Nand_Gate_1.A.t0 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1060 RingCounter_0.D_FlipFlop_4.Q' Nand_Gate_2.A.t11 VDD.t152 VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1061 a_68455_13083# RingCounter_0.D_FlipFlop_14.Inverter_0.Vout a_67841_13083# Vbias.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1062 Comparator_0.Vinm CDAC8_0.switch_7.Z.t47 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1063 VDD.t388 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1064 VDD.t747 VDD.t746 RingCounter_0.D_FlipFlop_10.Q' VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1065 a_134897_46849# D_FlipFlop_0.D.t27 a_134283_46849# Vbias.t577 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1066 Comparator_0.Vinm CDAC8_0.switch_7.Z.t46 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1067 Vbias.t612 Nand_Gate_7.B.t13 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout Vbias.t611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1068 VDD.t522 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 VDD.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1069 VDD.t263 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1070 a_90535_15797# Nand_Gate_6.B.t10 a_89921_15797# Vbias.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1071 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 a_65125_52572# Vbias.t492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1072 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout Nand_Gate_5.A.t13 Vbias.t825 Vbias.t824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1073 VDD.t1039 CLK.t75 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 VDD.t1038 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1074 D_FlipFlop_2.3-input-nand_2.Vout.t0 D_FlipFlop_2.3-input-nand_0.Vout VDD.t169 VDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1075 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD.t744 VDD.t745 VDD.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1076 a_123655_13083# RingCounter_0.D_FlipFlop_10.Inverter_0.Vout a_123041_13083# Vbias.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1077 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 VDD.t281 VDD.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1078 a_134897_30478# D_FlipFlop_0.D.t28 a_134283_30478# Vbias.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1079 VDD.t928 D_FlipFlop_7.Q' Q0.t2 VDD.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1080 a_84619_52572# VDD.t1143 Vbias.t195 Vbias.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1081 a_65869_13083# RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 Vbias.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1082 Comparator_0.Vinm CDAC8_0.switch_9.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1083 Vbias.t792 Nand_Gate_5.B.t10 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout Vbias.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1084 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout Nand_Gate_0.B.t7 VDD.t838 VDD.t837 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1085 Comparator_0.Vinm CDAC8_0.switch_7.Z.t45 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1086 Comparator_0.Vinm CDAC8_0.switch_7.Z.t44 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1087 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 a_120325_52572# Vbias.t454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1088 Comparator_0.Vinm CDAC8_0.switch_9.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1089 And_Gate_4.A.t0 Nand_Gate_0.B.t8 a_71017_47663# Vbias.t744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1090 Vbias.t294 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 a_74807_15797# Vbias.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1091 Comparator_0.Vinm CDAC8_0.switch_6.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1092 D_FlipFlop_6.3-input-nand_2.Vout.t2 D_FlipFlop_6.3-input-nand_0.Vout VDD.t900 VDD.t712 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1093 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 CLK.t76 a_74193_49858# Vbias.t500 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1094 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 EN.t76 VDD.t56 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1095 Vbias.t321 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 a_107927_13083# Vbias.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1096 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 VDD.t998 VDD.t660 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1097 VDD.t743 VDD.t742 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 VDD.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1098 a_121069_13083# RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 Vbias.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1099 Vbias.t349 D_FlipFlop_3.3-input-nand_2.Vout.t7 a_130209_43285# Vbias.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1100 Comparator_0.Vinm CDAC8_0.switch_6.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1101 Comparator_0.Vinm CDAC8_0.switch_8.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1102 Vbias.t512 FFCLR.t37 a_134897_43285# Vbias.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1103 Q0.t0 D_FlipFlop_7.Nand_Gate_0.Vout VDD.t473 VDD.t472 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1104 a_85233_52572# Nand_Gate_0.B.t9 a_84619_52572# Vbias.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1105 Comparator_0.Vinm CDAC8_0.switch_0.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1106 VDD.t1037 CLK.t77 And_Gate_1.Inverter_0.Vin VDD.t1036 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1107 a_132311_33443# D_FlipFlop_1.3-input-nand_2.Vout.t6 D_FlipFlop_1.3-input-nand_2.C.t2 Vbias.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1108 VDD.t284 D_FlipFlop_1.3-input-nand_2.C.t7 D_FlipFlop_1.3-input-nand_2.Vout.t1 VDD.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1109 Comparator_0.Vinm CDAC8_0.switch_8.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1110 VDD.t1105 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 VDD.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1111 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 a_89307_52572# Vbias.t413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1112 VDD.t573 Nand_Gate_0.A.t16 D_FlipFlop_2.3-input-nand_1.Vout VDD.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1113 a_30647_13083# RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 Vbias.t581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1114 Comparator_0.Vinm CDAC8_0.switch_6.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1115 VDD.t945 FFCLR.t38 D_FlipFlop_1.3-input-nand_2.Vout.t3 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1116 VDD.t175 D_FlipFlop_0.3-input-nand_2.C.t7 D_FlipFlop_0.3-input-nand_2.Vout.t0 VDD.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1117 Comparator_0.Vinm CDAC8_0.switch_6.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1118 a_35335_13083# RingCounter_0.D_FlipFlop_16.Inverter_0.Vout a_34721_13083# Vbias.t873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1119 Vbias.t841 FFCLR.t39 a_128851_36157# Vbias.t507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1120 VDD.t932 Nand_Gate_5.A.t14 D_FlipFlop_0.3-input-nand_2.Vout.t3 VDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1121 a_118353_49858# RingCounter_0.D_FlipFlop_6.Inverter_0.Vout a_117739_49858# Vbias.t439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1122 a_94915_15797# RingCounter_0.D_FlipFlop_11.Q' Nand_Gate_6.B.t2 Vbias.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1123 Vbias.t478 Nand_Gate_4.A.t9 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout Vbias.t477 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1124 VDD.t334 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1125 Vbias.t827 Nand_Gate_5.A.t15 a_128851_46849# Vbias.t826 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1126 Comparator_0.Vinm CDAC8_0.switch_7.Z.t43 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1127 a_99603_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 a_98989_15797# Vbias.t849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1128 VDD.t1035 CLK.t78 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 VDD.t1034 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1129 a_132925_33443# D_FlipFlop_1.3-input-nand_1.Vout a_132311_33443# Vbias.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1130 a_128237_26914# D_FlipFlop_5.Q' Q2.t1 Vbias.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1131 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 VDD.t277 VDD.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1132 a_51499_52572# VDD.t1144 Vbias.t197 Vbias.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1133 a_32749_13083# RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 Vbias.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1134 Vbias.t562 Nand_Gate_1.B.t15 a_128851_30478# Vbias.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1135 VDD.t820 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 VDD.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1136 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout FFCLR.t40 VDD.t947 VDD.t946 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1137 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 Nand_Gate_7.B.t14 VDD.t354 VDD.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1138 Vbias.t357 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 a_118967_15797# Vbias.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1139 Vbias.t572 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 a_41687_15797# Vbias.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1140 VDD.t741 VDD.t740 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1141 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 CLK.t79 a_118353_49858# Vbias.t861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1142 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 EN.t77 VDD.t54 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1143 VDD.t302 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 VDD.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1144 Vbias.t45 EN.t78 a_99603_15797# Vbias.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1145 Comparator_0.Vinm CDAC8_0.switch_7.Z.t42 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1146 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 VDD.t560 VDD.t527 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1147 VDD.t739 VDD.t738 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1148 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_5.Inverter_0.Vout VDD.t917 VDD.t843 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1149 And_Gate_0.Vout.t0 And_Gate_0.Inverter_0.Vin VDD.t577 VDD.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1150 a_128851_39721# D_FlipFlop_2.Nand_Gate_0.Vout a_128237_39721# Vbias.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1151 a_130209_24200# D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout Vbias.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1152 VDD.t671 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout VDD.t670 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1153 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK.t80 VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1154 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 Nand_Gate_5.B.t11 VDD.t902 VDD.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1155 a_100347_49858# RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 Vbias.t687 Vbias.t686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1156 Comparator_0.Vinm CDAC8_0.switch_6.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1157 a_52113_52572# FFCLR.t41 a_51499_52572# Vbias.t842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1158 a_41687_15797# RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout Vbias.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1159 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 a_87205_49858# Vbias.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1160 VDD.t622 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 VDD.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1161 a_75898_21528# Q1.t5 Vbias.t141 Vbias.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1162 VDD.t421 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 VDD.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1163 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 a_56187_52572# Vbias.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1164 a_46375_15797# Nand_Gate_4.B.t13 a_45761_15797# Vbias.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1165 Comparator_0.Vinm CDAC8_0.switch_7.Z.t41 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1166 Comparator_0.Vinm CDAC8_0.switch_8.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1167 VDD.t737 VDD.t736 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 VDD.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1168 VDD.t624 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 VDD.t377 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1169 a_39715_13083# Nand_Gate_4.A.t10 RingCounter_0.D_FlipFlop_8.Q' Vbias.t582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1170 VDD.t901 D_FlipFlop_4.Q' Q3.t2 VDD.t403 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1171 VDD.t52 EN.t79 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1172 a_128851_23350# D_FlipFlop_6.Nand_Gate_0.Vout a_128237_23350# Vbias.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1173 Comparator_0.Vinm CDAC8_0.switch_6.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1174 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout VDD.t632 VDD.t318 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1175 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 VDD.t857 VDD.t855 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1176 Vbias.t843 FFCLR.t42 a_132925_40571# Vbias.t726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1177 Comparator_0.Vinm CDAC8_0.switch_6.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1178 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 VDD.t639 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1179 Comparator_0.Vinm CDAC8_0.switch_7.Z.t40 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1180 Vbias.t597 D_FlipFlop_7.3-input-nand_2.Vout.t7 a_130209_19786# Vbias.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1181 VDD.t929 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 VDD.t423 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1182 a_61795_15797# RingCounter_0.D_FlipFlop_14.Q' Nand_Gate_7.A.t2 Vbias.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1183 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout RingCounter_0.D_FlipFlop_16.Q.t7 VDD.t346 VDD.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1184 VDD.t824 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 VDD.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1185 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 a_111387_52572# Vbias.t546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1186 a_101575_15797# Nand_Gate_1.A.t7 a_100961_15797# Vbias.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1187 Nand_Gate_0.B.t0 EN.t80 VDD.t50 VDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1188 a_56187_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 Vbias.t535 Vbias.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1189 Vbias.t844 FFCLR.t43 a_134897_19786# Vbias.t550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1190 VDD.t676 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout VDD.t675 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1191 And_Gate_6.Inverter_0.Vin CLK.t81 a_103765_47663# Vbias.t862 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1192 VDD.t356 Nand_Gate_7.B.t15 RingCounter_0.D_FlipFlop_13.Q' VDD.t355 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1193 VDD.t150 And_Gate_0.Vout.t7 D_FlipFlop_6.3-input-nand_1.Vout VDD.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1194 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout VDD.t647 VDD.t646 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1195 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 VDD.t657 VDD.t655 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1196 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 VDD.t427 VDD.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1197 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_6.3-input-nand_2.C.t7 VDD.t556 VDD.t555 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1198 Vbias.t864 CLK.t82 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 Vbias.t863 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1199 Comparator_0.Vinm CDAC8_0.switch_0.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1200 VDD.t292 Nand_Gate_6.B.t11 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout VDD.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1201 VDD.t570 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout Nand_Gate_3.B.t1 VDD.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1202 Q3.t3 D_FlipFlop_4.Nand_Gate_0.Vout VDD.t996 VDD.t887 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1203 And_Gate_0.B.t2 Nand_Gate_7.B.t16 VDD.t358 VDD.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1204 a_132311_44135# D_FlipFlop_0.3-input-nand_2.Vout.t6 D_FlipFlop_0.3-input-nand_2.C.t0 Vbias.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1205 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout Nand_Gate_4.A.t11 VDD.t693 VDD.t692 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1206 a_130209_20636# D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout Vbias.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1207 VDD.t891 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout VDD.t890 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1208 a_139496_37417.t2 Comparator_0.Vinm a_139696_27690# Vbias.t893 sky130_fd_pr__nfet_g5v0d10v5 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=1
X1209 D_FlipFlop_3.3-input-nand_2.C.t0 D_FlipFlop_3.3-input-nand_1.Vout VDD.t636 VDD.t635 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1210 VDD.t735 VDD.t734 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1211 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 EN.t81 VDD.t48 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1212 VDD.t173 Nand_Gate_0.B.t10 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1213 a_128237_17072# Q0.t6 D_FlipFlop_7.Q' Vbias.t694 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1214 Comparator_0.Vinm CDAC8_0.switch_7.Z.t39 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1215 Vbias.t19 EN.t82 a_66483_15797# Vbias.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1216 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 CLK.t83 VDD.t1031 VDD.t1030 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1217 Comparator_0.Vinm CDAC8_0.switch_9.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1218 VDD.t822 Nand_Gate_2.Vout.t4 And_Gate_6.Inverter_0.Vin VDD.t821 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1219 Comparator_0.Vinm CDAC8_0.switch_7.Z.t38 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1220 Comparator_0.Vinm CDAC8_0.switch_7.Z.t37 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1221 a_128237_27764# Q3.t8 D_FlipFlop_4.Q' Vbias.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1222 a_53471_49858# VDD.t1145 Vbias.t199 Vbias.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1223 Comparator_0.Vinm CDAC8_0.switch_9.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1224 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK.t84 VDD.t1029 VDD.t1028 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1225 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 a_54085_49858# Vbias.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1226 VDD.t683 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1227 a_132925_44135# D_FlipFlop_0.3-input-nand_1.Vout a_132311_44135# Vbias.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1228 a_86591_52572# EN.t83 Vbias.t23 Vbias.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1229 a_67841_13083# CLK.t85 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 Vbias.t865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1230 Nand_Gate_2.Vout.t1 Nand_Gate_2.B.t11 VDD.t569 VDD.t568 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1231 a_113359_49858# RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 a_112745_49858# Vbias.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1232 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 VDD.t732 VDD.t733 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1233 VDD.t948 FFCLR.t44 D_FlipFlop_1.3-input-nand_1.Vout VDD.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1234 a_105955_15797# RingCounter_0.D_FlipFlop_9.Q' Nand_Gate_1.A.t2 Vbias.t630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1235 a_54085_49858# RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 a_53471_49858# Vbias.t355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1236 RingCounter_0.D_FlipFlop_1.Q' Nand_Gate_3.B.t9 a_58159_49858# Vbias.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1237 a_123041_13083# CLK.t86 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 Vbias.t866 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1238 VDD.t536 Nand_Gate_1.B.t16 RingCounter_0.D_FlipFlop_10.Q' VDD.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1239 a_73449_13083# RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 a_72835_13083# Vbias.t706 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1240 a_87205_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_86591_52572# Vbias.t642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1241 VDD.t141 And_Gate_5.Vout.t6 D_FlipFlop_1.3-input-nand_0.Vout VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1242 VDD.t294 Nand_Gate_6.B.t12 Q2.t0 VDD.t293 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1243 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.3-input-nand_2.Vout.t7 VDD.t503 VDD.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1244 Comparator_0.Vinm CDAC8_0.switch_2.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1245 a_74193_49858# RingCounter_0.D_FlipFlop_3.Inverter_0.Vout a_73579_49858# Vbias.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1246 Comparator_0.Vinm CDAC8_0.switch_7.Z.t36 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1247 RingCounter_0.D_FlipFlop_7.Q' Nand_Gate_5.A.t16 a_113359_49858# Vbias.t828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1248 VDD.t413 And_Gate_7.Vout.t6 D_FlipFlop_0.3-input-nand_0.Vout VDD.t411 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1249 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.3-input-nand_2.Vout.t7 VDD.t674 VDD.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1250 VDD.t956 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 VDD.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1251 a_93097_47663# Nand_Gate_2.A.t12 Vbias.t136 Vbias.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1252 a_130209_37007# D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout Vbias.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1253 VDD.t134 And_Gate_2.Vout.t5 D_FlipFlop_5.Inverter_1.Vout VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1254 Vbias.t352 Nand_Gate_6.B.t13 a_132925_26914# Vbias.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1255 And_Gate_1.Inverter_0.Vin And_Gate_1.B.t4 a_48565_16975# Vbias.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1256 And_Gate_4.Inverter_0.Vin CLK.t87 VDD.t1027 VDD.t1026 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1257 Vbias.t201 VDD.t1146 a_73449_13083# Vbias.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1258 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 CLK.t88 VDD.t1025 VDD.t1024 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1259 a_134897_33443# D_FlipFlop_1.Inverter_0.Vout a_134283_33443# Vbias.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1260 a_78881_15797# CLK.t89 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 Vbias.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1261 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_2.Inverter_0.Vout VDD.t586 VDD.t585 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1262 a_78267_49858# RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 Vbias.t751 Vbias.t750 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1263 VDD.t575 Nand_Gate_0.A.t17 Q6.t1 VDD.t574 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1264 Comparator_0.Vinm CDAC8_0.switch_7.Z.t35 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1265 a_34721_13083# CLK.t90 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 Vbias.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1266 Vbias.t203 VDD.t1147 a_79495_15797# Vbias.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1267 Comparator_0.Vinm CDAC8_0.switch_7.Z.t34 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1268 D_FlipFlop_7.3-input-nand_2.C.t0 D_FlipFlop_7.3-input-nand_1.Vout VDD.t310 VDD.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1269 a_128851_36157# D_FlipFlop_1.Nand_Gate_0.Vout a_128237_36157# Vbias.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1270 Comparator_0.Vinm CDAC8_0.switch_7.Z.t33 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1271 Comparator_0.Vinm CDAC8_0.switch_7.Z.t32 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1272 VDD.t348 RingCounter_0.D_FlipFlop_16.Q.t8 RingCounter_0.D_FlipFlop_16.Q' VDD.t347 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1273 a_134283_43285# And_Gate_6.Vout.t5 D_FlipFlop_3.3-input-nand_0.Vout Vbias.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1274 Comparator_0.Vinm CDAC8_0.switch_9.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1275 a_117739_49858# EN.t84 Vbias.t43 Vbias.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1276 Comparator_0.Vinm CDAC8_0.switch_7.Z.t31 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1277 a_128851_46849# D_FlipFlop_0.Nand_Gate_0.Vout a_128237_46849# Vbias.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1278 a_104137_16975# Nand_Gate_1.A.t8 Vbias.t768 Vbias.t767 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1279 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK.t91 a_96273_52572# Vbias.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1280 a_98989_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 Vbias.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1281 VDD.t359 Nand_Gate_7.B.t17 Q1.t1 VDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1282 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 CLK.t92 Vbias.t396 Vbias.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1283 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 VDD.t664 VDD.t643 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1284 a_57545_52572# EN.t85 Vbias.t41 Vbias.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1285 a_40329_13083# RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 a_39715_13083# Vbias.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1286 Comparator_0.Vinm CDAC8_0.switch_5.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1287 Comparator_0.Vinm CDAC8_0.switch_6.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1288 a_128851_30478# D_FlipFlop_4.Nand_Gate_0.Vout a_128237_30478# Vbias.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1289 Comparator_0.Vinm CDAC8_0.switch_7.Z.t30 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1290 VDD.t1023 CLK.t93 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 VDD.t1022 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1291 Vbias.t398 CLK.t94 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 Vbias.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1292 And_Gate_2.Vout.t1 And_Gate_2.Inverter_0.Vin Vbias.t629 Vbias.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1293 RingCounter_0.D_FlipFlop_2.Q' VDD.t730 VDD.t731 VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1294 VDD.t267 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout VDD.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1295 VDD.t924 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 VDD.t548 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1296 VDD.t541 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout Nand_Gate_0.B.t1 VDD.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1297 Comparator_0.Vinm CDAC8_0.switch_7.Z.t29 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1298 Vbias.t281 D_FlipFlop_3.3-input-nand_2.C.t6 a_130209_40571# Vbias.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1299 VDD.t839 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 VDD.t295 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1300 a_112745_52572# EN.t86 Vbias.t39 Vbias.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1301 Vbias.t138 Nand_Gate_2.A.t13 a_134897_40571# Vbias.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1302 VDD.t649 FFCLR.t45 D_FlipFlop_3.3-input-nand_0.Vout VDD.t648 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1303 VDD.t1021 CLK.t95 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 VDD.t1020 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1304 a_75898_35820# Q7.t7 Vbias.t869 Vbias.t868 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1305 Vbias.t205 VDD.t1148 a_40329_13083# Vbias.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1306 RingCounter_0.D_FlipFlop_6.Q' VDD.t728 VDD.t729 VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1307 VDD.t934 Nand_Gate_5.A.t17 D_FlipFlop_0.3-input-nand_1.Vout VDD.t933 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1308 Nand_Gate_7.B.t1 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD.t494 VDD.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1309 VDD.t159 Q1.t6 CDAC8_0.switch_2.Z.t0 Vbias.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1310 a_45761_15797# CLK.t96 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 Vbias.t399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1311 a_45147_49858# RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 Vbias.t846 Vbias.t845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1312 Vbias.t37 EN.t87 a_128851_33443# Vbias.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1313 Vbias.t207 VDD.t1149 a_121683_13083# Vbias.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1314 Vbias.t209 VDD.t1150 a_46375_15797# Vbias.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1315 Nand_Gate_0.B.t2 RingCounter_0.D_FlipFlop_3.Q' VDD.t659 VDD.t658 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1316 VDD.t1019 CLK.t97 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 VDD.t1018 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1317 Vbias.t675 FFCLR.t46 a_132925_17072# Vbias.t674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1318 Comparator_0.Vinm CDAC8_0.switch_7.Z.t28 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1319 Comparator_0.Vinm CDAC8_0.switch_7.Z.t27 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1320 VDD.t609 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD.t607 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1321 Comparator_0.Vinm CDAC8_0.switch_7.Z.t26 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1322 Comparator_0.Vinm CDAC8_0.switch_9.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1323 VDD.t46 EN.t88 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1324 CDAC8_0.switch_2.Z.t3 a_75898_21528# Vbias.t595 Vbias.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1325 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 VDD.t726 VDD.t727 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1326 a_100961_15797# CLK.t98 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 Vbias.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1327 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK.t99 a_63153_52572# Vbias.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1328 Vbias.t676 FFCLR.t47 a_132925_27764# Vbias.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1329 Nand_Gate_6.Vout.t0 Nand_Gate_6.B.t14 a_82057_16975# Vbias.t820 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1330 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 EN.t89 VDD.t44 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1331 a_51369_15797# RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_50755_15797# Vbias.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1332 VDD.t42 EN.t90 Nand_Gate_7.B.t0 VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1333 Vbias.t211 VDD.t1151 a_101575_15797# Vbias.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1334 VDD.t1017 CLK.t100 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 VDD.t1016 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1335 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 CLK.t101 Vbias.t382 Vbias.t381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1336 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 VDD.t304 VDD.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1337 Comparator_0.Vinm CDAC8_0.switch_6.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1338 RingCounter_0.D_FlipFlop_14.Q' RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 VDD.t475 VDD.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1339 Comparator_0.Vinm CDAC8_0.switch_6.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1340 a_125845_47663# Nand_Gate_5.Vout.t4 Vbias.t701 Vbias.t700 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1341 a_48937_47663# FFCLR.t48 Vbias.t678 Vbias.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1342 Comparator_0.Vinm CDAC8_0.switch_5.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1343 VDD.t1015 CLK.t102 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD.t1014 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1344 Vbias.t384 CLK.t103 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 Vbias.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1345 a_134283_19786# And_Gate_1.Vout.t6 D_FlipFlop_7.3-input-nand_0.Vout Vbias.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1346 a_134897_44135# D_FlipFlop_0.Inverter_0.Vout a_134283_44135# Vbias.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1347 Comparator_0.Vinm CDAC8_0.switch_7.Z.t25 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1348 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD.t724 VDD.t725 VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1349 a_90535_13083# RingCounter_0.D_FlipFlop_12.Inverter_0.Vout a_89921_13083# Vbias.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1350 Comparator_0.Vinm CDAC8_0.switch_8.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1351 VDD.t249 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_5.B.t1 VDD.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1352 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 CLK.t104 Vbias.t386 Vbias.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1353 D_FlipFlop_4.3-input-nand_2.C.t2 D_FlipFlop_4.3-input-nand_1.Vout VDD.t691 VDD.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1354 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 VDD.t422 VDD.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1355 Vbias.t35 EN.t91 a_51369_15797# Vbias.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1356 Vbias.t822 Nand_Gate_6.B.t15 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout Vbias.t821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1357 VDD.t723 VDD.t722 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1358 Nand_Gate_0.A.t3 RingCounter_0.D_FlipFlop_2.Q' VDD.t312 VDD.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1359 a_107927_15797# RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout Vbias.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1360 a_75898_21528# Q1.t7 VDD.t161 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1361 Nand_Gate_1.B.t3 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD.t927 VDD.t897 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1362 Nand_Gate_4.A.t3 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD.t705 VDD.t704 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1363 Vbias.t672 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 a_74807_13083# Vbias.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1364 VDD.t179 And_Gate_4.Vout.t7 D_FlipFlop_2.Inverter_1.Vout VDD.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1365 VDD.t259 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout VDD.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1366 Comparator_0.Vinm CDAC8_0.switch_7.Z.t24 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1367 VDD.t425 D_FlipFlop_5.Q' Q2.t2 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1368 VDD.t977 D_FlipFlop_0.D.t29 D_FlipFlop_1.Inverter_0.Vout VDD.t976 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1369 VDD.t154 Nand_Gate_2.A.t14 Nand_Gate_2.Vout.t0 VDD.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1370 Comparator_0.Vinm CDAC8_0.switch_6.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1371 a_79625_49858# VDD.t1152 Vbias.t213 Vbias.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1372 Nand_Gate_5.B.t2 RingCounter_0.D_FlipFlop_6.Q' VDD.t493 VDD.t492 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1373 Comparator_0.Vinm CDAC8_0.switch_7.Z.t23 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1374 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 VDD.t833 VDD.t363 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1375 Comparator_0.Vinm CDAC8_0.switch_6.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1376 VDD.t651 FFCLR.t49 D_FlipFlop_7.3-input-nand_0.Vout VDD.t650 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1377 D_FlipFlop_1.3-input-nand_1.Vout D_FlipFlop_1.Inverter_0.Vout VDD.t227 VDD.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1378 VDD.t979 D_FlipFlop_0.D.t30 D_FlipFlop_0.Inverter_0.Vout VDD.t978 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1379 Comparator_0.Vinm CDAC8_0.switch_7.Z.t22 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1380 VDD.t40 EN.t92 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1381 a_110029_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 Vbias.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1382 VDD.t372 D_FlipFlop_5.3-input-nand_2.Vout.t6 D_FlipFlop_5.3-input-nand_2.C.t1 VDD.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1383 a_58159_49858# RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 a_57545_49858# Vbias.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1384 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 VDD.t374 VDD.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1385 VDD.t653 FFCLR.t50 D_FlipFlop_3.Q' VDD.t652 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1386 Vbias.t125 D_FlipFlop_5.3-input-nand_2.Vout.t7 a_130209_26914# Vbias.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1387 Comparator_0.Vinm CDAC8_0.switch_7.Z.t21 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1388 VDD.t38 EN.t93 Nand_Gate_4.A.t0 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1389 Comparator_0.Vinm CDAC8_0.switch_9.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1390 VDD.t654 FFCLR.t51 D_FlipFlop_5.3-input-nand_2.C.t3 VDD.t580 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1391 Vbias.t459 FFCLR.t52 a_134897_26914# Vbias.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1392 And_Gate_1.Vout.t0 And_Gate_1.Inverter_0.Vin VDD.t325 VDD.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1393 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 VDD.t12 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1394 VDD.t1013 CLK.t105 And_Gate_0.Inverter_0.Vin VDD.t1012 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1395 Q2.t3 D_FlipFlop_5.Nand_Gate_0.Vout VDD.t588 VDD.t587 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1396 Comparator_0.Vinm CDAC8_0.switch_6.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1397 VDD.t886 D_FlipFlop_2.Q' Q6.t2 VDD.t885 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1398 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 a_76165_52572# Vbias.t752 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1399 Vbias.t589 CLK.t106 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 Vbias.t588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1400 Vbias.t591 CLK.t107 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 Vbias.t590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1401 VDD.t1011 CLK.t108 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 VDD.t1010 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1402 a_94915_13083# Nand_Gate_6.B.t16 RingCounter_0.D_FlipFlop_11.Q' Vbias.t823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1403 RingCounter_0.D_FlipFlop_16.Q.t3 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD.t909 VDD.t633 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1404 Vbias.t461 FFCLR.t53 a_128851_44135# Vbias.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1405 a_99603_13083# RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 a_98989_13083# Vbias.t547 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1406 Comparator_0.Vinm CDAC8_0.switch_7.Z.t20 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1407 a_75898_39392# Q6.t7 VDD.t991 VDD.t990 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1408 Vbias.t876 D_FlipFlop_0.D.t31 D_FlipFlop_3.Inverter_0.Vout Vbias.t875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1409 Comparator_0.Vinm CDAC8_0.switch_5.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1410 a_119711_49858# VDD.t1153 Vbias.t215 Vbias.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1411 a_95659_52572# VDD.t1154 Vbias.t217 Vbias.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1412 a_128237_24200# Q2.t9 D_FlipFlop_5.Q' Vbias.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1413 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout Nand_Gate_2.A.t15 VDD.t156 VDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1414 Comparator_0.Vinm CDAC8_0.switch_7.Z.t19 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1415 VDD.t915 D_FlipFlop_6.Q' Q1.t2 VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1416 a_75898_18814# Q0.t7 VDD.t673 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1417 Vbias.t683 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 a_85847_15797# Vbias.t682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1418 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 CLK.t109 a_85233_49858# Vbias.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1419 Q6.t0 D_FlipFlop_2.Nand_Gate_0.Vout VDD.t314 VDD.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1420 Vbias.t808 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 a_41687_13083# Vbias.t807 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1421 Vbias.t803 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 a_118967_13083# Vbias.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1422 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 VDD.t430 VDD.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1423 VDD.t36 EN.t94 RingCounter_0.D_FlipFlop_16.Q.t0 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1424 a_46505_49858# EN.t95 Vbias.t33 Vbias.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1425 Vbias.t219 VDD.t1155 a_99603_13083# Vbias.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1426 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 Nand_Gate_6.B.t17 VDD.t931 VDD.t564 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1427 Vbias.t872 And_Gate_6.Vout.t6 D_FlipFlop_3.Inverter_1.Vout Vbias.t871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1428 Comparator_0.Vinm CDAC8_0.switch_7.Z.t18 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1429 And_Gate_5.Vout.t1 And_Gate_5.Inverter_0.Vin Vbias.t761 Vbias.t760 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1430 Comparator_0.Vinm CDAC8_0.switch_6.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1431 And_Gate_3.Inverter_0.Vin Nand_Gate_1.Vout.t4 VDD.t410 VDD.t409 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1432 a_96273_52572# Nand_Gate_2.A.t16 a_95659_52572# Vbias.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1433 Comparator_0.Vinm CDAC8_0.switch_7.Z.t17 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1434 Comparator_0.Vinm CDAC8_0.switch_6.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1435 Q1.t0 D_FlipFlop_6.Nand_Gate_0.Vout VDD.t663 VDD.t662 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1436 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout RingCounter_0.D_FlipFlop_16.Q.t9 Vbias.t689 Vbias.t688 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1437 a_41687_13083# RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 Vbias.t391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1438 a_130209_39721# D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout Vbias.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1439 a_46375_13083# RingCounter_0.D_FlipFlop_8.Inverter_0.Vout a_45761_13083# Vbias.t578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1440 a_101705_49858# VDD.t1156 Vbias.t221 Vbias.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1441 Comparator_0.Vinm CDAC8_0.switch_7.Z.t16 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1442 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 VDD.t235 VDD.t234 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1443 VDD.t1009 CLK.t110 And_Gate_3.Inverter_0.Vin VDD.t1008 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1444 Comparator_0.Vinm CDAC8_0.switch_9.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1445 Vbias.t157 Nand_Gate_4.B.t14 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout Vbias.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1446 a_128237_20636# Q1.t8 D_FlipFlop_6.Q' Vbias.t363 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1447 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 a_43045_52572# Vbias.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1448 VDD.t1007 CLK.t111 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 VDD.t1006 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1449 Comparator_0.Vinm CDAC8_0.switch_6.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1450 Vbias.t419 D_FlipFlop_7.3-input-nand_2.C.t6 a_130209_17072# Vbias.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1451 a_61795_13083# Nand_Gate_7.A.t10 RingCounter_0.D_FlipFlop_14.Q' Vbias.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1452 a_130209_23350# D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout Vbias.t693 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1453 a_101575_13083# RingCounter_0.D_FlipFlop_11.Inverter_0.Vout a_100961_13083# Vbias.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1454 VDD.t505 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout VDD.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1455 a_120325_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_119711_52572# Vbias.t474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1456 Vbias.t159 Nand_Gate_4.B.t15 a_134897_17072# Vbias.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1457 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_0.D.t32 VDD.t980 VDD.t316 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1458 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 VDD.t816 VDD.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1459 Comparator_0.Vinm CDAC8_0.switch_7.Z.t15 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1460 VDD.t431 FFCLR.t54 D_FlipFlop_7.Q' VDD.t331 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1461 Vbias.t412 D_FlipFlop_4.3-input-nand_2.C.t7 a_130209_27764# Vbias.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1462 a_62539_52572# VDD.t1157 Vbias.t223 Vbias.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1463 VDD.t974 Q7.t8 CDAC8_0.switch_7.Z.t3 Vbias.t870 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1464 Vbias.t773 Nand_Gate_1.A.t9 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout Vbias.t772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1465 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout Nand_Gate_3.B.t10 VDD.t210 VDD.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1466 Vbias.t563 Nand_Gate_1.B.t17 a_134897_27764# Vbias.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1467 VDD.t433 FFCLR.t55 D_FlipFlop_4.3-input-nand_0.Vout VDD.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1468 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_0.Inverter_0.Vout VDD.t336 VDD.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1469 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 Nand_Gate_6.A.t10 VDD.t907 VDD.t591 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1470 Vbias.t565 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 a_52727_15797# Vbias.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1471 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 CLK.t112 a_52113_49858# Vbias.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1472 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 EN.t96 VDD.t34 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1473 a_128851_33443# D_FlipFlop_1.Nand_Gate_1.Vout a_128237_33443# Vbias.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1474 VDD.t171 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 VDD.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1475 a_134283_40571# And_Gate_6.Vout.t7 D_FlipFlop_3.3-input-nand_1.Vout Vbias.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1476 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 VDD.t623 VDD.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1477 a_89307_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 Vbias.t405 Vbias.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1478 Vbias.t469 a_138318_16817# D_FlipFlop_0.D.t1 Vbias.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X1479 CDAC8_0.switch_7.Z.t1 a_75898_35820# Vbias.t423 Vbias.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1480 Vbias.t225 VDD.t1158 a_66483_13083# Vbias.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1481 Vbias.t878 D_FlipFlop_0.D.t33 D_FlipFlop_7.Inverter_0.Vout Vbias.t877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1482 a_111387_49858# RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 Vbias.t641 Vbias.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1483 a_63153_52572# Nand_Gate_3.B.t11 a_62539_52572# Vbias.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1484 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 a_98245_49858# Vbias.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1485 VDD.t497 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 VDD.t236 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1486 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 a_67227_52572# Vbias.t754 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1487 VDD.t143 And_Gate_5.Vout.t7 D_FlipFlop_1.Inverter_1.Vout VDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1488 Comparator_0.Vinm CDAC8_0.switch_7.Z.t14 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1489 And_Gate_6.Vout.t0 And_Gate_6.Inverter_0.Vin VDD.t638 VDD.t637 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1490 VDD.t32 EN.t97 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1491 a_132311_43285# D_FlipFlop_3.3-input-nand_2.C.t7 D_FlipFlop_3.3-input-nand_2.Vout.t1 Vbias.t282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1492 VDD.t255 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 VDD.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1493 VDD.t30 EN.t98 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1494 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 VDD.t972 VDD.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1495 VDD.t962 D_FlipFlop_2.3-input-nand_2.Vout.t7 D_FlipFlop_2.3-input-nand_2.C.t3 VDD.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1496 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 VDD.t306 VDD.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1497 a_72835_15797# RingCounter_0.D_FlipFlop_13.Q' Nand_Gate_7.B.t2 Vbias.t549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1498 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 a_122427_52572# Vbias.t804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1499 a_77523_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 a_76909_15797# Vbias.t777 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1500 VDD.t435 FFCLR.t56 D_FlipFlop_2.3-input-nand_2.C.t0 VDD.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1501 a_105955_13083# Nand_Gate_1.A.t10 RingCounter_0.D_FlipFlop_9.Q' Vbias.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1502 VDD.t908 Nand_Gate_6.A.t11 RingCounter_0.D_FlipFlop_12.Q' VDD.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1503 Comparator_0.Vinm CDAC8_0.switch_7.Z.t13 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1504 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 VDD.t452 VDD.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1505 Comparator_0.Vinm CDAC8_0.switch_7.Z.t12 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1506 VDD.t185 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout Nand_Gate_0.A.t1 VDD.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1507 Comparator_0.Vinm CDAC8_0.switch_7.Z.t11 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1508 a_132925_43285# D_FlipFlop_3.3-input-nand_0.Vout a_132311_43285# Vbias.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1509 a_128237_37007# Q6.t8 D_FlipFlop_2.Q' Vbias.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1510 VDD.t251 And_Gate_5.A.t4 And_Gate_5.Inverter_0.Vin VDD.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1511 Comparator_0.Vinm CDAC8_0.switch_7.Z.t10 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1512 Vbias.t364 Q1.t9 CDAC8_0.switch_2.Z.t1 VDD.t315 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1513 a_75898_28676# Q3.t9 Vbias.t747 Vbias.t746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1514 VDD.t896 Q5.t9 D_FlipFlop_3.Q' VDD.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1515 Comparator_0.Vinm CDAC8_0.switch_7.Z.t9 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1516 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 Nand_Gate_4.B.t16 VDD.t181 VDD.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1517 VDD.t135 And_Gate_2.Vout.t6 D_FlipFlop_5.3-input-nand_1.Vout VDD.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1518 RingCounter_0.D_FlipFlop_3.Q' Nand_Gate_0.B.t11 a_80239_49858# Vbias.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1519 VDD.t721 VDD.t720 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 VDD.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1520 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_5.3-input-nand_2.C.t7 VDD.t401 VDD.t369 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1521 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD.t718 VDD.t719 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1522 VDD.t399 Nand_Gate_2.A.t17 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD.t398 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1523 Vbias.t31 EN.t99 a_77523_15797# Vbias.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1524 Comparator_0.Vinm CDAC8_0.switch_6.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1525 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 VDD.t684 VDD.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1526 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 CLK.t113 VDD.t1005 VDD.t1004 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1527 Comparator_0.Vinm CDAC8_0.switch_9.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1528 Comparator_0.Vinm CDAC8_0.switch_7.Z.t8 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1529 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK.t114 VDD.t1003 VDD.t1002 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1530 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 Nand_Gate_1.A.t11 VDD.t884 VDD.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1531 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_0.D.t34 VDD.t981 VDD.t604 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1532 a_91279_52572# RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_90665_52572# Vbias.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1533 a_92725_16975# CLK.t115 Vbias.t486 Vbias.t485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1534 a_117609_15797# RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_116995_15797# Vbias.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1535 Vbias.t463 FFCLR.t57 a_132925_24200# Vbias.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1536 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 a_65125_49858# Vbias.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1537 Comparator_0.Vinm CDAC8_0.switch_7.Z.t7 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1538 VDD.t511 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 VDD.t510 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1539 Comparator_0.Vinm CDAC8_0.switch_6.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1540 D_FlipFlop_3.Q' D_FlipFlop_3.Nand_Gate_1.Vout VDD.t350 VDD.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1541 VDD.t666 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 VDD.t665 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1542 a_78881_13083# CLK.t116 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 Vbias.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1543 a_97631_52572# EN.t100 Vbias.t29 Vbias.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1544 D_FlipFlop_0.D.t35 Vbias.t567 sky130_fd_pr__cap_mim_m3_2 l=5.35 w=2
X1545 VDD.t28 EN.t101 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1546 VDD.t563 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1547 Comparator_0.Vinm CDAC8_0.switch_7.Z.t6 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1548 Comparator_0.Vinm CDAC8_0.switch_5.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1549 VDD.t437 FFCLR.t58 D_FlipFlop_4.Q' VDD.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1550 And_Gate_0.Inverter_0.Vin And_Gate_0.B.t4 a_70645_16975# Vbias.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1551 a_84619_49858# EN.t102 Vbias.t27 Vbias.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1552 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 VDD.t298 VDD.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1553 Vbias.t25 EN.t103 a_79495_13083# Vbias.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1554 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 a_120325_49858# Vbias.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1555 a_44403_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 a_43789_15797# Vbias.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1556 Nand_Gate_3.B.t0 EN.t104 VDD.t26 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1557 a_130209_36157# D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout Vbias.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1558 a_128851_44135# D_FlipFlop_0.Nand_Gate_1.Vout a_128237_44135# Vbias.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1559 a_98989_13083# RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 Vbias.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1560 Vbias.t884 Q6.t9 CDAC8_0.switch_6.Z.t3 VDD.t992 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1561 Vbias.t21 EN.t105 a_117609_15797# Vbias.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1562 VDD.t183 Nand_Gate_4.B.t17 RingCounter_0.D_FlipFlop_15.Q' VDD.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1563 a_134283_26914# And_Gate_2.Vout.t7 D_FlipFlop_5.3-input-nand_0.Vout Vbias.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1564 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 VDD.t342 VDD.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1565 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 VDD.t926 VDD.t925 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1566 a_130209_46849# D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_0.Vout Vbias.t650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1567 a_98245_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_97631_52572# Vbias.t531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1568 a_132311_19786# D_FlipFlop_7.3-input-nand_2.C.t7 D_FlipFlop_7.3-input-nand_2.Vout.t2 Vbias.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1569 Vbias.t695 Q0.t8 CDAC8_0.switch_1.Z.t3 VDD.t315 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1570 Comparator_0.Vinm CDAC8_0.switch_7.Z.t5 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1571 a_85233_49858# RingCounter_0.D_FlipFlop_4.Inverter_0.Vout a_84619_49858# Vbias.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1572 Nand_Gate_5.A.t0 EN.t106 VDD.t24 VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1573 VDD.t415 And_Gate_7.Vout.t7 D_FlipFlop_0.Inverter_1.Vout VDD.t414 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1574 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 a_89307_49858# Vbias.t736 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1575 VDD.t717 VDD.t716 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1576 a_29289_15797# RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_28675_15797# Vbias.t788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1577 VDD.t836 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 VDD.t685 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1578 Vbias.t891 FFCLR.t59 a_132925_20636# Vbias.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1579 a_130209_30478# D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_0.Vout Vbias.t467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1580 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 VDD.t919 VDD.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1581 Vbias.t17 EN.t107 a_44403_15797# Vbias.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1582 Vbias.t324 And_Gate_1.Vout.t7 D_FlipFlop_7.Inverter_1.Vout Vbias.t323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1583 VDD.t603 RingCounter_0.D_FlipFlop_9.Q' Nand_Gate_1.A.t3 VDD.t602 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1584 Comparator_0.Vinm CDAC8_0.switch_6.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1585 RingCounter_0.D_FlipFlop_4.Q' VDD.t714 VDD.t715 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1586 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 CLK.t117 VDD.t1001 VDD.t1000 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1587 a_132925_19786# D_FlipFlop_7.3-input-nand_0.Vout a_132311_19786# Vbias.t692 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1588 Comparator_0.Vinm CDAC8_0.switch_7.Z.t4 sky130_fd_pr__cap_mim_m3_2 l=2 w=22.7
X1589 a_59977_16975# Nand_Gate_7.A.t11 Vbias.t15 Vbias.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1590 Vbias.t451 And_Gate_3.Vout.t7 D_FlipFlop_4.Inverter_1.Vout Vbias.t450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1591 a_75898_35820# Q7.t9 VDD.t465 VDD.t464 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
X1592 a_28675_15797# RingCounter_0.D_FlipFlop_16.Q' RingCounter_0.D_FlipFlop_16.Q.t1 Vbias.t566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=1.44
X1593 VDD.t499 Q0.t9 D_FlipFlop_7.Q' VDD.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4176 pd=3.46 as=0.4176 ps=3.46 w=1.44 l=0.72
R0 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.t0 168.609
R1 CDAC8_0.switch_7.Z CDAC8_0.switch_7.Z.t2 168.565
R2 CDAC8_0.switch_7.Z.n0 CDAC8_0.switch_7.Z.t1 60.321
R3 CDAC8_0.switch_7.Z.n0 CDAC8_0.switch_7.Z.t3 60.321
R4 CDAC8_0.switch_7.Z.n237 CDAC8_0.switch_7.Z.n236 40.463
R5 CDAC8_0.switch_7.Z.n296 CDAC8_0.switch_7.Z.n2 20.4699
R6 CDAC8_0.switch_7.Z.n296 CDAC8_0.switch_7.Z.n295 19.9889
R7 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.n296 11.6479
R8 CDAC8_0.switch_7.Z.n48 CDAC8_0.switch_7.Z.n47 4.61363
R9 CDAC8_0.switch_7.Z.n46 CDAC8_0.switch_7.Z.n36 4.61363
R10 CDAC8_0.switch_7.Z.n53 CDAC8_0.switch_7.Z.n52 4.61363
R11 CDAC8_0.switch_7.Z.n34 CDAC8_0.switch_7.Z.n26 4.61363
R12 CDAC8_0.switch_7.Z.n56 CDAC8_0.switch_7.Z.n55 4.61363
R13 CDAC8_0.switch_7.Z.n32 CDAC8_0.switch_7.Z.n24 4.61363
R14 CDAC8_0.switch_7.Z.n61 CDAC8_0.switch_7.Z.n60 4.61363
R15 CDAC8_0.switch_7.Z.n30 CDAC8_0.switch_7.Z.n22 4.61363
R16 CDAC8_0.switch_7.Z.n65 CDAC8_0.switch_7.Z.n64 4.61363
R17 CDAC8_0.switch_7.Z.n28 CDAC8_0.switch_7.Z.n20 4.61363
R18 CDAC8_0.switch_7.Z.n69 CDAC8_0.switch_7.Z.n18 4.61363
R19 CDAC8_0.switch_7.Z.n70 CDAC8_0.switch_7.Z.n13 4.61363
R20 CDAC8_0.switch_7.Z.n74 CDAC8_0.switch_7.Z.n3 4.61363
R21 CDAC8_0.switch_7.Z.n75 CDAC8_0.switch_7.Z.n74 4.61363
R22 CDAC8_0.switch_7.Z.n15 CDAC8_0.switch_7.Z.n5 4.61363
R23 CDAC8_0.switch_7.Z.n293 CDAC8_0.switch_7.Z.n292 4.61363
R24 CDAC8_0.switch_7.Z.n287 CDAC8_0.switch_7.Z.n9 4.61363
R25 CDAC8_0.switch_7.Z.n288 CDAC8_0.switch_7.Z.n8 4.61363
R26 CDAC8_0.switch_7.Z.n283 CDAC8_0.switch_7.Z.n282 4.61363
R27 CDAC8_0.switch_7.Z.n239 CDAC8_0.switch_7.Z.n80 4.61363
R28 CDAC8_0.switch_7.Z.n280 CDAC8_0.switch_7.Z.n279 4.61363
R29 CDAC8_0.switch_7.Z.n241 CDAC8_0.switch_7.Z.n83 4.61363
R30 CDAC8_0.switch_7.Z.n275 CDAC8_0.switch_7.Z.n274 4.61363
R31 CDAC8_0.switch_7.Z.n243 CDAC8_0.switch_7.Z.n85 4.61363
R32 CDAC8_0.switch_7.Z.n272 CDAC8_0.switch_7.Z.n271 4.61363
R33 CDAC8_0.switch_7.Z.n245 CDAC8_0.switch_7.Z.n87 4.61363
R34 CDAC8_0.switch_7.Z.n247 CDAC8_0.switch_7.Z.n89 4.61363
R35 CDAC8_0.switch_7.Z.n267 CDAC8_0.switch_7.Z.n266 4.61363
R36 CDAC8_0.switch_7.Z.n264 CDAC8_0.switch_7.Z.n263 4.61363
R37 CDAC8_0.switch_7.Z.n261 CDAC8_0.switch_7.Z.n249 4.61363
R38 CDAC8_0.switch_7.Z.n221 CDAC8_0.switch_7.Z.n220 4.61363
R39 CDAC8_0.switch_7.Z.n159 CDAC8_0.switch_7.Z.n158 4.61363
R40 CDAC8_0.switch_7.Z.n156 CDAC8_0.switch_7.Z.n144 4.61363
R41 CDAC8_0.switch_7.Z.n162 CDAC8_0.switch_7.Z.n161 4.61363
R42 CDAC8_0.switch_7.Z.n142 CDAC8_0.switch_7.Z.n132 4.61363
R43 CDAC8_0.switch_7.Z.n167 CDAC8_0.switch_7.Z.n166 4.61363
R44 CDAC8_0.switch_7.Z.n140 CDAC8_0.switch_7.Z.n130 4.61363
R45 CDAC8_0.switch_7.Z.n170 CDAC8_0.switch_7.Z.n169 4.61363
R46 CDAC8_0.switch_7.Z.n138 CDAC8_0.switch_7.Z.n128 4.61363
R47 CDAC8_0.switch_7.Z.n175 CDAC8_0.switch_7.Z.n174 4.61363
R48 CDAC8_0.switch_7.Z.n136 CDAC8_0.switch_7.Z.n126 4.61363
R49 CDAC8_0.switch_7.Z.n179 CDAC8_0.switch_7.Z.n178 4.61363
R50 CDAC8_0.switch_7.Z.n134 CDAC8_0.switch_7.Z.n124 4.61363
R51 CDAC8_0.switch_7.Z.n183 CDAC8_0.switch_7.Z.n122 4.61363
R52 CDAC8_0.switch_7.Z.n184 CDAC8_0.switch_7.Z.n121 4.61363
R53 CDAC8_0.switch_7.Z.n192 CDAC8_0.switch_7.Z.n191 4.61363
R54 CDAC8_0.switch_7.Z.n188 CDAC8_0.switch_7.Z.n118 4.61363
R55 CDAC8_0.switch_7.Z.n196 CDAC8_0.switch_7.Z.n90 4.61363
R56 CDAC8_0.switch_7.Z.n197 CDAC8_0.switch_7.Z.n115 4.61363
R57 CDAC8_0.switch_7.Z.n234 CDAC8_0.switch_7.Z.n233 4.61363
R58 CDAC8_0.switch_7.Z.n113 CDAC8_0.switch_7.Z.n92 4.61363
R59 CDAC8_0.switch_7.Z.n229 CDAC8_0.switch_7.Z.n228 4.61363
R60 CDAC8_0.switch_7.Z.n111 CDAC8_0.switch_7.Z.n95 4.61363
R61 CDAC8_0.switch_7.Z.n226 CDAC8_0.switch_7.Z.n225 4.61363
R62 CDAC8_0.switch_7.Z.n109 CDAC8_0.switch_7.Z.n97 4.61363
R63 CDAC8_0.switch_7.Z.n107 CDAC8_0.switch_7.Z.n99 4.61363
R64 CDAC8_0.switch_7.Z.n218 CDAC8_0.switch_7.Z.n217 4.61363
R65 CDAC8_0.switch_7.Z.n105 CDAC8_0.switch_7.Z.n101 4.61363
R66 CDAC8_0.switch_7.Z.n211 CDAC8_0.switch_7.Z.n102 4.61363
R67 CDAC8_0.switch_7.Z.n213 CDAC8_0.switch_7.Z.n212 4.61363
R68 CDAC8_0.switch_7.Z.n48 CDAC8_0.switch_7.Z.n46 4.23363
R69 CDAC8_0.switch_7.Z.n52 CDAC8_0.switch_7.Z.n26 4.23363
R70 CDAC8_0.switch_7.Z.n56 CDAC8_0.switch_7.Z.n24 4.23363
R71 CDAC8_0.switch_7.Z.n60 CDAC8_0.switch_7.Z.n22 4.23363
R72 CDAC8_0.switch_7.Z.n65 CDAC8_0.switch_7.Z.n20 4.23363
R73 CDAC8_0.switch_7.Z.n70 CDAC8_0.switch_7.Z.n69 4.23363
R74 CDAC8_0.switch_7.Z.n292 CDAC8_0.switch_7.Z.n5 4.23363
R75 CDAC8_0.switch_7.Z.n288 CDAC8_0.switch_7.Z.n287 4.23363
R76 CDAC8_0.switch_7.Z.n283 CDAC8_0.switch_7.Z.n80 4.23363
R77 CDAC8_0.switch_7.Z.n279 CDAC8_0.switch_7.Z.n83 4.23363
R78 CDAC8_0.switch_7.Z.n275 CDAC8_0.switch_7.Z.n85 4.23363
R79 CDAC8_0.switch_7.Z.n271 CDAC8_0.switch_7.Z.n87 4.23363
R80 CDAC8_0.switch_7.Z.n267 CDAC8_0.switch_7.Z.n89 4.23363
R81 CDAC8_0.switch_7.Z.n263 CDAC8_0.switch_7.Z.n261 4.23363
R82 CDAC8_0.switch_7.Z.n158 CDAC8_0.switch_7.Z.n156 4.23363
R83 CDAC8_0.switch_7.Z.n162 CDAC8_0.switch_7.Z.n132 4.23363
R84 CDAC8_0.switch_7.Z.n166 CDAC8_0.switch_7.Z.n130 4.23363
R85 CDAC8_0.switch_7.Z.n170 CDAC8_0.switch_7.Z.n128 4.23363
R86 CDAC8_0.switch_7.Z.n174 CDAC8_0.switch_7.Z.n126 4.23363
R87 CDAC8_0.switch_7.Z.n179 CDAC8_0.switch_7.Z.n124 4.23363
R88 CDAC8_0.switch_7.Z.n184 CDAC8_0.switch_7.Z.n183 4.23363
R89 CDAC8_0.switch_7.Z.n192 CDAC8_0.switch_7.Z.n188 4.23363
R90 CDAC8_0.switch_7.Z.n197 CDAC8_0.switch_7.Z.n196 4.23363
R91 CDAC8_0.switch_7.Z.n233 CDAC8_0.switch_7.Z.n92 4.23363
R92 CDAC8_0.switch_7.Z.n229 CDAC8_0.switch_7.Z.n95 4.23363
R93 CDAC8_0.switch_7.Z.n225 CDAC8_0.switch_7.Z.n97 4.23363
R94 CDAC8_0.switch_7.Z.n221 CDAC8_0.switch_7.Z.n99 4.23363
R95 CDAC8_0.switch_7.Z.n217 CDAC8_0.switch_7.Z.n101 4.23363
R96 CDAC8_0.switch_7.Z.n213 CDAC8_0.switch_7.Z.n211 4.23363
R97 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z.n1 1.60376
R98 CDAC8_0.switch_7.Z.n262 CDAC8_0.switch_7.Z.t127 0.726216
R99 CDAC8_0.switch_7.Z.n260 CDAC8_0.switch_7.Z.t43 0.726216
R100 CDAC8_0.switch_7.Z.n264 CDAC8_0.switch_7.Z.t9 0.726216
R101 CDAC8_0.switch_7.Z.n249 CDAC8_0.switch_7.Z.t105 0.726216
R102 CDAC8_0.switch_7.Z.n210 CDAC8_0.switch_7.Z.t80 0.726216
R103 CDAC8_0.switch_7.Z.n214 CDAC8_0.switch_7.Z.t40 0.726216
R104 CDAC8_0.switch_7.Z.n102 CDAC8_0.switch_7.Z.t19 0.726216
R105 CDAC8_0.switch_7.Z.n212 CDAC8_0.switch_7.Z.t101 0.726216
R106 CDAC8_0.switch_7.Z.n159 CDAC8_0.switch_7.Z.t90 0.658247
R107 CDAC8_0.switch_7.Z.n36 CDAC8_0.switch_7.Z.t98 0.658247
R108 CDAC8_0.switch_7.Z.n47 CDAC8_0.switch_7.Z.t129 0.658247
R109 CDAC8_0.switch_7.Z.n45 CDAC8_0.switch_7.Z.t36 0.658247
R110 CDAC8_0.switch_7.Z.n49 CDAC8_0.switch_7.Z.t117 0.658247
R111 CDAC8_0.switch_7.Z.n144 CDAC8_0.switch_7.Z.t8 0.658247
R112 CDAC8_0.switch_7.Z.n157 CDAC8_0.switch_7.Z.t30 0.658247
R113 CDAC8_0.switch_7.Z.n155 CDAC8_0.switch_7.Z.t70 0.658247
R114 CDAC8_0.switch_7.Z.n160 CDAC8_0.switch_7.Z.t86 0.611304
R115 CDAC8_0.switch_7.Z.n129 CDAC8_0.switch_7.Z.t112 0.611304
R116 CDAC8_0.switch_7.Z.n168 CDAC8_0.switch_7.Z.t107 0.611304
R117 CDAC8_0.switch_7.Z.n125 CDAC8_0.switch_7.Z.t32 0.611304
R118 CDAC8_0.switch_7.Z.n176 CDAC8_0.switch_7.Z.t49 0.611304
R119 CDAC8_0.switch_7.Z.n177 CDAC8_0.switch_7.Z.t44 0.611304
R120 CDAC8_0.switch_7.Z.n189 CDAC8_0.switch_7.Z.t69 0.611304
R121 CDAC8_0.switch_7.Z.n190 CDAC8_0.switch_7.Z.t65 0.611304
R122 CDAC8_0.switch_7.Z.n35 CDAC8_0.switch_7.Z.t92 0.611304
R123 CDAC8_0.switch_7.Z.n33 CDAC8_0.switch_7.Z.t120 0.611304
R124 CDAC8_0.switch_7.Z.n31 CDAC8_0.switch_7.Z.t113 0.611304
R125 CDAC8_0.switch_7.Z.n29 CDAC8_0.switch_7.Z.t39 0.611304
R126 CDAC8_0.switch_7.Z.n27 CDAC8_0.switch_7.Z.t58 0.611304
R127 CDAC8_0.switch_7.Z.n12 CDAC8_0.switch_7.Z.t51 0.611304
R128 CDAC8_0.switch_7.Z.n294 CDAC8_0.switch_7.Z.t76 0.611304
R129 CDAC8_0.switch_7.Z.n4 CDAC8_0.switch_7.Z.t71 0.611304
R130 CDAC8_0.switch_7.Z.n238 CDAC8_0.switch_7.Z.t128 0.611304
R131 CDAC8_0.switch_7.Z.n240 CDAC8_0.switch_7.Z.t21 0.611304
R132 CDAC8_0.switch_7.Z.n242 CDAC8_0.switch_7.Z.t16 0.611304
R133 CDAC8_0.switch_7.Z.n244 CDAC8_0.switch_7.Z.t38 0.611304
R134 CDAC8_0.switch_7.Z.n246 CDAC8_0.switch_7.Z.t89 0.611304
R135 CDAC8_0.switch_7.Z.n248 CDAC8_0.switch_7.Z.t84 0.611304
R136 CDAC8_0.switch_7.Z.n25 CDAC8_0.switch_7.Z.t125 0.611304
R137 CDAC8_0.switch_7.Z.n54 CDAC8_0.switch_7.Z.t23 0.611304
R138 CDAC8_0.switch_7.Z.n21 CDAC8_0.switch_7.Z.t17 0.611304
R139 CDAC8_0.switch_7.Z.n62 CDAC8_0.switch_7.Z.t66 0.611304
R140 CDAC8_0.switch_7.Z.n63 CDAC8_0.switch_7.Z.t85 0.611304
R141 CDAC8_0.switch_7.Z.n17 CDAC8_0.switch_7.Z.t81 0.611304
R142 CDAC8_0.switch_7.Z.n16 CDAC8_0.switch_7.Z.t106 0.611304
R143 CDAC8_0.switch_7.Z.n14 CDAC8_0.switch_7.Z.t103 0.611304
R144 CDAC8_0.switch_7.Z.n81 CDAC8_0.switch_7.Z.t35 0.611304
R145 CDAC8_0.switch_7.Z.n281 CDAC8_0.switch_7.Z.t52 0.611304
R146 CDAC8_0.switch_7.Z.n82 CDAC8_0.switch_7.Z.t46 0.611304
R147 CDAC8_0.switch_7.Z.n273 CDAC8_0.switch_7.Z.t64 0.611304
R148 CDAC8_0.switch_7.Z.n86 CDAC8_0.switch_7.Z.t122 0.611304
R149 CDAC8_0.switch_7.Z.n44 CDAC8_0.switch_7.Z.t29 0.611304
R150 CDAC8_0.switch_7.Z.n42 CDAC8_0.switch_7.Z.t54 0.611304
R151 CDAC8_0.switch_7.Z.n40 CDAC8_0.switch_7.Z.t48 0.611304
R152 CDAC8_0.switch_7.Z.n38 CDAC8_0.switch_7.Z.t100 0.611304
R153 CDAC8_0.switch_7.Z.n11 CDAC8_0.switch_7.Z.t121 0.611304
R154 CDAC8_0.switch_7.Z.n72 CDAC8_0.switch_7.Z.t114 0.611304
R155 CDAC8_0.switch_7.Z.n6 CDAC8_0.switch_7.Z.t14 0.611304
R156 CDAC8_0.switch_7.Z.n290 CDAC8_0.switch_7.Z.t6 0.611304
R157 CDAC8_0.switch_7.Z.n7 CDAC8_0.switch_7.Z.t62 0.611304
R158 CDAC8_0.switch_7.Z.n251 CDAC8_0.switch_7.Z.t82 0.611304
R159 CDAC8_0.switch_7.Z.n253 CDAC8_0.switch_7.Z.t77 0.611304
R160 CDAC8_0.switch_7.Z.n255 CDAC8_0.switch_7.Z.t99 0.611304
R161 CDAC8_0.switch_7.Z.n50 CDAC8_0.switch_7.Z.t111 0.611304
R162 CDAC8_0.switch_7.Z.n23 CDAC8_0.switch_7.Z.t12 0.611304
R163 CDAC8_0.switch_7.Z.n58 CDAC8_0.switch_7.Z.t5 0.611304
R164 CDAC8_0.switch_7.Z.n19 CDAC8_0.switch_7.Z.t57 0.611304
R165 CDAC8_0.switch_7.Z.n67 CDAC8_0.switch_7.Z.t74 0.611304
R166 CDAC8_0.switch_7.Z.n10 CDAC8_0.switch_7.Z.t68 0.611304
R167 CDAC8_0.switch_7.Z.n76 CDAC8_0.switch_7.Z.t97 0.611304
R168 CDAC8_0.switch_7.Z.n78 CDAC8_0.switch_7.Z.t91 0.611304
R169 CDAC8_0.switch_7.Z.n285 CDAC8_0.switch_7.Z.t20 0.611304
R170 CDAC8_0.switch_7.Z.n79 CDAC8_0.switch_7.Z.t42 0.611304
R171 CDAC8_0.switch_7.Z.n277 CDAC8_0.switch_7.Z.t37 0.611304
R172 CDAC8_0.switch_7.Z.n84 CDAC8_0.switch_7.Z.t55 0.611304
R173 CDAC8_0.switch_7.Z.n269 CDAC8_0.switch_7.Z.t109 0.611304
R174 CDAC8_0.switch_7.Z.n88 CDAC8_0.switch_7.Z.t104 0.611304
R175 CDAC8_0.switch_7.Z.n257 CDAC8_0.switch_7.Z.t28 0.611304
R176 CDAC8_0.switch_7.Z.n259 CDAC8_0.switch_7.Z.t22 0.611304
R177 CDAC8_0.switch_7.Z.n265 CDAC8_0.switch_7.Z.t118 0.611304
R178 CDAC8_0.switch_7.Z.n235 CDAC8_0.switch_7.Z.t123 0.611304
R179 CDAC8_0.switch_7.Z.n91 CDAC8_0.switch_7.Z.t15 0.611304
R180 CDAC8_0.switch_7.Z.n227 CDAC8_0.switch_7.Z.t10 0.611304
R181 CDAC8_0.switch_7.Z.n96 CDAC8_0.switch_7.Z.t31 0.611304
R182 CDAC8_0.switch_7.Z.n219 CDAC8_0.switch_7.Z.t83 0.611304
R183 CDAC8_0.switch_7.Z.n100 CDAC8_0.switch_7.Z.t79 0.611304
R184 CDAC8_0.switch_7.Z.n143 CDAC8_0.switch_7.Z.t4 0.611304
R185 CDAC8_0.switch_7.Z.n141 CDAC8_0.switch_7.Z.t33 0.611304
R186 CDAC8_0.switch_7.Z.n139 CDAC8_0.switch_7.Z.t26 0.611304
R187 CDAC8_0.switch_7.Z.n137 CDAC8_0.switch_7.Z.t75 0.611304
R188 CDAC8_0.switch_7.Z.n135 CDAC8_0.switch_7.Z.t96 0.611304
R189 CDAC8_0.switch_7.Z.n133 CDAC8_0.switch_7.Z.t88 0.611304
R190 CDAC8_0.switch_7.Z.n120 CDAC8_0.switch_7.Z.t116 0.611304
R191 CDAC8_0.switch_7.Z.n117 CDAC8_0.switch_7.Z.t110 0.611304
R192 CDAC8_0.switch_7.Z.n114 CDAC8_0.switch_7.Z.t41 0.611304
R193 CDAC8_0.switch_7.Z.n112 CDAC8_0.switch_7.Z.t60 0.611304
R194 CDAC8_0.switch_7.Z.n110 CDAC8_0.switch_7.Z.t56 0.611304
R195 CDAC8_0.switch_7.Z.n108 CDAC8_0.switch_7.Z.t73 0.611304
R196 CDAC8_0.switch_7.Z.n106 CDAC8_0.switch_7.Z.t130 0.611304
R197 CDAC8_0.switch_7.Z.n131 CDAC8_0.switch_7.Z.t25 0.611304
R198 CDAC8_0.switch_7.Z.n164 CDAC8_0.switch_7.Z.t50 0.611304
R199 CDAC8_0.switch_7.Z.n127 CDAC8_0.switch_7.Z.t45 0.611304
R200 CDAC8_0.switch_7.Z.n172 CDAC8_0.switch_7.Z.t95 0.611304
R201 CDAC8_0.switch_7.Z.n123 CDAC8_0.switch_7.Z.t115 0.611304
R202 CDAC8_0.switch_7.Z.n181 CDAC8_0.switch_7.Z.t108 0.611304
R203 CDAC8_0.switch_7.Z.n116 CDAC8_0.switch_7.Z.t7 0.611304
R204 CDAC8_0.switch_7.Z.n194 CDAC8_0.switch_7.Z.t131 0.611304
R205 CDAC8_0.switch_7.Z.n93 CDAC8_0.switch_7.Z.t59 0.611304
R206 CDAC8_0.switch_7.Z.n231 CDAC8_0.switch_7.Z.t78 0.611304
R207 CDAC8_0.switch_7.Z.n94 CDAC8_0.switch_7.Z.t72 0.611304
R208 CDAC8_0.switch_7.Z.n223 CDAC8_0.switch_7.Z.t94 0.611304
R209 CDAC8_0.switch_7.Z.n154 CDAC8_0.switch_7.Z.t67 0.611304
R210 CDAC8_0.switch_7.Z.n152 CDAC8_0.switch_7.Z.t93 0.611304
R211 CDAC8_0.switch_7.Z.n150 CDAC8_0.switch_7.Z.t87 0.611304
R212 CDAC8_0.switch_7.Z.n148 CDAC8_0.switch_7.Z.t13 0.611304
R213 CDAC8_0.switch_7.Z.n146 CDAC8_0.switch_7.Z.t34 0.611304
R214 CDAC8_0.switch_7.Z.n119 CDAC8_0.switch_7.Z.t27 0.611304
R215 CDAC8_0.switch_7.Z.n186 CDAC8_0.switch_7.Z.t53 0.611304
R216 CDAC8_0.switch_7.Z.n103 CDAC8_0.switch_7.Z.t47 0.611304
R217 CDAC8_0.switch_7.Z.n199 CDAC8_0.switch_7.Z.t102 0.611304
R218 CDAC8_0.switch_7.Z.n201 CDAC8_0.switch_7.Z.t124 0.611304
R219 CDAC8_0.switch_7.Z.n203 CDAC8_0.switch_7.Z.t119 0.611304
R220 CDAC8_0.switch_7.Z.n205 CDAC8_0.switch_7.Z.t11 0.611304
R221 CDAC8_0.switch_7.Z.n207 CDAC8_0.switch_7.Z.t63 0.611304
R222 CDAC8_0.switch_7.Z.n209 CDAC8_0.switch_7.Z.t61 0.611304
R223 CDAC8_0.switch_7.Z.n98 CDAC8_0.switch_7.Z.t24 0.611304
R224 CDAC8_0.switch_7.Z.n215 CDAC8_0.switch_7.Z.t18 0.611304
R225 CDAC8_0.switch_7.Z.n104 CDAC8_0.switch_7.Z.t126 0.611304
R226 CDAC8_0.switch_7.Z.n276 CDAC8_0.switch_7.Z.n275 0.3805
R227 CDAC8_0.switch_7.Z.n279 CDAC8_0.switch_7.Z.n278 0.3805
R228 CDAC8_0.switch_7.Z.n284 CDAC8_0.switch_7.Z.n283 0.3805
R229 CDAC8_0.switch_7.Z.n287 CDAC8_0.switch_7.Z.n286 0.3805
R230 CDAC8_0.switch_7.Z.n77 CDAC8_0.switch_7.Z.n5 0.3805
R231 CDAC8_0.switch_7.Z.n69 CDAC8_0.switch_7.Z.n68 0.3805
R232 CDAC8_0.switch_7.Z.n66 CDAC8_0.switch_7.Z.n65 0.3805
R233 CDAC8_0.switch_7.Z.n60 CDAC8_0.switch_7.Z.n59 0.3805
R234 CDAC8_0.switch_7.Z.n57 CDAC8_0.switch_7.Z.n56 0.3805
R235 CDAC8_0.switch_7.Z.n52 CDAC8_0.switch_7.Z.n51 0.3805
R236 CDAC8_0.switch_7.Z.n49 CDAC8_0.switch_7.Z.n48 0.3805
R237 CDAC8_0.switch_7.Z.n271 CDAC8_0.switch_7.Z.n270 0.3805
R238 CDAC8_0.switch_7.Z.n256 CDAC8_0.switch_7.Z.n87 0.3805
R239 CDAC8_0.switch_7.Z.n254 CDAC8_0.switch_7.Z.n85 0.3805
R240 CDAC8_0.switch_7.Z.n252 CDAC8_0.switch_7.Z.n83 0.3805
R241 CDAC8_0.switch_7.Z.n250 CDAC8_0.switch_7.Z.n80 0.3805
R242 CDAC8_0.switch_7.Z.n289 CDAC8_0.switch_7.Z.n288 0.3805
R243 CDAC8_0.switch_7.Z.n292 CDAC8_0.switch_7.Z.n291 0.3805
R244 CDAC8_0.switch_7.Z.n74 CDAC8_0.switch_7.Z.n73 0.3805
R245 CDAC8_0.switch_7.Z.n71 CDAC8_0.switch_7.Z.n70 0.3805
R246 CDAC8_0.switch_7.Z.n37 CDAC8_0.switch_7.Z.n20 0.3805
R247 CDAC8_0.switch_7.Z.n39 CDAC8_0.switch_7.Z.n22 0.3805
R248 CDAC8_0.switch_7.Z.n41 CDAC8_0.switch_7.Z.n24 0.3805
R249 CDAC8_0.switch_7.Z.n43 CDAC8_0.switch_7.Z.n26 0.3805
R250 CDAC8_0.switch_7.Z.n46 CDAC8_0.switch_7.Z.n45 0.3805
R251 CDAC8_0.switch_7.Z.n258 CDAC8_0.switch_7.Z.n89 0.3805
R252 CDAC8_0.switch_7.Z.n268 CDAC8_0.switch_7.Z.n267 0.3805
R253 CDAC8_0.switch_7.Z.n263 CDAC8_0.switch_7.Z.n262 0.3805
R254 CDAC8_0.switch_7.Z.n261 CDAC8_0.switch_7.Z.n260 0.3805
R255 CDAC8_0.switch_7.Z.n204 CDAC8_0.switch_7.Z.n97 0.3805
R256 CDAC8_0.switch_7.Z.n202 CDAC8_0.switch_7.Z.n95 0.3805
R257 CDAC8_0.switch_7.Z.n200 CDAC8_0.switch_7.Z.n92 0.3805
R258 CDAC8_0.switch_7.Z.n198 CDAC8_0.switch_7.Z.n197 0.3805
R259 CDAC8_0.switch_7.Z.n188 CDAC8_0.switch_7.Z.n187 0.3805
R260 CDAC8_0.switch_7.Z.n185 CDAC8_0.switch_7.Z.n184 0.3805
R261 CDAC8_0.switch_7.Z.n145 CDAC8_0.switch_7.Z.n124 0.3805
R262 CDAC8_0.switch_7.Z.n147 CDAC8_0.switch_7.Z.n126 0.3805
R263 CDAC8_0.switch_7.Z.n149 CDAC8_0.switch_7.Z.n128 0.3805
R264 CDAC8_0.switch_7.Z.n151 CDAC8_0.switch_7.Z.n130 0.3805
R265 CDAC8_0.switch_7.Z.n153 CDAC8_0.switch_7.Z.n132 0.3805
R266 CDAC8_0.switch_7.Z.n156 CDAC8_0.switch_7.Z.n155 0.3805
R267 CDAC8_0.switch_7.Z.n206 CDAC8_0.switch_7.Z.n99 0.3805
R268 CDAC8_0.switch_7.Z.n222 CDAC8_0.switch_7.Z.n221 0.3805
R269 CDAC8_0.switch_7.Z.n225 CDAC8_0.switch_7.Z.n224 0.3805
R270 CDAC8_0.switch_7.Z.n230 CDAC8_0.switch_7.Z.n229 0.3805
R271 CDAC8_0.switch_7.Z.n233 CDAC8_0.switch_7.Z.n232 0.3805
R272 CDAC8_0.switch_7.Z.n196 CDAC8_0.switch_7.Z.n195 0.3805
R273 CDAC8_0.switch_7.Z.n193 CDAC8_0.switch_7.Z.n192 0.3805
R274 CDAC8_0.switch_7.Z.n183 CDAC8_0.switch_7.Z.n182 0.3805
R275 CDAC8_0.switch_7.Z.n180 CDAC8_0.switch_7.Z.n179 0.3805
R276 CDAC8_0.switch_7.Z.n174 CDAC8_0.switch_7.Z.n173 0.3805
R277 CDAC8_0.switch_7.Z.n171 CDAC8_0.switch_7.Z.n170 0.3805
R278 CDAC8_0.switch_7.Z.n166 CDAC8_0.switch_7.Z.n165 0.3805
R279 CDAC8_0.switch_7.Z.n163 CDAC8_0.switch_7.Z.n162 0.3805
R280 CDAC8_0.switch_7.Z.n158 CDAC8_0.switch_7.Z.n157 0.3805
R281 CDAC8_0.switch_7.Z.n217 CDAC8_0.switch_7.Z.n216 0.3805
R282 CDAC8_0.switch_7.Z.n208 CDAC8_0.switch_7.Z.n101 0.3805
R283 CDAC8_0.switch_7.Z.n211 CDAC8_0.switch_7.Z.n210 0.3805
R284 CDAC8_0.switch_7.Z.n214 CDAC8_0.switch_7.Z.n213 0.3805
R285 CDAC8_0.switch_7.Z.n1 CDAC8_0.switch_7.Z 0.259656
R286 CDAC8_0.switch_7.Z.n297 CDAC8_0.switch_7.Z 0.166261
R287 CDAC8_0.switch_7.Z.n17 CDAC8_0.switch_7.Z.n16 0.162356
R288 CDAC8_0.switch_7.Z.n50 CDAC8_0.switch_7.Z.n49 0.115412
R289 CDAC8_0.switch_7.Z.n51 CDAC8_0.switch_7.Z.n23 0.115412
R290 CDAC8_0.switch_7.Z.n58 CDAC8_0.switch_7.Z.n57 0.115412
R291 CDAC8_0.switch_7.Z.n59 CDAC8_0.switch_7.Z.n19 0.115412
R292 CDAC8_0.switch_7.Z.n67 CDAC8_0.switch_7.Z.n66 0.115412
R293 CDAC8_0.switch_7.Z.n68 CDAC8_0.switch_7.Z.n10 0.115412
R294 CDAC8_0.switch_7.Z.n76 CDAC8_0.switch_7.Z.n75 0.115412
R295 CDAC8_0.switch_7.Z.n78 CDAC8_0.switch_7.Z.n77 0.115412
R296 CDAC8_0.switch_7.Z.n286 CDAC8_0.switch_7.Z.n285 0.115412
R297 CDAC8_0.switch_7.Z.n284 CDAC8_0.switch_7.Z.n79 0.115412
R298 CDAC8_0.switch_7.Z.n278 CDAC8_0.switch_7.Z.n277 0.115412
R299 CDAC8_0.switch_7.Z.n276 CDAC8_0.switch_7.Z.n84 0.115412
R300 CDAC8_0.switch_7.Z.n270 CDAC8_0.switch_7.Z.n269 0.115412
R301 CDAC8_0.switch_7.Z.n268 CDAC8_0.switch_7.Z.n88 0.115412
R302 CDAC8_0.switch_7.Z.n45 CDAC8_0.switch_7.Z.n44 0.115412
R303 CDAC8_0.switch_7.Z.n43 CDAC8_0.switch_7.Z.n42 0.115412
R304 CDAC8_0.switch_7.Z.n41 CDAC8_0.switch_7.Z.n40 0.115412
R305 CDAC8_0.switch_7.Z.n39 CDAC8_0.switch_7.Z.n38 0.115412
R306 CDAC8_0.switch_7.Z.n37 CDAC8_0.switch_7.Z.n11 0.115412
R307 CDAC8_0.switch_7.Z.n72 CDAC8_0.switch_7.Z.n71 0.115412
R308 CDAC8_0.switch_7.Z.n73 CDAC8_0.switch_7.Z.n6 0.115412
R309 CDAC8_0.switch_7.Z.n291 CDAC8_0.switch_7.Z.n290 0.115412
R310 CDAC8_0.switch_7.Z.n289 CDAC8_0.switch_7.Z.n7 0.115412
R311 CDAC8_0.switch_7.Z.n251 CDAC8_0.switch_7.Z.n250 0.115412
R312 CDAC8_0.switch_7.Z.n253 CDAC8_0.switch_7.Z.n252 0.115412
R313 CDAC8_0.switch_7.Z.n255 CDAC8_0.switch_7.Z.n254 0.115412
R314 CDAC8_0.switch_7.Z.n257 CDAC8_0.switch_7.Z.n256 0.115412
R315 CDAC8_0.switch_7.Z.n259 CDAC8_0.switch_7.Z.n258 0.115412
R316 CDAC8_0.switch_7.Z.n47 CDAC8_0.switch_7.Z.n25 0.115412
R317 CDAC8_0.switch_7.Z.n54 CDAC8_0.switch_7.Z.n53 0.115412
R318 CDAC8_0.switch_7.Z.n55 CDAC8_0.switch_7.Z.n21 0.115412
R319 CDAC8_0.switch_7.Z.n62 CDAC8_0.switch_7.Z.n61 0.115412
R320 CDAC8_0.switch_7.Z.n64 CDAC8_0.switch_7.Z.n63 0.115412
R321 CDAC8_0.switch_7.Z.n18 CDAC8_0.switch_7.Z.n17 0.115412
R322 CDAC8_0.switch_7.Z.n15 CDAC8_0.switch_7.Z.n14 0.115412
R323 CDAC8_0.switch_7.Z.n81 CDAC8_0.switch_7.Z.n9 0.115412
R324 CDAC8_0.switch_7.Z.n282 CDAC8_0.switch_7.Z.n281 0.115412
R325 CDAC8_0.switch_7.Z.n280 CDAC8_0.switch_7.Z.n82 0.115412
R326 CDAC8_0.switch_7.Z.n274 CDAC8_0.switch_7.Z.n273 0.115412
R327 CDAC8_0.switch_7.Z.n272 CDAC8_0.switch_7.Z.n86 0.115412
R328 CDAC8_0.switch_7.Z.n266 CDAC8_0.switch_7.Z.n265 0.115412
R329 CDAC8_0.switch_7.Z.n36 CDAC8_0.switch_7.Z.n35 0.115412
R330 CDAC8_0.switch_7.Z.n34 CDAC8_0.switch_7.Z.n33 0.115412
R331 CDAC8_0.switch_7.Z.n32 CDAC8_0.switch_7.Z.n31 0.115412
R332 CDAC8_0.switch_7.Z.n30 CDAC8_0.switch_7.Z.n29 0.115412
R333 CDAC8_0.switch_7.Z.n28 CDAC8_0.switch_7.Z.n27 0.115412
R334 CDAC8_0.switch_7.Z.n13 CDAC8_0.switch_7.Z.n12 0.115412
R335 CDAC8_0.switch_7.Z.n293 CDAC8_0.switch_7.Z.n4 0.115412
R336 CDAC8_0.switch_7.Z.n240 CDAC8_0.switch_7.Z.n239 0.115412
R337 CDAC8_0.switch_7.Z.n242 CDAC8_0.switch_7.Z.n241 0.115412
R338 CDAC8_0.switch_7.Z.n244 CDAC8_0.switch_7.Z.n243 0.115412
R339 CDAC8_0.switch_7.Z.n246 CDAC8_0.switch_7.Z.n245 0.115412
R340 CDAC8_0.switch_7.Z.n248 CDAC8_0.switch_7.Z.n247 0.115412
R341 CDAC8_0.switch_7.Z.n155 CDAC8_0.switch_7.Z.n154 0.115412
R342 CDAC8_0.switch_7.Z.n153 CDAC8_0.switch_7.Z.n152 0.115412
R343 CDAC8_0.switch_7.Z.n151 CDAC8_0.switch_7.Z.n150 0.115412
R344 CDAC8_0.switch_7.Z.n149 CDAC8_0.switch_7.Z.n148 0.115412
R345 CDAC8_0.switch_7.Z.n147 CDAC8_0.switch_7.Z.n146 0.115412
R346 CDAC8_0.switch_7.Z.n145 CDAC8_0.switch_7.Z.n119 0.115412
R347 CDAC8_0.switch_7.Z.n186 CDAC8_0.switch_7.Z.n185 0.115412
R348 CDAC8_0.switch_7.Z.n187 CDAC8_0.switch_7.Z.n103 0.115412
R349 CDAC8_0.switch_7.Z.n199 CDAC8_0.switch_7.Z.n198 0.115412
R350 CDAC8_0.switch_7.Z.n201 CDAC8_0.switch_7.Z.n200 0.115412
R351 CDAC8_0.switch_7.Z.n203 CDAC8_0.switch_7.Z.n202 0.115412
R352 CDAC8_0.switch_7.Z.n205 CDAC8_0.switch_7.Z.n204 0.115412
R353 CDAC8_0.switch_7.Z.n207 CDAC8_0.switch_7.Z.n206 0.115412
R354 CDAC8_0.switch_7.Z.n209 CDAC8_0.switch_7.Z.n208 0.115412
R355 CDAC8_0.switch_7.Z.n157 CDAC8_0.switch_7.Z.n131 0.115412
R356 CDAC8_0.switch_7.Z.n164 CDAC8_0.switch_7.Z.n163 0.115412
R357 CDAC8_0.switch_7.Z.n165 CDAC8_0.switch_7.Z.n127 0.115412
R358 CDAC8_0.switch_7.Z.n172 CDAC8_0.switch_7.Z.n171 0.115412
R359 CDAC8_0.switch_7.Z.n173 CDAC8_0.switch_7.Z.n123 0.115412
R360 CDAC8_0.switch_7.Z.n181 CDAC8_0.switch_7.Z.n180 0.115412
R361 CDAC8_0.switch_7.Z.n182 CDAC8_0.switch_7.Z.n116 0.115412
R362 CDAC8_0.switch_7.Z.n194 CDAC8_0.switch_7.Z.n193 0.115412
R363 CDAC8_0.switch_7.Z.n195 CDAC8_0.switch_7.Z.n93 0.115412
R364 CDAC8_0.switch_7.Z.n232 CDAC8_0.switch_7.Z.n231 0.115412
R365 CDAC8_0.switch_7.Z.n230 CDAC8_0.switch_7.Z.n94 0.115412
R366 CDAC8_0.switch_7.Z.n224 CDAC8_0.switch_7.Z.n223 0.115412
R367 CDAC8_0.switch_7.Z.n222 CDAC8_0.switch_7.Z.n98 0.115412
R368 CDAC8_0.switch_7.Z.n216 CDAC8_0.switch_7.Z.n215 0.115412
R369 CDAC8_0.switch_7.Z.n144 CDAC8_0.switch_7.Z.n143 0.115412
R370 CDAC8_0.switch_7.Z.n142 CDAC8_0.switch_7.Z.n141 0.115412
R371 CDAC8_0.switch_7.Z.n140 CDAC8_0.switch_7.Z.n139 0.115412
R372 CDAC8_0.switch_7.Z.n138 CDAC8_0.switch_7.Z.n137 0.115412
R373 CDAC8_0.switch_7.Z.n136 CDAC8_0.switch_7.Z.n135 0.115412
R374 CDAC8_0.switch_7.Z.n134 CDAC8_0.switch_7.Z.n133 0.115412
R375 CDAC8_0.switch_7.Z.n121 CDAC8_0.switch_7.Z.n120 0.115412
R376 CDAC8_0.switch_7.Z.n118 CDAC8_0.switch_7.Z.n117 0.115412
R377 CDAC8_0.switch_7.Z.n115 CDAC8_0.switch_7.Z.n114 0.115412
R378 CDAC8_0.switch_7.Z.n113 CDAC8_0.switch_7.Z.n112 0.115412
R379 CDAC8_0.switch_7.Z.n111 CDAC8_0.switch_7.Z.n110 0.115412
R380 CDAC8_0.switch_7.Z.n109 CDAC8_0.switch_7.Z.n108 0.115412
R381 CDAC8_0.switch_7.Z.n107 CDAC8_0.switch_7.Z.n106 0.115412
R382 CDAC8_0.switch_7.Z.n105 CDAC8_0.switch_7.Z.n104 0.115412
R383 CDAC8_0.switch_7.Z.n160 CDAC8_0.switch_7.Z.n159 0.115412
R384 CDAC8_0.switch_7.Z.n161 CDAC8_0.switch_7.Z.n129 0.115412
R385 CDAC8_0.switch_7.Z.n168 CDAC8_0.switch_7.Z.n167 0.115412
R386 CDAC8_0.switch_7.Z.n169 CDAC8_0.switch_7.Z.n125 0.115412
R387 CDAC8_0.switch_7.Z.n176 CDAC8_0.switch_7.Z.n175 0.115412
R388 CDAC8_0.switch_7.Z.n178 CDAC8_0.switch_7.Z.n177 0.115412
R389 CDAC8_0.switch_7.Z.n191 CDAC8_0.switch_7.Z.n190 0.115412
R390 CDAC8_0.switch_7.Z.n234 CDAC8_0.switch_7.Z.n91 0.115412
R391 CDAC8_0.switch_7.Z.n228 CDAC8_0.switch_7.Z.n227 0.115412
R392 CDAC8_0.switch_7.Z.n226 CDAC8_0.switch_7.Z.n96 0.115412
R393 CDAC8_0.switch_7.Z.n220 CDAC8_0.switch_7.Z.n219 0.115412
R394 CDAC8_0.switch_7.Z.n218 CDAC8_0.switch_7.Z.n100 0.115412
R395 CDAC8_0.switch_7.Z.n295 CDAC8_0.switch_7.Z.n294 0.0845094
R396 CDAC8_0.switch_7.Z.n238 CDAC8_0.switch_7.Z.n237 0.0845094
R397 CDAC8_0.switch_7.Z.n189 CDAC8_0.switch_7.Z.n2 0.0845094
R398 CDAC8_0.switch_7.Z.n236 CDAC8_0.switch_7.Z.n235 0.0845094
R399 CDAC8_0.switch_7.Z.n51 CDAC8_0.switch_7.Z.n50 0.0474438
R400 CDAC8_0.switch_7.Z.n57 CDAC8_0.switch_7.Z.n23 0.0474438
R401 CDAC8_0.switch_7.Z.n59 CDAC8_0.switch_7.Z.n58 0.0474438
R402 CDAC8_0.switch_7.Z.n66 CDAC8_0.switch_7.Z.n19 0.0474438
R403 CDAC8_0.switch_7.Z.n68 CDAC8_0.switch_7.Z.n67 0.0474438
R404 CDAC8_0.switch_7.Z.n75 CDAC8_0.switch_7.Z.n10 0.0474438
R405 CDAC8_0.switch_7.Z.n77 CDAC8_0.switch_7.Z.n76 0.0474438
R406 CDAC8_0.switch_7.Z.n286 CDAC8_0.switch_7.Z.n78 0.0474438
R407 CDAC8_0.switch_7.Z.n285 CDAC8_0.switch_7.Z.n284 0.0474438
R408 CDAC8_0.switch_7.Z.n278 CDAC8_0.switch_7.Z.n79 0.0474438
R409 CDAC8_0.switch_7.Z.n277 CDAC8_0.switch_7.Z.n276 0.0474438
R410 CDAC8_0.switch_7.Z.n270 CDAC8_0.switch_7.Z.n84 0.0474438
R411 CDAC8_0.switch_7.Z.n269 CDAC8_0.switch_7.Z.n268 0.0474438
R412 CDAC8_0.switch_7.Z.n262 CDAC8_0.switch_7.Z.n88 0.0474438
R413 CDAC8_0.switch_7.Z.n44 CDAC8_0.switch_7.Z.n43 0.0474438
R414 CDAC8_0.switch_7.Z.n42 CDAC8_0.switch_7.Z.n41 0.0474438
R415 CDAC8_0.switch_7.Z.n40 CDAC8_0.switch_7.Z.n39 0.0474438
R416 CDAC8_0.switch_7.Z.n38 CDAC8_0.switch_7.Z.n37 0.0474438
R417 CDAC8_0.switch_7.Z.n71 CDAC8_0.switch_7.Z.n11 0.0474438
R418 CDAC8_0.switch_7.Z.n73 CDAC8_0.switch_7.Z.n72 0.0474438
R419 CDAC8_0.switch_7.Z.n291 CDAC8_0.switch_7.Z.n6 0.0474438
R420 CDAC8_0.switch_7.Z.n290 CDAC8_0.switch_7.Z.n289 0.0474438
R421 CDAC8_0.switch_7.Z.n250 CDAC8_0.switch_7.Z.n7 0.0474438
R422 CDAC8_0.switch_7.Z.n252 CDAC8_0.switch_7.Z.n251 0.0474438
R423 CDAC8_0.switch_7.Z.n254 CDAC8_0.switch_7.Z.n253 0.0474438
R424 CDAC8_0.switch_7.Z.n256 CDAC8_0.switch_7.Z.n255 0.0474438
R425 CDAC8_0.switch_7.Z.n258 CDAC8_0.switch_7.Z.n257 0.0474438
R426 CDAC8_0.switch_7.Z.n260 CDAC8_0.switch_7.Z.n259 0.0474438
R427 CDAC8_0.switch_7.Z.n53 CDAC8_0.switch_7.Z.n25 0.0474438
R428 CDAC8_0.switch_7.Z.n55 CDAC8_0.switch_7.Z.n54 0.0474438
R429 CDAC8_0.switch_7.Z.n61 CDAC8_0.switch_7.Z.n21 0.0474438
R430 CDAC8_0.switch_7.Z.n64 CDAC8_0.switch_7.Z.n62 0.0474438
R431 CDAC8_0.switch_7.Z.n63 CDAC8_0.switch_7.Z.n18 0.0474438
R432 CDAC8_0.switch_7.Z.n16 CDAC8_0.switch_7.Z.n15 0.0474438
R433 CDAC8_0.switch_7.Z.n14 CDAC8_0.switch_7.Z.n9 0.0474438
R434 CDAC8_0.switch_7.Z.n282 CDAC8_0.switch_7.Z.n81 0.0474438
R435 CDAC8_0.switch_7.Z.n281 CDAC8_0.switch_7.Z.n280 0.0474438
R436 CDAC8_0.switch_7.Z.n274 CDAC8_0.switch_7.Z.n82 0.0474438
R437 CDAC8_0.switch_7.Z.n273 CDAC8_0.switch_7.Z.n272 0.0474438
R438 CDAC8_0.switch_7.Z.n266 CDAC8_0.switch_7.Z.n86 0.0474438
R439 CDAC8_0.switch_7.Z.n265 CDAC8_0.switch_7.Z.n264 0.0474438
R440 CDAC8_0.switch_7.Z.n35 CDAC8_0.switch_7.Z.n34 0.0474438
R441 CDAC8_0.switch_7.Z.n33 CDAC8_0.switch_7.Z.n32 0.0474438
R442 CDAC8_0.switch_7.Z.n31 CDAC8_0.switch_7.Z.n30 0.0474438
R443 CDAC8_0.switch_7.Z.n29 CDAC8_0.switch_7.Z.n28 0.0474438
R444 CDAC8_0.switch_7.Z.n27 CDAC8_0.switch_7.Z.n13 0.0474438
R445 CDAC8_0.switch_7.Z.n12 CDAC8_0.switch_7.Z.n3 0.0474438
R446 CDAC8_0.switch_7.Z.n294 CDAC8_0.switch_7.Z.n293 0.0474438
R447 CDAC8_0.switch_7.Z.n8 CDAC8_0.switch_7.Z.n4 0.0474438
R448 CDAC8_0.switch_7.Z.n239 CDAC8_0.switch_7.Z.n238 0.0474438
R449 CDAC8_0.switch_7.Z.n241 CDAC8_0.switch_7.Z.n240 0.0474438
R450 CDAC8_0.switch_7.Z.n243 CDAC8_0.switch_7.Z.n242 0.0474438
R451 CDAC8_0.switch_7.Z.n245 CDAC8_0.switch_7.Z.n244 0.0474438
R452 CDAC8_0.switch_7.Z.n247 CDAC8_0.switch_7.Z.n246 0.0474438
R453 CDAC8_0.switch_7.Z.n249 CDAC8_0.switch_7.Z.n248 0.0474438
R454 CDAC8_0.switch_7.Z.n154 CDAC8_0.switch_7.Z.n153 0.0474438
R455 CDAC8_0.switch_7.Z.n152 CDAC8_0.switch_7.Z.n151 0.0474438
R456 CDAC8_0.switch_7.Z.n150 CDAC8_0.switch_7.Z.n149 0.0474438
R457 CDAC8_0.switch_7.Z.n148 CDAC8_0.switch_7.Z.n147 0.0474438
R458 CDAC8_0.switch_7.Z.n146 CDAC8_0.switch_7.Z.n145 0.0474438
R459 CDAC8_0.switch_7.Z.n185 CDAC8_0.switch_7.Z.n119 0.0474438
R460 CDAC8_0.switch_7.Z.n187 CDAC8_0.switch_7.Z.n186 0.0474438
R461 CDAC8_0.switch_7.Z.n198 CDAC8_0.switch_7.Z.n103 0.0474438
R462 CDAC8_0.switch_7.Z.n200 CDAC8_0.switch_7.Z.n199 0.0474438
R463 CDAC8_0.switch_7.Z.n202 CDAC8_0.switch_7.Z.n201 0.0474438
R464 CDAC8_0.switch_7.Z.n204 CDAC8_0.switch_7.Z.n203 0.0474438
R465 CDAC8_0.switch_7.Z.n206 CDAC8_0.switch_7.Z.n205 0.0474438
R466 CDAC8_0.switch_7.Z.n208 CDAC8_0.switch_7.Z.n207 0.0474438
R467 CDAC8_0.switch_7.Z.n210 CDAC8_0.switch_7.Z.n209 0.0474438
R468 CDAC8_0.switch_7.Z.n163 CDAC8_0.switch_7.Z.n131 0.0474438
R469 CDAC8_0.switch_7.Z.n165 CDAC8_0.switch_7.Z.n164 0.0474438
R470 CDAC8_0.switch_7.Z.n171 CDAC8_0.switch_7.Z.n127 0.0474438
R471 CDAC8_0.switch_7.Z.n173 CDAC8_0.switch_7.Z.n172 0.0474438
R472 CDAC8_0.switch_7.Z.n180 CDAC8_0.switch_7.Z.n123 0.0474438
R473 CDAC8_0.switch_7.Z.n182 CDAC8_0.switch_7.Z.n181 0.0474438
R474 CDAC8_0.switch_7.Z.n193 CDAC8_0.switch_7.Z.n116 0.0474438
R475 CDAC8_0.switch_7.Z.n195 CDAC8_0.switch_7.Z.n194 0.0474438
R476 CDAC8_0.switch_7.Z.n232 CDAC8_0.switch_7.Z.n93 0.0474438
R477 CDAC8_0.switch_7.Z.n231 CDAC8_0.switch_7.Z.n230 0.0474438
R478 CDAC8_0.switch_7.Z.n224 CDAC8_0.switch_7.Z.n94 0.0474438
R479 CDAC8_0.switch_7.Z.n223 CDAC8_0.switch_7.Z.n222 0.0474438
R480 CDAC8_0.switch_7.Z.n216 CDAC8_0.switch_7.Z.n98 0.0474438
R481 CDAC8_0.switch_7.Z.n215 CDAC8_0.switch_7.Z.n214 0.0474438
R482 CDAC8_0.switch_7.Z.n143 CDAC8_0.switch_7.Z.n142 0.0474438
R483 CDAC8_0.switch_7.Z.n141 CDAC8_0.switch_7.Z.n140 0.0474438
R484 CDAC8_0.switch_7.Z.n139 CDAC8_0.switch_7.Z.n138 0.0474438
R485 CDAC8_0.switch_7.Z.n137 CDAC8_0.switch_7.Z.n136 0.0474438
R486 CDAC8_0.switch_7.Z.n135 CDAC8_0.switch_7.Z.n134 0.0474438
R487 CDAC8_0.switch_7.Z.n133 CDAC8_0.switch_7.Z.n121 0.0474438
R488 CDAC8_0.switch_7.Z.n120 CDAC8_0.switch_7.Z.n118 0.0474438
R489 CDAC8_0.switch_7.Z.n117 CDAC8_0.switch_7.Z.n115 0.0474438
R490 CDAC8_0.switch_7.Z.n114 CDAC8_0.switch_7.Z.n113 0.0474438
R491 CDAC8_0.switch_7.Z.n112 CDAC8_0.switch_7.Z.n111 0.0474438
R492 CDAC8_0.switch_7.Z.n110 CDAC8_0.switch_7.Z.n109 0.0474438
R493 CDAC8_0.switch_7.Z.n108 CDAC8_0.switch_7.Z.n107 0.0474438
R494 CDAC8_0.switch_7.Z.n106 CDAC8_0.switch_7.Z.n105 0.0474438
R495 CDAC8_0.switch_7.Z.n104 CDAC8_0.switch_7.Z.n102 0.0474438
R496 CDAC8_0.switch_7.Z.n161 CDAC8_0.switch_7.Z.n160 0.0474438
R497 CDAC8_0.switch_7.Z.n167 CDAC8_0.switch_7.Z.n129 0.0474438
R498 CDAC8_0.switch_7.Z.n169 CDAC8_0.switch_7.Z.n168 0.0474438
R499 CDAC8_0.switch_7.Z.n175 CDAC8_0.switch_7.Z.n125 0.0474438
R500 CDAC8_0.switch_7.Z.n178 CDAC8_0.switch_7.Z.n176 0.0474438
R501 CDAC8_0.switch_7.Z.n177 CDAC8_0.switch_7.Z.n122 0.0474438
R502 CDAC8_0.switch_7.Z.n191 CDAC8_0.switch_7.Z.n189 0.0474438
R503 CDAC8_0.switch_7.Z.n190 CDAC8_0.switch_7.Z.n90 0.0474438
R504 CDAC8_0.switch_7.Z.n235 CDAC8_0.switch_7.Z.n234 0.0474438
R505 CDAC8_0.switch_7.Z.n228 CDAC8_0.switch_7.Z.n91 0.0474438
R506 CDAC8_0.switch_7.Z.n227 CDAC8_0.switch_7.Z.n226 0.0474438
R507 CDAC8_0.switch_7.Z.n220 CDAC8_0.switch_7.Z.n96 0.0474438
R508 CDAC8_0.switch_7.Z.n219 CDAC8_0.switch_7.Z.n218 0.0474438
R509 CDAC8_0.switch_7.Z.n212 CDAC8_0.switch_7.Z.n100 0.0474438
R510 CDAC8_0.switch_7.Z CDAC8_0.switch_7.Z.n297 0.0454219
R511 CDAC8_0.switch_7.Z.n295 CDAC8_0.switch_7.Z.n3 0.0314031
R512 CDAC8_0.switch_7.Z.n237 CDAC8_0.switch_7.Z.n8 0.0314031
R513 CDAC8_0.switch_7.Z.n122 CDAC8_0.switch_7.Z.n2 0.0314031
R514 CDAC8_0.switch_7.Z.n236 CDAC8_0.switch_7.Z.n90 0.0314031
R515 CDAC8_0.switch_7.Z.n1 CDAC8_0.switch_7.Z.n0 0.0188121
R516 EN.n61 EN.t56 158.988
R517 EN.n155 EN.t42 158.988
R518 EN EN.t13 158.581
R519 EN EN.t21 158.581
R520 EN EN.t88 158.581
R521 EN EN.t77 158.581
R522 EN EN.t9 158.581
R523 EN EN.t96 158.581
R524 EN EN.t36 158.581
R525 EN EN.t60 158.581
R526 EN EN.t35 158.581
R527 EN EN.t76 158.581
R528 EN EN.t39 158.581
R529 EN EN.t81 158.581
R530 EN EN.t79 158.581
R531 EN EN.t37 158.581
R532 EN EN.t40 158.581
R533 EN EN.t98 158.581
R534 EN.n69 EN.t6 150.293
R535 EN.n63 EN.t61 150.293
R536 EN.n145 EN.t10 150.293
R537 EN.n139 EN.t12 150.293
R538 EN.t13 EN.n181 150.293
R539 EN.t21 EN.n212 150.293
R540 EN.t88 EN.n221 150.293
R541 EN.t77 EN.n135 150.293
R542 EN.t9 EN.n244 150.293
R543 EN.t96 EN.n274 150.293
R544 EN.t36 EN.n284 150.293
R545 EN.t60 EN.n97 150.293
R546 EN.t35 EN.n106 150.293
R547 EN.t76 EN.n318 150.293
R548 EN.t39 EN.n327 150.293
R549 EN.t81 EN.n33 150.293
R550 EN.t79 EN.n350 150.293
R551 EN.t37 EN.n163 150.293
R552 EN.t40 EN.n52 150.293
R553 EN.t98 EN.n5 150.293
R554 EN.t56 EN.n60 150.273
R555 EN.t42 EN.n154 150.273
R556 EN.n186 EN.t50 150.273
R557 EN.n176 EN.t94 150.273
R558 EN.n205 EN.t71 150.273
R559 EN.n199 EN.t104 150.273
R560 EN.n226 EN.t23 150.273
R561 EN.n216 EN.t15 150.273
R562 EN.n128 EN.t89 150.273
R563 EN.n122 EN.t25 150.273
R564 EN.n249 EN.t47 150.273
R565 EN.n239 EN.t72 150.273
R566 EN.n267 EN.t46 150.273
R567 EN.n261 EN.t80 150.273
R568 EN.n289 EN.t97 150.273
R569 EN.n279 EN.t90 150.273
R570 EN.n90 EN.t66 150.273
R571 EN.n84 EN.t45 150.273
R572 EN.n111 EN.t18 150.273
R573 EN.n101 EN.t11 150.273
R574 EN.n311 EN.t17 150.273
R575 EN.n305 EN.t55 150.273
R576 EN.n332 EN.t92 150.273
R577 EN.n322 EN.t67 150.273
R578 EN.n26 EN.t29 150.273
R579 EN.n20 EN.t106 150.273
R580 EN.n355 EN.t14 150.273
R581 EN.n345 EN.t75 150.273
R582 EN.n168 EN.t101 150.273
R583 EN.n158 EN.t93 150.273
R584 EN.n45 EN.t49 150.273
R585 EN.n39 EN.t26 150.273
R586 EN.n10 EN.t38 150.273
R587 EN.n0 EN.t16 150.273
R588 EN.n194 EN.t1 115.191
R589 EN.n234 EN.t91 81.8568
R590 EN.n257 EN.t48 81.8568
R591 EN.n297 EN.t69 81.8568
R592 EN.n300 EN.t19 81.8568
R593 EN.n340 EN.t44 81.8568
R594 EN.n363 EN.t53 81.8568
R595 EN.n195 EN.t73 81.8568
R596 EN.t105 EN.n365 81.8568
R597 EN.n58 EN.t41 73.6406
R598 EN.n152 EN.t20 73.6406
R599 EN.n184 EN.t57 73.6406
R600 EN.t1 EN.n193 73.6406
R601 EN.n203 EN.t58 73.6406
R602 EN.n197 EN.t85 73.6406
R603 EN.n224 EN.t28 73.6406
R604 EN.t91 EN.n233 73.6406
R605 EN.n126 EN.t0 73.6406
R606 EN.n120 EN.t4 73.6406
R607 EN.n247 EN.t82 73.6406
R608 EN.t48 EN.n256 73.6406
R609 EN.n265 EN.t31 73.6406
R610 EN.n259 EN.t63 73.6406
R611 EN.n287 EN.t99 73.6406
R612 EN.t69 EN.n296 73.6406
R613 EN.n88 EN.t83 73.6406
R614 EN.n82 EN.t27 73.6406
R615 EN.n109 EN.t22 73.6406
R616 EN.t19 EN.n118 73.6406
R617 EN.n309 EN.t100 73.6406
R618 EN.n303 EN.t68 73.6406
R619 EN.n330 EN.t78 73.6406
R620 EN.t44 EN.n339 73.6406
R621 EN.n24 EN.t8 73.6406
R622 EN.n18 EN.t86 73.6406
R623 EN.n353 EN.t30 73.6406
R624 EN.t53 EN.n362 73.6406
R625 EN.n166 EN.t107 73.6406
R626 EN.t73 EN.n175 73.6406
R627 EN.n43 EN.t64 73.6406
R628 EN.n37 EN.t7 73.6406
R629 EN.n8 EN.t74 73.6406
R630 EN.n366 EN.t105 73.6406
R631 EN.n71 EN.t43 73.6304
R632 EN.n65 EN.t87 73.6304
R633 EN.n147 EN.t62 73.6304
R634 EN.n141 EN.t95 73.6304
R635 EN.n179 EN.t59 73.6304
R636 EN.n210 EN.t2 73.6304
R637 EN.n219 EN.t33 73.6304
R638 EN.n133 EN.t32 73.6304
R639 EN.n242 EN.t52 73.6304
R640 EN.n272 EN.t51 73.6304
R641 EN.n282 EN.t103 73.6304
R642 EN.n95 EN.t102 73.6304
R643 EN.n104 EN.t70 73.6304
R644 EN.n316 EN.t24 73.6304
R645 EN.n325 EN.t5 73.6304
R646 EN.n31 EN.t65 73.6304
R647 EN.n348 EN.t34 73.6304
R648 EN.n161 EN.t3 73.6304
R649 EN.n50 EN.t84 73.6304
R650 EN.n3 EN.t54 73.6304
R651 EN.n365 EN.n364 33.3344
R652 EN.n236 EN.n196 33.3344
R653 EN.n343 EN.n80 33.3344
R654 EN.n364 EN.n17 29.9244
R655 EN.n299 EN.n17 29.9244
R656 EN.n299 EN.n298 29.9244
R657 EN.n298 EN.n258 29.9244
R658 EN.n258 EN.n119 29.9244
R659 EN.n194 EN.n119 29.9244
R660 EN.n237 EN.n236 29.9244
R661 EN.n237 EN.n81 29.9244
R662 EN.n302 EN.n81 29.9244
R663 EN.n342 EN.n302 29.9244
R664 EN.n343 EN.n342 29.9244
R665 EN.n235 EN.n234 25.7228
R666 EN.n257 EN.n238 25.7228
R667 EN.n297 EN.n278 25.7228
R668 EN.n301 EN.n300 25.7228
R669 EN.n341 EN.n340 25.7228
R670 EN.n363 EN.n344 25.7228
R671 EN.n196 EN.n195 25.7228
R672 EN.n79 EN 23.3453
R673 EN.n77 EN.n76 20.9244
R674 EN.n75 EN.n68 15.5222
R675 EN.n151 EN.n144 15.5222
R676 EN.n191 EN.n190 15.5222
R677 EN.n209 EN.n202 15.5222
R678 EN.n231 EN.n230 15.5222
R679 EN.n132 EN.n125 15.5222
R680 EN.n254 EN.n253 15.5222
R681 EN.n271 EN.n264 15.5222
R682 EN.n294 EN.n293 15.5222
R683 EN.n94 EN.n87 15.5222
R684 EN.n116 EN.n115 15.5222
R685 EN.n315 EN.n308 15.5222
R686 EN.n337 EN.n336 15.5222
R687 EN.n30 EN.n23 15.5222
R688 EN.n360 EN.n359 15.5222
R689 EN.n173 EN.n172 15.5222
R690 EN.n49 EN.n42 15.5222
R691 EN.n15 EN.n14 15.5222
R692 EN.n78 EN 12.9568
R693 EN.n57 EN.n56 12.8934
R694 EN.n79 EN.n78 12.7234
R695 EN.n57 EN 10.1822
R696 EN.n190 EN.n183 8.26552
R697 EN.n230 EN.n223 8.26552
R698 EN.n253 EN.n246 8.26552
R699 EN.n293 EN.n286 8.26552
R700 EN.n115 EN.n108 8.26552
R701 EN.n336 EN.n329 8.26552
R702 EN.n359 EN.n352 8.26552
R703 EN.n172 EN.n165 8.26552
R704 EN.n14 EN.n7 8.26552
R705 EN.n76 EN.n75 7.83713
R706 EN.n235 EN.n215 5.58033
R707 EN.n238 EN.n138 5.58033
R708 EN.n278 EN.n277 5.58033
R709 EN.n301 EN.n100 5.58033
R710 EN.n341 EN.n321 5.58033
R711 EN.n344 EN.n36 5.58033
R712 EN.n80 EN.n55 5.58033
R713 EN.n75 EN.n74 4.5005
R714 EN.n151 EN.n150 4.5005
R715 EN.n190 EN.n189 4.5005
R716 EN.n209 EN.n208 4.5005
R717 EN.n230 EN.n229 4.5005
R718 EN.n132 EN.n131 4.5005
R719 EN.n253 EN.n252 4.5005
R720 EN.n271 EN.n270 4.5005
R721 EN.n293 EN.n292 4.5005
R722 EN.n94 EN.n93 4.5005
R723 EN.n115 EN.n114 4.5005
R724 EN.n315 EN.n314 4.5005
R725 EN.n336 EN.n335 4.5005
R726 EN.n30 EN.n29 4.5005
R727 EN.n359 EN.n358 4.5005
R728 EN.n172 EN.n171 4.5005
R729 EN.n49 EN.n48 4.5005
R730 EN.n14 EN.n13 4.5005
R731 EN.n196 EN.n157 4.31133
R732 EN.n215 EN.n214 4.20846
R733 EN.n138 EN.n137 4.20846
R734 EN.n277 EN.n276 4.20846
R735 EN.n100 EN.n99 4.20846
R736 EN.n321 EN.n320 4.20846
R737 EN.n36 EN.n35 4.20846
R738 EN.n55 EN.n54 4.20846
R739 EN.n157 EN.n151 3.98148
R740 EN.n215 EN.n209 3.98148
R741 EN.n138 EN.n132 3.98148
R742 EN.n277 EN.n271 3.98148
R743 EN.n100 EN.n94 3.98148
R744 EN.n321 EN.n315 3.98148
R745 EN.n36 EN.n30 3.98148
R746 EN.n55 EN.n49 3.98148
R747 EN.n157 EN 3.8
R748 EN.n364 EN.n363 3.4105
R749 EN.n340 EN.n17 3.4105
R750 EN.n300 EN.n299 3.4105
R751 EN.n298 EN.n297 3.4105
R752 EN.n258 EN.n257 3.4105
R753 EN.n234 EN.n119 3.4105
R754 EN.n195 EN.n194 3.4105
R755 EN.n236 EN.n235 3.4105
R756 EN.n238 EN.n237 3.4105
R757 EN.n278 EN.n81 3.4105
R758 EN.n302 EN.n301 3.4105
R759 EN.n342 EN.n341 3.4105
R760 EN.n344 EN.n343 3.4105
R761 EN.n59 EN.n58 1.19615
R762 EN.n153 EN.n152 1.19615
R763 EN.n181 EN.n180 1.19615
R764 EN.n212 EN.n211 1.19615
R765 EN.n221 EN.n220 1.19615
R766 EN.n135 EN.n134 1.19615
R767 EN.n244 EN.n243 1.19615
R768 EN.n274 EN.n273 1.19615
R769 EN.n284 EN.n283 1.19615
R770 EN.n97 EN.n96 1.19615
R771 EN.n106 EN.n105 1.19615
R772 EN.n318 EN.n317 1.19615
R773 EN.n327 EN.n326 1.19615
R774 EN.n33 EN.n32 1.19615
R775 EN.n350 EN.n349 1.19615
R776 EN.n163 EN.n162 1.19615
R777 EN.n52 EN.n51 1.19615
R778 EN.n5 EN.n4 1.19615
R779 EN.n70 EN 1.09561
R780 EN.n64 EN 1.09561
R781 EN.n146 EN 1.09561
R782 EN.n140 EN 1.09561
R783 EN.n73 EN.n72 0.796696
R784 EN.n67 EN.n66 0.796696
R785 EN.n149 EN.n148 0.796696
R786 EN.n143 EN.n142 0.796696
R787 EN.n185 EN.n184 0.796696
R788 EN.n193 EN.n192 0.796696
R789 EN.n204 EN.n203 0.796696
R790 EN.n198 EN.n197 0.796696
R791 EN.n225 EN.n224 0.796696
R792 EN.n233 EN.n232 0.796696
R793 EN.n127 EN.n126 0.796696
R794 EN.n121 EN.n120 0.796696
R795 EN.n248 EN.n247 0.796696
R796 EN.n256 EN.n255 0.796696
R797 EN.n266 EN.n265 0.796696
R798 EN.n260 EN.n259 0.796696
R799 EN.n288 EN.n287 0.796696
R800 EN.n296 EN.n295 0.796696
R801 EN.n89 EN.n88 0.796696
R802 EN.n83 EN.n82 0.796696
R803 EN.n110 EN.n109 0.796696
R804 EN.n118 EN.n117 0.796696
R805 EN.n310 EN.n309 0.796696
R806 EN.n304 EN.n303 0.796696
R807 EN.n331 EN.n330 0.796696
R808 EN.n339 EN.n338 0.796696
R809 EN.n25 EN.n24 0.796696
R810 EN.n19 EN.n18 0.796696
R811 EN.n354 EN.n353 0.796696
R812 EN.n362 EN.n361 0.796696
R813 EN.n167 EN.n166 0.796696
R814 EN.n175 EN.n174 0.796696
R815 EN.n44 EN.n43 0.796696
R816 EN.n38 EN.n37 0.796696
R817 EN.n9 EN.n8 0.796696
R818 EN.n366 EN.n16 0.796696
R819 EN.n62 EN.n61 0.783833
R820 EN.n156 EN.n155 0.783833
R821 EN.n183 EN.n182 0.783833
R822 EN.n214 EN.n213 0.783833
R823 EN.n223 EN.n222 0.783833
R824 EN.n137 EN.n136 0.783833
R825 EN.n246 EN.n245 0.783833
R826 EN.n276 EN.n275 0.783833
R827 EN.n286 EN.n285 0.783833
R828 EN.n99 EN.n98 0.783833
R829 EN.n108 EN.n107 0.783833
R830 EN.n320 EN.n319 0.783833
R831 EN.n329 EN.n328 0.783833
R832 EN.n35 EN.n34 0.783833
R833 EN.n352 EN.n351 0.783833
R834 EN.n165 EN.n164 0.783833
R835 EN.n54 EN.n53 0.783833
R836 EN.n7 EN.n6 0.783833
R837 EN.n61 EN 0.716182
R838 EN.n155 EN 0.716182
R839 EN.n183 EN 0.716182
R840 EN.n214 EN 0.716182
R841 EN.n223 EN 0.716182
R842 EN.n137 EN 0.716182
R843 EN.n246 EN 0.716182
R844 EN.n276 EN 0.716182
R845 EN.n286 EN 0.716182
R846 EN.n99 EN 0.716182
R847 EN.n108 EN 0.716182
R848 EN.n320 EN 0.716182
R849 EN.n329 EN 0.716182
R850 EN.n35 EN 0.716182
R851 EN.n352 EN 0.716182
R852 EN.n165 EN 0.716182
R853 EN.n54 EN 0.716182
R854 EN.n7 EN 0.716182
R855 EN.n73 EN 0.662609
R856 EN.n67 EN 0.662609
R857 EN.n149 EN 0.662609
R858 EN.n143 EN 0.662609
R859 EN.n185 EN 0.524957
R860 EN.n192 EN 0.524957
R861 EN.n204 EN 0.524957
R862 EN.n198 EN 0.524957
R863 EN.n225 EN 0.524957
R864 EN.n232 EN 0.524957
R865 EN.n127 EN 0.524957
R866 EN.n121 EN 0.524957
R867 EN.n248 EN 0.524957
R868 EN.n255 EN 0.524957
R869 EN.n266 EN 0.524957
R870 EN.n260 EN 0.524957
R871 EN.n288 EN 0.524957
R872 EN.n295 EN 0.524957
R873 EN.n89 EN 0.524957
R874 EN.n83 EN 0.524957
R875 EN.n110 EN 0.524957
R876 EN.n117 EN 0.524957
R877 EN.n310 EN 0.524957
R878 EN.n304 EN 0.524957
R879 EN.n331 EN 0.524957
R880 EN.n338 EN 0.524957
R881 EN.n25 EN 0.524957
R882 EN.n19 EN 0.524957
R883 EN.n354 EN 0.524957
R884 EN.n361 EN 0.524957
R885 EN.n167 EN 0.524957
R886 EN.n174 EN 0.524957
R887 EN.n44 EN 0.524957
R888 EN.n38 EN 0.524957
R889 EN.n9 EN 0.524957
R890 EN.n16 EN 0.524957
R891 EN.n69 EN 0.447191
R892 EN.n63 EN 0.447191
R893 EN.n145 EN 0.447191
R894 EN.n139 EN 0.447191
R895 EN.n181 EN 0.447191
R896 EN.n212 EN 0.447191
R897 EN.n221 EN 0.447191
R898 EN.n135 EN 0.447191
R899 EN.n244 EN 0.447191
R900 EN.n274 EN 0.447191
R901 EN.n284 EN 0.447191
R902 EN.n97 EN 0.447191
R903 EN.n106 EN 0.447191
R904 EN.n318 EN 0.447191
R905 EN.n327 EN 0.447191
R906 EN.n33 EN 0.447191
R907 EN.n350 EN 0.447191
R908 EN.n163 EN 0.447191
R909 EN.n52 EN 0.447191
R910 EN.n5 EN 0.447191
R911 EN.n188 EN 0.252453
R912 EN.n178 EN 0.252453
R913 EN.n207 EN 0.252453
R914 EN.n201 EN 0.252453
R915 EN.n228 EN 0.252453
R916 EN.n218 EN 0.252453
R917 EN.n130 EN 0.252453
R918 EN.n124 EN 0.252453
R919 EN.n251 EN 0.252453
R920 EN.n241 EN 0.252453
R921 EN.n269 EN 0.252453
R922 EN.n263 EN 0.252453
R923 EN.n291 EN 0.252453
R924 EN.n281 EN 0.252453
R925 EN.n92 EN 0.252453
R926 EN.n86 EN 0.252453
R927 EN.n113 EN 0.252453
R928 EN.n103 EN 0.252453
R929 EN.n313 EN 0.252453
R930 EN.n307 EN 0.252453
R931 EN.n334 EN 0.252453
R932 EN.n324 EN 0.252453
R933 EN.n28 EN 0.252453
R934 EN.n22 EN 0.252453
R935 EN.n357 EN 0.252453
R936 EN.n347 EN 0.252453
R937 EN.n170 EN 0.252453
R938 EN.n160 EN 0.252453
R939 EN.n47 EN 0.252453
R940 EN.n41 EN 0.252453
R941 EN.n12 EN 0.252453
R942 EN.n2 EN 0.252453
R943 EN.n70 EN.n69 0.226043
R944 EN.n64 EN.n63 0.226043
R945 EN.n146 EN.n145 0.226043
R946 EN.n140 EN.n139 0.226043
R947 EN.n188 EN.n187 0.226043
R948 EN.n178 EN.n177 0.226043
R949 EN.n207 EN.n206 0.226043
R950 EN.n201 EN.n200 0.226043
R951 EN.n228 EN.n227 0.226043
R952 EN.n218 EN.n217 0.226043
R953 EN.n130 EN.n129 0.226043
R954 EN.n124 EN.n123 0.226043
R955 EN.n251 EN.n250 0.226043
R956 EN.n241 EN.n240 0.226043
R957 EN.n269 EN.n268 0.226043
R958 EN.n263 EN.n262 0.226043
R959 EN.n291 EN.n290 0.226043
R960 EN.n281 EN.n280 0.226043
R961 EN.n92 EN.n91 0.226043
R962 EN.n86 EN.n85 0.226043
R963 EN.n113 EN.n112 0.226043
R964 EN.n103 EN.n102 0.226043
R965 EN.n313 EN.n312 0.226043
R966 EN.n307 EN.n306 0.226043
R967 EN.n334 EN.n333 0.226043
R968 EN.n324 EN.n323 0.226043
R969 EN.n28 EN.n27 0.226043
R970 EN.n22 EN.n21 0.226043
R971 EN.n357 EN.n356 0.226043
R972 EN.n347 EN.n346 0.226043
R973 EN.n170 EN.n169 0.226043
R974 EN.n160 EN.n159 0.226043
R975 EN.n47 EN.n46 0.226043
R976 EN.n41 EN.n40 0.226043
R977 EN.n12 EN.n11 0.226043
R978 EN.n2 EN.n1 0.226043
R979 EN.n58 EN 0.217464
R980 EN.n152 EN 0.217464
R981 EN.n184 EN 0.217464
R982 EN.n193 EN 0.217464
R983 EN.n203 EN 0.217464
R984 EN.n197 EN 0.217464
R985 EN.n224 EN 0.217464
R986 EN.n233 EN 0.217464
R987 EN.n126 EN 0.217464
R988 EN.n120 EN 0.217464
R989 EN.n247 EN 0.217464
R990 EN.n256 EN 0.217464
R991 EN.n265 EN 0.217464
R992 EN.n259 EN 0.217464
R993 EN.n287 EN 0.217464
R994 EN.n296 EN 0.217464
R995 EN.n88 EN 0.217464
R996 EN.n82 EN 0.217464
R997 EN.n109 EN 0.217464
R998 EN.n118 EN 0.217464
R999 EN.n309 EN 0.217464
R1000 EN.n303 EN 0.217464
R1001 EN.n330 EN 0.217464
R1002 EN.n339 EN 0.217464
R1003 EN.n24 EN 0.217464
R1004 EN.n18 EN 0.217464
R1005 EN.n353 EN 0.217464
R1006 EN.n362 EN 0.217464
R1007 EN.n166 EN 0.217464
R1008 EN.n175 EN 0.217464
R1009 EN.n43 EN 0.217464
R1010 EN.n37 EN 0.217464
R1011 EN.n8 EN 0.217464
R1012 EN EN.n366 0.217464
R1013 EN.n72 EN 0.1255
R1014 EN.n66 EN 0.1255
R1015 EN.n59 EN 0.1255
R1016 EN.n153 EN 0.1255
R1017 EN.n148 EN 0.1255
R1018 EN.n142 EN 0.1255
R1019 EN.n187 EN 0.1255
R1020 EN.n180 EN 0.1255
R1021 EN.n177 EN 0.1255
R1022 EN.n211 EN 0.1255
R1023 EN.n206 EN 0.1255
R1024 EN.n200 EN 0.1255
R1025 EN.n227 EN 0.1255
R1026 EN.n220 EN 0.1255
R1027 EN.n217 EN 0.1255
R1028 EN.n134 EN 0.1255
R1029 EN.n129 EN 0.1255
R1030 EN.n123 EN 0.1255
R1031 EN.n250 EN 0.1255
R1032 EN.n243 EN 0.1255
R1033 EN.n240 EN 0.1255
R1034 EN.n273 EN 0.1255
R1035 EN.n268 EN 0.1255
R1036 EN.n262 EN 0.1255
R1037 EN.n290 EN 0.1255
R1038 EN.n283 EN 0.1255
R1039 EN.n280 EN 0.1255
R1040 EN.n96 EN 0.1255
R1041 EN.n91 EN 0.1255
R1042 EN.n85 EN 0.1255
R1043 EN.n112 EN 0.1255
R1044 EN.n105 EN 0.1255
R1045 EN.n102 EN 0.1255
R1046 EN.n317 EN 0.1255
R1047 EN.n312 EN 0.1255
R1048 EN.n306 EN 0.1255
R1049 EN.n333 EN 0.1255
R1050 EN.n326 EN 0.1255
R1051 EN.n323 EN 0.1255
R1052 EN.n32 EN 0.1255
R1053 EN.n27 EN 0.1255
R1054 EN.n21 EN 0.1255
R1055 EN.n356 EN 0.1255
R1056 EN.n349 EN 0.1255
R1057 EN.n346 EN 0.1255
R1058 EN.n169 EN 0.1255
R1059 EN.n162 EN 0.1255
R1060 EN.n159 EN 0.1255
R1061 EN.n51 EN 0.1255
R1062 EN.n46 EN 0.1255
R1063 EN.n40 EN 0.1255
R1064 EN.n11 EN 0.1255
R1065 EN.n4 EN 0.1255
R1066 EN.n1 EN 0.1255
R1067 EN.n74 EN.n70 0.063
R1068 EN.n74 EN.n73 0.063
R1069 EN.n68 EN.n64 0.063
R1070 EN.n68 EN.n67 0.063
R1071 EN.n150 EN.n146 0.063
R1072 EN.n150 EN.n149 0.063
R1073 EN.n144 EN.n140 0.063
R1074 EN.n144 EN.n143 0.063
R1075 EN.n189 EN.n185 0.063
R1076 EN.n189 EN.n188 0.063
R1077 EN.n192 EN.n191 0.063
R1078 EN.n191 EN.n178 0.063
R1079 EN.n208 EN.n204 0.063
R1080 EN.n208 EN.n207 0.063
R1081 EN.n202 EN.n198 0.063
R1082 EN.n202 EN.n201 0.063
R1083 EN.n229 EN.n225 0.063
R1084 EN.n229 EN.n228 0.063
R1085 EN.n232 EN.n231 0.063
R1086 EN.n231 EN.n218 0.063
R1087 EN.n131 EN.n127 0.063
R1088 EN.n131 EN.n130 0.063
R1089 EN.n125 EN.n121 0.063
R1090 EN.n125 EN.n124 0.063
R1091 EN.n252 EN.n248 0.063
R1092 EN.n252 EN.n251 0.063
R1093 EN.n255 EN.n254 0.063
R1094 EN.n254 EN.n241 0.063
R1095 EN.n270 EN.n266 0.063
R1096 EN.n270 EN.n269 0.063
R1097 EN.n264 EN.n260 0.063
R1098 EN.n264 EN.n263 0.063
R1099 EN.n292 EN.n288 0.063
R1100 EN.n292 EN.n291 0.063
R1101 EN.n295 EN.n294 0.063
R1102 EN.n294 EN.n281 0.063
R1103 EN.n93 EN.n89 0.063
R1104 EN.n93 EN.n92 0.063
R1105 EN.n87 EN.n83 0.063
R1106 EN.n87 EN.n86 0.063
R1107 EN.n114 EN.n110 0.063
R1108 EN.n114 EN.n113 0.063
R1109 EN.n117 EN.n116 0.063
R1110 EN.n116 EN.n103 0.063
R1111 EN.n314 EN.n310 0.063
R1112 EN.n314 EN.n313 0.063
R1113 EN.n308 EN.n304 0.063
R1114 EN.n308 EN.n307 0.063
R1115 EN.n335 EN.n331 0.063
R1116 EN.n335 EN.n334 0.063
R1117 EN.n338 EN.n337 0.063
R1118 EN.n337 EN.n324 0.063
R1119 EN.n29 EN.n25 0.063
R1120 EN.n29 EN.n28 0.063
R1121 EN.n23 EN.n19 0.063
R1122 EN.n23 EN.n22 0.063
R1123 EN.n358 EN.n354 0.063
R1124 EN.n358 EN.n357 0.063
R1125 EN.n361 EN.n360 0.063
R1126 EN.n360 EN.n347 0.063
R1127 EN.n171 EN.n167 0.063
R1128 EN.n171 EN.n170 0.063
R1129 EN.n174 EN.n173 0.063
R1130 EN.n173 EN.n160 0.063
R1131 EN.n48 EN.n44 0.063
R1132 EN.n48 EN.n47 0.063
R1133 EN.n42 EN.n38 0.063
R1134 EN.n42 EN.n41 0.063
R1135 EN.n13 EN.n9 0.063
R1136 EN.n13 EN.n12 0.063
R1137 EN.n16 EN.n15 0.063
R1138 EN.n15 EN.n2 0.063
R1139 EN.n80 EN.n79 0.024
R1140 EN.n78 EN.n77 0.024
R1141 EN.n77 EN.n57 0.024
R1142 EN.n60 EN.n59 0.0216397
R1143 EN.n60 EN 0.0216397
R1144 EN.n154 EN.n153 0.0216397
R1145 EN.n154 EN 0.0216397
R1146 EN.n187 EN.n186 0.0216397
R1147 EN.n186 EN 0.0216397
R1148 EN.n177 EN.n176 0.0216397
R1149 EN.n176 EN 0.0216397
R1150 EN.n206 EN.n205 0.0216397
R1151 EN.n205 EN 0.0216397
R1152 EN.n200 EN.n199 0.0216397
R1153 EN.n199 EN 0.0216397
R1154 EN.n227 EN.n226 0.0216397
R1155 EN.n226 EN 0.0216397
R1156 EN.n217 EN.n216 0.0216397
R1157 EN.n216 EN 0.0216397
R1158 EN.n129 EN.n128 0.0216397
R1159 EN.n128 EN 0.0216397
R1160 EN.n123 EN.n122 0.0216397
R1161 EN.n122 EN 0.0216397
R1162 EN.n250 EN.n249 0.0216397
R1163 EN.n249 EN 0.0216397
R1164 EN.n240 EN.n239 0.0216397
R1165 EN.n239 EN 0.0216397
R1166 EN.n268 EN.n267 0.0216397
R1167 EN.n267 EN 0.0216397
R1168 EN.n262 EN.n261 0.0216397
R1169 EN.n261 EN 0.0216397
R1170 EN.n290 EN.n289 0.0216397
R1171 EN.n289 EN 0.0216397
R1172 EN.n280 EN.n279 0.0216397
R1173 EN.n279 EN 0.0216397
R1174 EN.n91 EN.n90 0.0216397
R1175 EN.n90 EN 0.0216397
R1176 EN.n85 EN.n84 0.0216397
R1177 EN.n84 EN 0.0216397
R1178 EN.n112 EN.n111 0.0216397
R1179 EN.n111 EN 0.0216397
R1180 EN.n102 EN.n101 0.0216397
R1181 EN.n101 EN 0.0216397
R1182 EN.n312 EN.n311 0.0216397
R1183 EN.n311 EN 0.0216397
R1184 EN.n306 EN.n305 0.0216397
R1185 EN.n305 EN 0.0216397
R1186 EN.n333 EN.n332 0.0216397
R1187 EN.n332 EN 0.0216397
R1188 EN.n323 EN.n322 0.0216397
R1189 EN.n322 EN 0.0216397
R1190 EN.n27 EN.n26 0.0216397
R1191 EN.n26 EN 0.0216397
R1192 EN.n21 EN.n20 0.0216397
R1193 EN.n20 EN 0.0216397
R1194 EN.n356 EN.n355 0.0216397
R1195 EN.n355 EN 0.0216397
R1196 EN.n346 EN.n345 0.0216397
R1197 EN.n345 EN 0.0216397
R1198 EN.n169 EN.n168 0.0216397
R1199 EN.n168 EN 0.0216397
R1200 EN.n159 EN.n158 0.0216397
R1201 EN.n158 EN 0.0216397
R1202 EN.n46 EN.n45 0.0216397
R1203 EN.n45 EN 0.0216397
R1204 EN.n40 EN.n39 0.0216397
R1205 EN.n39 EN 0.0216397
R1206 EN.n11 EN.n10 0.0216397
R1207 EN.n10 EN 0.0216397
R1208 EN.n1 EN.n0 0.0216397
R1209 EN.n0 EN 0.0216397
R1210 EN.n76 EN 0.0204394
R1211 EN.n365 EN 0.0204394
R1212 EN.n72 EN.n71 0.0107679
R1213 EN.n71 EN 0.0107679
R1214 EN.n66 EN.n65 0.0107679
R1215 EN.n65 EN 0.0107679
R1216 EN.n148 EN.n147 0.0107679
R1217 EN.n147 EN 0.0107679
R1218 EN.n142 EN.n141 0.0107679
R1219 EN.n141 EN 0.0107679
R1220 EN.n180 EN.n179 0.0107679
R1221 EN.n179 EN 0.0107679
R1222 EN.n211 EN.n210 0.0107679
R1223 EN.n210 EN 0.0107679
R1224 EN.n220 EN.n219 0.0107679
R1225 EN.n219 EN 0.0107679
R1226 EN.n134 EN.n133 0.0107679
R1227 EN.n133 EN 0.0107679
R1228 EN.n243 EN.n242 0.0107679
R1229 EN.n242 EN 0.0107679
R1230 EN.n273 EN.n272 0.0107679
R1231 EN.n272 EN 0.0107679
R1232 EN.n283 EN.n282 0.0107679
R1233 EN.n282 EN 0.0107679
R1234 EN.n96 EN.n95 0.0107679
R1235 EN.n95 EN 0.0107679
R1236 EN.n105 EN.n104 0.0107679
R1237 EN.n104 EN 0.0107679
R1238 EN.n317 EN.n316 0.0107679
R1239 EN.n316 EN 0.0107679
R1240 EN.n326 EN.n325 0.0107679
R1241 EN.n325 EN 0.0107679
R1242 EN.n32 EN.n31 0.0107679
R1243 EN.n31 EN 0.0107679
R1244 EN.n349 EN.n348 0.0107679
R1245 EN.n348 EN 0.0107679
R1246 EN.n162 EN.n161 0.0107679
R1247 EN.n161 EN 0.0107679
R1248 EN.n51 EN.n50 0.0107679
R1249 EN.n50 EN 0.0107679
R1250 EN.n4 EN.n3 0.0107679
R1251 EN.n3 EN 0.0107679
R1252 EN.n62 EN 0.00441667
R1253 EN.n156 EN 0.00441667
R1254 EN.n182 EN 0.00441667
R1255 EN.n213 EN 0.00441667
R1256 EN.n222 EN 0.00441667
R1257 EN.n136 EN 0.00441667
R1258 EN.n245 EN 0.00441667
R1259 EN.n275 EN 0.00441667
R1260 EN.n285 EN 0.00441667
R1261 EN.n98 EN 0.00441667
R1262 EN.n107 EN 0.00441667
R1263 EN.n319 EN 0.00441667
R1264 EN.n328 EN 0.00441667
R1265 EN.n34 EN 0.00441667
R1266 EN.n351 EN 0.00441667
R1267 EN.n164 EN 0.00441667
R1268 EN.n53 EN 0.00441667
R1269 EN.n56 EN 0.00441667
R1270 EN.n6 EN 0.00441667
R1271 EN EN.n62 0.00406061
R1272 EN EN.n156 0.00406061
R1273 EN.n182 EN 0.00406061
R1274 EN.n213 EN 0.00406061
R1275 EN.n222 EN 0.00406061
R1276 EN.n136 EN 0.00406061
R1277 EN.n245 EN 0.00406061
R1278 EN.n275 EN 0.00406061
R1279 EN.n285 EN 0.00406061
R1280 EN.n98 EN 0.00406061
R1281 EN.n107 EN 0.00406061
R1282 EN.n319 EN 0.00406061
R1283 EN.n328 EN 0.00406061
R1284 EN.n34 EN 0.00406061
R1285 EN.n351 EN 0.00406061
R1286 EN.n164 EN 0.00406061
R1287 EN.n53 EN 0.00406061
R1288 EN.n6 EN 0.00406061
R1289 EN.n56 EN 0.00406061
R1290 Vbias.n4899 Vbias.n4846 93853.1
R1291 Vbias.n4899 Vbias.n4893 93853.1
R1292 Vbias.n4895 Vbias.n4846 93853.1
R1293 Vbias.n7802 Vbias.n7801 49144.5
R1294 Vbias.n7937 Vbias.n7936 49144.5
R1295 Vbias.n7822 Vbias.n7821 45562.9
R1296 Vbias.n350 Vbias.n349 45562.9
R1297 Vbias.n7016 Vbias.n1339 45562.9
R1298 Vbias.n7015 Vbias.n1340 45562.9
R1299 Vbias.n5919 Vbias.n1638 45562.9
R1300 Vbias.n5918 Vbias.n1639 45562.9
R1301 Vbias.n5122 Vbias.n2370 45562.9
R1302 Vbias.n5121 Vbias.n2371 45562.9
R1303 Vbias.n4682 Vbias.n4550 45562.9
R1304 Vbias.n7225 Vbias.n7224 18472.2
R1305 Vbias.n4902 Vbias.n4901 17553.4
R1306 Vbias.n7871 Vbias.n7870 12551.1
R1307 Vbias.n7736 Vbias.n7735 12551.1
R1308 Vbias.n4685 Vbias.n4682 8982.04
R1309 Vbias.n7753 Vbias.n7752 8969.43
R1310 Vbias.n7888 Vbias.n7887 8969.43
R1311 Vbias.n7121 Vbias.n1152 8969.43
R1312 Vbias.n7121 Vbias.n7120 8969.43
R1313 Vbias.n6045 Vbias.n1557 8969.43
R1314 Vbias.n6045 Vbias.n6044 8969.43
R1315 Vbias.n5278 Vbias.n2288 8969.43
R1316 Vbias.n5263 Vbias.n2288 8969.43
R1317 Vbias.n2446 Vbias.n2433 8969.43
R1318 Vbias.n4491 Vbias.n2433 8969.43
R1319 Vbias.n4883 Vbias.n4854 7992.36
R1320 Vbias.n4884 Vbias.n4854 7992.36
R1321 Vbias.n4889 Vbias.n4849 7992.36
R1322 Vbias.n4889 Vbias.n4848 7992.36
R1323 Vbias.n4880 Vbias.n4879 7126.28
R1324 Vbias.n4879 Vbias.n4853 7126.28
R1325 Vbias.n4873 Vbias.n4872 6345.81
R1326 Vbias.n4872 Vbias.n4867 6345.81
R1327 Vbias.n4857 Vbias.n4856 6345.81
R1328 Vbias.n4877 Vbias.n4857 6345.81
R1329 Vbias.n4898 Vbias.n4894 6098.07
R1330 Vbias.n4896 Vbias.n4894 6098.07
R1331 Vbias.n4898 Vbias.n4897 5915.51
R1332 Vbias.n4897 Vbias.n4896 5915.51
R1333 Vbias.n8008 Vbias.n86 5897.47
R1334 Vbias.n7544 Vbias.n917 5734.32
R1335 Vbias.n6531 Vbias.n6504 5734.32
R1336 Vbias.n6598 Vbias.n6226 5734.32
R1337 Vbias.n7668 Vbias.n755 5734.32
R1338 Vbias.n4862 Vbias.n4858 5479.72
R1339 Vbias.n4863 Vbias.n4862 5479.72
R1340 Vbias.n2663 Vbias.n5 4900.92
R1341 Vbias.n4845 Vbias.n2663 4900.92
R1342 Vbias.n4903 Vbias.n4845 4900.92
R1343 Vbias.n4869 Vbias.n4 4699.26
R1344 Vbias.n8079 Vbias.n4 4699.26
R1345 Vbias.n8079 Vbias.n2 4699.26
R1346 Vbias.n4869 Vbias.n2 4699.26
R1347 Vbias.n1203 Vbias.n1190 4207.44
R1348 Vbias.n6936 Vbias.n6923 4207.44
R1349 Vbias.n6847 Vbias.n6846 4207.44
R1350 Vbias.n5989 Vbias.n5988 4207.44
R1351 Vbias.n5307 Vbias.n5294 4207.44
R1352 Vbias.n5216 Vbias.n5215 4207.44
R1353 Vbias.n2475 Vbias.n2462 4207.44
R1354 Vbias.n4452 Vbias.n4434 4207.44
R1355 Vbias.n7225 Vbias.n1071 3443.83
R1356 Vbias.n4903 Vbias.n4902 3201.12
R1357 Vbias.n7122 Vbias.n7121 3097.63
R1358 Vbias.n6075 Vbias.n6045 3097.63
R1359 Vbias.n5485 Vbias.n2288 3097.63
R1360 Vbias.n5037 Vbias.n2433 3097.63
R1361 Vbias.n7122 Vbias.n1151 2528.02
R1362 Vbias.n6076 Vbias.n6075 2528.02
R1363 Vbias.n5486 Vbias.n5485 2528.02
R1364 Vbias.n5037 Vbias.n5036 2528.02
R1365 Vbias.n7016 Vbias.n7015 2291.01
R1366 Vbias.n5919 Vbias.n5918 2291.01
R1367 Vbias.n5122 Vbias.n5121 2291.01
R1368 Vbias.n2905 Vbias.n2663 2200
R1369 Vbias.n4845 Vbias.n4844 2200
R1370 Vbias.n4261 Vbias.n5 2200
R1371 Vbias.n7545 Vbias.n7544 2152.7
R1372 Vbias.n6532 Vbias.n6531 2152.7
R1373 Vbias.n6599 Vbias.n6598 2152.7
R1374 Vbias.n7669 Vbias.n7668 2152.7
R1375 Vbias.n4901 Vbias.t702 2033.91
R1376 Vbias.n4405 Vbias.n2778 2025.26
R1377 Vbias.n4405 Vbias.n2779 2025.26
R1378 Vbias.n4366 Vbias.n2798 2025.26
R1379 Vbias.n4369 Vbias.n4366 2025.26
R1380 Vbias.n4363 Vbias.n2803 2025.26
R1381 Vbias.n4363 Vbias.n2804 2025.26
R1382 Vbias.n4342 Vbias.n2811 2025.26
R1383 Vbias.n4342 Vbias.n4339 2025.26
R1384 Vbias.n4337 Vbias.n2820 2025.26
R1385 Vbias.n4337 Vbias.n2821 2025.26
R1386 Vbias.n2832 Vbias.n2821 2025.26
R1387 Vbias.n2832 Vbias.n2820 2025.26
R1388 Vbias.n4329 Vbias.n2829 2025.26
R1389 Vbias.n4330 Vbias.n2829 2025.26
R1390 Vbias.n2854 Vbias.n2853 2025.26
R1391 Vbias.n4306 Vbias.n2854 2025.26
R1392 Vbias.n4296 Vbias.n2865 2025.26
R1393 Vbias.n4297 Vbias.n2865 2025.26
R1394 Vbias.n2888 Vbias.n2887 2025.26
R1395 Vbias.n4273 Vbias.n2888 2025.26
R1396 Vbias.n2787 Vbias.n2777 2025.26
R1397 Vbias.n4400 Vbias.n2777 2025.26
R1398 Vbias.n4370 Vbias.n2801 2025.26
R1399 Vbias.n2801 Vbias.n2799 2025.26
R1400 Vbias.n2808 Vbias.n2802 2025.26
R1401 Vbias.n4347 Vbias.n2802 2025.26
R1402 Vbias.n4345 Vbias.n4344 2025.26
R1403 Vbias.n4344 Vbias.n2812 2025.26
R1404 Vbias.n4311 Vbias.n2826 2025.26
R1405 Vbias.n4311 Vbias.n2831 2025.26
R1406 Vbias.n4307 Vbias.n2847 2025.26
R1407 Vbias.n2852 Vbias.n2847 2025.26
R1408 Vbias.n4278 Vbias.n2862 2025.26
R1409 Vbias.n4278 Vbias.n2867 2025.26
R1410 Vbias.n4274 Vbias.n2881 2025.26
R1411 Vbias.n2886 Vbias.n2881 2025.26
R1412 Vbias.n4263 Vbias.n4257 2025.26
R1413 Vbias.n4263 Vbias.n4259 2025.26
R1414 Vbias.n4260 Vbias.n4259 2025.26
R1415 Vbias.n4260 Vbias.n4257 2025.26
R1416 Vbias.n5864 Vbias.n5861 2025.26
R1417 Vbias.n5861 Vbias.n5860 2025.26
R1418 Vbias.n1690 Vbias.n1682 2025.26
R1419 Vbias.n1692 Vbias.n1690 2025.26
R1420 Vbias.n1687 Vbias.n1675 2025.26
R1421 Vbias.n1687 Vbias.n1676 2025.26
R1422 Vbias.n5875 Vbias.n1676 2025.26
R1423 Vbias.n5875 Vbias.n1675 2025.26
R1424 Vbias.n5524 Vbias.n5517 2025.26
R1425 Vbias.n5525 Vbias.n5517 2025.26
R1426 Vbias.n5531 Vbias.n5510 2025.26
R1427 Vbias.n5531 Vbias.n5509 2025.26
R1428 Vbias.n5540 Vbias.n5537 2025.26
R1429 Vbias.n5537 Vbias.n5536 2025.26
R1430 Vbias.n2243 Vbias.n2235 2025.26
R1431 Vbias.n2245 Vbias.n2243 2025.26
R1432 Vbias.n2240 Vbias.n2229 2025.26
R1433 Vbias.n2240 Vbias.n2230 2025.26
R1434 Vbias.n5551 Vbias.n2230 2025.26
R1435 Vbias.n5551 Vbias.n2229 2025.26
R1436 Vbias.n5021 Vbias.n5018 2025.26
R1437 Vbias.n5018 Vbias.n5017 2025.26
R1438 Vbias.n5013 Vbias.n2587 2025.26
R1439 Vbias.n5015 Vbias.n5013 2025.26
R1440 Vbias.n5008 Vbias.n2593 2025.26
R1441 Vbias.n5008 Vbias.n2594 2025.26
R1442 Vbias.n5001 Vbias.n2598 2025.26
R1443 Vbias.n5000 Vbias.n2598 2025.26
R1444 Vbias.n4991 Vbias.n2600 2025.26
R1445 Vbias.n4991 Vbias.n2601 2025.26
R1446 Vbias.n4683 Vbias.n2601 2025.26
R1447 Vbias.n4683 Vbias.n2600 2025.26
R1448 Vbias.n7949 Vbias.n164 2025.26
R1449 Vbias.n7950 Vbias.n164 2025.26
R1450 Vbias.n158 Vbias.n156 2025.26
R1451 Vbias.n156 Vbias.n146 2025.26
R1452 Vbias.n7963 Vbias.n136 2025.26
R1453 Vbias.n7964 Vbias.n136 2025.26
R1454 Vbias.n7969 Vbias.n131 2025.26
R1455 Vbias.n7969 Vbias.n130 2025.26
R1456 Vbias.n7974 Vbias.n129 2025.26
R1457 Vbias.n7973 Vbias.n129 2025.26
R1458 Vbias.n7984 Vbias.n110 2025.26
R1459 Vbias.n7984 Vbias.n109 2025.26
R1460 Vbias.n7989 Vbias.n108 2025.26
R1461 Vbias.n7988 Vbias.n108 2025.26
R1462 Vbias.n7999 Vbias.n91 2025.26
R1463 Vbias.n7999 Vbias.n90 2025.26
R1464 Vbias.n8002 Vbias.n87 2025.26
R1465 Vbias.n8002 Vbias.n88 2025.26
R1466 Vbias.n8006 Vbias.n88 2025.26
R1467 Vbias.n8006 Vbias.n87 2025.26
R1468 Vbias.n8012 Vbias.n85 2025.26
R1469 Vbias.n8011 Vbias.n85 2025.26
R1470 Vbias.n8023 Vbias.n67 2025.26
R1471 Vbias.n8023 Vbias.n66 2025.26
R1472 Vbias.n8031 Vbias.n64 2025.26
R1473 Vbias.n8032 Vbias.n64 2025.26
R1474 Vbias.n8038 Vbias.n58 2025.26
R1475 Vbias.n8038 Vbias.n57 2025.26
R1476 Vbias.n8041 Vbias.n54 2025.26
R1477 Vbias.n8041 Vbias.n52 2025.26
R1478 Vbias.n55 Vbias.n52 2025.26
R1479 Vbias.n55 Vbias.n54 2025.26
R1480 Vbias.n8049 Vbias.n46 2025.26
R1481 Vbias.n8048 Vbias.n46 2025.26
R1482 Vbias.n38 Vbias.n32 2025.26
R1483 Vbias.n40 Vbias.n38 2025.26
R1484 Vbias.n8064 Vbias.n28 2025.26
R1485 Vbias.n8063 Vbias.n28 2025.26
R1486 Vbias.n8074 Vbias.n11 2025.26
R1487 Vbias.n8074 Vbias.n10 2025.26
R1488 Vbias.n6711 Vbias.n6700 2025.26
R1489 Vbias.n6711 Vbias.n6698 2025.26
R1490 Vbias.n6702 Vbias.n6696 2025.26
R1491 Vbias.n6705 Vbias.n6702 2025.26
R1492 Vbias.n6738 Vbias.n6724 2025.26
R1493 Vbias.n6738 Vbias.n6722 2025.26
R1494 Vbias.n6728 Vbias.n6720 2025.26
R1495 Vbias.n6731 Vbias.n6728 2025.26
R1496 Vbias.n6725 Vbias.n1445 2025.26
R1497 Vbias.n6725 Vbias.n1446 2025.26
R1498 Vbias.n6748 Vbias.n1446 2025.26
R1499 Vbias.n6748 Vbias.n1445 2025.26
R1500 Vbias.n2038 Vbias.n2037 2025.26
R1501 Vbias.n2037 Vbias.n1733 2025.26
R1502 Vbias.n1742 Vbias.n1739 2025.26
R1503 Vbias.n1739 Vbias.n1738 2025.26
R1504 Vbias.n5853 Vbias.n1703 2025.26
R1505 Vbias.n5852 Vbias.n1703 2025.26
R1506 Vbias.n5846 Vbias.n2065 2025.26
R1507 Vbias.n5845 Vbias.n2065 2025.26
R1508 Vbias.n5838 Vbias.n5833 2025.26
R1509 Vbias.n5838 Vbias.n5836 2025.26
R1510 Vbias.n5836 Vbias.n5835 2025.26
R1511 Vbias.n5835 Vbias.n5833 2025.26
R1512 Vbias.n7743 Vbias.n676 2025.26
R1513 Vbias.n7744 Vbias.n676 2025.26
R1514 Vbias.n7750 Vbias.n669 2025.26
R1515 Vbias.n7750 Vbias.n668 2025.26
R1516 Vbias.n5824 Vbias.n2073 2025.26
R1517 Vbias.n5823 Vbias.n2073 2025.26
R1518 Vbias.n5794 Vbias.n5793 2025.26
R1519 Vbias.n5794 Vbias.n2085 2025.26
R1520 Vbias.n5810 Vbias.n5790 2025.26
R1521 Vbias.n5809 Vbias.n5790 2025.26
R1522 Vbias.n5805 Vbias.n5801 2025.26
R1523 Vbias.n5804 Vbias.n5801 2025.26
R1524 Vbias.n5782 Vbias.n5781 2025.26
R1525 Vbias.n5781 Vbias.n5780 2025.26
R1526 Vbias.n2110 Vbias.n2109 2025.26
R1527 Vbias.n2110 Vbias.n2101 2025.26
R1528 Vbias.n5767 Vbias.n2106 2025.26
R1529 Vbias.n5766 Vbias.n2106 2025.26
R1530 Vbias.n5749 Vbias.n5748 2025.26
R1531 Vbias.n5749 Vbias.n2123 2025.26
R1532 Vbias.n5752 Vbias.n5743 2025.26
R1533 Vbias.n5752 Vbias.n5746 2025.26
R1534 Vbias.n5746 Vbias.n5745 2025.26
R1535 Vbias.n5745 Vbias.n5743 2025.26
R1536 Vbias.n7808 Vbias.n7805 2025.26
R1537 Vbias.n7805 Vbias.n7804 2025.26
R1538 Vbias.n568 Vbias.n560 2025.26
R1539 Vbias.n570 Vbias.n568 2025.26
R1540 Vbias.n565 Vbias.n554 2025.26
R1541 Vbias.n565 Vbias.n555 2025.26
R1542 Vbias.n7819 Vbias.n555 2025.26
R1543 Vbias.n7819 Vbias.n554 2025.26
R1544 Vbias.n5735 Vbias.n2128 2025.26
R1545 Vbias.n5734 Vbias.n2128 2025.26
R1546 Vbias.n2149 Vbias.n2148 2025.26
R1547 Vbias.n2149 Vbias.n2140 2025.26
R1548 Vbias.n5721 Vbias.n2145 2025.26
R1549 Vbias.n5720 Vbias.n2145 2025.26
R1550 Vbias.n5716 Vbias.n2156 2025.26
R1551 Vbias.n5715 Vbias.n2156 2025.26
R1552 Vbias.n5711 Vbias.n2157 2025.26
R1553 Vbias.n5711 Vbias.n2158 2025.26
R1554 Vbias.n5696 Vbias.n2174 2025.26
R1555 Vbias.n5697 Vbias.n2174 2025.26
R1556 Vbias.n5692 Vbias.n2175 2025.26
R1557 Vbias.n5692 Vbias.n2176 2025.26
R1558 Vbias.n5678 Vbias.n2192 2025.26
R1559 Vbias.n5679 Vbias.n2192 2025.26
R1560 Vbias.n5674 Vbias.n2193 2025.26
R1561 Vbias.n5674 Vbias.n2194 2025.26
R1562 Vbias.n5670 Vbias.n2194 2025.26
R1563 Vbias.n5670 Vbias.n2193 2025.26
R1564 Vbias.n7878 Vbias.n455 2025.26
R1565 Vbias.n7879 Vbias.n455 2025.26
R1566 Vbias.n7885 Vbias.n449 2025.26
R1567 Vbias.n7885 Vbias.n448 2025.26
R1568 Vbias.n5661 Vbias.n2199 2025.26
R1569 Vbias.n5660 Vbias.n2199 2025.26
R1570 Vbias.n2220 Vbias.n2219 2025.26
R1571 Vbias.n2220 Vbias.n2211 2025.26
R1572 Vbias.n5647 Vbias.n2216 2025.26
R1573 Vbias.n5646 Vbias.n2216 2025.26
R1574 Vbias.n5642 Vbias.n2227 2025.26
R1575 Vbias.n5641 Vbias.n2227 2025.26
R1576 Vbias.n5637 Vbias.n5554 2025.26
R1577 Vbias.n5637 Vbias.n5555 2025.26
R1578 Vbias.n5622 Vbias.n5571 2025.26
R1579 Vbias.n5623 Vbias.n5571 2025.26
R1580 Vbias.n5618 Vbias.n5572 2025.26
R1581 Vbias.n5618 Vbias.n5573 2025.26
R1582 Vbias.n5604 Vbias.n5589 2025.26
R1583 Vbias.n5605 Vbias.n5589 2025.26
R1584 Vbias.n5600 Vbias.n5590 2025.26
R1585 Vbias.n5600 Vbias.n5591 2025.26
R1586 Vbias.n5596 Vbias.n5591 2025.26
R1587 Vbias.n5596 Vbias.n5590 2025.26
R1588 Vbias.n7939 Vbias.n173 2025.26
R1589 Vbias.n7939 Vbias.n171 2025.26
R1590 Vbias.n340 Vbias.n329 2025.26
R1591 Vbias.n340 Vbias.n328 2025.26
R1592 Vbias.n343 Vbias.n324 2025.26
R1593 Vbias.n343 Vbias.n325 2025.26
R1594 Vbias.n347 Vbias.n325 2025.26
R1595 Vbias.n347 Vbias.n324 2025.26
R1596 Vbias.n1025 Vbias.n1024 2025.26
R1597 Vbias.n1025 Vbias.n922 2025.26
R1598 Vbias.n1016 Vbias.n1013 2025.26
R1599 Vbias.n1016 Vbias.n1012 2025.26
R1600 Vbias.n7532 Vbias.n928 2025.26
R1601 Vbias.n7532 Vbias.n926 2025.26
R1602 Vbias.n6521 Vbias.n6520 2025.26
R1603 Vbias.n6530 Vbias.n6521 2025.26
R1604 Vbias.n6516 Vbias.n6505 2025.26
R1605 Vbias.n6516 Vbias.n6506 2025.26
R1606 Vbias.n6509 Vbias.n6506 2025.26
R1607 Vbias.n6509 Vbias.n6505 2025.26
R1608 Vbias.n7653 Vbias.n777 2025.26
R1609 Vbias.n7653 Vbias.n775 2025.26
R1610 Vbias.n6591 Vbias.n773 2025.26
R1611 Vbias.n6594 Vbias.n6591 2025.26
R1612 Vbias.n7663 Vbias.n764 2025.26
R1613 Vbias.n7662 Vbias.n764 2025.26
R1614 Vbias.n759 Vbias.n758 2025.26
R1615 Vbias.n7667 Vbias.n759 2025.26
R1616 Vbias.n7264 Vbias.n7261 2025.26
R1617 Vbias.n7255 Vbias.n7253 2025.26
R1618 Vbias.n7253 Vbias.n7243 2025.26
R1619 Vbias.n7279 Vbias.n7233 2025.26
R1620 Vbias.n7280 Vbias.n7233 2025.26
R1621 Vbias.n7285 Vbias.n7228 2025.26
R1622 Vbias.n7285 Vbias.n7227 2025.26
R1623 Vbias.n7290 Vbias.n1070 2025.26
R1624 Vbias.n7289 Vbias.n1070 2025.26
R1625 Vbias.n7300 Vbias.n1051 2025.26
R1626 Vbias.n7300 Vbias.n1050 2025.26
R1627 Vbias.n7305 Vbias.n1049 2025.26
R1628 Vbias.n7304 Vbias.n1049 2025.26
R1629 Vbias.n7315 Vbias.n1030 2025.26
R1630 Vbias.n7315 Vbias.n1029 2025.26
R1631 Vbias.n7318 Vbias.n1020 2025.26
R1632 Vbias.n7318 Vbias.n1022 2025.26
R1633 Vbias.n1027 Vbias.n1022 2025.26
R1634 Vbias.n1027 Vbias.n1020 2025.26
R1635 Vbias.n7471 Vbias.n1011 2025.26
R1636 Vbias.n7472 Vbias.n1011 2025.26
R1637 Vbias.n1005 Vbias.n1003 2025.26
R1638 Vbias.n1003 Vbias.n993 2025.26
R1639 Vbias.n7485 Vbias.n983 2025.26
R1640 Vbias.n7486 Vbias.n983 2025.26
R1641 Vbias.n7491 Vbias.n978 2025.26
R1642 Vbias.n7491 Vbias.n977 2025.26
R1643 Vbias.n7497 Vbias.n975 2025.26
R1644 Vbias.n7496 Vbias.n975 2025.26
R1645 Vbias.n7507 Vbias.n956 2025.26
R1646 Vbias.n7507 Vbias.n955 2025.26
R1647 Vbias.n7512 Vbias.n954 2025.26
R1648 Vbias.n7511 Vbias.n954 2025.26
R1649 Vbias.n7522 Vbias.n933 2025.26
R1650 Vbias.n7522 Vbias.n932 2025.26
R1651 Vbias.n7525 Vbias.n929 2025.26
R1652 Vbias.n7525 Vbias.n930 2025.26
R1653 Vbias.n7529 Vbias.n930 2025.26
R1654 Vbias.n7529 Vbias.n929 2025.26
R1655 Vbias.n7593 Vbias.n856 2025.26
R1656 Vbias.n7594 Vbias.n856 2025.26
R1657 Vbias.n850 Vbias.n848 2025.26
R1658 Vbias.n848 Vbias.n838 2025.26
R1659 Vbias.n7607 Vbias.n828 2025.26
R1660 Vbias.n7608 Vbias.n828 2025.26
R1661 Vbias.n7613 Vbias.n823 2025.26
R1662 Vbias.n7613 Vbias.n822 2025.26
R1663 Vbias.n7618 Vbias.n820 2025.26
R1664 Vbias.n7617 Vbias.n820 2025.26
R1665 Vbias.n7628 Vbias.n801 2025.26
R1666 Vbias.n7628 Vbias.n800 2025.26
R1667 Vbias.n7633 Vbias.n799 2025.26
R1668 Vbias.n7632 Vbias.n799 2025.26
R1669 Vbias.n7643 Vbias.n782 2025.26
R1670 Vbias.n7643 Vbias.n781 2025.26
R1671 Vbias.n7646 Vbias.n778 2025.26
R1672 Vbias.n7646 Vbias.n779 2025.26
R1673 Vbias.n7650 Vbias.n779 2025.26
R1674 Vbias.n7650 Vbias.n778 2025.26
R1675 Vbias.n6588 Vbias.n6227 2025.26
R1676 Vbias.n6588 Vbias.n6228 2025.26
R1677 Vbias.n6355 Vbias.n6244 2025.26
R1678 Vbias.n6356 Vbias.n6244 2025.26
R1679 Vbias.n6351 Vbias.n6245 2025.26
R1680 Vbias.n6351 Vbias.n6246 2025.26
R1681 Vbias.n6346 Vbias.n6250 2025.26
R1682 Vbias.n6345 Vbias.n6250 2025.26
R1683 Vbias.n6338 Vbias.n6262 2025.26
R1684 Vbias.n6337 Vbias.n6262 2025.26
R1685 Vbias.n6283 Vbias.n6282 2025.26
R1686 Vbias.n6283 Vbias.n6274 2025.26
R1687 Vbias.n6324 Vbias.n6279 2025.26
R1688 Vbias.n6323 Vbias.n6279 2025.26
R1689 Vbias.n6306 Vbias.n6305 2025.26
R1690 Vbias.n6306 Vbias.n6296 2025.26
R1691 Vbias.n6309 Vbias.n6299 2025.26
R1692 Vbias.n6309 Vbias.n6301 2025.26
R1693 Vbias.n6302 Vbias.n6301 2025.26
R1694 Vbias.n6302 Vbias.n6299 2025.26
R1695 Vbias.n6654 Vbias.n1500 2025.26
R1696 Vbias.n6655 Vbias.n1500 2025.26
R1697 Vbias.n1494 Vbias.n1493 2025.26
R1698 Vbias.n1493 Vbias.n1483 2025.26
R1699 Vbias.n6668 Vbias.n1474 2025.26
R1700 Vbias.n6669 Vbias.n1474 2025.26
R1701 Vbias.n6674 Vbias.n1469 2025.26
R1702 Vbias.n6674 Vbias.n1468 2025.26
R1703 Vbias.n7672 Vbias.n754 2025.26
R1704 Vbias.n7671 Vbias.n754 2025.26
R1705 Vbias.n7683 Vbias.n736 2025.26
R1706 Vbias.n7683 Vbias.n735 2025.26
R1707 Vbias.n7691 Vbias.n733 2025.26
R1708 Vbias.n7692 Vbias.n733 2025.26
R1709 Vbias.n7698 Vbias.n727 2025.26
R1710 Vbias.n7698 Vbias.n726 2025.26
R1711 Vbias.n7701 Vbias.n723 2025.26
R1712 Vbias.n7701 Vbias.n721 2025.26
R1713 Vbias.n724 Vbias.n721 2025.26
R1714 Vbias.n724 Vbias.n723 2025.26
R1715 Vbias.n7709 Vbias.n715 2025.26
R1716 Vbias.n7708 Vbias.n715 2025.26
R1717 Vbias.n707 Vbias.n701 2025.26
R1718 Vbias.n709 Vbias.n707 2025.26
R1719 Vbias.n7724 Vbias.n697 2025.26
R1720 Vbias.n7723 Vbias.n697 2025.26
R1721 Vbias.n7734 Vbias.n680 2025.26
R1722 Vbias.n7734 Vbias.n679 2025.26
R1723 Vbias.n7754 Vbias.n653 2025.26
R1724 Vbias.n7754 Vbias.n651 2025.26
R1725 Vbias.n7763 Vbias.n644 2025.26
R1726 Vbias.n7763 Vbias.n643 2025.26
R1727 Vbias.n7766 Vbias.n631 2025.26
R1728 Vbias.n7766 Vbias.n629 2025.26
R1729 Vbias.n635 Vbias.n627 2025.26
R1730 Vbias.n638 Vbias.n635 2025.26
R1731 Vbias.n632 Vbias.n620 2025.26
R1732 Vbias.n632 Vbias.n621 2025.26
R1733 Vbias.n7776 Vbias.n621 2025.26
R1734 Vbias.n7776 Vbias.n620 2025.26
R1735 Vbias.n7779 Vbias.n606 2025.26
R1736 Vbias.n7779 Vbias.n604 2025.26
R1737 Vbias.n7788 Vbias.n597 2025.26
R1738 Vbias.n7788 Vbias.n596 2025.26
R1739 Vbias.n7800 Vbias.n572 2025.26
R1740 Vbias.n7800 Vbias.n573 2025.26
R1741 Vbias.n7791 Vbias.n582 2025.26
R1742 Vbias.n7791 Vbias.n580 2025.26
R1743 Vbias.n7823 Vbias.n539 2025.26
R1744 Vbias.n7823 Vbias.n537 2025.26
R1745 Vbias.n7832 Vbias.n530 2025.26
R1746 Vbias.n7832 Vbias.n529 2025.26
R1747 Vbias.n7835 Vbias.n517 2025.26
R1748 Vbias.n7835 Vbias.n515 2025.26
R1749 Vbias.n521 Vbias.n513 2025.26
R1750 Vbias.n524 Vbias.n521 2025.26
R1751 Vbias.n518 Vbias.n506 2025.26
R1752 Vbias.n518 Vbias.n507 2025.26
R1753 Vbias.n7845 Vbias.n507 2025.26
R1754 Vbias.n7845 Vbias.n506 2025.26
R1755 Vbias.n7848 Vbias.n492 2025.26
R1756 Vbias.n7848 Vbias.n490 2025.26
R1757 Vbias.n7857 Vbias.n483 2025.26
R1758 Vbias.n7857 Vbias.n482 2025.26
R1759 Vbias.n7869 Vbias.n458 2025.26
R1760 Vbias.n7869 Vbias.n459 2025.26
R1761 Vbias.n7860 Vbias.n468 2025.26
R1762 Vbias.n7860 Vbias.n466 2025.26
R1763 Vbias.n7889 Vbias.n433 2025.26
R1764 Vbias.n7889 Vbias.n431 2025.26
R1765 Vbias.n7898 Vbias.n424 2025.26
R1766 Vbias.n7898 Vbias.n423 2025.26
R1767 Vbias.n7901 Vbias.n411 2025.26
R1768 Vbias.n7901 Vbias.n409 2025.26
R1769 Vbias.n415 Vbias.n407 2025.26
R1770 Vbias.n418 Vbias.n415 2025.26
R1771 Vbias.n412 Vbias.n400 2025.26
R1772 Vbias.n412 Vbias.n401 2025.26
R1773 Vbias.n7911 Vbias.n401 2025.26
R1774 Vbias.n7911 Vbias.n400 2025.26
R1775 Vbias.n7914 Vbias.n386 2025.26
R1776 Vbias.n7914 Vbias.n384 2025.26
R1777 Vbias.n7923 Vbias.n377 2025.26
R1778 Vbias.n7923 Vbias.n376 2025.26
R1779 Vbias.n7935 Vbias.n175 2025.26
R1780 Vbias.n7935 Vbias.n176 2025.26
R1781 Vbias.n7926 Vbias.n362 2025.26
R1782 Vbias.n7926 Vbias.n360 2025.26
R1783 Vbias.n351 Vbias.n183 2025.26
R1784 Vbias.n351 Vbias.n181 2025.26
R1785 Vbias.n315 Vbias.n188 2025.26
R1786 Vbias.n316 Vbias.n188 2025.26
R1787 Vbias.n308 Vbias.n202 2025.26
R1788 Vbias.n308 Vbias.n200 2025.26
R1789 Vbias.n300 Vbias.n207 2025.26
R1790 Vbias.n301 Vbias.n300 2025.26
R1791 Vbias.n297 Vbias.n208 2025.26
R1792 Vbias.n297 Vbias.n209 2025.26
R1793 Vbias.n285 Vbias.n209 2025.26
R1794 Vbias.n285 Vbias.n208 2025.26
R1795 Vbias.n288 Vbias.n216 2025.26
R1796 Vbias.n288 Vbias.n214 2025.26
R1797 Vbias.n276 Vbias.n221 2025.26
R1798 Vbias.n277 Vbias.n221 2025.26
R1799 Vbias.n260 Vbias.n240 2025.26
R1800 Vbias.n259 Vbias.n240 2025.26
R1801 Vbias.n269 Vbias.n235 2025.26
R1802 Vbias.n269 Vbias.n233 2025.26
R1803 Vbias.n5035 Vbias.n2434 2025.26
R1804 Vbias.n5035 Vbias.n2435 2025.26
R1805 Vbias.n4611 Vbias.n4602 2025.26
R1806 Vbias.n4634 Vbias.n4611 2025.26
R1807 Vbias.n4631 Vbias.n4630 2025.26
R1808 Vbias.n4631 Vbias.n4599 2025.26
R1809 Vbias.n4619 Vbias.n4595 2025.26
R1810 Vbias.n4621 Vbias.n4619 2025.26
R1811 Vbias.n4616 Vbias.n4589 2025.26
R1812 Vbias.n4616 Vbias.n4590 2025.26
R1813 Vbias.n4659 Vbias.n4590 2025.26
R1814 Vbias.n4659 Vbias.n4589 2025.26
R1815 Vbias.n4662 Vbias.n4582 2025.26
R1816 Vbias.n4662 Vbias.n4580 2025.26
R1817 Vbias.n4669 Vbias.n4575 2025.26
R1818 Vbias.n4669 Vbias.n4574 2025.26
R1819 Vbias.n4492 Vbias.n4486 2025.26
R1820 Vbias.n4492 Vbias.n4488 2025.26
R1821 Vbias.n4489 Vbias.n4488 2025.26
R1822 Vbias.n4489 Vbias.n4486 2025.26
R1823 Vbias.n4499 Vbias.n4481 2025.26
R1824 Vbias.n4500 Vbias.n4481 2025.26
R1825 Vbias.n4475 Vbias.n4473 2025.26
R1826 Vbias.n4473 Vbias.n4463 2025.26
R1827 Vbias.n4513 Vbias.n4459 2025.26
R1828 Vbias.n4514 Vbias.n4459 2025.26
R1829 Vbias.n4453 Vbias.n4451 2025.26
R1830 Vbias.n4451 Vbias.n4441 2025.26
R1831 Vbias.n4527 Vbias.n4432 2025.26
R1832 Vbias.n4528 Vbias.n4432 2025.26
R1833 Vbias.n4533 Vbias.n4427 2025.26
R1834 Vbias.n4533 Vbias.n4426 2025.26
R1835 Vbias.n4538 Vbias.n4425 2025.26
R1836 Vbias.n4537 Vbias.n4425 2025.26
R1837 Vbias.n4549 Vbias.n4408 2025.26
R1838 Vbias.n4549 Vbias.n4407 2025.26
R1839 Vbias.n5119 Vbias.n2372 2025.26
R1840 Vbias.n5119 Vbias.n2373 2025.26
R1841 Vbias.n5103 Vbias.n2387 2025.26
R1842 Vbias.n5104 Vbias.n2387 2025.26
R1843 Vbias.n5099 Vbias.n2388 2025.26
R1844 Vbias.n5099 Vbias.n2389 2025.26
R1845 Vbias.n5083 Vbias.n5081 2025.26
R1846 Vbias.n5084 Vbias.n5081 2025.26
R1847 Vbias.n5078 Vbias.n2403 2025.26
R1848 Vbias.n5078 Vbias.n2404 2025.26
R1849 Vbias.n5066 Vbias.n2404 2025.26
R1850 Vbias.n5066 Vbias.n2403 2025.26
R1851 Vbias.n5069 Vbias.n2411 2025.26
R1852 Vbias.n5069 Vbias.n2409 2025.26
R1853 Vbias.n5059 Vbias.n2416 2025.26
R1854 Vbias.n5060 Vbias.n5059 2025.26
R1855 Vbias.n5487 Vbias.n2274 2025.26
R1856 Vbias.n5487 Vbias.n2272 2025.26
R1857 Vbias.n5496 Vbias.n2266 2025.26
R1858 Vbias.n5496 Vbias.n2265 2025.26
R1859 Vbias.n5499 Vbias.n2256 2025.26
R1860 Vbias.n5499 Vbias.n2254 2025.26
R1861 Vbias.n5156 Vbias.n5153 2025.26
R1862 Vbias.n5156 Vbias.n5152 2025.26
R1863 Vbias.n5159 Vbias.n5149 2025.26
R1864 Vbias.n5159 Vbias.n5150 2025.26
R1865 Vbias.n5166 Vbias.n5150 2025.26
R1866 Vbias.n5166 Vbias.n5149 2025.26
R1867 Vbias.n5169 Vbias.n2363 2025.26
R1868 Vbias.n5169 Vbias.n2361 2025.26
R1869 Vbias.n5141 Vbias.n2359 2025.26
R1870 Vbias.n5144 Vbias.n5141 2025.26
R1871 Vbias.n5138 Vbias.n5137 2025.26
R1872 Vbias.n5138 Vbias.n2355 2025.26
R1873 Vbias.n5124 Vbias.n2351 2025.26
R1874 Vbias.n5126 Vbias.n5124 2025.26
R1875 Vbias.n5916 Vbias.n1640 2025.26
R1876 Vbias.n5916 Vbias.n1641 2025.26
R1877 Vbias.n5900 Vbias.n1655 2025.26
R1878 Vbias.n5901 Vbias.n1655 2025.26
R1879 Vbias.n5896 Vbias.n1656 2025.26
R1880 Vbias.n5896 Vbias.n1657 2025.26
R1881 Vbias.n5880 Vbias.n1671 2025.26
R1882 Vbias.n5881 Vbias.n1671 2025.26
R1883 Vbias.n5455 Vbias.n5451 2025.26
R1884 Vbias.n5455 Vbias.n5452 2025.26
R1885 Vbias.n5461 Vbias.n5452 2025.26
R1886 Vbias.n5461 Vbias.n5451 2025.26
R1887 Vbias.n5464 Vbias.n5444 2025.26
R1888 Vbias.n5464 Vbias.n5442 2025.26
R1889 Vbias.n5471 Vbias.n5437 2025.26
R1890 Vbias.n5471 Vbias.n5436 2025.26
R1891 Vbias.n5474 Vbias.n5422 2025.26
R1892 Vbias.n5474 Vbias.n5420 2025.26
R1893 Vbias.n5483 Vbias.n2290 2025.26
R1894 Vbias.n5483 Vbias.n2289 2025.26
R1895 Vbias.n5942 Vbias.n5941 2025.26
R1896 Vbias.n5942 Vbias.n1625 2025.26
R1897 Vbias.n5934 Vbias.n1623 2025.26
R1898 Vbias.n5937 Vbias.n5934 2025.26
R1899 Vbias.n5931 Vbias.n5930 2025.26
R1900 Vbias.n5931 Vbias.n1618 2025.26
R1901 Vbias.n1634 Vbias.n1614 2025.26
R1902 Vbias.n5921 Vbias.n1634 2025.26
R1903 Vbias.n1805 Vbias.n1533 2025.26
R1904 Vbias.n1805 Vbias.n1534 2025.26
R1905 Vbias.n6099 Vbias.n1534 2025.26
R1906 Vbias.n6099 Vbias.n1533 2025.26
R1907 Vbias.n1818 Vbias.n1758 2025.26
R1908 Vbias.n1817 Vbias.n1758 2025.26
R1909 Vbias.n1809 Vbias.n1803 2025.26
R1910 Vbias.n1810 Vbias.n1803 2025.26
R1911 Vbias.n1872 Vbias.n1868 2025.26
R1912 Vbias.n1873 Vbias.n1868 2025.26
R1913 Vbias.n1862 Vbias.n1860 2025.26
R1914 Vbias.n1861 Vbias.n1860 2025.26
R1915 Vbias.n1938 Vbias.n1934 2025.26
R1916 Vbias.n1939 Vbias.n1934 2025.26
R1917 Vbias.n1930 Vbias.n1928 2025.26
R1918 Vbias.n1929 Vbias.n1928 2025.26
R1919 Vbias.n2012 Vbias.n1986 2025.26
R1920 Vbias.n2012 Vbias.n2011 2025.26
R1921 Vbias.n2003 Vbias.n1992 2025.26
R1922 Vbias.n2002 Vbias.n1992 2025.26
R1923 Vbias.n6112 Vbias.n6108 2025.26
R1924 Vbias.n6113 Vbias.n6108 2025.26
R1925 Vbias.n6104 Vbias.n1522 2025.26
R1926 Vbias.n6103 Vbias.n1522 2025.26
R1927 Vbias.n1972 Vbias.n1968 2025.26
R1928 Vbias.n1973 Vbias.n1968 2025.26
R1929 Vbias.n1964 Vbias.n1962 2025.26
R1930 Vbias.n1963 Vbias.n1962 2025.26
R1931 Vbias.n1904 Vbias.n1895 2025.26
R1932 Vbias.n1903 Vbias.n1895 2025.26
R1933 Vbias.n1911 Vbias.n1885 2025.26
R1934 Vbias.n1912 Vbias.n1885 2025.26
R1935 Vbias.n6077 Vbias.n1553 2025.26
R1936 Vbias.n6077 Vbias.n1551 2025.26
R1937 Vbias.n1788 Vbias.n1547 2025.26
R1938 Vbias.n1788 Vbias.n1787 2025.26
R1939 Vbias.n1793 Vbias.n1791 2025.26
R1940 Vbias.n1791 Vbias.n1543 2025.26
R1941 Vbias.n1768 Vbias.n1539 2025.26
R1942 Vbias.n1799 Vbias.n1768 2025.26
R1943 Vbias.n7013 Vbias.n1341 2025.26
R1944 Vbias.n7013 Vbias.n1342 2025.26
R1945 Vbias.n1439 Vbias.n1430 2025.26
R1946 Vbias.n6772 Vbias.n1439 2025.26
R1947 Vbias.n6769 Vbias.n6768 2025.26
R1948 Vbias.n6769 Vbias.n1427 2025.26
R1949 Vbias.n6755 Vbias.n1423 2025.26
R1950 Vbias.n6757 Vbias.n6755 2025.26
R1951 Vbias.n6752 Vbias.n1416 2025.26
R1952 Vbias.n6752 Vbias.n1417 2025.26
R1953 Vbias.n6797 Vbias.n1417 2025.26
R1954 Vbias.n6797 Vbias.n1416 2025.26
R1955 Vbias.n6800 Vbias.n1415 2025.26
R1956 Vbias.n6800 Vbias.n1413 2025.26
R1957 Vbias.n6059 Vbias.n1411 2025.26
R1958 Vbias.n6059 Vbias.n6058 2025.26
R1959 Vbias.n6064 Vbias.n6062 2025.26
R1960 Vbias.n6062 Vbias.n1407 2025.26
R1961 Vbias.n6073 Vbias.n1403 2025.26
R1962 Vbias.n6073 Vbias.n6072 2025.26
R1963 Vbias.n7091 Vbias.n7090 2025.26
R1964 Vbias.n7091 Vbias.n1276 2025.26
R1965 Vbias.n7081 Vbias.n1282 2025.26
R1966 Vbias.n7082 Vbias.n1282 2025.26
R1967 Vbias.n7074 Vbias.n1296 2025.26
R1968 Vbias.n7074 Vbias.n1294 2025.26
R1969 Vbias.n7064 Vbias.n1301 2025.26
R1970 Vbias.n7065 Vbias.n1301 2025.26
R1971 Vbias.n7057 Vbias.n1315 2025.26
R1972 Vbias.n7057 Vbias.n1313 2025.26
R1973 Vbias.n7054 Vbias.n1313 2025.26
R1974 Vbias.n7054 Vbias.n1315 2025.26
R1975 Vbias.n7052 Vbias.n1316 2025.26
R1976 Vbias.n7052 Vbias.n1317 2025.26
R1977 Vbias.n7045 Vbias.n1321 2025.26
R1978 Vbias.n7044 Vbias.n1321 2025.26
R1979 Vbias.n7035 Vbias.n1323 2025.26
R1980 Vbias.n7035 Vbias.n1324 2025.26
R1981 Vbias.n7019 Vbias.n1338 2025.26
R1982 Vbias.n7020 Vbias.n1338 2025.26
R1983 Vbias.n7197 Vbias.n7196 2025.26
R1984 Vbias.n7197 Vbias.n1089 2025.26
R1985 Vbias.n7187 Vbias.n1095 2025.26
R1986 Vbias.n7188 Vbias.n1095 2025.26
R1987 Vbias.n7180 Vbias.n1109 2025.26
R1988 Vbias.n7180 Vbias.n1107 2025.26
R1989 Vbias.n7170 Vbias.n1114 2025.26
R1990 Vbias.n7171 Vbias.n1114 2025.26
R1991 Vbias.n7163 Vbias.n1127 2025.26
R1992 Vbias.n7163 Vbias.n1125 2025.26
R1993 Vbias.n7160 Vbias.n1125 2025.26
R1994 Vbias.n7160 Vbias.n1127 2025.26
R1995 Vbias.n7158 Vbias.n1128 2025.26
R1996 Vbias.n7158 Vbias.n1129 2025.26
R1997 Vbias.n7151 Vbias.n1133 2025.26
R1998 Vbias.n7150 Vbias.n1133 2025.26
R1999 Vbias.n7141 Vbias.n1135 2025.26
R2000 Vbias.n7141 Vbias.n1136 2025.26
R2001 Vbias.n7125 Vbias.n1150 2025.26
R2002 Vbias.n7126 Vbias.n1150 2025.26
R2003 Vbias.n7219 Vbias.n1072 2025.26
R2004 Vbias.n7223 Vbias.n1072 2025.26
R2005 Vbias.n7223 Vbias.n1073 2025.26
R2006 Vbias.n7219 Vbias.n1073 2025.26
R2007 Vbias.n7216 Vbias.n1075 2025.26
R2008 Vbias.n7216 Vbias.n1076 2025.26
R2009 Vbias.n1223 Vbias.n1215 2025.26
R2010 Vbias.n1223 Vbias.n1214 2025.26
R2011 Vbias.n1234 Vbias.n1210 2025.26
R2012 Vbias.n1233 Vbias.n1210 2025.26
R2013 Vbias.n1206 Vbias.n1204 2025.26
R2014 Vbias.n1204 Vbias.n1198 2025.26
R2015 Vbias.n1247 Vbias.n1192 2025.26
R2016 Vbias.n1192 Vbias.n1191 2025.26
R2017 Vbias.n1254 Vbias.n1184 2025.26
R2018 Vbias.n1254 Vbias.n1183 2025.26
R2019 Vbias.n1265 Vbias.n1181 2025.26
R2020 Vbias.n1264 Vbias.n1181 2025.26
R2021 Vbias.n1177 Vbias.n1175 2025.26
R2022 Vbias.n1175 Vbias.n1170 2025.26
R2023 Vbias.n7119 Vbias.n1153 2025.26
R2024 Vbias.n7119 Vbias.n1154 2025.26
R2025 Vbias.n7115 Vbias.n1154 2025.26
R2026 Vbias.n7115 Vbias.n1153 2025.26
R2027 Vbias.n7112 Vbias.n1156 2025.26
R2028 Vbias.n7112 Vbias.n1157 2025.26
R2029 Vbias.n6956 Vbias.n6948 2025.26
R2030 Vbias.n6956 Vbias.n6947 2025.26
R2031 Vbias.n6967 Vbias.n6943 2025.26
R2032 Vbias.n6966 Vbias.n6943 2025.26
R2033 Vbias.n6939 Vbias.n6937 2025.26
R2034 Vbias.n6937 Vbias.n6931 2025.26
R2035 Vbias.n6980 Vbias.n6925 2025.26
R2036 Vbias.n6925 Vbias.n6924 2025.26
R2037 Vbias.n6987 Vbias.n6917 2025.26
R2038 Vbias.n6987 Vbias.n6916 2025.26
R2039 Vbias.n6998 Vbias.n6914 2025.26
R2040 Vbias.n6997 Vbias.n6914 2025.26
R2041 Vbias.n6910 Vbias.n6908 2025.26
R2042 Vbias.n6908 Vbias.n6903 2025.26
R2043 Vbias.n6896 Vbias.n1349 2025.26
R2044 Vbias.n6895 Vbias.n1349 2025.26
R2045 Vbias.n6895 Vbias.n1348 2025.26
R2046 Vbias.n6896 Vbias.n1348 2025.26
R2047 Vbias.n6891 Vbias.n1350 2025.26
R2048 Vbias.n6891 Vbias.n1351 2025.26
R2049 Vbias.n6876 Vbias.n1362 2025.26
R2050 Vbias.n6877 Vbias.n1362 2025.26
R2051 Vbias.n6868 Vbias.n1363 2025.26
R2052 Vbias.n6868 Vbias.n1364 2025.26
R2053 Vbias.n6853 Vbias.n1375 2025.26
R2054 Vbias.n6854 Vbias.n1375 2025.26
R2055 Vbias.n6845 Vbias.n1376 2025.26
R2056 Vbias.n6845 Vbias.n1377 2025.26
R2057 Vbias.n1385 Vbias.n1384 2025.26
R2058 Vbias.n6838 Vbias.n1385 2025.26
R2059 Vbias.n6830 Vbias.n1391 2025.26
R2060 Vbias.n6829 Vbias.n1391 2025.26
R2061 Vbias.n1556 Vbias.n1555 2025.26
R2062 Vbias.n1556 Vbias.n1400 2025.26
R2063 Vbias.n6043 Vbias.n1558 2025.26
R2064 Vbias.n6043 Vbias.n1559 2025.26
R2065 Vbias.n6039 Vbias.n1559 2025.26
R2066 Vbias.n6039 Vbias.n1558 2025.26
R2067 Vbias.n6036 Vbias.n1561 2025.26
R2068 Vbias.n6036 Vbias.n1562 2025.26
R2069 Vbias.n6018 Vbias.n1573 2025.26
R2070 Vbias.n6019 Vbias.n1573 2025.26
R2071 Vbias.n6010 Vbias.n1574 2025.26
R2072 Vbias.n6010 Vbias.n1575 2025.26
R2073 Vbias.n5995 Vbias.n1586 2025.26
R2074 Vbias.n5996 Vbias.n1586 2025.26
R2075 Vbias.n5987 Vbias.n1587 2025.26
R2076 Vbias.n5987 Vbias.n1588 2025.26
R2077 Vbias.n1596 Vbias.n1595 2025.26
R2078 Vbias.n5980 Vbias.n1596 2025.26
R2079 Vbias.n5972 Vbias.n1602 2025.26
R2080 Vbias.n5971 Vbias.n1602 2025.26
R2081 Vbias.n1637 Vbias.n1636 2025.26
R2082 Vbias.n1637 Vbias.n1611 2025.26
R2083 Vbias.n5344 Vbias.n5338 2025.26
R2084 Vbias.n5344 Vbias.n5339 2025.26
R2085 Vbias.n5348 Vbias.n5339 2025.26
R2086 Vbias.n5348 Vbias.n5338 2025.26
R2087 Vbias.n5353 Vbias.n5337 2025.26
R2088 Vbias.n5352 Vbias.n5337 2025.26
R2089 Vbias.n5364 Vbias.n5317 2025.26
R2090 Vbias.n5364 Vbias.n5316 2025.26
R2091 Vbias.n5375 Vbias.n5314 2025.26
R2092 Vbias.n5374 Vbias.n5314 2025.26
R2093 Vbias.n5310 Vbias.n5308 2025.26
R2094 Vbias.n5308 Vbias.n5302 2025.26
R2095 Vbias.n5388 Vbias.n5296 2025.26
R2096 Vbias.n5296 Vbias.n5295 2025.26
R2097 Vbias.n5395 Vbias.n5288 2025.26
R2098 Vbias.n5395 Vbias.n5287 2025.26
R2099 Vbias.n5406 Vbias.n5285 2025.26
R2100 Vbias.n5405 Vbias.n5285 2025.26
R2101 Vbias.n5281 Vbias.n5279 2025.26
R2102 Vbias.n5279 Vbias.n5273 2025.26
R2103 Vbias.n5266 Vbias.n2297 2025.26
R2104 Vbias.n5265 Vbias.n2297 2025.26
R2105 Vbias.n5265 Vbias.n2296 2025.26
R2106 Vbias.n5266 Vbias.n2296 2025.26
R2107 Vbias.n5260 Vbias.n2298 2025.26
R2108 Vbias.n5260 Vbias.n2299 2025.26
R2109 Vbias.n5245 Vbias.n2310 2025.26
R2110 Vbias.n5246 Vbias.n2310 2025.26
R2111 Vbias.n5237 Vbias.n2311 2025.26
R2112 Vbias.n5237 Vbias.n2312 2025.26
R2113 Vbias.n5222 Vbias.n2323 2025.26
R2114 Vbias.n5223 Vbias.n2323 2025.26
R2115 Vbias.n5214 Vbias.n2324 2025.26
R2116 Vbias.n5214 Vbias.n2325 2025.26
R2117 Vbias.n2333 Vbias.n2332 2025.26
R2118 Vbias.n5207 Vbias.n2333 2025.26
R2119 Vbias.n5199 Vbias.n2339 2025.26
R2120 Vbias.n5198 Vbias.n2339 2025.26
R2121 Vbias.n2369 Vbias.n2368 2025.26
R2122 Vbias.n2369 Vbias.n2348 2025.26
R2123 Vbias.n2512 Vbias.n2506 2025.26
R2124 Vbias.n2512 Vbias.n2507 2025.26
R2125 Vbias.n2516 Vbias.n2507 2025.26
R2126 Vbias.n2516 Vbias.n2506 2025.26
R2127 Vbias.n2521 Vbias.n2505 2025.26
R2128 Vbias.n2520 Vbias.n2505 2025.26
R2129 Vbias.n2532 Vbias.n2485 2025.26
R2130 Vbias.n2532 Vbias.n2484 2025.26
R2131 Vbias.n2543 Vbias.n2482 2025.26
R2132 Vbias.n2542 Vbias.n2482 2025.26
R2133 Vbias.n2478 Vbias.n2476 2025.26
R2134 Vbias.n2476 Vbias.n2470 2025.26
R2135 Vbias.n2556 Vbias.n2464 2025.26
R2136 Vbias.n2464 Vbias.n2463 2025.26
R2137 Vbias.n2563 Vbias.n2456 2025.26
R2138 Vbias.n2563 Vbias.n2455 2025.26
R2139 Vbias.n2574 Vbias.n2453 2025.26
R2140 Vbias.n2573 Vbias.n2453 2025.26
R2141 Vbias.n2449 Vbias.n2447 2025.26
R2142 Vbias.n2447 Vbias.n2441 2025.26
R2143 Vbias.n5041 Vbias.n2432 2025.26
R2144 Vbias.n5040 Vbias.n2432 2025.26
R2145 Vbias.n5056 Vbias.n2417 2025.26
R2146 Vbias.n5056 Vbias.n2418 2025.26
R2147 Vbias.n3842 Vbias.n3816 2025.26
R2148 Vbias.n3841 Vbias.n3816 2025.26
R2149 Vbias.n3854 Vbias.n3792 2025.26
R2150 Vbias.n3854 Vbias.n3791 2025.26
R2151 Vbias.n3880 Vbias.n3858 2025.26
R2152 Vbias.n3858 Vbias.n3857 2025.26
R2153 Vbias.n3866 Vbias.n3779 2025.26
R2154 Vbias.n3866 Vbias.n3863 2025.26
R2155 Vbias.n3861 Vbias.n3772 2025.26
R2156 Vbias.n3861 Vbias.n3773 2025.26
R2157 Vbias.n3892 Vbias.n3773 2025.26
R2158 Vbias.n3892 Vbias.n3772 2025.26
R2159 Vbias.n3918 Vbias.n3769 2025.26
R2160 Vbias.n3917 Vbias.n3769 2025.26
R2161 Vbias.n3930 Vbias.n3745 2025.26
R2162 Vbias.n3930 Vbias.n3744 2025.26
R2163 Vbias.n3956 Vbias.n3740 2025.26
R2164 Vbias.n3955 Vbias.n3740 2025.26
R2165 Vbias.n3968 Vbias.n3716 2025.26
R2166 Vbias.n3968 Vbias.n3715 2025.26
R2167 Vbias.n3837 Vbias.n3817 2025.26
R2168 Vbias.n3837 Vbias.n3818 2025.26
R2169 Vbias.n3826 Vbias.n3790 2025.26
R2170 Vbias.n3795 Vbias.n3790 2025.26
R2171 Vbias.n3874 Vbias.n3788 2025.26
R2172 Vbias.n3874 Vbias.n3789 2025.26
R2173 Vbias.n3870 Vbias.n3868 2025.26
R2174 Vbias.n3868 Vbias.n3780 2025.26
R2175 Vbias.n3913 Vbias.n3770 2025.26
R2176 Vbias.n3913 Vbias.n3771 2025.26
R2177 Vbias.n3902 Vbias.n3743 2025.26
R2178 Vbias.n3748 Vbias.n3743 2025.26
R2179 Vbias.n3951 Vbias.n3741 2025.26
R2180 Vbias.n3951 Vbias.n3742 2025.26
R2181 Vbias.n3940 Vbias.n3714 2025.26
R2182 Vbias.n3719 Vbias.n3714 2025.26
R2183 Vbias.n3973 Vbias.n3713 2025.26
R2184 Vbias.n3972 Vbias.n3713 2025.26
R2185 Vbias.n3972 Vbias.n3712 2025.26
R2186 Vbias.n3973 Vbias.n3712 2025.26
R2187 Vbias.n3304 Vbias.n3278 2025.26
R2188 Vbias.n3303 Vbias.n3278 2025.26
R2189 Vbias.n3316 Vbias.n3254 2025.26
R2190 Vbias.n3316 Vbias.n3253 2025.26
R2191 Vbias.n3342 Vbias.n3320 2025.26
R2192 Vbias.n3320 Vbias.n3319 2025.26
R2193 Vbias.n3328 Vbias.n3241 2025.26
R2194 Vbias.n3328 Vbias.n3325 2025.26
R2195 Vbias.n3323 Vbias.n3234 2025.26
R2196 Vbias.n3323 Vbias.n3235 2025.26
R2197 Vbias.n3354 Vbias.n3235 2025.26
R2198 Vbias.n3354 Vbias.n3234 2025.26
R2199 Vbias.n3380 Vbias.n3231 2025.26
R2200 Vbias.n3379 Vbias.n3231 2025.26
R2201 Vbias.n3392 Vbias.n3207 2025.26
R2202 Vbias.n3392 Vbias.n3206 2025.26
R2203 Vbias.n3418 Vbias.n3202 2025.26
R2204 Vbias.n3417 Vbias.n3202 2025.26
R2205 Vbias.n3430 Vbias.n3178 2025.26
R2206 Vbias.n3430 Vbias.n3177 2025.26
R2207 Vbias.n3299 Vbias.n3279 2025.26
R2208 Vbias.n3299 Vbias.n3280 2025.26
R2209 Vbias.n3288 Vbias.n3252 2025.26
R2210 Vbias.n3257 Vbias.n3252 2025.26
R2211 Vbias.n3336 Vbias.n3250 2025.26
R2212 Vbias.n3336 Vbias.n3251 2025.26
R2213 Vbias.n3332 Vbias.n3330 2025.26
R2214 Vbias.n3330 Vbias.n3242 2025.26
R2215 Vbias.n3375 Vbias.n3232 2025.26
R2216 Vbias.n3375 Vbias.n3233 2025.26
R2217 Vbias.n3364 Vbias.n3205 2025.26
R2218 Vbias.n3210 Vbias.n3205 2025.26
R2219 Vbias.n3413 Vbias.n3203 2025.26
R2220 Vbias.n3413 Vbias.n3204 2025.26
R2221 Vbias.n3402 Vbias.n3176 2025.26
R2222 Vbias.n3181 Vbias.n3176 2025.26
R2223 Vbias.n3435 Vbias.n3175 2025.26
R2224 Vbias.n3434 Vbias.n3175 2025.26
R2225 Vbias.n3434 Vbias.n3174 2025.26
R2226 Vbias.n3435 Vbias.n3174 2025.26
R2227 Vbias.n3573 Vbias.n3547 2025.26
R2228 Vbias.n3572 Vbias.n3547 2025.26
R2229 Vbias.n3585 Vbias.n3523 2025.26
R2230 Vbias.n3585 Vbias.n3522 2025.26
R2231 Vbias.n3611 Vbias.n3589 2025.26
R2232 Vbias.n3589 Vbias.n3588 2025.26
R2233 Vbias.n3597 Vbias.n3510 2025.26
R2234 Vbias.n3597 Vbias.n3594 2025.26
R2235 Vbias.n3592 Vbias.n3503 2025.26
R2236 Vbias.n3592 Vbias.n3504 2025.26
R2237 Vbias.n3623 Vbias.n3504 2025.26
R2238 Vbias.n3623 Vbias.n3503 2025.26
R2239 Vbias.n3649 Vbias.n3500 2025.26
R2240 Vbias.n3648 Vbias.n3500 2025.26
R2241 Vbias.n3661 Vbias.n3476 2025.26
R2242 Vbias.n3661 Vbias.n3475 2025.26
R2243 Vbias.n3687 Vbias.n3471 2025.26
R2244 Vbias.n3686 Vbias.n3471 2025.26
R2245 Vbias.n3699 Vbias.n3447 2025.26
R2246 Vbias.n3699 Vbias.n3446 2025.26
R2247 Vbias.n3568 Vbias.n3548 2025.26
R2248 Vbias.n3568 Vbias.n3549 2025.26
R2249 Vbias.n3557 Vbias.n3521 2025.26
R2250 Vbias.n3526 Vbias.n3521 2025.26
R2251 Vbias.n3605 Vbias.n3519 2025.26
R2252 Vbias.n3605 Vbias.n3520 2025.26
R2253 Vbias.n3601 Vbias.n3599 2025.26
R2254 Vbias.n3599 Vbias.n3511 2025.26
R2255 Vbias.n3644 Vbias.n3501 2025.26
R2256 Vbias.n3644 Vbias.n3502 2025.26
R2257 Vbias.n3633 Vbias.n3474 2025.26
R2258 Vbias.n3479 Vbias.n3474 2025.26
R2259 Vbias.n3682 Vbias.n3472 2025.26
R2260 Vbias.n3682 Vbias.n3473 2025.26
R2261 Vbias.n3671 Vbias.n3445 2025.26
R2262 Vbias.n3450 Vbias.n3445 2025.26
R2263 Vbias.n3704 Vbias.n3444 2025.26
R2264 Vbias.n3703 Vbias.n3444 2025.26
R2265 Vbias.n3703 Vbias.n3443 2025.26
R2266 Vbias.n3704 Vbias.n3443 2025.26
R2267 Vbias.n4188 Vbias.n4070 2025.26
R2268 Vbias.n4187 Vbias.n4070 2025.26
R2269 Vbias.n4199 Vbias.n4050 2025.26
R2270 Vbias.n4199 Vbias.n4049 2025.26
R2271 Vbias.n4206 Vbias.n4203 2025.26
R2272 Vbias.n4203 Vbias.n4202 2025.26
R2273 Vbias.n4154 Vbias.n4039 2025.26
R2274 Vbias.n4154 Vbias.n4153 2025.26
R2275 Vbias.n4150 Vbias.n4032 2025.26
R2276 Vbias.n4150 Vbias.n4033 2025.26
R2277 Vbias.n4217 Vbias.n4033 2025.26
R2278 Vbias.n4217 Vbias.n4032 2025.26
R2279 Vbias.n4222 Vbias.n4028 2025.26
R2280 Vbias.n4221 Vbias.n4028 2025.26
R2281 Vbias.n4233 Vbias.n4008 2025.26
R2282 Vbias.n4233 Vbias.n4007 2025.26
R2283 Vbias.n4237 Vbias.n4002 2025.26
R2284 Vbias.n4238 Vbias.n4002 2025.26
R2285 Vbias.n4248 Vbias.n3983 2025.26
R2286 Vbias.n4247 Vbias.n3983 2025.26
R2287 Vbias.n4073 Vbias.n4071 2025.26
R2288 Vbias.n4185 Vbias.n4073 2025.26
R2289 Vbias.n4172 Vbias.n4048 2025.26
R2290 Vbias.n4176 Vbias.n4048 2025.26
R2291 Vbias.n4047 Vbias.n4045 2025.26
R2292 Vbias.n4047 Vbias.n4046 2025.26
R2293 Vbias.n4158 Vbias.n4156 2025.26
R2294 Vbias.n4156 Vbias.n4149 2025.26
R2295 Vbias.n4031 Vbias.n4029 2025.26
R2296 Vbias.n4031 Vbias.n4030 2025.26
R2297 Vbias.n4133 Vbias.n4006 2025.26
R2298 Vbias.n4129 Vbias.n4006 2025.26
R2299 Vbias.n4005 Vbias.n4003 2025.26
R2300 Vbias.n4005 Vbias.n4004 2025.26
R2301 Vbias.n4116 Vbias.n3987 2025.26
R2302 Vbias.n4116 Vbias.n3986 2025.26
R2303 Vbias.n4110 Vbias.n4106 2025.26
R2304 Vbias.n4109 Vbias.n4106 2025.26
R2305 Vbias.n4109 Vbias.n4105 2025.26
R2306 Vbias.n4110 Vbias.n4105 2025.26
R2307 Vbias.n4984 Vbias.n2608 2025.26
R2308 Vbias.n4983 Vbias.n2608 2025.26
R2309 Vbias.n2626 Vbias.n2625 2025.26
R2310 Vbias.n2626 Vbias.n2617 2025.26
R2311 Vbias.n4966 Vbias.n2622 2025.26
R2312 Vbias.n4965 Vbias.n2622 2025.26
R2313 Vbias.n4959 Vbias.n2631 2025.26
R2314 Vbias.n4958 Vbias.n2631 2025.26
R2315 Vbias.n4954 Vbias.n2632 2025.26
R2316 Vbias.n4954 Vbias.n2633 2025.26
R2317 Vbias.n4939 Vbias.n2645 2025.26
R2318 Vbias.n4940 Vbias.n2645 2025.26
R2319 Vbias.n4931 Vbias.n2646 2025.26
R2320 Vbias.n4931 Vbias.n2647 2025.26
R2321 Vbias.n4917 Vbias.n2659 2025.26
R2322 Vbias.n4918 Vbias.n2659 2025.26
R2323 Vbias.n4909 Vbias.n2660 2025.26
R2324 Vbias.n4909 Vbias.n2661 2025.26
R2325 Vbias.n4905 Vbias.n2661 2025.26
R2326 Vbias.n4905 Vbias.n2660 2025.26
R2327 Vbias.n3034 Vbias.n3008 2025.26
R2328 Vbias.n3033 Vbias.n3008 2025.26
R2329 Vbias.n3046 Vbias.n2984 2025.26
R2330 Vbias.n3046 Vbias.n2983 2025.26
R2331 Vbias.n3072 Vbias.n3050 2025.26
R2332 Vbias.n3050 Vbias.n3049 2025.26
R2333 Vbias.n3058 Vbias.n2971 2025.26
R2334 Vbias.n3058 Vbias.n3055 2025.26
R2335 Vbias.n3053 Vbias.n2964 2025.26
R2336 Vbias.n3053 Vbias.n2965 2025.26
R2337 Vbias.n3084 Vbias.n2965 2025.26
R2338 Vbias.n3084 Vbias.n2964 2025.26
R2339 Vbias.n3110 Vbias.n2961 2025.26
R2340 Vbias.n3109 Vbias.n2961 2025.26
R2341 Vbias.n3122 Vbias.n2937 2025.26
R2342 Vbias.n3122 Vbias.n2936 2025.26
R2343 Vbias.n3148 Vbias.n2932 2025.26
R2344 Vbias.n3147 Vbias.n2932 2025.26
R2345 Vbias.n3160 Vbias.n2908 2025.26
R2346 Vbias.n3160 Vbias.n2907 2025.26
R2347 Vbias.n3029 Vbias.n3009 2025.26
R2348 Vbias.n3029 Vbias.n3010 2025.26
R2349 Vbias.n3018 Vbias.n2982 2025.26
R2350 Vbias.n2987 Vbias.n2982 2025.26
R2351 Vbias.n3066 Vbias.n2980 2025.26
R2352 Vbias.n3066 Vbias.n2981 2025.26
R2353 Vbias.n3062 Vbias.n3060 2025.26
R2354 Vbias.n3060 Vbias.n2972 2025.26
R2355 Vbias.n3105 Vbias.n2962 2025.26
R2356 Vbias.n3105 Vbias.n2963 2025.26
R2357 Vbias.n3094 Vbias.n2935 2025.26
R2358 Vbias.n2940 Vbias.n2935 2025.26
R2359 Vbias.n3143 Vbias.n2933 2025.26
R2360 Vbias.n3143 Vbias.n2934 2025.26
R2361 Vbias.n3132 Vbias.n2906 2025.26
R2362 Vbias.n2911 Vbias.n2906 2025.26
R2363 Vbias.n3165 Vbias.n2904 2025.26
R2364 Vbias.n3164 Vbias.n2904 2025.26
R2365 Vbias.n3164 Vbias.n2903 2025.26
R2366 Vbias.n3165 Vbias.n2903 2025.26
R2367 Vbias.n4710 Vbias.n2769 2025.26
R2368 Vbias.n4709 Vbias.n2769 2025.26
R2369 Vbias.n4722 Vbias.n2745 2025.26
R2370 Vbias.n4722 Vbias.n2744 2025.26
R2371 Vbias.n4748 Vbias.n4726 2025.26
R2372 Vbias.n4726 Vbias.n4725 2025.26
R2373 Vbias.n4734 Vbias.n2732 2025.26
R2374 Vbias.n4734 Vbias.n4731 2025.26
R2375 Vbias.n4729 Vbias.n2725 2025.26
R2376 Vbias.n4729 Vbias.n2726 2025.26
R2377 Vbias.n4760 Vbias.n2726 2025.26
R2378 Vbias.n4760 Vbias.n2725 2025.26
R2379 Vbias.n4786 Vbias.n2722 2025.26
R2380 Vbias.n4785 Vbias.n2722 2025.26
R2381 Vbias.n4798 Vbias.n2698 2025.26
R2382 Vbias.n4798 Vbias.n2697 2025.26
R2383 Vbias.n4824 Vbias.n2693 2025.26
R2384 Vbias.n4823 Vbias.n2693 2025.26
R2385 Vbias.n4836 Vbias.n2669 2025.26
R2386 Vbias.n4836 Vbias.n2668 2025.26
R2387 Vbias.n4705 Vbias.n2770 2025.26
R2388 Vbias.n4705 Vbias.n2771 2025.26
R2389 Vbias.n4694 Vbias.n2743 2025.26
R2390 Vbias.n2748 Vbias.n2743 2025.26
R2391 Vbias.n4742 Vbias.n2741 2025.26
R2392 Vbias.n4742 Vbias.n2742 2025.26
R2393 Vbias.n4738 Vbias.n4736 2025.26
R2394 Vbias.n4736 Vbias.n2733 2025.26
R2395 Vbias.n4781 Vbias.n2723 2025.26
R2396 Vbias.n4781 Vbias.n2724 2025.26
R2397 Vbias.n4770 Vbias.n2696 2025.26
R2398 Vbias.n2701 Vbias.n2696 2025.26
R2399 Vbias.n4819 Vbias.n2694 2025.26
R2400 Vbias.n4819 Vbias.n2695 2025.26
R2401 Vbias.n4808 Vbias.n2667 2025.26
R2402 Vbias.n2672 Vbias.n2667 2025.26
R2403 Vbias.n4839 Vbias.n2664 2025.26
R2404 Vbias.n4839 Vbias.n2665 2025.26
R2405 Vbias.n4843 Vbias.n2665 2025.26
R2406 Vbias.n4843 Vbias.n2664 2025.26
R2407 Vbias.n4680 Vbias.n4551 2025.26
R2408 Vbias.n4680 Vbias.n4552 2025.26
R2409 Vbias.n4672 Vbias.n4560 2025.26
R2410 Vbias.n4672 Vbias.n4558 2025.26
R2411 Vbias.n6600 Vbias.n6212 2025.26
R2412 Vbias.n6600 Vbias.n6210 2025.26
R2413 Vbias.n6609 Vbias.n6203 2025.26
R2414 Vbias.n6609 Vbias.n6202 2025.26
R2415 Vbias.n6612 Vbias.n6195 2025.26
R2416 Vbias.n6612 Vbias.n6193 2025.26
R2417 Vbias.n6619 Vbias.n6189 2025.26
R2418 Vbias.n6619 Vbias.n6188 2025.26
R2419 Vbias.n6622 Vbias.n6165 2025.26
R2420 Vbias.n6622 Vbias.n6163 2025.26
R2421 Vbias.n6186 Vbias.n6163 2025.26
R2422 Vbias.n6186 Vbias.n6165 2025.26
R2423 Vbias.n6184 Vbias.n6183 2025.26
R2424 Vbias.n6184 Vbias.n6160 2025.26
R2425 Vbias.n6170 Vbias.n6156 2025.26
R2426 Vbias.n6172 Vbias.n6170 2025.26
R2427 Vbias.n6533 Vbias.n6449 2025.26
R2428 Vbias.n6533 Vbias.n6447 2025.26
R2429 Vbias.n6542 Vbias.n6440 2025.26
R2430 Vbias.n6542 Vbias.n6439 2025.26
R2431 Vbias.n6545 Vbias.n6432 2025.26
R2432 Vbias.n6545 Vbias.n6430 2025.26
R2433 Vbias.n6552 Vbias.n6426 2025.26
R2434 Vbias.n6552 Vbias.n6425 2025.26
R2435 Vbias.n6555 Vbias.n6383 2025.26
R2436 Vbias.n6555 Vbias.n6381 2025.26
R2437 Vbias.n6423 Vbias.n6381 2025.26
R2438 Vbias.n6423 Vbias.n6383 2025.26
R2439 Vbias.n6421 Vbias.n6420 2025.26
R2440 Vbias.n6421 Vbias.n6378 2025.26
R2441 Vbias.n6407 Vbias.n6374 2025.26
R2442 Vbias.n6409 Vbias.n6407 2025.26
R2443 Vbias.n6404 Vbias.n6403 2025.26
R2444 Vbias.n6404 Vbias.n6370 2025.26
R2445 Vbias.n6390 Vbias.n6366 2025.26
R2446 Vbias.n6392 Vbias.n6390 2025.26
R2447 Vbias.n7546 Vbias.n903 2025.26
R2448 Vbias.n7546 Vbias.n901 2025.26
R2449 Vbias.n7555 Vbias.n894 2025.26
R2450 Vbias.n7555 Vbias.n893 2025.26
R2451 Vbias.n7558 Vbias.n886 2025.26
R2452 Vbias.n7558 Vbias.n884 2025.26
R2453 Vbias.n7565 Vbias.n880 2025.26
R2454 Vbias.n7565 Vbias.n879 2025.26
R2455 Vbias.n7568 Vbias.n878 2025.26
R2456 Vbias.n7568 Vbias.n876 2025.26
R2457 Vbias.n6475 Vbias.n876 2025.26
R2458 Vbias.n6475 Vbias.n878 2025.26
R2459 Vbias.n6480 Vbias.n6478 2025.26
R2460 Vbias.n6478 Vbias.n873 2025.26
R2461 Vbias.n6489 Vbias.n869 2025.26
R2462 Vbias.n6489 Vbias.n6488 2025.26
R2463 Vbias.n6494 Vbias.n6492 2025.26
R2464 Vbias.n6492 Vbias.n865 2025.26
R2465 Vbias.n6503 Vbias.n861 2025.26
R2466 Vbias.n6503 Vbias.n6502 2025.26
R2467 Vbias.n7403 Vbias.n7399 2025.26
R2468 Vbias.n7414 Vbias.n7381 2025.26
R2469 Vbias.n7414 Vbias.n7380 2025.26
R2470 Vbias.n7421 Vbias.n7418 2025.26
R2471 Vbias.n7418 Vbias.n7417 2025.26
R2472 Vbias.n7377 Vbias.n7369 2025.26
R2473 Vbias.n7379 Vbias.n7377 2025.26
R2474 Vbias.n7374 Vbias.n7362 2025.26
R2475 Vbias.n7374 Vbias.n7363 2025.26
R2476 Vbias.n7432 Vbias.n7363 2025.26
R2477 Vbias.n7432 Vbias.n7362 2025.26
R2478 Vbias.n7437 Vbias.n7361 2025.26
R2479 Vbias.n7436 Vbias.n7361 2025.26
R2480 Vbias.n7448 Vbias.n7343 2025.26
R2481 Vbias.n7448 Vbias.n7342 2025.26
R2482 Vbias.n7452 Vbias.n7341 2025.26
R2483 Vbias.n7453 Vbias.n7341 2025.26
R2484 Vbias.n7463 Vbias.n7327 2025.26
R2485 Vbias.n7462 Vbias.n7327 2025.26
R2486 Vbias.n6143 Vbias.n6141 2025.26
R2487 Vbias.n6141 Vbias.n6136 2025.26
R2488 Vbias.n6638 Vbias.n6149 2025.26
R2489 Vbias.n6637 Vbias.n6149 2025.26
R2490 Vbias.n6130 Vbias.n1501 2025.26
R2491 Vbias.n1505 Vbias.n1501 2025.26
R2492 Vbias.n6130 Vbias.n1502 2025.26
R2493 Vbias.n1505 Vbias.n1502 2025.26
R2494 Vbias.n2058 Vbias.n1704 2025.26
R2495 Vbias.n2047 Vbias.n1720 2025.26
R2496 Vbias.n2046 Vbias.n1720 2025.26
R2497 Vbias.n2058 Vbias.n1705 2025.26
R2498 Vbias.n6681 Vbias.n6680 2025.26
R2499 Vbias.n6680 Vbias.n1457 2025.26
R2500 Vbias.n6688 Vbias.n6687 2025.26
R2501 Vbias.n6688 Vbias.n1451 2025.26
R2502 Vbias.n8008 Vbias.n8007 1937.25
R2503 Vbias.n6261 Vbias.n6252 1847.07
R2504 Vbias.n7615 Vbias.n7614 1847.07
R2505 Vbias.n7493 Vbias.n7492 1847.07
R2506 Vbias.n7287 Vbias.n7286 1847.07
R2507 Vbias.n7015 Vbias.n7014 1797.97
R2508 Vbias.n5918 Vbias.n5917 1797.97
R2509 Vbias.n5121 Vbias.n5120 1797.97
R2510 Vbias.n8077 Vbias.n5 1711.26
R2511 Vbias.n7801 Vbias.t50 1477.9
R2512 Vbias.n585 Vbias.t50 1477.9
R2513 Vbias.n585 Vbias.t600 1477.9
R2514 Vbias.n595 Vbias.t600 1477.9
R2515 Vbias.t441 Vbias.n595 1477.9
R2516 Vbias.n7790 Vbias.t441 1477.9
R2517 Vbias.n7789 Vbias.t275 1477.9
R2518 Vbias.n609 Vbias.t275 1477.9
R2519 Vbias.n609 Vbias.t614 1477.9
R2520 Vbias.n619 Vbias.t614 1477.9
R2521 Vbias.t681 Vbias.n619 1477.9
R2522 Vbias.n7778 Vbias.t681 1477.9
R2523 Vbias.n7777 Vbias.t817 1477.9
R2524 Vbias.n633 Vbias.t817 1477.9
R2525 Vbias.n634 Vbias.t855 1477.9
R2526 Vbias.n642 Vbias.t855 1477.9
R2527 Vbias.t848 Vbias.n642 1477.9
R2528 Vbias.n7765 Vbias.t848 1477.9
R2529 Vbias.n7764 Vbias.t273 1477.9
R2530 Vbias.n656 Vbias.t273 1477.9
R2531 Vbias.n656 Vbias.t721 1477.9
R2532 Vbias.n666 Vbias.t721 1477.9
R2533 Vbias.t786 Vbias.n666 1477.9
R2534 Vbias.n7753 Vbias.t786 1477.9
R2535 Vbias.n7870 Vbias.t112 1477.9
R2536 Vbias.n471 Vbias.t112 1477.9
R2537 Vbias.n471 Vbias.t161 1477.9
R2538 Vbias.n481 Vbias.t161 1477.9
R2539 Vbias.t327 Vbias.n481 1477.9
R2540 Vbias.n7859 Vbias.t327 1477.9
R2541 Vbias.n7858 Vbias.t218 1477.9
R2542 Vbias.n495 Vbias.t218 1477.9
R2543 Vbias.n495 Vbias.t547 1477.9
R2544 Vbias.n505 Vbias.t547 1477.9
R2545 Vbias.t153 Vbias.n505 1477.9
R2546 Vbias.n7847 Vbias.t153 1477.9
R2547 Vbias.n7846 Vbias.t397 1477.9
R2548 Vbias.n519 Vbias.t397 1477.9
R2549 Vbias.n520 Vbias.t889 1477.9
R2550 Vbias.n528 Vbias.t889 1477.9
R2551 Vbias.t741 Vbias.n528 1477.9
R2552 Vbias.n7834 Vbias.t741 1477.9
R2553 Vbias.n7833 Vbias.t184 1477.9
R2554 Vbias.n542 Vbias.t184 1477.9
R2555 Vbias.n542 Vbias.t505 1477.9
R2556 Vbias.n552 Vbias.t505 1477.9
R2557 Vbias.t823 Vbias.n552 1477.9
R2558 Vbias.n7822 Vbias.t823 1477.9
R2559 Vbias.n7936 Vbias.t86 1477.9
R2560 Vbias.n365 Vbias.t86 1477.9
R2561 Vbias.n365 Vbias.t673 1477.9
R2562 Vbias.n375 Vbias.t673 1477.9
R2563 Vbias.t443 Vbias.n375 1477.9
R2564 Vbias.n7925 Vbias.t443 1477.9
R2565 Vbias.n7924 Vbias.t172 1477.9
R2566 Vbias.n389 Vbias.t172 1477.9
R2567 Vbias.n389 Vbias.t797 1477.9
R2568 Vbias.n399 Vbias.t797 1477.9
R2569 Vbias.t430 Vbias.n399 1477.9
R2570 Vbias.n7913 Vbias.t430 1477.9
R2571 Vbias.n7912 Vbias.t590 1477.9
R2572 Vbias.n413 Vbias.t590 1477.9
R2573 Vbias.n414 Vbias.t320 1477.9
R2574 Vbias.n422 Vbias.t320 1477.9
R2575 Vbias.t633 Vbias.n422 1477.9
R2576 Vbias.n7900 Vbias.t633 1477.9
R2577 Vbias.n7899 Vbias.t190 1477.9
R2578 Vbias.n436 Vbias.t190 1477.9
R2579 Vbias.n436 Vbias.t886 1477.9
R2580 Vbias.n446 Vbias.t886 1477.9
R2581 Vbias.t774 Vbias.n446 1477.9
R2582 Vbias.n7888 Vbias.t774 1477.9
R2583 Vbias.t70 Vbias.n86 1477.9
R2584 Vbias.t70 Vbias.n242 1477.9
R2585 Vbias.n242 Vbias.t495 1477.9
R2586 Vbias.n267 Vbias.t495 1477.9
R2587 Vbias.t866 Vbias.n267 1477.9
R2588 Vbias.n268 Vbias.t866 1477.9
R2589 Vbias.t206 Vbias.n223 1477.9
R2590 Vbias.t206 Vbias.n224 1477.9
R2591 Vbias.n224 Vbias.t309 1477.9
R2592 Vbias.n284 Vbias.t309 1477.9
R2593 Vbias.t455 Vbias.n284 1477.9
R2594 Vbias.n287 Vbias.t455 1477.9
R2595 Vbias.n286 Vbias.t863 1477.9
R2596 Vbias.n298 Vbias.t863 1477.9
R2597 Vbias.n299 Vbias.t802 1477.9
R2598 Vbias.n306 Vbias.t802 1477.9
R2599 Vbias.t859 Vbias.n306 1477.9
R2600 Vbias.n307 Vbias.t859 1477.9
R2601 Vbias.t247 Vbias.n190 1477.9
R2602 Vbias.t247 Vbias.n191 1477.9
R2603 Vbias.n191 Vbias.t780 1477.9
R2604 Vbias.n323 Vbias.t780 1477.9
R2605 Vbias.t4 Vbias.n323 1477.9
R2606 Vbias.n350 Vbias.t4 1477.9
R2607 Vbias.t796 Vbias.n1152 1477.9
R2608 Vbias.n1268 Vbias.t796 1477.9
R2609 Vbias.n1268 Vbias.t704 1477.9
R2610 Vbias.t704 Vbias.n1178 1477.9
R2611 Vbias.t188 Vbias.n1178 1477.9
R2612 Vbias.t188 Vbias.n1256 1477.9
R2613 Vbias.n1255 Vbias.t429 1477.9
R2614 Vbias.n1248 Vbias.t429 1477.9
R2615 Vbias.n1248 Vbias.t315 1477.9
R2616 Vbias.t315 Vbias.n1190 1477.9
R2617 Vbias.t126 Vbias.n1203 1477.9
R2618 Vbias.n1237 Vbias.t126 1477.9
R2619 Vbias.n1237 Vbias.t874 1477.9
R2620 Vbias.t874 Vbias.n1207 1477.9
R2621 Vbias.t255 Vbias.n1207 1477.9
R2622 Vbias.t255 Vbias.n1225 1477.9
R2623 Vbias.n1224 Vbias.t336 1477.9
R2624 Vbias.t336 Vbias.n1082 1477.9
R2625 Vbias.t298 Vbias.n1082 1477.9
R2626 Vbias.n7210 Vbias.t298 1477.9
R2627 Vbias.n7210 Vbias.t104 1477.9
R2628 Vbias.n7217 Vbias.t104 1477.9
R2629 Vbias.n7218 Vbias.t688 1477.9
R2630 Vbias.n7224 Vbias.t688 1477.9
R2631 Vbias.t885 Vbias.n1339 1477.9
R2632 Vbias.n7001 Vbias.t885 1477.9
R2633 Vbias.n7001 Vbias.t606 1477.9
R2634 Vbias.t606 Vbias.n6911 1477.9
R2635 Vbias.t40 Vbias.n6911 1477.9
R2636 Vbias.t40 Vbias.n6989 1477.9
R2637 Vbias.n6988 Vbias.t145 1477.9
R2638 Vbias.n6981 Vbias.t145 1477.9
R2639 Vbias.n6981 Vbias.t534 1477.9
R2640 Vbias.t534 Vbias.n6923 1477.9
R2641 Vbias.t544 Vbias.n6936 1477.9
R2642 Vbias.n6970 Vbias.t544 1477.9
R2643 Vbias.n6970 Vbias.t378 1477.9
R2644 Vbias.t378 Vbias.n6940 1477.9
R2645 Vbias.t66 Vbias.n6940 1477.9
R2646 Vbias.t66 Vbias.n6958 1477.9
R2647 Vbias.n6957 Vbias.t497 1477.9
R2648 Vbias.t497 Vbias.n1163 1477.9
R2649 Vbias.t842 Vbias.n1163 1477.9
R2650 Vbias.n7106 Vbias.t842 1477.9
R2651 Vbias.n7106 Vbias.t196 1477.9
R2652 Vbias.n7113 Vbias.t196 1477.9
R2653 Vbias.n7114 Vbias.t509 1477.9
R2654 Vbias.n7120 Vbias.t509 1477.9
R2655 Vbias.n1557 Vbias.t361 1477.9
R2656 Vbias.t361 Vbias.n1397 1477.9
R2657 Vbias.t160 Vbias.n1397 1477.9
R2658 Vbias.t160 Vbias.n1392 1477.9
R2659 Vbias.t118 Vbias.n1392 1477.9
R2660 Vbias.t118 Vbias.n1393 1477.9
R2661 Vbias.t754 Vbias.n1383 1477.9
R2662 Vbias.n6839 Vbias.t754 1477.9
R2663 Vbias.n6839 Vbias.t488 1477.9
R2664 Vbias.n6846 Vbias.t488 1477.9
R2665 Vbias.t492 Vbias.n6847 1477.9
R2666 Vbias.t492 Vbias.n1370 1477.9
R2667 Vbias.t579 Vbias.n1370 1477.9
R2668 Vbias.n6862 Vbias.t579 1477.9
R2669 Vbias.n6862 Vbias.t122 1477.9
R2670 Vbias.n6869 Vbias.t122 1477.9
R2671 Vbias.t380 Vbias.n6870 1477.9
R2672 Vbias.t380 Vbias.n1357 1477.9
R2673 Vbias.t1 Vbias.n1357 1477.9
R2674 Vbias.n6885 Vbias.t1 1477.9
R2675 Vbias.n6885 Vbias.t222 1477.9
R2676 Vbias.n6892 Vbias.t222 1477.9
R2677 Vbias.t420 Vbias.n6893 1477.9
R2678 Vbias.t420 Vbias.n1340 1477.9
R2679 Vbias.n1638 Vbias.t680 1477.9
R2680 Vbias.t680 Vbias.n1608 1477.9
R2681 Vbias.t569 Vbias.n1608 1477.9
R2682 Vbias.t569 Vbias.n1603 1477.9
R2683 Vbias.t60 Vbias.n1603 1477.9
R2684 Vbias.t60 Vbias.n1604 1477.9
R2685 Vbias.t456 Vbias.n1594 1477.9
R2686 Vbias.n5981 Vbias.t456 1477.9
R2687 Vbias.n5981 Vbias.t318 1477.9
R2688 Vbias.n5988 Vbias.t318 1477.9
R2689 Vbias.t752 Vbias.n5989 1477.9
R2690 Vbias.t752 Vbias.n1581 1477.9
R2691 Vbias.t852 Vbias.n1581 1477.9
R2692 Vbias.n6004 Vbias.t852 1477.9
R2693 Vbias.n6004 Vbias.t94 1477.9
R2694 Vbias.n6011 Vbias.t94 1477.9
R2695 Vbias.t660 Vbias.n6012 1477.9
R2696 Vbias.t660 Vbias.n1568 1477.9
R2697 Vbias.t732 Vbias.n1568 1477.9
R2698 Vbias.n6030 Vbias.t732 1477.9
R2699 Vbias.n6030 Vbias.t243 1477.9
R2700 Vbias.n6037 Vbias.t243 1477.9
R2701 Vbias.n6038 Vbias.t728 1477.9
R2702 Vbias.n6044 Vbias.t728 1477.9
R2703 Vbias.t532 Vbias.n5278 1477.9
R2704 Vbias.n5409 Vbias.t532 1477.9
R2705 Vbias.n5409 Vbias.t635 1477.9
R2706 Vbias.t635 Vbias.n5282 1477.9
R2707 Vbias.t98 Vbias.n5282 1477.9
R2708 Vbias.t98 Vbias.n5397 1477.9
R2709 Vbias.n5396 Vbias.t413 1477.9
R2710 Vbias.n5389 Vbias.t413 1477.9
R2711 Vbias.n5389 Vbias.t404 1477.9
R2712 Vbias.t404 Vbias.n5294 1477.9
R2713 Vbias.t13 Vbias.n5307 1477.9
R2714 Vbias.n5378 Vbias.t13 1477.9
R2715 Vbias.n5378 Vbias.t642 1477.9
R2716 Vbias.t642 Vbias.n5311 1477.9
R2717 Vbias.t22 Vbias.n5311 1477.9
R2718 Vbias.t22 Vbias.n5366 1477.9
R2719 Vbias.n5365 Vbias.t814 1477.9
R2720 Vbias.n5323 Vbias.t814 1477.9
R2721 Vbias.t154 Vbias.n5323 1477.9
R2722 Vbias.t154 Vbias.n5324 1477.9
R2723 Vbias.t194 Vbias.n5324 1477.9
R2724 Vbias.t194 Vbias.n5350 1477.9
R2725 Vbias.n5349 Vbias.t742 1477.9
R2726 Vbias.t742 Vbias.n1639 1477.9
R2727 Vbias.n2370 Vbias.t765 1477.9
R2728 Vbias.t765 Vbias.n2345 1477.9
R2729 Vbias.t347 Vbias.n2345 1477.9
R2730 Vbias.t347 Vbias.n2340 1477.9
R2731 Vbias.t54 Vbias.n2340 1477.9
R2732 Vbias.t54 Vbias.n2341 1477.9
R2733 Vbias.t711 Vbias.n2331 1477.9
R2734 Vbias.n5208 Vbias.t711 1477.9
R2735 Vbias.n5208 Vbias.t664 1477.9
R2736 Vbias.n5215 Vbias.t664 1477.9
R2737 Vbias.t685 Vbias.n5216 1477.9
R2738 Vbias.t685 Vbias.n2318 1477.9
R2739 Vbias.t531 Vbias.n2318 1477.9
R2740 Vbias.n5231 Vbias.t531 1477.9
R2741 Vbias.n5231 Vbias.t28 1477.9
R2742 Vbias.n5238 Vbias.t28 1477.9
R2743 Vbias.t394 Vbias.n5239 1477.9
R2744 Vbias.t394 Vbias.n2305 1477.9
R2745 Vbias.t139 Vbias.n2305 1477.9
R2746 Vbias.n5254 Vbias.t139 1477.9
R2747 Vbias.n5254 Vbias.t216 1477.9
R2748 Vbias.n5261 Vbias.t216 1477.9
R2749 Vbias.t707 Vbias.n5262 1477.9
R2750 Vbias.t707 Vbias.n5263 1477.9
R2751 Vbias.t851 Vbias.n2446 1477.9
R2752 Vbias.n2577 Vbias.t851 1477.9
R2753 Vbias.n2577 Vbias.t762 1477.9
R2754 Vbias.t762 Vbias.n2450 1477.9
R2755 Vbias.t38 Vbias.n2450 1477.9
R2756 Vbias.t38 Vbias.n2565 1477.9
R2757 Vbias.n2564 Vbias.t546 1477.9
R2758 Vbias.n2557 Vbias.t546 1477.9
R2759 Vbias.n2557 Vbias.t690 1477.9
R2760 Vbias.t690 Vbias.n2462 1477.9
R2761 Vbias.t9 Vbias.n2475 1477.9
R2762 Vbias.n2546 Vbias.t9 1477.9
R2763 Vbias.n2546 Vbias.t598 1477.9
R2764 Vbias.t598 Vbias.n2479 1477.9
R2765 Vbias.t108 Vbias.n2479 1477.9
R2766 Vbias.t108 Vbias.n2534 1477.9
R2767 Vbias.n2533 Vbias.t480 1477.9
R2768 Vbias.n2491 Vbias.t480 1477.9
R2769 Vbias.t603 Vbias.n2491 1477.9
R2770 Vbias.t603 Vbias.n2492 1477.9
R2771 Vbias.t263 Vbias.n2492 1477.9
R2772 Vbias.t263 Vbias.n2518 1477.9
R2773 Vbias.n2517 Vbias.t601 1477.9
R2774 Vbias.t601 Vbias.n2371 1477.9
R2775 Vbias.n4550 Vbias.t536 1477.9
R2776 Vbias.n4414 Vbias.t536 1477.9
R2777 Vbias.t303 Vbias.n4414 1477.9
R2778 Vbias.t303 Vbias.n4415 1477.9
R2779 Vbias.t110 Vbias.n4415 1477.9
R2780 Vbias.t110 Vbias.n4535 1477.9
R2781 Vbias.n4534 Vbias.t804 1477.9
R2782 Vbias.n4433 Vbias.t804 1477.9
R2783 Vbias.t300 Vbias.n4433 1477.9
R2784 Vbias.t300 Vbias.n4434 1477.9
R2785 Vbias.t454 Vbias.n4452 1477.9
R2786 Vbias.t454 Vbias.n4446 1477.9
R2787 Vbias.t474 Vbias.n4446 1477.9
R2788 Vbias.t474 Vbias.n4447 1477.9
R2789 Vbias.t58 Vbias.n4447 1477.9
R2790 Vbias.t58 Vbias.n4460 1477.9
R2791 Vbias.t408 Vbias.n4474 1477.9
R2792 Vbias.t408 Vbias.n4468 1477.9
R2793 Vbias.t226 Vbias.n4468 1477.9
R2794 Vbias.t226 Vbias.n4469 1477.9
R2795 Vbias.t180 Vbias.n4469 1477.9
R2796 Vbias.t180 Vbias.n4482 1477.9
R2797 Vbias.t824 Vbias.n4490 1477.9
R2798 Vbias.n4491 Vbias.t824 1477.9
R2799 Vbias.t64 Vbias.n917 1477.9
R2800 Vbias.t64 Vbias.n7329 1477.9
R2801 Vbias.t873 Vbias.n7329 1477.9
R2802 Vbias.t873 Vbias.n7335 1477.9
R2803 Vbias.t393 Vbias.n7335 1477.9
R2804 Vbias.t393 Vbias.n7450 1477.9
R2805 Vbias.n7449 Vbias.t192 1477.9
R2806 Vbias.n7351 Vbias.t192 1477.9
R2807 Vbias.t146 Vbias.n7351 1477.9
R2808 Vbias.t146 Vbias.n7352 1477.9
R2809 Vbias.t302 Vbias.n7352 1477.9
R2810 Vbias.t302 Vbias.n7434 1477.9
R2811 Vbias.n7433 Vbias.t588 1477.9
R2812 Vbias.n7375 Vbias.t588 1477.9
R2813 Vbias.t667 Vbias.n7376 1477.9
R2814 Vbias.n7422 Vbias.t667 1477.9
R2815 Vbias.n7422 Vbias.t581 1477.9
R2816 Vbias.t581 Vbias.n7416 1477.9
R2817 Vbias.n7415 Vbias.t251 1477.9
R2818 Vbias.n7389 Vbias.t251 1477.9
R2819 Vbias.t705 Vbias.n7389 1477.9
R2820 Vbias.t705 Vbias.n7390 1477.9
R2821 Vbias.t299 Vbias.n7390 1477.9
R2822 Vbias.n6504 Vbias.t120 1477.9
R2823 Vbias.n6468 Vbias.t120 1477.9
R2824 Vbias.t578 Vbias.n6468 1477.9
R2825 Vbias.t578 Vbias.n6497 1477.9
R2826 Vbias.n6497 Vbias.t326 1477.9
R2827 Vbias.t326 Vbias.n6491 1477.9
R2828 Vbias.n6490 Vbias.t249 1477.9
R2829 Vbias.n6474 Vbias.t249 1477.9
R2830 Vbias.t476 Vbias.n6474 1477.9
R2831 Vbias.t476 Vbias.n6483 1477.9
R2832 Vbias.n6483 Vbias.t570 1477.9
R2833 Vbias.t570 Vbias.n6477 1477.9
R2834 Vbias.n6476 Vbias.t337 1477.9
R2835 Vbias.n7567 Vbias.t337 1477.9
R2836 Vbias.n7566 Vbias.t807 1477.9
R2837 Vbias.n892 Vbias.t807 1477.9
R2838 Vbias.t391 Vbias.n892 1477.9
R2839 Vbias.n7557 Vbias.t391 1477.9
R2840 Vbias.n7556 Vbias.t204 1477.9
R2841 Vbias.n906 Vbias.t204 1477.9
R2842 Vbias.n906 Vbias.t506 1477.9
R2843 Vbias.n916 Vbias.t506 1477.9
R2844 Vbias.t582 Vbias.n916 1477.9
R2845 Vbias.n7545 Vbias.t582 1477.9
R2846 Vbias.t88 Vbias.n6226 1477.9
R2847 Vbias.n6395 Vbias.t88 1477.9
R2848 Vbias.t654 Vbias.n6395 1477.9
R2849 Vbias.t654 Vbias.n6398 1477.9
R2850 Vbias.n6398 Vbias.t442 1477.9
R2851 Vbias.n6405 Vbias.t442 1477.9
R2852 Vbias.t277 Vbias.n6406 1477.9
R2853 Vbias.n6412 Vbias.t277 1477.9
R2854 Vbias.t800 Vbias.n6412 1477.9
R2855 Vbias.t800 Vbias.n6415 1477.9
R2856 Vbias.n6415 Vbias.t555 1477.9
R2857 Vbias.n6422 Vbias.t555 1477.9
R2858 Vbias.t483 Vbias.n6424 1477.9
R2859 Vbias.n6554 Vbias.t483 1477.9
R2860 Vbias.n6553 Vbias.t344 1477.9
R2861 Vbias.n6438 Vbias.t344 1477.9
R2862 Vbias.t745 Vbias.n6438 1477.9
R2863 Vbias.n6544 Vbias.t745 1477.9
R2864 Vbias.n6543 Vbias.t231 1477.9
R2865 Vbias.n6452 Vbias.t231 1477.9
R2866 Vbias.n6452 Vbias.t753 1477.9
R2867 Vbias.n6462 Vbias.t753 1477.9
R2868 Vbias.t373 Vbias.n6462 1477.9
R2869 Vbias.n6532 Vbias.t373 1477.9
R2870 Vbias.t74 Vbias.n755 1477.9
R2871 Vbias.n6643 Vbias.t74 1477.9
R2872 Vbias.n6643 Vbias.t625 1477.9
R2873 Vbias.t625 Vbias.n6144 1477.9
R2874 Vbias.t865 Vbias.n6144 1477.9
R2875 Vbias.t865 Vbias.n6150 1477.9
R2876 Vbias.t224 Vbias.n6169 1477.9
R2877 Vbias.n6175 Vbias.t224 1477.9
R2878 Vbias.t860 Vbias.n6175 1477.9
R2879 Vbias.t860 Vbias.n6178 1477.9
R2880 Vbias.n6178 Vbias.t132 1477.9
R2881 Vbias.n6185 Vbias.t132 1477.9
R2882 Vbias.t383 Vbias.n6187 1477.9
R2883 Vbias.n6621 Vbias.t383 1477.9
R2884 Vbias.n6620 Vbias.t733 1477.9
R2885 Vbias.n6201 Vbias.t733 1477.9
R2886 Vbias.t749 Vbias.n6201 1477.9
R2887 Vbias.n6611 Vbias.t749 1477.9
R2888 Vbias.n6610 Vbias.t186 1477.9
R2889 Vbias.n6215 Vbias.t186 1477.9
R2890 Vbias.n6215 Vbias.t515 1477.9
R2891 Vbias.n6225 Vbias.t515 1477.9
R2892 Vbias.t770 Vbias.n6225 1477.9
R2893 Vbias.n6599 Vbias.t770 1477.9
R2894 Vbias.n7735 Vbias.t24 1477.9
R2895 Vbias.n688 Vbias.t24 1477.9
R2896 Vbias.t623 Vbias.n688 1477.9
R2897 Vbias.t623 Vbias.n689 1477.9
R2898 Vbias.t487 Vbias.n689 1477.9
R2899 Vbias.t487 Vbias.n698 1477.9
R2900 Vbias.t245 Vbias.n706 1477.9
R2901 Vbias.n7714 Vbias.t245 1477.9
R2902 Vbias.n7714 Vbias.t778 1477.9
R2903 Vbias.t778 Vbias.n710 1477.9
R2904 Vbias.t292 Vbias.n710 1477.9
R2905 Vbias.t292 Vbias.n716 1477.9
R2906 Vbias.t332 Vbias.n725 1477.9
R2907 Vbias.n7700 Vbias.t332 1477.9
R2908 Vbias.n7699 Vbias.t671 1477.9
R2909 Vbias.n734 Vbias.t671 1477.9
R2910 Vbias.t540 Vbias.n734 1477.9
R2911 Vbias.t540 Vbias.n7685 1477.9
R2912 Vbias.n7684 Vbias.t200 1477.9
R2913 Vbias.n744 Vbias.t200 1477.9
R2914 Vbias.t706 Vbias.n744 1477.9
R2915 Vbias.t706 Vbias.n745 1477.9
R2916 Vbias.t552 Vbias.n745 1477.9
R2917 Vbias.t552 Vbias.n7669 1477.9
R2918 Vbias.n5639 Vbias.n5638 1297.44
R2919 Vbias.n5713 Vbias.n5712 1297.44
R2920 Vbias.n5802 Vbias.n1674 1297.44
R2921 Vbias.n7971 Vbias.n7970 1297.44
R2922 Vbias.n6590 Vbias.n6589 1246.88
R2923 Vbias.n7652 Vbias.n7651 1246.88
R2924 Vbias.n1018 Vbias.n1017 1246.88
R2925 Vbias.n1028 Vbias.n1026 1246.88
R2926 Vbias.n7226 Vbias.n7225 1235.69
R2927 Vbias.n7123 Vbias.n7122 1036.63
R2928 Vbias.n6075 Vbias.n6074 1036.63
R2929 Vbias.n5485 Vbias.n5484 1036.63
R2930 Vbias.n5038 Vbias.n5037 1036.63
R2931 Vbias.n8009 Vbias.n8008 1017.54
R2932 Vbias.n4378 Vbias.n2792 1014.28
R2933 Vbias.n4378 Vbias.n4377 1014.28
R2934 Vbias.n4393 Vbias.n2793 1014.28
R2935 Vbias.n4393 Vbias.n4392 1014.28
R2936 Vbias.n4353 Vbias.n2815 1014.28
R2937 Vbias.n4353 Vbias.n2816 1014.28
R2938 Vbias.n2856 Vbias.n2839 1014.28
R2939 Vbias.n2856 Vbias.n2843 1014.28
R2940 Vbias.n2836 Vbias.n2835 1014.28
R2941 Vbias.n2836 Vbias.n2828 1014.28
R2942 Vbias.n2890 Vbias.n2873 1014.28
R2943 Vbias.n2890 Vbias.n2877 1014.28
R2944 Vbias.n2870 Vbias.n2869 1014.28
R2945 Vbias.n2870 Vbias.n2864 1014.28
R2946 Vbias.n4374 Vbias.n4373 1014.28
R2947 Vbias.n4374 Vbias.n2784 1014.28
R2948 Vbias.n2788 Vbias.n2783 1014.28
R2949 Vbias.n4399 Vbias.n2783 1014.28
R2950 Vbias.n4351 Vbias.n2817 1014.28
R2951 Vbias.n4351 Vbias.n2818 1014.28
R2952 Vbias.n2851 Vbias.n2850 1014.28
R2953 Vbias.n2850 Vbias.n2848 1014.28
R2954 Vbias.n4317 Vbias.n4315 1014.28
R2955 Vbias.n4317 Vbias.n4316 1014.28
R2956 Vbias.n2885 Vbias.n2884 1014.28
R2957 Vbias.n2884 Vbias.n2882 1014.28
R2958 Vbias.n4284 Vbias.n4282 1014.28
R2959 Vbias.n4284 Vbias.n4283 1014.28
R2960 Vbias.n5866 Vbias.n1685 1014.28
R2961 Vbias.n5866 Vbias.n1686 1014.28
R2962 Vbias.n5520 Vbias.n5519 1014.28
R2963 Vbias.n5520 Vbias.n5516 1014.28
R2964 Vbias.n5542 Vbias.n2238 1014.28
R2965 Vbias.n5542 Vbias.n2239 1014.28
R2966 Vbias.n5023 Vbias.n2590 1014.28
R2967 Vbias.n5023 Vbias.n2591 1014.28
R2968 Vbias.n4996 Vbias.n4995 1014.28
R2969 Vbias.n4996 Vbias.n2599 1014.28
R2970 Vbias.n153 Vbias.n149 1014.28
R2971 Vbias.n154 Vbias.n153 1014.28
R2972 Vbias.n161 Vbias.n150 1014.28
R2973 Vbias.n161 Vbias.n155 1014.28
R2974 Vbias.n140 Vbias.n139 1014.28
R2975 Vbias.n139 Vbias.n135 1014.28
R2976 Vbias.n119 Vbias.n118 1014.28
R2977 Vbias.n118 Vbias.n114 1014.28
R2978 Vbias.n125 Vbias.n120 1014.28
R2979 Vbias.n125 Vbias.n115 1014.28
R2980 Vbias.n100 Vbias.n99 1014.28
R2981 Vbias.n99 Vbias.n95 1014.28
R2982 Vbias.n104 Vbias.n101 1014.28
R2983 Vbias.n104 Vbias.n96 1014.28
R2984 Vbias.n79 Vbias.n77 1014.28
R2985 Vbias.n79 Vbias.n73 1014.28
R2986 Vbias.n82 Vbias.n78 1014.28
R2987 Vbias.n82 Vbias.n74 1014.28
R2988 Vbias.n8027 Vbias.n8026 1014.28
R2989 Vbias.n8027 Vbias.n63 1014.28
R2990 Vbias.n8055 Vbias.n35 1014.28
R2991 Vbias.n8055 Vbias.n36 1014.28
R2992 Vbias.n48 Vbias.n43 1014.28
R2993 Vbias.n49 Vbias.n48 1014.28
R2994 Vbias.n22 Vbias.n21 1014.28
R2995 Vbias.n21 Vbias.n17 1014.28
R2996 Vbias.n25 Vbias.n23 1014.28
R2997 Vbias.n25 Vbias.n18 1014.28
R2998 Vbias.n6708 Vbias.n6706 1014.28
R2999 Vbias.n6708 Vbias.n6707 1014.28
R3000 Vbias.n6734 Vbias.n6732 1014.28
R3001 Vbias.n6734 Vbias.n6733 1014.28
R3002 Vbias.n1740 Vbias.n1727 1014.28
R3003 Vbias.n1741 Vbias.n1740 1014.28
R3004 Vbias.n2040 Vbias.n1728 1014.28
R3005 Vbias.n2040 Vbias.n1732 1014.28
R3006 Vbias.n2066 Vbias.n1696 1014.28
R3007 Vbias.n2067 Vbias.n2066 1014.28
R3008 Vbias.n2061 Vbias.n1697 1014.28
R3009 Vbias.n2062 Vbias.n2061 1014.28
R3010 Vbias.n7739 Vbias.n7738 1014.28
R3011 Vbias.n7739 Vbias.n675 1014.28
R3012 Vbias.n2082 Vbias.n2081 1014.28
R3013 Vbias.n2082 Vbias.n2079 1014.28
R3014 Vbias.n2076 Vbias.n2072 1014.28
R3015 Vbias.n2076 Vbias.n2075 1014.28
R3016 Vbias.n5798 Vbias.n5789 1014.28
R3017 Vbias.n5798 Vbias.n5797 1014.28
R3018 Vbias.n2098 Vbias.n2097 1014.28
R3019 Vbias.n2098 Vbias.n2093 1014.28
R3020 Vbias.n2095 Vbias.n2089 1014.28
R3021 Vbias.n2095 Vbias.n2090 1014.28
R3022 Vbias.n2120 Vbias.n2119 1014.28
R3023 Vbias.n2120 Vbias.n2117 1014.28
R3024 Vbias.n2114 Vbias.n2105 1014.28
R3025 Vbias.n2114 Vbias.n2113 1014.28
R3026 Vbias.n7810 Vbias.n563 1014.28
R3027 Vbias.n7810 Vbias.n564 1014.28
R3028 Vbias.n2137 Vbias.n2136 1014.28
R3029 Vbias.n2137 Vbias.n2134 1014.28
R3030 Vbias.n2131 Vbias.n2127 1014.28
R3031 Vbias.n2131 Vbias.n2130 1014.28
R3032 Vbias.n2153 Vbias.n2144 1014.28
R3033 Vbias.n2153 Vbias.n2152 1014.28
R3034 Vbias.n2169 Vbias.n2166 1014.28
R3035 Vbias.n2169 Vbias.n2162 1014.28
R3036 Vbias.n2168 Vbias.n2167 1014.28
R3037 Vbias.n2167 Vbias.n2163 1014.28
R3038 Vbias.n2187 Vbias.n2184 1014.28
R3039 Vbias.n2187 Vbias.n2180 1014.28
R3040 Vbias.n2186 Vbias.n2185 1014.28
R3041 Vbias.n2185 Vbias.n2181 1014.28
R3042 Vbias.n7874 Vbias.n7873 1014.28
R3043 Vbias.n7874 Vbias.n454 1014.28
R3044 Vbias.n2208 Vbias.n2207 1014.28
R3045 Vbias.n2208 Vbias.n2205 1014.28
R3046 Vbias.n2202 Vbias.n2198 1014.28
R3047 Vbias.n2202 Vbias.n2201 1014.28
R3048 Vbias.n2224 Vbias.n2215 1014.28
R3049 Vbias.n2224 Vbias.n2223 1014.28
R3050 Vbias.n5566 Vbias.n5563 1014.28
R3051 Vbias.n5566 Vbias.n5559 1014.28
R3052 Vbias.n5565 Vbias.n5564 1014.28
R3053 Vbias.n5564 Vbias.n5560 1014.28
R3054 Vbias.n5584 Vbias.n5581 1014.28
R3055 Vbias.n5584 Vbias.n5577 1014.28
R3056 Vbias.n5583 Vbias.n5582 1014.28
R3057 Vbias.n5582 Vbias.n5578 1014.28
R3058 Vbias.n333 Vbias.n330 1014.28
R3059 Vbias.n333 Vbias.n331 1014.28
R3060 Vbias.n7543 Vbias.n918 1014.28
R3061 Vbias.n7543 Vbias.n919 1014.28
R3062 Vbias.n6526 Vbias.n6522 1014.28
R3063 Vbias.n6526 Vbias.n6525 1014.28
R3064 Vbias.n6597 Vbias.n6595 1014.28
R3065 Vbias.n6597 Vbias.n6596 1014.28
R3066 Vbias.n766 Vbias.n760 1014.28
R3067 Vbias.n767 Vbias.n766 1014.28
R3068 Vbias.n7250 Vbias.n7246 1014.28
R3069 Vbias.n7251 Vbias.n7250 1014.28
R3070 Vbias.n7258 Vbias.n7247 1014.28
R3071 Vbias.n7258 Vbias.n7252 1014.28
R3072 Vbias.n7237 Vbias.n7236 1014.28
R3073 Vbias.n7236 Vbias.n7232 1014.28
R3074 Vbias.n1060 Vbias.n1059 1014.28
R3075 Vbias.n1059 Vbias.n1055 1014.28
R3076 Vbias.n1066 Vbias.n1061 1014.28
R3077 Vbias.n1066 Vbias.n1056 1014.28
R3078 Vbias.n1039 Vbias.n1038 1014.28
R3079 Vbias.n1038 Vbias.n1034 1014.28
R3080 Vbias.n1045 Vbias.n1040 1014.28
R3081 Vbias.n1045 Vbias.n1035 1014.28
R3082 Vbias.n1000 Vbias.n996 1014.28
R3083 Vbias.n1001 Vbias.n1000 1014.28
R3084 Vbias.n1008 Vbias.n997 1014.28
R3085 Vbias.n1008 Vbias.n1002 1014.28
R3086 Vbias.n987 Vbias.n986 1014.28
R3087 Vbias.n986 Vbias.n982 1014.28
R3088 Vbias.n965 Vbias.n964 1014.28
R3089 Vbias.n964 Vbias.n960 1014.28
R3090 Vbias.n971 Vbias.n966 1014.28
R3091 Vbias.n971 Vbias.n961 1014.28
R3092 Vbias.n942 Vbias.n941 1014.28
R3093 Vbias.n941 Vbias.n937 1014.28
R3094 Vbias.n950 Vbias.n943 1014.28
R3095 Vbias.n950 Vbias.n938 1014.28
R3096 Vbias.n845 Vbias.n841 1014.28
R3097 Vbias.n846 Vbias.n845 1014.28
R3098 Vbias.n853 Vbias.n842 1014.28
R3099 Vbias.n853 Vbias.n847 1014.28
R3100 Vbias.n832 Vbias.n831 1014.28
R3101 Vbias.n831 Vbias.n827 1014.28
R3102 Vbias.n810 Vbias.n809 1014.28
R3103 Vbias.n809 Vbias.n805 1014.28
R3104 Vbias.n816 Vbias.n811 1014.28
R3105 Vbias.n816 Vbias.n806 1014.28
R3106 Vbias.n791 Vbias.n790 1014.28
R3107 Vbias.n790 Vbias.n786 1014.28
R3108 Vbias.n795 Vbias.n792 1014.28
R3109 Vbias.n795 Vbias.n787 1014.28
R3110 Vbias.n6239 Vbias.n6236 1014.28
R3111 Vbias.n6239 Vbias.n6232 1014.28
R3112 Vbias.n6238 Vbias.n6237 1014.28
R3113 Vbias.n6237 Vbias.n6233 1014.28
R3114 Vbias.n6255 Vbias.n6254 1014.28
R3115 Vbias.n6254 Vbias.n6251 1014.28
R3116 Vbias.n6271 Vbias.n6270 1014.28
R3117 Vbias.n6271 Vbias.n6268 1014.28
R3118 Vbias.n6265 Vbias.n6260 1014.28
R3119 Vbias.n6265 Vbias.n6264 1014.28
R3120 Vbias.n6293 Vbias.n6292 1014.28
R3121 Vbias.n6293 Vbias.n6290 1014.28
R3122 Vbias.n6287 Vbias.n6278 1014.28
R3123 Vbias.n6287 Vbias.n6286 1014.28
R3124 Vbias.n1490 Vbias.n1486 1014.28
R3125 Vbias.n1491 Vbias.n1490 1014.28
R3126 Vbias.n1497 Vbias.n1487 1014.28
R3127 Vbias.n1497 Vbias.n1492 1014.28
R3128 Vbias.n1478 Vbias.n1477 1014.28
R3129 Vbias.n1477 Vbias.n1473 1014.28
R3130 Vbias.n748 Vbias.n746 1014.28
R3131 Vbias.n748 Vbias.n742 1014.28
R3132 Vbias.n751 Vbias.n747 1014.28
R3133 Vbias.n751 Vbias.n743 1014.28
R3134 Vbias.n7687 Vbias.n7686 1014.28
R3135 Vbias.n7687 Vbias.n732 1014.28
R3136 Vbias.n7715 Vbias.n704 1014.28
R3137 Vbias.n7715 Vbias.n705 1014.28
R3138 Vbias.n717 Vbias.n712 1014.28
R3139 Vbias.n718 Vbias.n717 1014.28
R3140 Vbias.n691 Vbias.n690 1014.28
R3141 Vbias.n690 Vbias.n686 1014.28
R3142 Vbias.n694 Vbias.n692 1014.28
R3143 Vbias.n694 Vbias.n687 1014.28
R3144 Vbias.n657 Vbias.n654 1014.28
R3145 Vbias.n657 Vbias.n655 1014.28
R3146 Vbias.n665 Vbias.n663 1014.28
R3147 Vbias.n665 Vbias.n664 1014.28
R3148 Vbias.n641 Vbias.n639 1014.28
R3149 Vbias.n641 Vbias.n640 1014.28
R3150 Vbias.n610 Vbias.n607 1014.28
R3151 Vbias.n610 Vbias.n608 1014.28
R3152 Vbias.n618 Vbias.n616 1014.28
R3153 Vbias.n618 Vbias.n617 1014.28
R3154 Vbias.n586 Vbias.n583 1014.28
R3155 Vbias.n586 Vbias.n584 1014.28
R3156 Vbias.n594 Vbias.n592 1014.28
R3157 Vbias.n594 Vbias.n593 1014.28
R3158 Vbias.n543 Vbias.n540 1014.28
R3159 Vbias.n543 Vbias.n541 1014.28
R3160 Vbias.n551 Vbias.n549 1014.28
R3161 Vbias.n551 Vbias.n550 1014.28
R3162 Vbias.n527 Vbias.n525 1014.28
R3163 Vbias.n527 Vbias.n526 1014.28
R3164 Vbias.n496 Vbias.n493 1014.28
R3165 Vbias.n496 Vbias.n494 1014.28
R3166 Vbias.n504 Vbias.n502 1014.28
R3167 Vbias.n504 Vbias.n503 1014.28
R3168 Vbias.n472 Vbias.n469 1014.28
R3169 Vbias.n472 Vbias.n470 1014.28
R3170 Vbias.n480 Vbias.n478 1014.28
R3171 Vbias.n480 Vbias.n479 1014.28
R3172 Vbias.n437 Vbias.n434 1014.28
R3173 Vbias.n437 Vbias.n435 1014.28
R3174 Vbias.n445 Vbias.n443 1014.28
R3175 Vbias.n445 Vbias.n444 1014.28
R3176 Vbias.n421 Vbias.n419 1014.28
R3177 Vbias.n421 Vbias.n420 1014.28
R3178 Vbias.n390 Vbias.n387 1014.28
R3179 Vbias.n390 Vbias.n388 1014.28
R3180 Vbias.n398 Vbias.n396 1014.28
R3181 Vbias.n398 Vbias.n397 1014.28
R3182 Vbias.n366 Vbias.n363 1014.28
R3183 Vbias.n366 Vbias.n364 1014.28
R3184 Vbias.n374 Vbias.n372 1014.28
R3185 Vbias.n374 Vbias.n373 1014.28
R3186 Vbias.n317 Vbias.n187 1014.28
R3187 Vbias.n192 Vbias.n187 1014.28
R3188 Vbias.n322 Vbias.n184 1014.28
R3189 Vbias.n322 Vbias.n185 1014.28
R3190 Vbias.n305 Vbias.n203 1014.28
R3191 Vbias.n305 Vbias.n204 1014.28
R3192 Vbias.n278 Vbias.n220 1014.28
R3193 Vbias.n225 Vbias.n220 1014.28
R3194 Vbias.n283 Vbias.n217 1014.28
R3195 Vbias.n283 Vbias.n218 1014.28
R3196 Vbias.n261 Vbias.n239 1014.28
R3197 Vbias.n243 Vbias.n239 1014.28
R3198 Vbias.n266 Vbias.n236 1014.28
R3199 Vbias.n266 Vbias.n237 1014.28
R3200 Vbias.n4609 Vbias.n4608 1014.28
R3201 Vbias.n4608 Vbias.n4604 1014.28
R3202 Vbias.n4637 Vbias.n4610 1014.28
R3203 Vbias.n4637 Vbias.n4605 1014.28
R3204 Vbias.n4622 Vbias.n4615 1014.28
R3205 Vbias.n4615 Vbias.n4614 1014.28
R3206 Vbias.n4624 Vbias.n4612 1014.28
R3207 Vbias.n4624 Vbias.n4623 1014.28
R3208 Vbias.n4587 Vbias.n4583 1014.28
R3209 Vbias.n4587 Vbias.n4584 1014.28
R3210 Vbias.n4470 Vbias.n4466 1014.28
R3211 Vbias.n4471 Vbias.n4470 1014.28
R3212 Vbias.n4478 Vbias.n4467 1014.28
R3213 Vbias.n4478 Vbias.n4472 1014.28
R3214 Vbias.n4448 Vbias.n4444 1014.28
R3215 Vbias.n4449 Vbias.n4448 1014.28
R3216 Vbias.n4456 Vbias.n4445 1014.28
R3217 Vbias.n4456 Vbias.n4450 1014.28
R3218 Vbias.n4436 Vbias.n4435 1014.28
R3219 Vbias.n4435 Vbias.n4431 1014.28
R3220 Vbias.n4417 Vbias.n4416 1014.28
R3221 Vbias.n4416 Vbias.n4412 1014.28
R3222 Vbias.n4420 Vbias.n4418 1014.28
R3223 Vbias.n4420 Vbias.n4413 1014.28
R3224 Vbias.n2384 Vbias.n2382 1014.28
R3225 Vbias.n2384 Vbias.n2378 1014.28
R3226 Vbias.n5107 Vbias.n2383 1014.28
R3227 Vbias.n5107 Vbias.n2379 1014.28
R3228 Vbias.n2400 Vbias.n2398 1014.28
R3229 Vbias.n2400 Vbias.n2394 1014.28
R3230 Vbias.n5087 Vbias.n2399 1014.28
R3231 Vbias.n5087 Vbias.n2395 1014.28
R3232 Vbias.n5064 Vbias.n2412 1014.28
R3233 Vbias.n5064 Vbias.n2413 1014.28
R3234 Vbias.n2278 Vbias.n2275 1014.28
R3235 Vbias.n2278 Vbias.n2276 1014.28
R3236 Vbias.n2286 Vbias.n2284 1014.28
R3237 Vbias.n2286 Vbias.n2285 1014.28
R3238 Vbias.n5507 Vbias.n2246 1014.28
R3239 Vbias.n5507 Vbias.n2247 1014.28
R3240 Vbias.n2263 Vbias.n2257 1014.28
R3241 Vbias.n2263 Vbias.n2258 1014.28
R3242 Vbias.n5147 Vbias.n5145 1014.28
R3243 Vbias.n5147 Vbias.n5146 1014.28
R3244 Vbias.n5128 Vbias.n2366 1014.28
R3245 Vbias.n5128 Vbias.n5127 1014.28
R3246 Vbias.n5131 Vbias.n2364 1014.28
R3247 Vbias.n5131 Vbias.n5130 1014.28
R3248 Vbias.n1652 Vbias.n1650 1014.28
R3249 Vbias.n1652 Vbias.n1646 1014.28
R3250 Vbias.n5904 Vbias.n1651 1014.28
R3251 Vbias.n5904 Vbias.n1647 1014.28
R3252 Vbias.n1668 Vbias.n1666 1014.28
R3253 Vbias.n1668 Vbias.n1662 1014.28
R3254 Vbias.n5884 Vbias.n1667 1014.28
R3255 Vbias.n5884 Vbias.n1663 1014.28
R3256 Vbias.n5449 Vbias.n5445 1014.28
R3257 Vbias.n5449 Vbias.n5446 1014.28
R3258 Vbias.n5426 Vbias.n5423 1014.28
R3259 Vbias.n5426 Vbias.n5424 1014.28
R3260 Vbias.n5434 Vbias.n5432 1014.28
R3261 Vbias.n5434 Vbias.n5433 1014.28
R3262 Vbias.n5939 Vbias.n1627 1014.28
R3263 Vbias.n5939 Vbias.n5938 1014.28
R3264 Vbias.n1633 Vbias.n1632 1014.28
R3265 Vbias.n1632 Vbias.n1631 1014.28
R3266 Vbias.n5928 Vbias.n1628 1014.28
R3267 Vbias.n5928 Vbias.n5927 1014.28
R3268 Vbias.n1811 Vbias.n1802 1014.28
R3269 Vbias.n1802 Vbias.n1764 1014.28
R3270 Vbias.n1766 Vbias.n1757 1014.28
R3271 Vbias.n1766 Vbias.n1761 1014.28
R3272 Vbias.n1857 Vbias.n1851 1014.28
R3273 Vbias.n1857 Vbias.n1855 1014.28
R3274 Vbias.n1865 Vbias.n1852 1014.28
R3275 Vbias.n1865 Vbias.n1856 1014.28
R3276 Vbias.n1925 Vbias.n1919 1014.28
R3277 Vbias.n1925 Vbias.n1923 1014.28
R3278 Vbias.n1941 Vbias.n1920 1014.28
R3279 Vbias.n1941 Vbias.n1924 1014.28
R3280 Vbias.n1995 Vbias.n1991 1014.28
R3281 Vbias.n2004 Vbias.n1991 1014.28
R3282 Vbias.n2009 Vbias.n1989 1014.28
R3283 Vbias.n2009 Vbias.n1988 1014.28
R3284 Vbias.n1519 Vbias.n1513 1014.28
R3285 Vbias.n1519 Vbias.n1517 1014.28
R3286 Vbias.n6115 Vbias.n1514 1014.28
R3287 Vbias.n6115 Vbias.n1518 1014.28
R3288 Vbias.n1959 Vbias.n1953 1014.28
R3289 Vbias.n1959 Vbias.n1957 1014.28
R3290 Vbias.n1975 Vbias.n1954 1014.28
R3291 Vbias.n1975 Vbias.n1958 1014.28
R3292 Vbias.n1889 Vbias.n1886 1014.28
R3293 Vbias.n1889 Vbias.n1888 1014.28
R3294 Vbias.n1905 Vbias.n1894 1014.28
R3295 Vbias.n1894 Vbias.n1892 1014.28
R3296 Vbias.n1778 Vbias.n1777 1014.28
R3297 Vbias.n1777 Vbias.n1775 1014.28
R3298 Vbias.n1782 Vbias.n1781 1014.28
R3299 Vbias.n1781 Vbias.n1780 1014.28
R3300 Vbias.n1771 Vbias.n1770 1014.28
R3301 Vbias.n1770 Vbias.n1769 1014.28
R3302 Vbias.n1794 Vbias.n1774 1014.28
R3303 Vbias.n1774 Vbias.n1773 1014.28
R3304 Vbias.n1437 Vbias.n1436 1014.28
R3305 Vbias.n1436 Vbias.n1432 1014.28
R3306 Vbias.n6775 Vbias.n1438 1014.28
R3307 Vbias.n6775 Vbias.n1433 1014.28
R3308 Vbias.n6759 Vbias.n1442 1014.28
R3309 Vbias.n6759 Vbias.n6758 1014.28
R3310 Vbias.n6762 Vbias.n1440 1014.28
R3311 Vbias.n6762 Vbias.n6761 1014.28
R3312 Vbias.n6055 Vbias.n6054 1014.28
R3313 Vbias.n6054 Vbias.n6052 1014.28
R3314 Vbias.n6050 Vbias.n6046 1014.28
R3315 Vbias.n6050 Vbias.n6049 1014.28
R3316 Vbias.n6066 Vbias.n6048 1014.28
R3317 Vbias.n6066 Vbias.n6065 1014.28
R3318 Vbias.n7083 Vbias.n1281 1014.28
R3319 Vbias.n1286 Vbias.n1281 1014.28
R3320 Vbias.n7088 Vbias.n1278 1014.28
R3321 Vbias.n7088 Vbias.n1279 1014.28
R3322 Vbias.n7066 Vbias.n1300 1014.28
R3323 Vbias.n1306 Vbias.n1300 1014.28
R3324 Vbias.n7071 Vbias.n1297 1014.28
R3325 Vbias.n7071 Vbias.n1298 1014.28
R3326 Vbias.n7040 Vbias.n7039 1014.28
R3327 Vbias.n7040 Vbias.n1322 1014.28
R3328 Vbias.n1335 Vbias.n1333 1014.28
R3329 Vbias.n1335 Vbias.n1329 1014.28
R3330 Vbias.n7023 Vbias.n1334 1014.28
R3331 Vbias.n7023 Vbias.n1330 1014.28
R3332 Vbias.n7189 Vbias.n1094 1014.28
R3333 Vbias.n1099 Vbias.n1094 1014.28
R3334 Vbias.n7194 Vbias.n1091 1014.28
R3335 Vbias.n7194 Vbias.n1092 1014.28
R3336 Vbias.n7172 Vbias.n1113 1014.28
R3337 Vbias.n1118 Vbias.n1113 1014.28
R3338 Vbias.n7177 Vbias.n1110 1014.28
R3339 Vbias.n7177 Vbias.n1111 1014.28
R3340 Vbias.n7146 Vbias.n7145 1014.28
R3341 Vbias.n7146 Vbias.n1134 1014.28
R3342 Vbias.n1147 Vbias.n1145 1014.28
R3343 Vbias.n1147 Vbias.n1141 1014.28
R3344 Vbias.n7129 Vbias.n1146 1014.28
R3345 Vbias.n7129 Vbias.n1142 1014.28
R3346 Vbias.n1218 Vbias.n1084 1014.28
R3347 Vbias.n1218 Vbias.n1217 1014.28
R3348 Vbias.n7211 Vbias.n1080 1014.28
R3349 Vbias.n7211 Vbias.n1081 1014.28
R3350 Vbias.n1238 Vbias.n1201 1014.28
R3351 Vbias.n1238 Vbias.n1202 1014.28
R3352 Vbias.n1235 Vbias.n1209 1014.28
R3353 Vbias.n1226 Vbias.n1209 1014.28
R3354 Vbias.n1249 Vbias.n1188 1014.28
R3355 Vbias.n1249 Vbias.n1189 1014.28
R3356 Vbias.n1269 Vbias.n1173 1014.28
R3357 Vbias.n1269 Vbias.n1174 1014.28
R3358 Vbias.n1266 Vbias.n1180 1014.28
R3359 Vbias.n1257 Vbias.n1180 1014.28
R3360 Vbias.n6951 Vbias.n1165 1014.28
R3361 Vbias.n6951 Vbias.n6950 1014.28
R3362 Vbias.n7107 Vbias.n1161 1014.28
R3363 Vbias.n7107 Vbias.n1162 1014.28
R3364 Vbias.n6971 Vbias.n6934 1014.28
R3365 Vbias.n6971 Vbias.n6935 1014.28
R3366 Vbias.n6968 Vbias.n6942 1014.28
R3367 Vbias.n6959 Vbias.n6942 1014.28
R3368 Vbias.n6982 Vbias.n6921 1014.28
R3369 Vbias.n6982 Vbias.n6922 1014.28
R3370 Vbias.n7002 Vbias.n6906 1014.28
R3371 Vbias.n7002 Vbias.n6907 1014.28
R3372 Vbias.n6999 Vbias.n6913 1014.28
R3373 Vbias.n6990 Vbias.n6913 1014.28
R3374 Vbias.n6872 Vbias.n1359 1014.28
R3375 Vbias.n6872 Vbias.n6871 1014.28
R3376 Vbias.n6886 Vbias.n1355 1014.28
R3377 Vbias.n6886 Vbias.n1356 1014.28
R3378 Vbias.n6849 Vbias.n1372 1014.28
R3379 Vbias.n6849 Vbias.n6848 1014.28
R3380 Vbias.n6863 Vbias.n1368 1014.28
R3381 Vbias.n6863 Vbias.n1369 1014.28
R3382 Vbias.n6840 Vbias.n1381 1014.28
R3383 Vbias.n6840 Vbias.n1382 1014.28
R3384 Vbias.n6818 Vbias.n1398 1014.28
R3385 Vbias.n6818 Vbias.n1396 1014.28
R3386 Vbias.n6825 Vbias.n1390 1014.28
R3387 Vbias.n6825 Vbias.n1394 1014.28
R3388 Vbias.n6014 Vbias.n1570 1014.28
R3389 Vbias.n6014 Vbias.n6013 1014.28
R3390 Vbias.n6031 Vbias.n1566 1014.28
R3391 Vbias.n6031 Vbias.n1567 1014.28
R3392 Vbias.n5991 Vbias.n1583 1014.28
R3393 Vbias.n5991 Vbias.n5990 1014.28
R3394 Vbias.n6005 Vbias.n1579 1014.28
R3395 Vbias.n6005 Vbias.n1580 1014.28
R3396 Vbias.n5982 Vbias.n1592 1014.28
R3397 Vbias.n5982 Vbias.n1593 1014.28
R3398 Vbias.n5960 Vbias.n1609 1014.28
R3399 Vbias.n5960 Vbias.n1607 1014.28
R3400 Vbias.n5967 Vbias.n1601 1014.28
R3401 Vbias.n5967 Vbias.n1605 1014.28
R3402 Vbias.n5326 Vbias.n5325 1014.28
R3403 Vbias.n5325 Vbias.n5321 1014.28
R3404 Vbias.n5329 Vbias.n5327 1014.28
R3405 Vbias.n5329 Vbias.n5322 1014.28
R3406 Vbias.n5379 Vbias.n5305 1014.28
R3407 Vbias.n5379 Vbias.n5306 1014.28
R3408 Vbias.n5376 Vbias.n5313 1014.28
R3409 Vbias.n5367 Vbias.n5313 1014.28
R3410 Vbias.n5390 Vbias.n5292 1014.28
R3411 Vbias.n5390 Vbias.n5293 1014.28
R3412 Vbias.n5410 Vbias.n5276 1014.28
R3413 Vbias.n5410 Vbias.n5277 1014.28
R3414 Vbias.n5407 Vbias.n5284 1014.28
R3415 Vbias.n5398 Vbias.n5284 1014.28
R3416 Vbias.n5241 Vbias.n2307 1014.28
R3417 Vbias.n5241 Vbias.n5240 1014.28
R3418 Vbias.n5255 Vbias.n2303 1014.28
R3419 Vbias.n5255 Vbias.n2304 1014.28
R3420 Vbias.n5218 Vbias.n2320 1014.28
R3421 Vbias.n5218 Vbias.n5217 1014.28
R3422 Vbias.n5232 Vbias.n2316 1014.28
R3423 Vbias.n5232 Vbias.n2317 1014.28
R3424 Vbias.n5209 Vbias.n2329 1014.28
R3425 Vbias.n5209 Vbias.n2330 1014.28
R3426 Vbias.n5187 Vbias.n2346 1014.28
R3427 Vbias.n5187 Vbias.n2344 1014.28
R3428 Vbias.n5194 Vbias.n2338 1014.28
R3429 Vbias.n5194 Vbias.n2342 1014.28
R3430 Vbias.n2494 Vbias.n2493 1014.28
R3431 Vbias.n2493 Vbias.n2489 1014.28
R3432 Vbias.n2497 Vbias.n2495 1014.28
R3433 Vbias.n2497 Vbias.n2490 1014.28
R3434 Vbias.n2547 Vbias.n2473 1014.28
R3435 Vbias.n2547 Vbias.n2474 1014.28
R3436 Vbias.n2544 Vbias.n2481 1014.28
R3437 Vbias.n2535 Vbias.n2481 1014.28
R3438 Vbias.n2558 Vbias.n2460 1014.28
R3439 Vbias.n2558 Vbias.n2461 1014.28
R3440 Vbias.n2578 Vbias.n2444 1014.28
R3441 Vbias.n2578 Vbias.n2445 1014.28
R3442 Vbias.n2575 Vbias.n2452 1014.28
R3443 Vbias.n2566 Vbias.n2452 1014.28
R3444 Vbias.n2429 Vbias.n2427 1014.28
R3445 Vbias.n2429 Vbias.n2423 1014.28
R3446 Vbias.n5044 Vbias.n2428 1014.28
R3447 Vbias.n5044 Vbias.n2424 1014.28
R3448 Vbias.n3810 Vbias.n3807 1014.28
R3449 Vbias.n3810 Vbias.n3802 1014.28
R3450 Vbias.n3813 Vbias.n3808 1014.28
R3451 Vbias.n3813 Vbias.n3803 1014.28
R3452 Vbias.n3882 Vbias.n3784 1014.28
R3453 Vbias.n3882 Vbias.n3785 1014.28
R3454 Vbias.n3763 Vbias.n3760 1014.28
R3455 Vbias.n3763 Vbias.n3755 1014.28
R3456 Vbias.n3766 Vbias.n3761 1014.28
R3457 Vbias.n3766 Vbias.n3756 1014.28
R3458 Vbias.n3734 Vbias.n3731 1014.28
R3459 Vbias.n3734 Vbias.n3726 1014.28
R3460 Vbias.n3737 Vbias.n3732 1014.28
R3461 Vbias.n3737 Vbias.n3727 1014.28
R3462 Vbias.n3824 Vbias.n3823 1014.28
R3463 Vbias.n3825 Vbias.n3824 1014.28
R3464 Vbias.n3833 Vbias.n3831 1014.28
R3465 Vbias.n3833 Vbias.n3832 1014.28
R3466 Vbias.n3787 Vbias.n3786 1014.28
R3467 Vbias.n3869 Vbias.n3786 1014.28
R3468 Vbias.n3900 Vbias.n3899 1014.28
R3469 Vbias.n3901 Vbias.n3900 1014.28
R3470 Vbias.n3909 Vbias.n3907 1014.28
R3471 Vbias.n3909 Vbias.n3908 1014.28
R3472 Vbias.n3938 Vbias.n3937 1014.28
R3473 Vbias.n3939 Vbias.n3938 1014.28
R3474 Vbias.n3947 Vbias.n3945 1014.28
R3475 Vbias.n3947 Vbias.n3946 1014.28
R3476 Vbias.n3272 Vbias.n3269 1014.28
R3477 Vbias.n3272 Vbias.n3264 1014.28
R3478 Vbias.n3275 Vbias.n3270 1014.28
R3479 Vbias.n3275 Vbias.n3265 1014.28
R3480 Vbias.n3344 Vbias.n3246 1014.28
R3481 Vbias.n3344 Vbias.n3247 1014.28
R3482 Vbias.n3225 Vbias.n3222 1014.28
R3483 Vbias.n3225 Vbias.n3217 1014.28
R3484 Vbias.n3228 Vbias.n3223 1014.28
R3485 Vbias.n3228 Vbias.n3218 1014.28
R3486 Vbias.n3196 Vbias.n3193 1014.28
R3487 Vbias.n3196 Vbias.n3188 1014.28
R3488 Vbias.n3199 Vbias.n3194 1014.28
R3489 Vbias.n3199 Vbias.n3189 1014.28
R3490 Vbias.n3286 Vbias.n3285 1014.28
R3491 Vbias.n3287 Vbias.n3286 1014.28
R3492 Vbias.n3295 Vbias.n3293 1014.28
R3493 Vbias.n3295 Vbias.n3294 1014.28
R3494 Vbias.n3249 Vbias.n3248 1014.28
R3495 Vbias.n3331 Vbias.n3248 1014.28
R3496 Vbias.n3362 Vbias.n3361 1014.28
R3497 Vbias.n3363 Vbias.n3362 1014.28
R3498 Vbias.n3371 Vbias.n3369 1014.28
R3499 Vbias.n3371 Vbias.n3370 1014.28
R3500 Vbias.n3400 Vbias.n3399 1014.28
R3501 Vbias.n3401 Vbias.n3400 1014.28
R3502 Vbias.n3409 Vbias.n3407 1014.28
R3503 Vbias.n3409 Vbias.n3408 1014.28
R3504 Vbias.n3541 Vbias.n3538 1014.28
R3505 Vbias.n3541 Vbias.n3533 1014.28
R3506 Vbias.n3544 Vbias.n3539 1014.28
R3507 Vbias.n3544 Vbias.n3534 1014.28
R3508 Vbias.n3613 Vbias.n3515 1014.28
R3509 Vbias.n3613 Vbias.n3516 1014.28
R3510 Vbias.n3494 Vbias.n3491 1014.28
R3511 Vbias.n3494 Vbias.n3486 1014.28
R3512 Vbias.n3497 Vbias.n3492 1014.28
R3513 Vbias.n3497 Vbias.n3487 1014.28
R3514 Vbias.n3465 Vbias.n3462 1014.28
R3515 Vbias.n3465 Vbias.n3457 1014.28
R3516 Vbias.n3468 Vbias.n3463 1014.28
R3517 Vbias.n3468 Vbias.n3458 1014.28
R3518 Vbias.n3555 Vbias.n3554 1014.28
R3519 Vbias.n3556 Vbias.n3555 1014.28
R3520 Vbias.n3564 Vbias.n3562 1014.28
R3521 Vbias.n3564 Vbias.n3563 1014.28
R3522 Vbias.n3518 Vbias.n3517 1014.28
R3523 Vbias.n3600 Vbias.n3517 1014.28
R3524 Vbias.n3631 Vbias.n3630 1014.28
R3525 Vbias.n3632 Vbias.n3631 1014.28
R3526 Vbias.n3640 Vbias.n3638 1014.28
R3527 Vbias.n3640 Vbias.n3639 1014.28
R3528 Vbias.n3669 Vbias.n3668 1014.28
R3529 Vbias.n3670 Vbias.n3669 1014.28
R3530 Vbias.n3678 Vbias.n3676 1014.28
R3531 Vbias.n3678 Vbias.n3677 1014.28
R3532 Vbias.n4064 Vbias.n4062 1014.28
R3533 Vbias.n4064 Vbias.n4056 1014.28
R3534 Vbias.n4067 Vbias.n4063 1014.28
R3535 Vbias.n4067 Vbias.n4057 1014.28
R3536 Vbias.n4208 Vbias.n4042 1014.28
R3537 Vbias.n4208 Vbias.n4043 1014.28
R3538 Vbias.n4022 Vbias.n4020 1014.28
R3539 Vbias.n4022 Vbias.n4014 1014.28
R3540 Vbias.n4025 Vbias.n4021 1014.28
R3541 Vbias.n4025 Vbias.n4015 1014.28
R3542 Vbias.n3990 Vbias.n3989 1014.28
R3543 Vbias.n3990 Vbias.n3984 1014.28
R3544 Vbias.n3998 Vbias.n3993 1014.28
R3545 Vbias.n3998 Vbias.n3997 1014.28
R3546 Vbias.n4175 Vbias.n4174 1014.28
R3547 Vbias.n4174 Vbias.n4173 1014.28
R3548 Vbias.n4076 Vbias.n4075 1014.28
R3549 Vbias.n4076 Vbias.n4072 1014.28
R3550 Vbias.n4147 Vbias.n4044 1014.28
R3551 Vbias.n4157 Vbias.n4044 1014.28
R3552 Vbias.n4131 Vbias.n4130 1014.28
R3553 Vbias.n4132 Vbias.n4131 1014.28
R3554 Vbias.n4083 Vbias.n4081 1014.28
R3555 Vbias.n4083 Vbias.n4082 1014.28
R3556 Vbias.n4097 Vbias.n4095 1014.28
R3557 Vbias.n4097 Vbias.n4096 1014.28
R3558 Vbias.n4093 Vbias.n4091 1014.28
R3559 Vbias.n4093 Vbias.n4092 1014.28
R3560 Vbias.n4972 Vbias.n2615 1014.28
R3561 Vbias.n4972 Vbias.n2613 1014.28
R3562 Vbias.n4979 Vbias.n2607 1014.28
R3563 Vbias.n4979 Vbias.n2611 1014.28
R3564 Vbias.n4961 Vbias.n2621 1014.28
R3565 Vbias.n4961 Vbias.n2629 1014.28
R3566 Vbias.n4935 Vbias.n2641 1014.28
R3567 Vbias.n4935 Vbias.n4934 1014.28
R3568 Vbias.n4949 Vbias.n2637 1014.28
R3569 Vbias.n4949 Vbias.n2638 1014.28
R3570 Vbias.n4913 Vbias.n2655 1014.28
R3571 Vbias.n4913 Vbias.n4912 1014.28
R3572 Vbias.n4926 Vbias.n2651 1014.28
R3573 Vbias.n4926 Vbias.n2652 1014.28
R3574 Vbias.n3002 Vbias.n2999 1014.28
R3575 Vbias.n3002 Vbias.n2994 1014.28
R3576 Vbias.n3005 Vbias.n3000 1014.28
R3577 Vbias.n3005 Vbias.n2995 1014.28
R3578 Vbias.n3074 Vbias.n2976 1014.28
R3579 Vbias.n3074 Vbias.n2977 1014.28
R3580 Vbias.n2955 Vbias.n2952 1014.28
R3581 Vbias.n2955 Vbias.n2947 1014.28
R3582 Vbias.n2958 Vbias.n2953 1014.28
R3583 Vbias.n2958 Vbias.n2948 1014.28
R3584 Vbias.n2926 Vbias.n2923 1014.28
R3585 Vbias.n2926 Vbias.n2918 1014.28
R3586 Vbias.n2929 Vbias.n2924 1014.28
R3587 Vbias.n2929 Vbias.n2919 1014.28
R3588 Vbias.n3016 Vbias.n3015 1014.28
R3589 Vbias.n3017 Vbias.n3016 1014.28
R3590 Vbias.n3025 Vbias.n3023 1014.28
R3591 Vbias.n3025 Vbias.n3024 1014.28
R3592 Vbias.n2979 Vbias.n2978 1014.28
R3593 Vbias.n3061 Vbias.n2978 1014.28
R3594 Vbias.n3092 Vbias.n3091 1014.28
R3595 Vbias.n3093 Vbias.n3092 1014.28
R3596 Vbias.n3101 Vbias.n3099 1014.28
R3597 Vbias.n3101 Vbias.n3100 1014.28
R3598 Vbias.n3130 Vbias.n3129 1014.28
R3599 Vbias.n3131 Vbias.n3130 1014.28
R3600 Vbias.n3139 Vbias.n3137 1014.28
R3601 Vbias.n3139 Vbias.n3138 1014.28
R3602 Vbias.n2763 Vbias.n2760 1014.28
R3603 Vbias.n2763 Vbias.n2755 1014.28
R3604 Vbias.n2766 Vbias.n2761 1014.28
R3605 Vbias.n2766 Vbias.n2756 1014.28
R3606 Vbias.n4750 Vbias.n2737 1014.28
R3607 Vbias.n4750 Vbias.n2738 1014.28
R3608 Vbias.n2716 Vbias.n2713 1014.28
R3609 Vbias.n2716 Vbias.n2708 1014.28
R3610 Vbias.n2719 Vbias.n2714 1014.28
R3611 Vbias.n2719 Vbias.n2709 1014.28
R3612 Vbias.n2687 Vbias.n2684 1014.28
R3613 Vbias.n2687 Vbias.n2679 1014.28
R3614 Vbias.n2690 Vbias.n2685 1014.28
R3615 Vbias.n2690 Vbias.n2680 1014.28
R3616 Vbias.n4692 Vbias.n4691 1014.28
R3617 Vbias.n4693 Vbias.n4692 1014.28
R3618 Vbias.n4701 Vbias.n4699 1014.28
R3619 Vbias.n4701 Vbias.n4700 1014.28
R3620 Vbias.n2740 Vbias.n2739 1014.28
R3621 Vbias.n4737 Vbias.n2739 1014.28
R3622 Vbias.n4768 Vbias.n4767 1014.28
R3623 Vbias.n4769 Vbias.n4768 1014.28
R3624 Vbias.n4777 Vbias.n4775 1014.28
R3625 Vbias.n4777 Vbias.n4776 1014.28
R3626 Vbias.n4806 Vbias.n4805 1014.28
R3627 Vbias.n4807 Vbias.n4806 1014.28
R3628 Vbias.n4815 Vbias.n4813 1014.28
R3629 Vbias.n4815 Vbias.n4814 1014.28
R3630 Vbias.n4564 Vbias.n4561 1014.28
R3631 Vbias.n4564 Vbias.n4562 1014.28
R3632 Vbias.n4572 Vbias.n4570 1014.28
R3633 Vbias.n4572 Vbias.n4571 1014.28
R3634 Vbias.n6216 Vbias.n6213 1014.28
R3635 Vbias.n6216 Vbias.n6214 1014.28
R3636 Vbias.n6224 Vbias.n6222 1014.28
R3637 Vbias.n6224 Vbias.n6223 1014.28
R3638 Vbias.n6200 Vbias.n6196 1014.28
R3639 Vbias.n6200 Vbias.n6197 1014.28
R3640 Vbias.n6174 Vbias.n6168 1014.28
R3641 Vbias.n6174 Vbias.n6173 1014.28
R3642 Vbias.n6177 Vbias.n6166 1014.28
R3643 Vbias.n6177 Vbias.n6176 1014.28
R3644 Vbias.n6453 Vbias.n6450 1014.28
R3645 Vbias.n6453 Vbias.n6451 1014.28
R3646 Vbias.n6461 Vbias.n6459 1014.28
R3647 Vbias.n6461 Vbias.n6460 1014.28
R3648 Vbias.n6437 Vbias.n6433 1014.28
R3649 Vbias.n6437 Vbias.n6434 1014.28
R3650 Vbias.n6411 Vbias.n6386 1014.28
R3651 Vbias.n6411 Vbias.n6410 1014.28
R3652 Vbias.n6414 Vbias.n6384 1014.28
R3653 Vbias.n6414 Vbias.n6413 1014.28
R3654 Vbias.n6394 Vbias.n6389 1014.28
R3655 Vbias.n6394 Vbias.n6393 1014.28
R3656 Vbias.n6397 Vbias.n6387 1014.28
R3657 Vbias.n6397 Vbias.n6396 1014.28
R3658 Vbias.n907 Vbias.n904 1014.28
R3659 Vbias.n907 Vbias.n905 1014.28
R3660 Vbias.n915 Vbias.n913 1014.28
R3661 Vbias.n915 Vbias.n914 1014.28
R3662 Vbias.n891 Vbias.n887 1014.28
R3663 Vbias.n891 Vbias.n888 1014.28
R3664 Vbias.n6473 Vbias.n6469 1014.28
R3665 Vbias.n6473 Vbias.n6472 1014.28
R3666 Vbias.n6482 Vbias.n6471 1014.28
R3667 Vbias.n6482 Vbias.n6481 1014.28
R3668 Vbias.n6467 Vbias.n6463 1014.28
R3669 Vbias.n6467 Vbias.n6466 1014.28
R3670 Vbias.n6496 Vbias.n6465 1014.28
R3671 Vbias.n6496 Vbias.n6495 1014.28
R3672 Vbias.n7393 Vbias.n7391 1014.28
R3673 Vbias.n7393 Vbias.n7387 1014.28
R3674 Vbias.n7396 Vbias.n7392 1014.28
R3675 Vbias.n7396 Vbias.n7388 1014.28
R3676 Vbias.n7423 Vbias.n7372 1014.28
R3677 Vbias.n7423 Vbias.n7373 1014.28
R3678 Vbias.n7355 Vbias.n7353 1014.28
R3679 Vbias.n7355 Vbias.n7349 1014.28
R3680 Vbias.n7358 Vbias.n7354 1014.28
R3681 Vbias.n7358 Vbias.n7350 1014.28
R3682 Vbias.n7331 Vbias.n7330 1014.28
R3683 Vbias.n7331 Vbias.n7328 1014.28
R3684 Vbias.n7337 Vbias.n7334 1014.28
R3685 Vbias.n7337 Vbias.n7336 1014.28
R3686 Vbias.n6644 Vbias.n6139 1014.28
R3687 Vbias.n6644 Vbias.n6140 1014.28
R3688 Vbias.n6151 Vbias.n6146 1014.28
R3689 Vbias.n6152 Vbias.n6151 1014.28
R3690 Vbias.n1722 Vbias.n1713 1014.28
R3691 Vbias.n1722 Vbias.n1710 1014.28
R3692 Vbias.n1712 Vbias.n1711 1014.28
R3693 Vbias.n1711 Vbias.n1709 1014.28
R3694 Vbias.n6685 Vbias.n1453 1014.28
R3695 Vbias.n6685 Vbias.n1454 1014.28
R3696 Vbias.n4377 Vbias.n2798 1010.98
R3697 Vbias.n4377 Vbias.n2791 1010.98
R3698 Vbias.n4392 Vbias.n2791 1010.98
R3699 Vbias.n4392 Vbias.n2779 1010.98
R3700 Vbias.n4369 Vbias.n2792 1010.98
R3701 Vbias.n4397 Vbias.n2792 1010.98
R3702 Vbias.n4397 Vbias.n2793 1010.98
R3703 Vbias.n2793 Vbias.n2778 1010.98
R3704 Vbias.n2816 Vbias.n2811 1010.98
R3705 Vbias.n2816 Vbias.n2804 1010.98
R3706 Vbias.n4339 Vbias.n2815 1010.98
R3707 Vbias.n2815 Vbias.n2803 1010.98
R3708 Vbias.n2853 Vbias.n2843 1010.98
R3709 Vbias.n4323 Vbias.n2843 1010.98
R3710 Vbias.n4323 Vbias.n2828 1010.98
R3711 Vbias.n4330 Vbias.n2828 1010.98
R3712 Vbias.n4306 Vbias.n2839 1010.98
R3713 Vbias.n4324 Vbias.n2839 1010.98
R3714 Vbias.n4324 Vbias.n2835 1010.98
R3715 Vbias.n4329 Vbias.n2835 1010.98
R3716 Vbias.n2887 Vbias.n2877 1010.98
R3717 Vbias.n4290 Vbias.n2877 1010.98
R3718 Vbias.n4290 Vbias.n2864 1010.98
R3719 Vbias.n4297 Vbias.n2864 1010.98
R3720 Vbias.n4273 Vbias.n2873 1010.98
R3721 Vbias.n4291 Vbias.n2873 1010.98
R3722 Vbias.n4291 Vbias.n2869 1010.98
R3723 Vbias.n4296 Vbias.n2869 1010.98
R3724 Vbias.n4370 Vbias.n2784 1010.98
R3725 Vbias.n4398 Vbias.n2784 1010.98
R3726 Vbias.n4399 Vbias.n4398 1010.98
R3727 Vbias.n4400 Vbias.n4399 1010.98
R3728 Vbias.n4373 Vbias.n2799 1010.98
R3729 Vbias.n4373 Vbias.n2789 1010.98
R3730 Vbias.n2789 Vbias.n2788 1010.98
R3731 Vbias.n2788 Vbias.n2787 1010.98
R3732 Vbias.n4345 Vbias.n2818 1010.98
R3733 Vbias.n4347 Vbias.n2818 1010.98
R3734 Vbias.n2817 Vbias.n2812 1010.98
R3735 Vbias.n2817 Vbias.n2808 1010.98
R3736 Vbias.n4307 Vbias.n2848 1010.98
R3737 Vbias.n2848 Vbias.n2842 1010.98
R3738 Vbias.n4316 Vbias.n2842 1010.98
R3739 Vbias.n4316 Vbias.n2831 1010.98
R3740 Vbias.n2852 Vbias.n2851 1010.98
R3741 Vbias.n2851 Vbias.n2841 1010.98
R3742 Vbias.n4315 Vbias.n2841 1010.98
R3743 Vbias.n4315 Vbias.n2826 1010.98
R3744 Vbias.n4274 Vbias.n2882 1010.98
R3745 Vbias.n2882 Vbias.n2876 1010.98
R3746 Vbias.n4283 Vbias.n2876 1010.98
R3747 Vbias.n4283 Vbias.n2867 1010.98
R3748 Vbias.n2886 Vbias.n2885 1010.98
R3749 Vbias.n2885 Vbias.n2875 1010.98
R3750 Vbias.n4282 Vbias.n2875 1010.98
R3751 Vbias.n4282 Vbias.n2862 1010.98
R3752 Vbias.n1686 Vbias.n1682 1010.98
R3753 Vbias.n5860 Vbias.n1686 1010.98
R3754 Vbias.n1692 Vbias.n1685 1010.98
R3755 Vbias.n5864 Vbias.n1685 1010.98
R3756 Vbias.n5516 Vbias.n5510 1010.98
R3757 Vbias.n5525 Vbias.n5516 1010.98
R3758 Vbias.n5519 Vbias.n5509 1010.98
R3759 Vbias.n5524 Vbias.n5519 1010.98
R3760 Vbias.n2239 Vbias.n2235 1010.98
R3761 Vbias.n5536 Vbias.n2239 1010.98
R3762 Vbias.n2245 Vbias.n2238 1010.98
R3763 Vbias.n5540 Vbias.n2238 1010.98
R3764 Vbias.n2591 Vbias.n2587 1010.98
R3765 Vbias.n5017 Vbias.n2591 1010.98
R3766 Vbias.n5015 Vbias.n2590 1010.98
R3767 Vbias.n5021 Vbias.n2590 1010.98
R3768 Vbias.n5001 Vbias.n2599 1010.98
R3769 Vbias.n2599 Vbias.n2594 1010.98
R3770 Vbias.n5000 Vbias.n4995 1010.98
R3771 Vbias.n4995 Vbias.n2593 1010.98
R3772 Vbias.n158 Vbias.n154 1010.98
R3773 Vbias.n7954 Vbias.n154 1010.98
R3774 Vbias.n7954 Vbias.n155 1010.98
R3775 Vbias.n7950 Vbias.n155 1010.98
R3776 Vbias.n149 Vbias.n146 1010.98
R3777 Vbias.n7955 Vbias.n149 1010.98
R3778 Vbias.n7955 Vbias.n150 1010.98
R3779 Vbias.n7949 Vbias.n150 1010.98
R3780 Vbias.n135 Vbias.n131 1010.98
R3781 Vbias.n7964 Vbias.n135 1010.98
R3782 Vbias.n140 Vbias.n130 1010.98
R3783 Vbias.n7963 Vbias.n140 1010.98
R3784 Vbias.n114 Vbias.n110 1010.98
R3785 Vbias.n7979 Vbias.n114 1010.98
R3786 Vbias.n7979 Vbias.n115 1010.98
R3787 Vbias.n7973 Vbias.n115 1010.98
R3788 Vbias.n119 Vbias.n109 1010.98
R3789 Vbias.n7978 Vbias.n119 1010.98
R3790 Vbias.n7978 Vbias.n120 1010.98
R3791 Vbias.n7974 Vbias.n120 1010.98
R3792 Vbias.n95 Vbias.n91 1010.98
R3793 Vbias.n7994 Vbias.n95 1010.98
R3794 Vbias.n7994 Vbias.n96 1010.98
R3795 Vbias.n7988 Vbias.n96 1010.98
R3796 Vbias.n100 Vbias.n90 1010.98
R3797 Vbias.n7993 Vbias.n100 1010.98
R3798 Vbias.n7993 Vbias.n101 1010.98
R3799 Vbias.n7989 Vbias.n101 1010.98
R3800 Vbias.n73 Vbias.n67 1010.98
R3801 Vbias.n8017 Vbias.n73 1010.98
R3802 Vbias.n8017 Vbias.n74 1010.98
R3803 Vbias.n8011 Vbias.n74 1010.98
R3804 Vbias.n77 Vbias.n66 1010.98
R3805 Vbias.n8016 Vbias.n77 1010.98
R3806 Vbias.n8016 Vbias.n78 1010.98
R3807 Vbias.n8012 Vbias.n78 1010.98
R3808 Vbias.n63 Vbias.n58 1010.98
R3809 Vbias.n8032 Vbias.n63 1010.98
R3810 Vbias.n8026 Vbias.n57 1010.98
R3811 Vbias.n8031 Vbias.n8026 1010.98
R3812 Vbias.n36 Vbias.n32 1010.98
R3813 Vbias.n42 Vbias.n36 1010.98
R3814 Vbias.n49 Vbias.n42 1010.98
R3815 Vbias.n8048 Vbias.n49 1010.98
R3816 Vbias.n40 Vbias.n35 1010.98
R3817 Vbias.n8053 Vbias.n35 1010.98
R3818 Vbias.n8053 Vbias.n43 1010.98
R3819 Vbias.n8049 Vbias.n43 1010.98
R3820 Vbias.n17 Vbias.n11 1010.98
R3821 Vbias.n8069 Vbias.n17 1010.98
R3822 Vbias.n8069 Vbias.n18 1010.98
R3823 Vbias.n8063 Vbias.n18 1010.98
R3824 Vbias.n22 Vbias.n10 1010.98
R3825 Vbias.n8068 Vbias.n22 1010.98
R3826 Vbias.n8068 Vbias.n23 1010.98
R3827 Vbias.n8064 Vbias.n23 1010.98
R3828 Vbias.n6707 Vbias.n6696 1010.98
R3829 Vbias.n6707 Vbias.n6698 1010.98
R3830 Vbias.n6706 Vbias.n6705 1010.98
R3831 Vbias.n6706 Vbias.n6700 1010.98
R3832 Vbias.n6733 Vbias.n6720 1010.98
R3833 Vbias.n6733 Vbias.n6722 1010.98
R3834 Vbias.n6732 Vbias.n6731 1010.98
R3835 Vbias.n6732 Vbias.n6724 1010.98
R3836 Vbias.n1742 Vbias.n1741 1010.98
R3837 Vbias.n1741 Vbias.n1726 1010.98
R3838 Vbias.n1732 Vbias.n1726 1010.98
R3839 Vbias.n1733 Vbias.n1732 1010.98
R3840 Vbias.n1738 Vbias.n1727 1010.98
R3841 Vbias.n2044 Vbias.n1727 1010.98
R3842 Vbias.n2044 Vbias.n1728 1010.98
R3843 Vbias.n2038 Vbias.n1728 1010.98
R3844 Vbias.n5846 Vbias.n2067 1010.98
R3845 Vbias.n2067 Vbias.n1695 1010.98
R3846 Vbias.n2062 Vbias.n1695 1010.98
R3847 Vbias.n5852 Vbias.n2062 1010.98
R3848 Vbias.n5845 Vbias.n1696 1010.98
R3849 Vbias.n5857 Vbias.n1696 1010.98
R3850 Vbias.n5857 Vbias.n1697 1010.98
R3851 Vbias.n5853 Vbias.n1697 1010.98
R3852 Vbias.n675 Vbias.n669 1010.98
R3853 Vbias.n7744 Vbias.n675 1010.98
R3854 Vbias.n7738 Vbias.n668 1010.98
R3855 Vbias.n7743 Vbias.n7738 1010.98
R3856 Vbias.n5793 Vbias.n2079 1010.98
R3857 Vbias.n5819 Vbias.n2079 1010.98
R3858 Vbias.n5819 Vbias.n2075 1010.98
R3859 Vbias.n5823 Vbias.n2075 1010.98
R3860 Vbias.n2085 Vbias.n2081 1010.98
R3861 Vbias.n5818 Vbias.n2081 1010.98
R3862 Vbias.n5818 Vbias.n2072 1010.98
R3863 Vbias.n5824 Vbias.n2072 1010.98
R3864 Vbias.n5805 Vbias.n5797 1010.98
R3865 Vbias.n5809 Vbias.n5797 1010.98
R3866 Vbias.n5804 Vbias.n5789 1010.98
R3867 Vbias.n5810 Vbias.n5789 1010.98
R3868 Vbias.n2109 Vbias.n2093 1010.98
R3869 Vbias.n5776 Vbias.n2093 1010.98
R3870 Vbias.n5776 Vbias.n2090 1010.98
R3871 Vbias.n5780 Vbias.n2090 1010.98
R3872 Vbias.n2101 Vbias.n2097 1010.98
R3873 Vbias.n5775 Vbias.n2097 1010.98
R3874 Vbias.n5775 Vbias.n2089 1010.98
R3875 Vbias.n5782 Vbias.n2089 1010.98
R3876 Vbias.n5748 Vbias.n2117 1010.98
R3877 Vbias.n5762 Vbias.n2117 1010.98
R3878 Vbias.n5762 Vbias.n2113 1010.98
R3879 Vbias.n5766 Vbias.n2113 1010.98
R3880 Vbias.n2123 Vbias.n2119 1010.98
R3881 Vbias.n5761 Vbias.n2119 1010.98
R3882 Vbias.n5761 Vbias.n2105 1010.98
R3883 Vbias.n5767 Vbias.n2105 1010.98
R3884 Vbias.n564 Vbias.n560 1010.98
R3885 Vbias.n7804 Vbias.n564 1010.98
R3886 Vbias.n570 Vbias.n563 1010.98
R3887 Vbias.n7808 Vbias.n563 1010.98
R3888 Vbias.n2148 Vbias.n2134 1010.98
R3889 Vbias.n5730 Vbias.n2134 1010.98
R3890 Vbias.n5730 Vbias.n2130 1010.98
R3891 Vbias.n5734 Vbias.n2130 1010.98
R3892 Vbias.n2140 Vbias.n2136 1010.98
R3893 Vbias.n5729 Vbias.n2136 1010.98
R3894 Vbias.n5729 Vbias.n2127 1010.98
R3895 Vbias.n5735 Vbias.n2127 1010.98
R3896 Vbias.n5716 Vbias.n2152 1010.98
R3897 Vbias.n5720 Vbias.n2152 1010.98
R3898 Vbias.n5715 Vbias.n2144 1010.98
R3899 Vbias.n5721 Vbias.n2144 1010.98
R3900 Vbias.n5696 Vbias.n2162 1010.98
R3901 Vbias.n5706 Vbias.n2162 1010.98
R3902 Vbias.n5706 Vbias.n2163 1010.98
R3903 Vbias.n2163 Vbias.n2158 1010.98
R3904 Vbias.n5697 Vbias.n2166 1010.98
R3905 Vbias.n5705 Vbias.n2166 1010.98
R3906 Vbias.n5705 Vbias.n2168 1010.98
R3907 Vbias.n2168 Vbias.n2157 1010.98
R3908 Vbias.n5678 Vbias.n2180 1010.98
R3909 Vbias.n5687 Vbias.n2180 1010.98
R3910 Vbias.n5687 Vbias.n2181 1010.98
R3911 Vbias.n2181 Vbias.n2176 1010.98
R3912 Vbias.n5679 Vbias.n2184 1010.98
R3913 Vbias.n5686 Vbias.n2184 1010.98
R3914 Vbias.n5686 Vbias.n2186 1010.98
R3915 Vbias.n2186 Vbias.n2175 1010.98
R3916 Vbias.n454 Vbias.n449 1010.98
R3917 Vbias.n7879 Vbias.n454 1010.98
R3918 Vbias.n7873 Vbias.n448 1010.98
R3919 Vbias.n7878 Vbias.n7873 1010.98
R3920 Vbias.n2219 Vbias.n2205 1010.98
R3921 Vbias.n5656 Vbias.n2205 1010.98
R3922 Vbias.n5656 Vbias.n2201 1010.98
R3923 Vbias.n5660 Vbias.n2201 1010.98
R3924 Vbias.n2211 Vbias.n2207 1010.98
R3925 Vbias.n5655 Vbias.n2207 1010.98
R3926 Vbias.n5655 Vbias.n2198 1010.98
R3927 Vbias.n5661 Vbias.n2198 1010.98
R3928 Vbias.n5642 Vbias.n2223 1010.98
R3929 Vbias.n5646 Vbias.n2223 1010.98
R3930 Vbias.n5641 Vbias.n2215 1010.98
R3931 Vbias.n5647 Vbias.n2215 1010.98
R3932 Vbias.n5622 Vbias.n5559 1010.98
R3933 Vbias.n5632 Vbias.n5559 1010.98
R3934 Vbias.n5632 Vbias.n5560 1010.98
R3935 Vbias.n5560 Vbias.n5555 1010.98
R3936 Vbias.n5623 Vbias.n5563 1010.98
R3937 Vbias.n5631 Vbias.n5563 1010.98
R3938 Vbias.n5631 Vbias.n5565 1010.98
R3939 Vbias.n5565 Vbias.n5554 1010.98
R3940 Vbias.n5604 Vbias.n5577 1010.98
R3941 Vbias.n5613 Vbias.n5577 1010.98
R3942 Vbias.n5613 Vbias.n5578 1010.98
R3943 Vbias.n5578 Vbias.n5573 1010.98
R3944 Vbias.n5605 Vbias.n5581 1010.98
R3945 Vbias.n5612 Vbias.n5581 1010.98
R3946 Vbias.n5612 Vbias.n5583 1010.98
R3947 Vbias.n5583 Vbias.n5572 1010.98
R3948 Vbias.n331 Vbias.n329 1010.98
R3949 Vbias.n331 Vbias.n171 1010.98
R3950 Vbias.n330 Vbias.n328 1010.98
R3951 Vbias.n330 Vbias.n173 1010.98
R3952 Vbias.n1013 Vbias.n919 1010.98
R3953 Vbias.n922 Vbias.n919 1010.98
R3954 Vbias.n1012 Vbias.n918 1010.98
R3955 Vbias.n1024 Vbias.n918 1010.98
R3956 Vbias.n6525 Vbias.n6520 1010.98
R3957 Vbias.n6525 Vbias.n926 1010.98
R3958 Vbias.n6530 Vbias.n6522 1010.98
R3959 Vbias.n6522 Vbias.n928 1010.98
R3960 Vbias.n6596 Vbias.n773 1010.98
R3961 Vbias.n6596 Vbias.n775 1010.98
R3962 Vbias.n6595 Vbias.n6594 1010.98
R3963 Vbias.n6595 Vbias.n777 1010.98
R3964 Vbias.n767 Vbias.n758 1010.98
R3965 Vbias.n7662 Vbias.n767 1010.98
R3966 Vbias.n7667 Vbias.n760 1010.98
R3967 Vbias.n7663 Vbias.n760 1010.98
R3968 Vbias.n7255 Vbias.n7251 1010.98
R3969 Vbias.n7270 Vbias.n7251 1010.98
R3970 Vbias.n7270 Vbias.n7252 1010.98
R3971 Vbias.n7266 Vbias.n7252 1010.98
R3972 Vbias.n7246 Vbias.n7243 1010.98
R3973 Vbias.n7271 Vbias.n7246 1010.98
R3974 Vbias.n7271 Vbias.n7247 1010.98
R3975 Vbias.n7264 Vbias.n7247 1010.98
R3976 Vbias.n7232 Vbias.n7228 1010.98
R3977 Vbias.n7280 Vbias.n7232 1010.98
R3978 Vbias.n7237 Vbias.n7227 1010.98
R3979 Vbias.n7279 Vbias.n7237 1010.98
R3980 Vbias.n1055 Vbias.n1051 1010.98
R3981 Vbias.n7295 Vbias.n1055 1010.98
R3982 Vbias.n7295 Vbias.n1056 1010.98
R3983 Vbias.n7289 Vbias.n1056 1010.98
R3984 Vbias.n1060 Vbias.n1050 1010.98
R3985 Vbias.n7294 Vbias.n1060 1010.98
R3986 Vbias.n7294 Vbias.n1061 1010.98
R3987 Vbias.n7290 Vbias.n1061 1010.98
R3988 Vbias.n1034 Vbias.n1030 1010.98
R3989 Vbias.n7310 Vbias.n1034 1010.98
R3990 Vbias.n7310 Vbias.n1035 1010.98
R3991 Vbias.n7304 Vbias.n1035 1010.98
R3992 Vbias.n1039 Vbias.n1029 1010.98
R3993 Vbias.n7309 Vbias.n1039 1010.98
R3994 Vbias.n7309 Vbias.n1040 1010.98
R3995 Vbias.n7305 Vbias.n1040 1010.98
R3996 Vbias.n1005 Vbias.n1001 1010.98
R3997 Vbias.n7476 Vbias.n1001 1010.98
R3998 Vbias.n7476 Vbias.n1002 1010.98
R3999 Vbias.n7472 Vbias.n1002 1010.98
R4000 Vbias.n996 Vbias.n993 1010.98
R4001 Vbias.n7477 Vbias.n996 1010.98
R4002 Vbias.n7477 Vbias.n997 1010.98
R4003 Vbias.n7471 Vbias.n997 1010.98
R4004 Vbias.n982 Vbias.n978 1010.98
R4005 Vbias.n7486 Vbias.n982 1010.98
R4006 Vbias.n987 Vbias.n977 1010.98
R4007 Vbias.n7485 Vbias.n987 1010.98
R4008 Vbias.n960 Vbias.n956 1010.98
R4009 Vbias.n7502 Vbias.n960 1010.98
R4010 Vbias.n7502 Vbias.n961 1010.98
R4011 Vbias.n7496 Vbias.n961 1010.98
R4012 Vbias.n965 Vbias.n955 1010.98
R4013 Vbias.n7501 Vbias.n965 1010.98
R4014 Vbias.n7501 Vbias.n966 1010.98
R4015 Vbias.n7497 Vbias.n966 1010.98
R4016 Vbias.n937 Vbias.n933 1010.98
R4017 Vbias.n7517 Vbias.n937 1010.98
R4018 Vbias.n7517 Vbias.n938 1010.98
R4019 Vbias.n7511 Vbias.n938 1010.98
R4020 Vbias.n942 Vbias.n932 1010.98
R4021 Vbias.n7516 Vbias.n942 1010.98
R4022 Vbias.n7516 Vbias.n943 1010.98
R4023 Vbias.n7512 Vbias.n943 1010.98
R4024 Vbias.n850 Vbias.n846 1010.98
R4025 Vbias.n7598 Vbias.n846 1010.98
R4026 Vbias.n7598 Vbias.n847 1010.98
R4027 Vbias.n7594 Vbias.n847 1010.98
R4028 Vbias.n841 Vbias.n838 1010.98
R4029 Vbias.n7599 Vbias.n841 1010.98
R4030 Vbias.n7599 Vbias.n842 1010.98
R4031 Vbias.n7593 Vbias.n842 1010.98
R4032 Vbias.n827 Vbias.n823 1010.98
R4033 Vbias.n7608 Vbias.n827 1010.98
R4034 Vbias.n832 Vbias.n822 1010.98
R4035 Vbias.n7607 Vbias.n832 1010.98
R4036 Vbias.n805 Vbias.n801 1010.98
R4037 Vbias.n7623 Vbias.n805 1010.98
R4038 Vbias.n7623 Vbias.n806 1010.98
R4039 Vbias.n7617 Vbias.n806 1010.98
R4040 Vbias.n810 Vbias.n800 1010.98
R4041 Vbias.n7622 Vbias.n810 1010.98
R4042 Vbias.n7622 Vbias.n811 1010.98
R4043 Vbias.n7618 Vbias.n811 1010.98
R4044 Vbias.n786 Vbias.n782 1010.98
R4045 Vbias.n7638 Vbias.n786 1010.98
R4046 Vbias.n7638 Vbias.n787 1010.98
R4047 Vbias.n7632 Vbias.n787 1010.98
R4048 Vbias.n791 Vbias.n781 1010.98
R4049 Vbias.n7637 Vbias.n791 1010.98
R4050 Vbias.n7637 Vbias.n792 1010.98
R4051 Vbias.n7633 Vbias.n792 1010.98
R4052 Vbias.n6355 Vbias.n6232 1010.98
R4053 Vbias.n6583 Vbias.n6232 1010.98
R4054 Vbias.n6583 Vbias.n6233 1010.98
R4055 Vbias.n6233 Vbias.n6228 1010.98
R4056 Vbias.n6356 Vbias.n6236 1010.98
R4057 Vbias.n6582 Vbias.n6236 1010.98
R4058 Vbias.n6582 Vbias.n6238 1010.98
R4059 Vbias.n6238 Vbias.n6227 1010.98
R4060 Vbias.n6346 Vbias.n6251 1010.98
R4061 Vbias.n6251 Vbias.n6246 1010.98
R4062 Vbias.n6345 Vbias.n6255 1010.98
R4063 Vbias.n6255 Vbias.n6245 1010.98
R4064 Vbias.n6282 Vbias.n6268 1010.98
R4065 Vbias.n6333 Vbias.n6268 1010.98
R4066 Vbias.n6333 Vbias.n6264 1010.98
R4067 Vbias.n6337 Vbias.n6264 1010.98
R4068 Vbias.n6274 Vbias.n6270 1010.98
R4069 Vbias.n6332 Vbias.n6270 1010.98
R4070 Vbias.n6332 Vbias.n6260 1010.98
R4071 Vbias.n6338 Vbias.n6260 1010.98
R4072 Vbias.n6305 Vbias.n6290 1010.98
R4073 Vbias.n6319 Vbias.n6290 1010.98
R4074 Vbias.n6319 Vbias.n6286 1010.98
R4075 Vbias.n6323 Vbias.n6286 1010.98
R4076 Vbias.n6296 Vbias.n6292 1010.98
R4077 Vbias.n6318 Vbias.n6292 1010.98
R4078 Vbias.n6318 Vbias.n6278 1010.98
R4079 Vbias.n6324 Vbias.n6278 1010.98
R4080 Vbias.n1494 Vbias.n1491 1010.98
R4081 Vbias.n6659 Vbias.n1491 1010.98
R4082 Vbias.n6659 Vbias.n1492 1010.98
R4083 Vbias.n6655 Vbias.n1492 1010.98
R4084 Vbias.n1486 Vbias.n1483 1010.98
R4085 Vbias.n6660 Vbias.n1486 1010.98
R4086 Vbias.n6660 Vbias.n1487 1010.98
R4087 Vbias.n6654 Vbias.n1487 1010.98
R4088 Vbias.n1473 Vbias.n1469 1010.98
R4089 Vbias.n6669 Vbias.n1473 1010.98
R4090 Vbias.n1478 Vbias.n1468 1010.98
R4091 Vbias.n6668 Vbias.n1478 1010.98
R4092 Vbias.n742 Vbias.n736 1010.98
R4093 Vbias.n7677 Vbias.n742 1010.98
R4094 Vbias.n7677 Vbias.n743 1010.98
R4095 Vbias.n7671 Vbias.n743 1010.98
R4096 Vbias.n746 Vbias.n735 1010.98
R4097 Vbias.n7676 Vbias.n746 1010.98
R4098 Vbias.n7676 Vbias.n747 1010.98
R4099 Vbias.n7672 Vbias.n747 1010.98
R4100 Vbias.n732 Vbias.n727 1010.98
R4101 Vbias.n7692 Vbias.n732 1010.98
R4102 Vbias.n7686 Vbias.n726 1010.98
R4103 Vbias.n7691 Vbias.n7686 1010.98
R4104 Vbias.n705 Vbias.n701 1010.98
R4105 Vbias.n711 Vbias.n705 1010.98
R4106 Vbias.n718 Vbias.n711 1010.98
R4107 Vbias.n7708 Vbias.n718 1010.98
R4108 Vbias.n709 Vbias.n704 1010.98
R4109 Vbias.n7713 Vbias.n704 1010.98
R4110 Vbias.n7713 Vbias.n712 1010.98
R4111 Vbias.n7709 Vbias.n712 1010.98
R4112 Vbias.n686 Vbias.n680 1010.98
R4113 Vbias.n7729 Vbias.n686 1010.98
R4114 Vbias.n7729 Vbias.n687 1010.98
R4115 Vbias.n7723 Vbias.n687 1010.98
R4116 Vbias.n691 Vbias.n679 1010.98
R4117 Vbias.n7728 Vbias.n691 1010.98
R4118 Vbias.n7728 Vbias.n692 1010.98
R4119 Vbias.n7724 Vbias.n692 1010.98
R4120 Vbias.n655 Vbias.n644 1010.98
R4121 Vbias.n655 Vbias.n649 1010.98
R4122 Vbias.n664 Vbias.n649 1010.98
R4123 Vbias.n664 Vbias.n651 1010.98
R4124 Vbias.n654 Vbias.n643 1010.98
R4125 Vbias.n662 Vbias.n654 1010.98
R4126 Vbias.n663 Vbias.n662 1010.98
R4127 Vbias.n663 Vbias.n653 1010.98
R4128 Vbias.n640 Vbias.n627 1010.98
R4129 Vbias.n640 Vbias.n629 1010.98
R4130 Vbias.n639 Vbias.n638 1010.98
R4131 Vbias.n639 Vbias.n631 1010.98
R4132 Vbias.n608 Vbias.n597 1010.98
R4133 Vbias.n608 Vbias.n602 1010.98
R4134 Vbias.n617 Vbias.n602 1010.98
R4135 Vbias.n617 Vbias.n604 1010.98
R4136 Vbias.n607 Vbias.n596 1010.98
R4137 Vbias.n615 Vbias.n607 1010.98
R4138 Vbias.n616 Vbias.n615 1010.98
R4139 Vbias.n616 Vbias.n606 1010.98
R4140 Vbias.n583 Vbias.n572 1010.98
R4141 Vbias.n591 Vbias.n583 1010.98
R4142 Vbias.n592 Vbias.n591 1010.98
R4143 Vbias.n592 Vbias.n582 1010.98
R4144 Vbias.n584 Vbias.n573 1010.98
R4145 Vbias.n584 Vbias.n578 1010.98
R4146 Vbias.n593 Vbias.n578 1010.98
R4147 Vbias.n593 Vbias.n580 1010.98
R4148 Vbias.n541 Vbias.n530 1010.98
R4149 Vbias.n541 Vbias.n535 1010.98
R4150 Vbias.n550 Vbias.n535 1010.98
R4151 Vbias.n550 Vbias.n537 1010.98
R4152 Vbias.n540 Vbias.n529 1010.98
R4153 Vbias.n548 Vbias.n540 1010.98
R4154 Vbias.n549 Vbias.n548 1010.98
R4155 Vbias.n549 Vbias.n539 1010.98
R4156 Vbias.n526 Vbias.n513 1010.98
R4157 Vbias.n526 Vbias.n515 1010.98
R4158 Vbias.n525 Vbias.n524 1010.98
R4159 Vbias.n525 Vbias.n517 1010.98
R4160 Vbias.n494 Vbias.n483 1010.98
R4161 Vbias.n494 Vbias.n488 1010.98
R4162 Vbias.n503 Vbias.n488 1010.98
R4163 Vbias.n503 Vbias.n490 1010.98
R4164 Vbias.n493 Vbias.n482 1010.98
R4165 Vbias.n501 Vbias.n493 1010.98
R4166 Vbias.n502 Vbias.n501 1010.98
R4167 Vbias.n502 Vbias.n492 1010.98
R4168 Vbias.n469 Vbias.n458 1010.98
R4169 Vbias.n477 Vbias.n469 1010.98
R4170 Vbias.n478 Vbias.n477 1010.98
R4171 Vbias.n478 Vbias.n468 1010.98
R4172 Vbias.n470 Vbias.n459 1010.98
R4173 Vbias.n470 Vbias.n464 1010.98
R4174 Vbias.n479 Vbias.n464 1010.98
R4175 Vbias.n479 Vbias.n466 1010.98
R4176 Vbias.n435 Vbias.n424 1010.98
R4177 Vbias.n435 Vbias.n429 1010.98
R4178 Vbias.n444 Vbias.n429 1010.98
R4179 Vbias.n444 Vbias.n431 1010.98
R4180 Vbias.n434 Vbias.n423 1010.98
R4181 Vbias.n442 Vbias.n434 1010.98
R4182 Vbias.n443 Vbias.n442 1010.98
R4183 Vbias.n443 Vbias.n433 1010.98
R4184 Vbias.n420 Vbias.n407 1010.98
R4185 Vbias.n420 Vbias.n409 1010.98
R4186 Vbias.n419 Vbias.n418 1010.98
R4187 Vbias.n419 Vbias.n411 1010.98
R4188 Vbias.n388 Vbias.n377 1010.98
R4189 Vbias.n388 Vbias.n382 1010.98
R4190 Vbias.n397 Vbias.n382 1010.98
R4191 Vbias.n397 Vbias.n384 1010.98
R4192 Vbias.n387 Vbias.n376 1010.98
R4193 Vbias.n395 Vbias.n387 1010.98
R4194 Vbias.n396 Vbias.n395 1010.98
R4195 Vbias.n396 Vbias.n386 1010.98
R4196 Vbias.n363 Vbias.n175 1010.98
R4197 Vbias.n371 Vbias.n363 1010.98
R4198 Vbias.n372 Vbias.n371 1010.98
R4199 Vbias.n372 Vbias.n362 1010.98
R4200 Vbias.n364 Vbias.n176 1010.98
R4201 Vbias.n364 Vbias.n358 1010.98
R4202 Vbias.n373 Vbias.n358 1010.98
R4203 Vbias.n373 Vbias.n360 1010.98
R4204 Vbias.n315 Vbias.n192 1010.98
R4205 Vbias.n195 Vbias.n192 1010.98
R4206 Vbias.n195 Vbias.n185 1010.98
R4207 Vbias.n185 Vbias.n181 1010.98
R4208 Vbias.n317 Vbias.n316 1010.98
R4209 Vbias.n318 Vbias.n317 1010.98
R4210 Vbias.n318 Vbias.n184 1010.98
R4211 Vbias.n184 Vbias.n183 1010.98
R4212 Vbias.n207 Vbias.n204 1010.98
R4213 Vbias.n204 Vbias.n200 1010.98
R4214 Vbias.n301 Vbias.n203 1010.98
R4215 Vbias.n203 Vbias.n202 1010.98
R4216 Vbias.n276 Vbias.n225 1010.98
R4217 Vbias.n228 Vbias.n225 1010.98
R4218 Vbias.n228 Vbias.n218 1010.98
R4219 Vbias.n218 Vbias.n214 1010.98
R4220 Vbias.n278 Vbias.n277 1010.98
R4221 Vbias.n279 Vbias.n278 1010.98
R4222 Vbias.n279 Vbias.n217 1010.98
R4223 Vbias.n217 Vbias.n216 1010.98
R4224 Vbias.n261 Vbias.n260 1010.98
R4225 Vbias.n262 Vbias.n261 1010.98
R4226 Vbias.n262 Vbias.n236 1010.98
R4227 Vbias.n236 Vbias.n235 1010.98
R4228 Vbias.n259 Vbias.n243 1010.98
R4229 Vbias.n245 Vbias.n243 1010.98
R4230 Vbias.n245 Vbias.n237 1010.98
R4231 Vbias.n237 Vbias.n233 1010.98
R4232 Vbias.n4604 Vbias.n4602 1010.98
R4233 Vbias.n4642 Vbias.n4604 1010.98
R4234 Vbias.n4642 Vbias.n4605 1010.98
R4235 Vbias.n4605 Vbias.n2435 1010.98
R4236 Vbias.n4634 Vbias.n4609 1010.98
R4237 Vbias.n4641 Vbias.n4609 1010.98
R4238 Vbias.n4641 Vbias.n4610 1010.98
R4239 Vbias.n4610 Vbias.n2434 1010.98
R4240 Vbias.n4614 Vbias.n4595 1010.98
R4241 Vbias.n4614 Vbias.n4597 1010.98
R4242 Vbias.n4623 Vbias.n4597 1010.98
R4243 Vbias.n4623 Vbias.n4599 1010.98
R4244 Vbias.n4622 Vbias.n4621 1010.98
R4245 Vbias.n4626 Vbias.n4622 1010.98
R4246 Vbias.n4626 Vbias.n4612 1010.98
R4247 Vbias.n4630 Vbias.n4612 1010.98
R4248 Vbias.n4584 Vbias.n4575 1010.98
R4249 Vbias.n4584 Vbias.n4580 1010.98
R4250 Vbias.n4583 Vbias.n4574 1010.98
R4251 Vbias.n4583 Vbias.n4582 1010.98
R4252 Vbias.n4475 Vbias.n4471 1010.98
R4253 Vbias.n4504 Vbias.n4471 1010.98
R4254 Vbias.n4504 Vbias.n4472 1010.98
R4255 Vbias.n4500 Vbias.n4472 1010.98
R4256 Vbias.n4466 Vbias.n4463 1010.98
R4257 Vbias.n4505 Vbias.n4466 1010.98
R4258 Vbias.n4505 Vbias.n4467 1010.98
R4259 Vbias.n4499 Vbias.n4467 1010.98
R4260 Vbias.n4453 Vbias.n4449 1010.98
R4261 Vbias.n4518 Vbias.n4449 1010.98
R4262 Vbias.n4518 Vbias.n4450 1010.98
R4263 Vbias.n4514 Vbias.n4450 1010.98
R4264 Vbias.n4444 Vbias.n4441 1010.98
R4265 Vbias.n4519 Vbias.n4444 1010.98
R4266 Vbias.n4519 Vbias.n4445 1010.98
R4267 Vbias.n4513 Vbias.n4445 1010.98
R4268 Vbias.n4431 Vbias.n4427 1010.98
R4269 Vbias.n4528 Vbias.n4431 1010.98
R4270 Vbias.n4436 Vbias.n4426 1010.98
R4271 Vbias.n4527 Vbias.n4436 1010.98
R4272 Vbias.n4412 Vbias.n4408 1010.98
R4273 Vbias.n4544 Vbias.n4412 1010.98
R4274 Vbias.n4544 Vbias.n4413 1010.98
R4275 Vbias.n4537 Vbias.n4413 1010.98
R4276 Vbias.n4417 Vbias.n4407 1010.98
R4277 Vbias.n4543 Vbias.n4417 1010.98
R4278 Vbias.n4543 Vbias.n4418 1010.98
R4279 Vbias.n4538 Vbias.n4418 1010.98
R4280 Vbias.n5103 Vbias.n2378 1010.98
R4281 Vbias.n5112 Vbias.n2378 1010.98
R4282 Vbias.n5112 Vbias.n2379 1010.98
R4283 Vbias.n2379 Vbias.n2373 1010.98
R4284 Vbias.n5104 Vbias.n2382 1010.98
R4285 Vbias.n5111 Vbias.n2382 1010.98
R4286 Vbias.n5111 Vbias.n2383 1010.98
R4287 Vbias.n2383 Vbias.n2372 1010.98
R4288 Vbias.n5083 Vbias.n2394 1010.98
R4289 Vbias.n5092 Vbias.n2394 1010.98
R4290 Vbias.n5092 Vbias.n2395 1010.98
R4291 Vbias.n2395 Vbias.n2389 1010.98
R4292 Vbias.n5084 Vbias.n2398 1010.98
R4293 Vbias.n5091 Vbias.n2398 1010.98
R4294 Vbias.n5091 Vbias.n2399 1010.98
R4295 Vbias.n2399 Vbias.n2388 1010.98
R4296 Vbias.n2416 Vbias.n2413 1010.98
R4297 Vbias.n2413 Vbias.n2409 1010.98
R4298 Vbias.n5060 Vbias.n2412 1010.98
R4299 Vbias.n2412 Vbias.n2411 1010.98
R4300 Vbias.n2276 Vbias.n2266 1010.98
R4301 Vbias.n2276 Vbias.n2270 1010.98
R4302 Vbias.n2285 Vbias.n2270 1010.98
R4303 Vbias.n2285 Vbias.n2272 1010.98
R4304 Vbias.n2275 Vbias.n2265 1010.98
R4305 Vbias.n2283 Vbias.n2275 1010.98
R4306 Vbias.n2284 Vbias.n2283 1010.98
R4307 Vbias.n2284 Vbias.n2274 1010.98
R4308 Vbias.n5153 Vbias.n2247 1010.98
R4309 Vbias.n2250 Vbias.n2247 1010.98
R4310 Vbias.n2258 Vbias.n2250 1010.98
R4311 Vbias.n2258 Vbias.n2254 1010.98
R4312 Vbias.n5152 Vbias.n2246 1010.98
R4313 Vbias.n2259 Vbias.n2246 1010.98
R4314 Vbias.n2259 Vbias.n2257 1010.98
R4315 Vbias.n2257 Vbias.n2256 1010.98
R4316 Vbias.n5146 Vbias.n2359 1010.98
R4317 Vbias.n5146 Vbias.n2361 1010.98
R4318 Vbias.n5145 Vbias.n5144 1010.98
R4319 Vbias.n5145 Vbias.n2363 1010.98
R4320 Vbias.n5127 Vbias.n2351 1010.98
R4321 Vbias.n5127 Vbias.n2353 1010.98
R4322 Vbias.n5130 Vbias.n2353 1010.98
R4323 Vbias.n5130 Vbias.n2355 1010.98
R4324 Vbias.n5126 Vbias.n2366 1010.98
R4325 Vbias.n5133 Vbias.n2366 1010.98
R4326 Vbias.n5133 Vbias.n2364 1010.98
R4327 Vbias.n5137 Vbias.n2364 1010.98
R4328 Vbias.n5900 Vbias.n1646 1010.98
R4329 Vbias.n5909 Vbias.n1646 1010.98
R4330 Vbias.n5909 Vbias.n1647 1010.98
R4331 Vbias.n1647 Vbias.n1641 1010.98
R4332 Vbias.n5901 Vbias.n1650 1010.98
R4333 Vbias.n5908 Vbias.n1650 1010.98
R4334 Vbias.n5908 Vbias.n1651 1010.98
R4335 Vbias.n1651 Vbias.n1640 1010.98
R4336 Vbias.n5880 Vbias.n1662 1010.98
R4337 Vbias.n5889 Vbias.n1662 1010.98
R4338 Vbias.n5889 Vbias.n1663 1010.98
R4339 Vbias.n1663 Vbias.n1657 1010.98
R4340 Vbias.n5881 Vbias.n1666 1010.98
R4341 Vbias.n5888 Vbias.n1666 1010.98
R4342 Vbias.n5888 Vbias.n1667 1010.98
R4343 Vbias.n1667 Vbias.n1656 1010.98
R4344 Vbias.n5446 Vbias.n5437 1010.98
R4345 Vbias.n5446 Vbias.n5442 1010.98
R4346 Vbias.n5445 Vbias.n5436 1010.98
R4347 Vbias.n5445 Vbias.n5444 1010.98
R4348 Vbias.n5424 Vbias.n2290 1010.98
R4349 Vbias.n5424 Vbias.n5418 1010.98
R4350 Vbias.n5433 Vbias.n5418 1010.98
R4351 Vbias.n5433 Vbias.n5420 1010.98
R4352 Vbias.n5423 Vbias.n2289 1010.98
R4353 Vbias.n5431 Vbias.n5423 1010.98
R4354 Vbias.n5432 Vbias.n5431 1010.98
R4355 Vbias.n5432 Vbias.n5422 1010.98
R4356 Vbias.n5938 Vbias.n1623 1010.98
R4357 Vbias.n5938 Vbias.n1625 1010.98
R4358 Vbias.n5937 Vbias.n1627 1010.98
R4359 Vbias.n5941 Vbias.n1627 1010.98
R4360 Vbias.n1631 Vbias.n1614 1010.98
R4361 Vbias.n1631 Vbias.n1616 1010.98
R4362 Vbias.n5927 Vbias.n1616 1010.98
R4363 Vbias.n5927 Vbias.n1618 1010.98
R4364 Vbias.n5921 Vbias.n1633 1010.98
R4365 Vbias.n5926 Vbias.n1633 1010.98
R4366 Vbias.n5926 Vbias.n1628 1010.98
R4367 Vbias.n5930 Vbias.n1628 1010.98
R4368 Vbias.n1809 Vbias.n1764 1010.98
R4369 Vbias.n1813 Vbias.n1764 1010.98
R4370 Vbias.n1813 Vbias.n1761 1010.98
R4371 Vbias.n1817 Vbias.n1761 1010.98
R4372 Vbias.n1811 Vbias.n1810 1010.98
R4373 Vbias.n1812 Vbias.n1811 1010.98
R4374 Vbias.n1812 Vbias.n1757 1010.98
R4375 Vbias.n1818 Vbias.n1757 1010.98
R4376 Vbias.n1862 Vbias.n1855 1010.98
R4377 Vbias.n1877 Vbias.n1855 1010.98
R4378 Vbias.n1877 Vbias.n1856 1010.98
R4379 Vbias.n1873 Vbias.n1856 1010.98
R4380 Vbias.n1861 Vbias.n1851 1010.98
R4381 Vbias.n1878 Vbias.n1851 1010.98
R4382 Vbias.n1878 Vbias.n1852 1010.98
R4383 Vbias.n1872 Vbias.n1852 1010.98
R4384 Vbias.n1930 Vbias.n1923 1010.98
R4385 Vbias.n1945 Vbias.n1923 1010.98
R4386 Vbias.n1945 Vbias.n1924 1010.98
R4387 Vbias.n1939 Vbias.n1924 1010.98
R4388 Vbias.n1929 Vbias.n1919 1010.98
R4389 Vbias.n1946 Vbias.n1919 1010.98
R4390 Vbias.n1946 Vbias.n1920 1010.98
R4391 Vbias.n1938 Vbias.n1920 1010.98
R4392 Vbias.n2004 Vbias.n2003 1010.98
R4393 Vbias.n2005 Vbias.n2004 1010.98
R4394 Vbias.n2005 Vbias.n1988 1010.98
R4395 Vbias.n2011 Vbias.n1988 1010.98
R4396 Vbias.n2002 Vbias.n1995 1010.98
R4397 Vbias.n1997 Vbias.n1995 1010.98
R4398 Vbias.n1997 Vbias.n1989 1010.98
R4399 Vbias.n1989 Vbias.n1986 1010.98
R4400 Vbias.n6104 Vbias.n1517 1010.98
R4401 Vbias.n6119 Vbias.n1517 1010.98
R4402 Vbias.n6119 Vbias.n1518 1010.98
R4403 Vbias.n6113 Vbias.n1518 1010.98
R4404 Vbias.n6103 Vbias.n1513 1010.98
R4405 Vbias.n6120 Vbias.n1513 1010.98
R4406 Vbias.n6120 Vbias.n1514 1010.98
R4407 Vbias.n6112 Vbias.n1514 1010.98
R4408 Vbias.n1964 Vbias.n1957 1010.98
R4409 Vbias.n1979 Vbias.n1957 1010.98
R4410 Vbias.n1979 Vbias.n1958 1010.98
R4411 Vbias.n1973 Vbias.n1958 1010.98
R4412 Vbias.n1963 Vbias.n1953 1010.98
R4413 Vbias.n1980 Vbias.n1953 1010.98
R4414 Vbias.n1980 Vbias.n1954 1010.98
R4415 Vbias.n1972 Vbias.n1954 1010.98
R4416 Vbias.n1911 Vbias.n1888 1010.98
R4417 Vbias.n1907 Vbias.n1888 1010.98
R4418 Vbias.n1907 Vbias.n1892 1010.98
R4419 Vbias.n1903 Vbias.n1892 1010.98
R4420 Vbias.n1912 Vbias.n1886 1010.98
R4421 Vbias.n1906 Vbias.n1886 1010.98
R4422 Vbias.n1906 Vbias.n1905 1010.98
R4423 Vbias.n1905 Vbias.n1904 1010.98
R4424 Vbias.n1775 Vbias.n1547 1010.98
R4425 Vbias.n1775 Vbias.n1549 1010.98
R4426 Vbias.n1780 Vbias.n1549 1010.98
R4427 Vbias.n1780 Vbias.n1551 1010.98
R4428 Vbias.n1787 Vbias.n1778 1010.98
R4429 Vbias.n1783 Vbias.n1778 1010.98
R4430 Vbias.n1783 Vbias.n1782 1010.98
R4431 Vbias.n1782 Vbias.n1553 1010.98
R4432 Vbias.n1769 Vbias.n1539 1010.98
R4433 Vbias.n1769 Vbias.n1541 1010.98
R4434 Vbias.n1773 Vbias.n1541 1010.98
R4435 Vbias.n1773 Vbias.n1543 1010.98
R4436 Vbias.n1799 Vbias.n1771 1010.98
R4437 Vbias.n1795 Vbias.n1771 1010.98
R4438 Vbias.n1795 Vbias.n1794 1010.98
R4439 Vbias.n1794 Vbias.n1793 1010.98
R4440 Vbias.n1432 Vbias.n1430 1010.98
R4441 Vbias.n6780 Vbias.n1432 1010.98
R4442 Vbias.n6780 Vbias.n1433 1010.98
R4443 Vbias.n1433 Vbias.n1342 1010.98
R4444 Vbias.n6772 Vbias.n1437 1010.98
R4445 Vbias.n6779 Vbias.n1437 1010.98
R4446 Vbias.n6779 Vbias.n1438 1010.98
R4447 Vbias.n1438 Vbias.n1341 1010.98
R4448 Vbias.n6758 Vbias.n1423 1010.98
R4449 Vbias.n6758 Vbias.n1425 1010.98
R4450 Vbias.n6761 Vbias.n1425 1010.98
R4451 Vbias.n6761 Vbias.n1427 1010.98
R4452 Vbias.n6757 Vbias.n1442 1010.98
R4453 Vbias.n6764 Vbias.n1442 1010.98
R4454 Vbias.n6764 Vbias.n1440 1010.98
R4455 Vbias.n6768 Vbias.n1440 1010.98
R4456 Vbias.n6052 Vbias.n1411 1010.98
R4457 Vbias.n6052 Vbias.n1413 1010.98
R4458 Vbias.n6058 Vbias.n6055 1010.98
R4459 Vbias.n6055 Vbias.n1415 1010.98
R4460 Vbias.n6049 Vbias.n1403 1010.98
R4461 Vbias.n6049 Vbias.n1405 1010.98
R4462 Vbias.n6065 Vbias.n1405 1010.98
R4463 Vbias.n6065 Vbias.n1407 1010.98
R4464 Vbias.n6072 Vbias.n6046 1010.98
R4465 Vbias.n6068 Vbias.n6046 1010.98
R4466 Vbias.n6068 Vbias.n6048 1010.98
R4467 Vbias.n6064 Vbias.n6048 1010.98
R4468 Vbias.n7081 Vbias.n1286 1010.98
R4469 Vbias.n1289 Vbias.n1286 1010.98
R4470 Vbias.n1289 Vbias.n1279 1010.98
R4471 Vbias.n1279 Vbias.n1276 1010.98
R4472 Vbias.n7083 Vbias.n7082 1010.98
R4473 Vbias.n7084 Vbias.n7083 1010.98
R4474 Vbias.n7084 Vbias.n1278 1010.98
R4475 Vbias.n7090 Vbias.n1278 1010.98
R4476 Vbias.n7064 Vbias.n1306 1010.98
R4477 Vbias.n1309 Vbias.n1306 1010.98
R4478 Vbias.n1309 Vbias.n1298 1010.98
R4479 Vbias.n1298 Vbias.n1294 1010.98
R4480 Vbias.n7066 Vbias.n7065 1010.98
R4481 Vbias.n7067 Vbias.n7066 1010.98
R4482 Vbias.n7067 Vbias.n1297 1010.98
R4483 Vbias.n1297 Vbias.n1296 1010.98
R4484 Vbias.n7045 Vbias.n1322 1010.98
R4485 Vbias.n1322 Vbias.n1317 1010.98
R4486 Vbias.n7044 Vbias.n7039 1010.98
R4487 Vbias.n7039 Vbias.n1316 1010.98
R4488 Vbias.n7019 Vbias.n1329 1010.98
R4489 Vbias.n7028 Vbias.n1329 1010.98
R4490 Vbias.n7028 Vbias.n1330 1010.98
R4491 Vbias.n1330 Vbias.n1324 1010.98
R4492 Vbias.n7020 Vbias.n1333 1010.98
R4493 Vbias.n7027 Vbias.n1333 1010.98
R4494 Vbias.n7027 Vbias.n1334 1010.98
R4495 Vbias.n1334 Vbias.n1323 1010.98
R4496 Vbias.n7187 Vbias.n1099 1010.98
R4497 Vbias.n1102 Vbias.n1099 1010.98
R4498 Vbias.n1102 Vbias.n1092 1010.98
R4499 Vbias.n1092 Vbias.n1089 1010.98
R4500 Vbias.n7189 Vbias.n7188 1010.98
R4501 Vbias.n7190 Vbias.n7189 1010.98
R4502 Vbias.n7190 Vbias.n1091 1010.98
R4503 Vbias.n7196 Vbias.n1091 1010.98
R4504 Vbias.n7170 Vbias.n1118 1010.98
R4505 Vbias.n1121 Vbias.n1118 1010.98
R4506 Vbias.n1121 Vbias.n1111 1010.98
R4507 Vbias.n1111 Vbias.n1107 1010.98
R4508 Vbias.n7172 Vbias.n7171 1010.98
R4509 Vbias.n7173 Vbias.n7172 1010.98
R4510 Vbias.n7173 Vbias.n1110 1010.98
R4511 Vbias.n1110 Vbias.n1109 1010.98
R4512 Vbias.n7151 Vbias.n1134 1010.98
R4513 Vbias.n1134 Vbias.n1129 1010.98
R4514 Vbias.n7150 Vbias.n7145 1010.98
R4515 Vbias.n7145 Vbias.n1128 1010.98
R4516 Vbias.n7125 Vbias.n1141 1010.98
R4517 Vbias.n7134 Vbias.n1141 1010.98
R4518 Vbias.n7134 Vbias.n1142 1010.98
R4519 Vbias.n1142 Vbias.n1136 1010.98
R4520 Vbias.n7126 Vbias.n1145 1010.98
R4521 Vbias.n7133 Vbias.n1145 1010.98
R4522 Vbias.n7133 Vbias.n1146 1010.98
R4523 Vbias.n1146 Vbias.n1135 1010.98
R4524 Vbias.n1217 Vbias.n1215 1010.98
R4525 Vbias.n1217 Vbias.n1083 1010.98
R4526 Vbias.n1083 Vbias.n1081 1010.98
R4527 Vbias.n1081 Vbias.n1076 1010.98
R4528 Vbias.n1214 Vbias.n1084 1010.98
R4529 Vbias.n7209 Vbias.n1084 1010.98
R4530 Vbias.n7209 Vbias.n1080 1010.98
R4531 Vbias.n1080 Vbias.n1075 1010.98
R4532 Vbias.n1206 Vbias.n1202 1010.98
R4533 Vbias.n1208 Vbias.n1202 1010.98
R4534 Vbias.n1226 Vbias.n1208 1010.98
R4535 Vbias.n1233 Vbias.n1226 1010.98
R4536 Vbias.n1201 Vbias.n1198 1010.98
R4537 Vbias.n1236 Vbias.n1201 1010.98
R4538 Vbias.n1236 Vbias.n1235 1010.98
R4539 Vbias.n1235 Vbias.n1234 1010.98
R4540 Vbias.n1189 Vbias.n1184 1010.98
R4541 Vbias.n1191 Vbias.n1189 1010.98
R4542 Vbias.n1188 Vbias.n1183 1010.98
R4543 Vbias.n1247 Vbias.n1188 1010.98
R4544 Vbias.n1177 Vbias.n1174 1010.98
R4545 Vbias.n1179 Vbias.n1174 1010.98
R4546 Vbias.n1257 Vbias.n1179 1010.98
R4547 Vbias.n1264 Vbias.n1257 1010.98
R4548 Vbias.n1173 Vbias.n1170 1010.98
R4549 Vbias.n1267 Vbias.n1173 1010.98
R4550 Vbias.n1267 Vbias.n1266 1010.98
R4551 Vbias.n1266 Vbias.n1265 1010.98
R4552 Vbias.n6950 Vbias.n6948 1010.98
R4553 Vbias.n6950 Vbias.n1164 1010.98
R4554 Vbias.n1164 Vbias.n1162 1010.98
R4555 Vbias.n1162 Vbias.n1157 1010.98
R4556 Vbias.n6947 Vbias.n1165 1010.98
R4557 Vbias.n7105 Vbias.n1165 1010.98
R4558 Vbias.n7105 Vbias.n1161 1010.98
R4559 Vbias.n1161 Vbias.n1156 1010.98
R4560 Vbias.n6939 Vbias.n6935 1010.98
R4561 Vbias.n6941 Vbias.n6935 1010.98
R4562 Vbias.n6959 Vbias.n6941 1010.98
R4563 Vbias.n6966 Vbias.n6959 1010.98
R4564 Vbias.n6934 Vbias.n6931 1010.98
R4565 Vbias.n6969 Vbias.n6934 1010.98
R4566 Vbias.n6969 Vbias.n6968 1010.98
R4567 Vbias.n6968 Vbias.n6967 1010.98
R4568 Vbias.n6922 Vbias.n6917 1010.98
R4569 Vbias.n6924 Vbias.n6922 1010.98
R4570 Vbias.n6921 Vbias.n6916 1010.98
R4571 Vbias.n6980 Vbias.n6921 1010.98
R4572 Vbias.n6910 Vbias.n6907 1010.98
R4573 Vbias.n6912 Vbias.n6907 1010.98
R4574 Vbias.n6990 Vbias.n6912 1010.98
R4575 Vbias.n6997 Vbias.n6990 1010.98
R4576 Vbias.n6906 Vbias.n6903 1010.98
R4577 Vbias.n7000 Vbias.n6906 1010.98
R4578 Vbias.n7000 Vbias.n6999 1010.98
R4579 Vbias.n6999 Vbias.n6998 1010.98
R4580 Vbias.n6876 Vbias.n6871 1010.98
R4581 Vbias.n6871 Vbias.n1358 1010.98
R4582 Vbias.n1358 Vbias.n1356 1010.98
R4583 Vbias.n1356 Vbias.n1351 1010.98
R4584 Vbias.n6877 Vbias.n1359 1010.98
R4585 Vbias.n6884 Vbias.n1359 1010.98
R4586 Vbias.n6884 Vbias.n1355 1010.98
R4587 Vbias.n1355 Vbias.n1350 1010.98
R4588 Vbias.n6853 Vbias.n6848 1010.98
R4589 Vbias.n6848 Vbias.n1371 1010.98
R4590 Vbias.n1371 Vbias.n1369 1010.98
R4591 Vbias.n1369 Vbias.n1364 1010.98
R4592 Vbias.n6854 Vbias.n1372 1010.98
R4593 Vbias.n6861 Vbias.n1372 1010.98
R4594 Vbias.n6861 Vbias.n1368 1010.98
R4595 Vbias.n1368 Vbias.n1363 1010.98
R4596 Vbias.n1384 Vbias.n1382 1010.98
R4597 Vbias.n1382 Vbias.n1377 1010.98
R4598 Vbias.n6838 Vbias.n1381 1010.98
R4599 Vbias.n1381 Vbias.n1376 1010.98
R4600 Vbias.n1555 Vbias.n1396 1010.98
R4601 Vbias.n6823 Vbias.n1396 1010.98
R4602 Vbias.n6823 Vbias.n1394 1010.98
R4603 Vbias.n6829 Vbias.n1394 1010.98
R4604 Vbias.n1400 Vbias.n1398 1010.98
R4605 Vbias.n6822 Vbias.n1398 1010.98
R4606 Vbias.n6822 Vbias.n1390 1010.98
R4607 Vbias.n6830 Vbias.n1390 1010.98
R4608 Vbias.n6018 Vbias.n6013 1010.98
R4609 Vbias.n6013 Vbias.n1569 1010.98
R4610 Vbias.n1569 Vbias.n1567 1010.98
R4611 Vbias.n1567 Vbias.n1562 1010.98
R4612 Vbias.n6019 Vbias.n1570 1010.98
R4613 Vbias.n6029 Vbias.n1570 1010.98
R4614 Vbias.n6029 Vbias.n1566 1010.98
R4615 Vbias.n1566 Vbias.n1561 1010.98
R4616 Vbias.n5995 Vbias.n5990 1010.98
R4617 Vbias.n5990 Vbias.n1582 1010.98
R4618 Vbias.n1582 Vbias.n1580 1010.98
R4619 Vbias.n1580 Vbias.n1575 1010.98
R4620 Vbias.n5996 Vbias.n1583 1010.98
R4621 Vbias.n6003 Vbias.n1583 1010.98
R4622 Vbias.n6003 Vbias.n1579 1010.98
R4623 Vbias.n1579 Vbias.n1574 1010.98
R4624 Vbias.n1595 Vbias.n1593 1010.98
R4625 Vbias.n1593 Vbias.n1588 1010.98
R4626 Vbias.n5980 Vbias.n1592 1010.98
R4627 Vbias.n1592 Vbias.n1587 1010.98
R4628 Vbias.n1636 Vbias.n1607 1010.98
R4629 Vbias.n5965 Vbias.n1607 1010.98
R4630 Vbias.n5965 Vbias.n1605 1010.98
R4631 Vbias.n5971 Vbias.n1605 1010.98
R4632 Vbias.n1611 Vbias.n1609 1010.98
R4633 Vbias.n5964 Vbias.n1609 1010.98
R4634 Vbias.n5964 Vbias.n1601 1010.98
R4635 Vbias.n5972 Vbias.n1601 1010.98
R4636 Vbias.n5321 Vbias.n5317 1010.98
R4637 Vbias.n5359 Vbias.n5321 1010.98
R4638 Vbias.n5359 Vbias.n5322 1010.98
R4639 Vbias.n5352 Vbias.n5322 1010.98
R4640 Vbias.n5326 Vbias.n5316 1010.98
R4641 Vbias.n5358 Vbias.n5326 1010.98
R4642 Vbias.n5358 Vbias.n5327 1010.98
R4643 Vbias.n5353 Vbias.n5327 1010.98
R4644 Vbias.n5310 Vbias.n5306 1010.98
R4645 Vbias.n5312 Vbias.n5306 1010.98
R4646 Vbias.n5367 Vbias.n5312 1010.98
R4647 Vbias.n5374 Vbias.n5367 1010.98
R4648 Vbias.n5305 Vbias.n5302 1010.98
R4649 Vbias.n5377 Vbias.n5305 1010.98
R4650 Vbias.n5377 Vbias.n5376 1010.98
R4651 Vbias.n5376 Vbias.n5375 1010.98
R4652 Vbias.n5293 Vbias.n5288 1010.98
R4653 Vbias.n5295 Vbias.n5293 1010.98
R4654 Vbias.n5292 Vbias.n5287 1010.98
R4655 Vbias.n5388 Vbias.n5292 1010.98
R4656 Vbias.n5281 Vbias.n5277 1010.98
R4657 Vbias.n5283 Vbias.n5277 1010.98
R4658 Vbias.n5398 Vbias.n5283 1010.98
R4659 Vbias.n5405 Vbias.n5398 1010.98
R4660 Vbias.n5276 Vbias.n5273 1010.98
R4661 Vbias.n5408 Vbias.n5276 1010.98
R4662 Vbias.n5408 Vbias.n5407 1010.98
R4663 Vbias.n5407 Vbias.n5406 1010.98
R4664 Vbias.n5245 Vbias.n5240 1010.98
R4665 Vbias.n5240 Vbias.n2306 1010.98
R4666 Vbias.n2306 Vbias.n2304 1010.98
R4667 Vbias.n2304 Vbias.n2299 1010.98
R4668 Vbias.n5246 Vbias.n2307 1010.98
R4669 Vbias.n5253 Vbias.n2307 1010.98
R4670 Vbias.n5253 Vbias.n2303 1010.98
R4671 Vbias.n2303 Vbias.n2298 1010.98
R4672 Vbias.n5222 Vbias.n5217 1010.98
R4673 Vbias.n5217 Vbias.n2319 1010.98
R4674 Vbias.n2319 Vbias.n2317 1010.98
R4675 Vbias.n2317 Vbias.n2312 1010.98
R4676 Vbias.n5223 Vbias.n2320 1010.98
R4677 Vbias.n5230 Vbias.n2320 1010.98
R4678 Vbias.n5230 Vbias.n2316 1010.98
R4679 Vbias.n2316 Vbias.n2311 1010.98
R4680 Vbias.n2332 Vbias.n2330 1010.98
R4681 Vbias.n2330 Vbias.n2325 1010.98
R4682 Vbias.n5207 Vbias.n2329 1010.98
R4683 Vbias.n2329 Vbias.n2324 1010.98
R4684 Vbias.n2368 Vbias.n2344 1010.98
R4685 Vbias.n5192 Vbias.n2344 1010.98
R4686 Vbias.n5192 Vbias.n2342 1010.98
R4687 Vbias.n5198 Vbias.n2342 1010.98
R4688 Vbias.n2348 Vbias.n2346 1010.98
R4689 Vbias.n5191 Vbias.n2346 1010.98
R4690 Vbias.n5191 Vbias.n2338 1010.98
R4691 Vbias.n5199 Vbias.n2338 1010.98
R4692 Vbias.n2489 Vbias.n2485 1010.98
R4693 Vbias.n2527 Vbias.n2489 1010.98
R4694 Vbias.n2527 Vbias.n2490 1010.98
R4695 Vbias.n2520 Vbias.n2490 1010.98
R4696 Vbias.n2494 Vbias.n2484 1010.98
R4697 Vbias.n2526 Vbias.n2494 1010.98
R4698 Vbias.n2526 Vbias.n2495 1010.98
R4699 Vbias.n2521 Vbias.n2495 1010.98
R4700 Vbias.n2478 Vbias.n2474 1010.98
R4701 Vbias.n2480 Vbias.n2474 1010.98
R4702 Vbias.n2535 Vbias.n2480 1010.98
R4703 Vbias.n2542 Vbias.n2535 1010.98
R4704 Vbias.n2473 Vbias.n2470 1010.98
R4705 Vbias.n2545 Vbias.n2473 1010.98
R4706 Vbias.n2545 Vbias.n2544 1010.98
R4707 Vbias.n2544 Vbias.n2543 1010.98
R4708 Vbias.n2461 Vbias.n2456 1010.98
R4709 Vbias.n2463 Vbias.n2461 1010.98
R4710 Vbias.n2460 Vbias.n2455 1010.98
R4711 Vbias.n2556 Vbias.n2460 1010.98
R4712 Vbias.n2449 Vbias.n2445 1010.98
R4713 Vbias.n2451 Vbias.n2445 1010.98
R4714 Vbias.n2566 Vbias.n2451 1010.98
R4715 Vbias.n2573 Vbias.n2566 1010.98
R4716 Vbias.n2444 Vbias.n2441 1010.98
R4717 Vbias.n2576 Vbias.n2444 1010.98
R4718 Vbias.n2576 Vbias.n2575 1010.98
R4719 Vbias.n2575 Vbias.n2574 1010.98
R4720 Vbias.n5041 Vbias.n2427 1010.98
R4721 Vbias.n5048 Vbias.n2427 1010.98
R4722 Vbias.n5048 Vbias.n2428 1010.98
R4723 Vbias.n2428 Vbias.n2417 1010.98
R4724 Vbias.n5040 Vbias.n2423 1010.98
R4725 Vbias.n5049 Vbias.n2423 1010.98
R4726 Vbias.n5049 Vbias.n2424 1010.98
R4727 Vbias.n2424 Vbias.n2418 1010.98
R4728 Vbias.n3802 Vbias.n3792 1010.98
R4729 Vbias.n3847 Vbias.n3802 1010.98
R4730 Vbias.n3847 Vbias.n3803 1010.98
R4731 Vbias.n3841 Vbias.n3803 1010.98
R4732 Vbias.n3807 Vbias.n3791 1010.98
R4733 Vbias.n3846 Vbias.n3807 1010.98
R4734 Vbias.n3846 Vbias.n3808 1010.98
R4735 Vbias.n3842 Vbias.n3808 1010.98
R4736 Vbias.n3785 Vbias.n3779 1010.98
R4737 Vbias.n3857 Vbias.n3785 1010.98
R4738 Vbias.n3863 Vbias.n3784 1010.98
R4739 Vbias.n3880 Vbias.n3784 1010.98
R4740 Vbias.n3755 Vbias.n3745 1010.98
R4741 Vbias.n3923 Vbias.n3755 1010.98
R4742 Vbias.n3923 Vbias.n3756 1010.98
R4743 Vbias.n3917 Vbias.n3756 1010.98
R4744 Vbias.n3760 Vbias.n3744 1010.98
R4745 Vbias.n3922 Vbias.n3760 1010.98
R4746 Vbias.n3922 Vbias.n3761 1010.98
R4747 Vbias.n3918 Vbias.n3761 1010.98
R4748 Vbias.n3726 Vbias.n3716 1010.98
R4749 Vbias.n3961 Vbias.n3726 1010.98
R4750 Vbias.n3961 Vbias.n3727 1010.98
R4751 Vbias.n3955 Vbias.n3727 1010.98
R4752 Vbias.n3731 Vbias.n3715 1010.98
R4753 Vbias.n3960 Vbias.n3731 1010.98
R4754 Vbias.n3960 Vbias.n3732 1010.98
R4755 Vbias.n3956 Vbias.n3732 1010.98
R4756 Vbias.n3826 Vbias.n3825 1010.98
R4757 Vbias.n3825 Vbias.n3805 1010.98
R4758 Vbias.n3832 Vbias.n3805 1010.98
R4759 Vbias.n3832 Vbias.n3818 1010.98
R4760 Vbias.n3823 Vbias.n3795 1010.98
R4761 Vbias.n3823 Vbias.n3800 1010.98
R4762 Vbias.n3831 Vbias.n3800 1010.98
R4763 Vbias.n3831 Vbias.n3817 1010.98
R4764 Vbias.n3870 Vbias.n3869 1010.98
R4765 Vbias.n3869 Vbias.n3789 1010.98
R4766 Vbias.n3787 Vbias.n3780 1010.98
R4767 Vbias.n3788 Vbias.n3787 1010.98
R4768 Vbias.n3902 Vbias.n3901 1010.98
R4769 Vbias.n3901 Vbias.n3758 1010.98
R4770 Vbias.n3908 Vbias.n3758 1010.98
R4771 Vbias.n3908 Vbias.n3771 1010.98
R4772 Vbias.n3899 Vbias.n3748 1010.98
R4773 Vbias.n3899 Vbias.n3753 1010.98
R4774 Vbias.n3907 Vbias.n3753 1010.98
R4775 Vbias.n3907 Vbias.n3770 1010.98
R4776 Vbias.n3940 Vbias.n3939 1010.98
R4777 Vbias.n3939 Vbias.n3729 1010.98
R4778 Vbias.n3946 Vbias.n3729 1010.98
R4779 Vbias.n3946 Vbias.n3742 1010.98
R4780 Vbias.n3937 Vbias.n3719 1010.98
R4781 Vbias.n3937 Vbias.n3724 1010.98
R4782 Vbias.n3945 Vbias.n3724 1010.98
R4783 Vbias.n3945 Vbias.n3741 1010.98
R4784 Vbias.n3264 Vbias.n3254 1010.98
R4785 Vbias.n3309 Vbias.n3264 1010.98
R4786 Vbias.n3309 Vbias.n3265 1010.98
R4787 Vbias.n3303 Vbias.n3265 1010.98
R4788 Vbias.n3269 Vbias.n3253 1010.98
R4789 Vbias.n3308 Vbias.n3269 1010.98
R4790 Vbias.n3308 Vbias.n3270 1010.98
R4791 Vbias.n3304 Vbias.n3270 1010.98
R4792 Vbias.n3247 Vbias.n3241 1010.98
R4793 Vbias.n3319 Vbias.n3247 1010.98
R4794 Vbias.n3325 Vbias.n3246 1010.98
R4795 Vbias.n3342 Vbias.n3246 1010.98
R4796 Vbias.n3217 Vbias.n3207 1010.98
R4797 Vbias.n3385 Vbias.n3217 1010.98
R4798 Vbias.n3385 Vbias.n3218 1010.98
R4799 Vbias.n3379 Vbias.n3218 1010.98
R4800 Vbias.n3222 Vbias.n3206 1010.98
R4801 Vbias.n3384 Vbias.n3222 1010.98
R4802 Vbias.n3384 Vbias.n3223 1010.98
R4803 Vbias.n3380 Vbias.n3223 1010.98
R4804 Vbias.n3188 Vbias.n3178 1010.98
R4805 Vbias.n3423 Vbias.n3188 1010.98
R4806 Vbias.n3423 Vbias.n3189 1010.98
R4807 Vbias.n3417 Vbias.n3189 1010.98
R4808 Vbias.n3193 Vbias.n3177 1010.98
R4809 Vbias.n3422 Vbias.n3193 1010.98
R4810 Vbias.n3422 Vbias.n3194 1010.98
R4811 Vbias.n3418 Vbias.n3194 1010.98
R4812 Vbias.n3288 Vbias.n3287 1010.98
R4813 Vbias.n3287 Vbias.n3267 1010.98
R4814 Vbias.n3294 Vbias.n3267 1010.98
R4815 Vbias.n3294 Vbias.n3280 1010.98
R4816 Vbias.n3285 Vbias.n3257 1010.98
R4817 Vbias.n3285 Vbias.n3262 1010.98
R4818 Vbias.n3293 Vbias.n3262 1010.98
R4819 Vbias.n3293 Vbias.n3279 1010.98
R4820 Vbias.n3332 Vbias.n3331 1010.98
R4821 Vbias.n3331 Vbias.n3251 1010.98
R4822 Vbias.n3249 Vbias.n3242 1010.98
R4823 Vbias.n3250 Vbias.n3249 1010.98
R4824 Vbias.n3364 Vbias.n3363 1010.98
R4825 Vbias.n3363 Vbias.n3220 1010.98
R4826 Vbias.n3370 Vbias.n3220 1010.98
R4827 Vbias.n3370 Vbias.n3233 1010.98
R4828 Vbias.n3361 Vbias.n3210 1010.98
R4829 Vbias.n3361 Vbias.n3215 1010.98
R4830 Vbias.n3369 Vbias.n3215 1010.98
R4831 Vbias.n3369 Vbias.n3232 1010.98
R4832 Vbias.n3402 Vbias.n3401 1010.98
R4833 Vbias.n3401 Vbias.n3191 1010.98
R4834 Vbias.n3408 Vbias.n3191 1010.98
R4835 Vbias.n3408 Vbias.n3204 1010.98
R4836 Vbias.n3399 Vbias.n3181 1010.98
R4837 Vbias.n3399 Vbias.n3186 1010.98
R4838 Vbias.n3407 Vbias.n3186 1010.98
R4839 Vbias.n3407 Vbias.n3203 1010.98
R4840 Vbias.n3533 Vbias.n3523 1010.98
R4841 Vbias.n3578 Vbias.n3533 1010.98
R4842 Vbias.n3578 Vbias.n3534 1010.98
R4843 Vbias.n3572 Vbias.n3534 1010.98
R4844 Vbias.n3538 Vbias.n3522 1010.98
R4845 Vbias.n3577 Vbias.n3538 1010.98
R4846 Vbias.n3577 Vbias.n3539 1010.98
R4847 Vbias.n3573 Vbias.n3539 1010.98
R4848 Vbias.n3516 Vbias.n3510 1010.98
R4849 Vbias.n3588 Vbias.n3516 1010.98
R4850 Vbias.n3594 Vbias.n3515 1010.98
R4851 Vbias.n3611 Vbias.n3515 1010.98
R4852 Vbias.n3486 Vbias.n3476 1010.98
R4853 Vbias.n3654 Vbias.n3486 1010.98
R4854 Vbias.n3654 Vbias.n3487 1010.98
R4855 Vbias.n3648 Vbias.n3487 1010.98
R4856 Vbias.n3491 Vbias.n3475 1010.98
R4857 Vbias.n3653 Vbias.n3491 1010.98
R4858 Vbias.n3653 Vbias.n3492 1010.98
R4859 Vbias.n3649 Vbias.n3492 1010.98
R4860 Vbias.n3457 Vbias.n3447 1010.98
R4861 Vbias.n3692 Vbias.n3457 1010.98
R4862 Vbias.n3692 Vbias.n3458 1010.98
R4863 Vbias.n3686 Vbias.n3458 1010.98
R4864 Vbias.n3462 Vbias.n3446 1010.98
R4865 Vbias.n3691 Vbias.n3462 1010.98
R4866 Vbias.n3691 Vbias.n3463 1010.98
R4867 Vbias.n3687 Vbias.n3463 1010.98
R4868 Vbias.n3557 Vbias.n3556 1010.98
R4869 Vbias.n3556 Vbias.n3536 1010.98
R4870 Vbias.n3563 Vbias.n3536 1010.98
R4871 Vbias.n3563 Vbias.n3549 1010.98
R4872 Vbias.n3554 Vbias.n3526 1010.98
R4873 Vbias.n3554 Vbias.n3531 1010.98
R4874 Vbias.n3562 Vbias.n3531 1010.98
R4875 Vbias.n3562 Vbias.n3548 1010.98
R4876 Vbias.n3601 Vbias.n3600 1010.98
R4877 Vbias.n3600 Vbias.n3520 1010.98
R4878 Vbias.n3518 Vbias.n3511 1010.98
R4879 Vbias.n3519 Vbias.n3518 1010.98
R4880 Vbias.n3633 Vbias.n3632 1010.98
R4881 Vbias.n3632 Vbias.n3489 1010.98
R4882 Vbias.n3639 Vbias.n3489 1010.98
R4883 Vbias.n3639 Vbias.n3502 1010.98
R4884 Vbias.n3630 Vbias.n3479 1010.98
R4885 Vbias.n3630 Vbias.n3484 1010.98
R4886 Vbias.n3638 Vbias.n3484 1010.98
R4887 Vbias.n3638 Vbias.n3501 1010.98
R4888 Vbias.n3671 Vbias.n3670 1010.98
R4889 Vbias.n3670 Vbias.n3460 1010.98
R4890 Vbias.n3677 Vbias.n3460 1010.98
R4891 Vbias.n3677 Vbias.n3473 1010.98
R4892 Vbias.n3668 Vbias.n3450 1010.98
R4893 Vbias.n3668 Vbias.n3455 1010.98
R4894 Vbias.n3676 Vbias.n3455 1010.98
R4895 Vbias.n3676 Vbias.n3472 1010.98
R4896 Vbias.n4056 Vbias.n4050 1010.98
R4897 Vbias.n4193 Vbias.n4056 1010.98
R4898 Vbias.n4193 Vbias.n4057 1010.98
R4899 Vbias.n4187 Vbias.n4057 1010.98
R4900 Vbias.n4062 Vbias.n4049 1010.98
R4901 Vbias.n4192 Vbias.n4062 1010.98
R4902 Vbias.n4192 Vbias.n4063 1010.98
R4903 Vbias.n4188 Vbias.n4063 1010.98
R4904 Vbias.n4043 Vbias.n4039 1010.98
R4905 Vbias.n4202 Vbias.n4043 1010.98
R4906 Vbias.n4153 Vbias.n4042 1010.98
R4907 Vbias.n4206 Vbias.n4042 1010.98
R4908 Vbias.n4014 Vbias.n4008 1010.98
R4909 Vbias.n4227 Vbias.n4014 1010.98
R4910 Vbias.n4227 Vbias.n4015 1010.98
R4911 Vbias.n4221 Vbias.n4015 1010.98
R4912 Vbias.n4020 Vbias.n4007 1010.98
R4913 Vbias.n4226 Vbias.n4020 1010.98
R4914 Vbias.n4226 Vbias.n4021 1010.98
R4915 Vbias.n4222 Vbias.n4021 1010.98
R4916 Vbias.n4248 Vbias.n3984 1010.98
R4917 Vbias.n4242 Vbias.n3984 1010.98
R4918 Vbias.n4242 Vbias.n3997 1010.98
R4919 Vbias.n4238 Vbias.n3997 1010.98
R4920 Vbias.n4247 Vbias.n3989 1010.98
R4921 Vbias.n4243 Vbias.n3989 1010.98
R4922 Vbias.n4243 Vbias.n3993 1010.98
R4923 Vbias.n4237 Vbias.n3993 1010.98
R4924 Vbias.n4173 Vbias.n4172 1010.98
R4925 Vbias.n4173 Vbias.n4060 1010.98
R4926 Vbias.n4072 Vbias.n4060 1010.98
R4927 Vbias.n4185 Vbias.n4072 1010.98
R4928 Vbias.n4176 Vbias.n4175 1010.98
R4929 Vbias.n4175 Vbias.n4059 1010.98
R4930 Vbias.n4075 Vbias.n4059 1010.98
R4931 Vbias.n4075 Vbias.n4071 1010.98
R4932 Vbias.n4158 Vbias.n4157 1010.98
R4933 Vbias.n4157 Vbias.n4046 1010.98
R4934 Vbias.n4149 Vbias.n4147 1010.98
R4935 Vbias.n4147 Vbias.n4045 1010.98
R4936 Vbias.n4133 Vbias.n4132 1010.98
R4937 Vbias.n4132 Vbias.n4018 1010.98
R4938 Vbias.n4082 Vbias.n4018 1010.98
R4939 Vbias.n4082 Vbias.n4030 1010.98
R4940 Vbias.n4130 Vbias.n4129 1010.98
R4941 Vbias.n4130 Vbias.n4017 1010.98
R4942 Vbias.n4081 Vbias.n4017 1010.98
R4943 Vbias.n4081 Vbias.n4029 1010.98
R4944 Vbias.n4096 Vbias.n3987 1010.98
R4945 Vbias.n4096 Vbias.n3995 1010.98
R4946 Vbias.n4092 Vbias.n3995 1010.98
R4947 Vbias.n4092 Vbias.n4004 1010.98
R4948 Vbias.n4095 Vbias.n3986 1010.98
R4949 Vbias.n4095 Vbias.n3994 1010.98
R4950 Vbias.n4091 Vbias.n3994 1010.98
R4951 Vbias.n4091 Vbias.n4003 1010.98
R4952 Vbias.n2625 Vbias.n2613 1010.98
R4953 Vbias.n4977 Vbias.n2613 1010.98
R4954 Vbias.n4977 Vbias.n2611 1010.98
R4955 Vbias.n4983 Vbias.n2611 1010.98
R4956 Vbias.n2617 Vbias.n2615 1010.98
R4957 Vbias.n4976 Vbias.n2615 1010.98
R4958 Vbias.n4976 Vbias.n2607 1010.98
R4959 Vbias.n4984 Vbias.n2607 1010.98
R4960 Vbias.n4959 Vbias.n2629 1010.98
R4961 Vbias.n4965 Vbias.n2629 1010.98
R4962 Vbias.n4958 Vbias.n2621 1010.98
R4963 Vbias.n4966 Vbias.n2621 1010.98
R4964 Vbias.n4939 Vbias.n4934 1010.98
R4965 Vbias.n4934 Vbias.n2640 1010.98
R4966 Vbias.n2640 Vbias.n2638 1010.98
R4967 Vbias.n2638 Vbias.n2633 1010.98
R4968 Vbias.n4940 Vbias.n2641 1010.98
R4969 Vbias.n4947 Vbias.n2641 1010.98
R4970 Vbias.n4947 Vbias.n2637 1010.98
R4971 Vbias.n2637 Vbias.n2632 1010.98
R4972 Vbias.n4917 Vbias.n4912 1010.98
R4973 Vbias.n4912 Vbias.n2654 1010.98
R4974 Vbias.n2654 Vbias.n2652 1010.98
R4975 Vbias.n2652 Vbias.n2647 1010.98
R4976 Vbias.n4918 Vbias.n2655 1010.98
R4977 Vbias.n4924 Vbias.n2655 1010.98
R4978 Vbias.n4924 Vbias.n2651 1010.98
R4979 Vbias.n2651 Vbias.n2646 1010.98
R4980 Vbias.n2994 Vbias.n2984 1010.98
R4981 Vbias.n3039 Vbias.n2994 1010.98
R4982 Vbias.n3039 Vbias.n2995 1010.98
R4983 Vbias.n3033 Vbias.n2995 1010.98
R4984 Vbias.n2999 Vbias.n2983 1010.98
R4985 Vbias.n3038 Vbias.n2999 1010.98
R4986 Vbias.n3038 Vbias.n3000 1010.98
R4987 Vbias.n3034 Vbias.n3000 1010.98
R4988 Vbias.n2977 Vbias.n2971 1010.98
R4989 Vbias.n3049 Vbias.n2977 1010.98
R4990 Vbias.n3055 Vbias.n2976 1010.98
R4991 Vbias.n3072 Vbias.n2976 1010.98
R4992 Vbias.n2947 Vbias.n2937 1010.98
R4993 Vbias.n3115 Vbias.n2947 1010.98
R4994 Vbias.n3115 Vbias.n2948 1010.98
R4995 Vbias.n3109 Vbias.n2948 1010.98
R4996 Vbias.n2952 Vbias.n2936 1010.98
R4997 Vbias.n3114 Vbias.n2952 1010.98
R4998 Vbias.n3114 Vbias.n2953 1010.98
R4999 Vbias.n3110 Vbias.n2953 1010.98
R5000 Vbias.n2918 Vbias.n2908 1010.98
R5001 Vbias.n3153 Vbias.n2918 1010.98
R5002 Vbias.n3153 Vbias.n2919 1010.98
R5003 Vbias.n3147 Vbias.n2919 1010.98
R5004 Vbias.n2923 Vbias.n2907 1010.98
R5005 Vbias.n3152 Vbias.n2923 1010.98
R5006 Vbias.n3152 Vbias.n2924 1010.98
R5007 Vbias.n3148 Vbias.n2924 1010.98
R5008 Vbias.n3018 Vbias.n3017 1010.98
R5009 Vbias.n3017 Vbias.n2997 1010.98
R5010 Vbias.n3024 Vbias.n2997 1010.98
R5011 Vbias.n3024 Vbias.n3010 1010.98
R5012 Vbias.n3015 Vbias.n2987 1010.98
R5013 Vbias.n3015 Vbias.n2992 1010.98
R5014 Vbias.n3023 Vbias.n2992 1010.98
R5015 Vbias.n3023 Vbias.n3009 1010.98
R5016 Vbias.n3062 Vbias.n3061 1010.98
R5017 Vbias.n3061 Vbias.n2981 1010.98
R5018 Vbias.n2979 Vbias.n2972 1010.98
R5019 Vbias.n2980 Vbias.n2979 1010.98
R5020 Vbias.n3094 Vbias.n3093 1010.98
R5021 Vbias.n3093 Vbias.n2950 1010.98
R5022 Vbias.n3100 Vbias.n2950 1010.98
R5023 Vbias.n3100 Vbias.n2963 1010.98
R5024 Vbias.n3091 Vbias.n2940 1010.98
R5025 Vbias.n3091 Vbias.n2945 1010.98
R5026 Vbias.n3099 Vbias.n2945 1010.98
R5027 Vbias.n3099 Vbias.n2962 1010.98
R5028 Vbias.n3132 Vbias.n3131 1010.98
R5029 Vbias.n3131 Vbias.n2921 1010.98
R5030 Vbias.n3138 Vbias.n2921 1010.98
R5031 Vbias.n3138 Vbias.n2934 1010.98
R5032 Vbias.n3129 Vbias.n2911 1010.98
R5033 Vbias.n3129 Vbias.n2916 1010.98
R5034 Vbias.n3137 Vbias.n2916 1010.98
R5035 Vbias.n3137 Vbias.n2933 1010.98
R5036 Vbias.n2755 Vbias.n2745 1010.98
R5037 Vbias.n4715 Vbias.n2755 1010.98
R5038 Vbias.n4715 Vbias.n2756 1010.98
R5039 Vbias.n4709 Vbias.n2756 1010.98
R5040 Vbias.n2760 Vbias.n2744 1010.98
R5041 Vbias.n4714 Vbias.n2760 1010.98
R5042 Vbias.n4714 Vbias.n2761 1010.98
R5043 Vbias.n4710 Vbias.n2761 1010.98
R5044 Vbias.n2738 Vbias.n2732 1010.98
R5045 Vbias.n4725 Vbias.n2738 1010.98
R5046 Vbias.n4731 Vbias.n2737 1010.98
R5047 Vbias.n4748 Vbias.n2737 1010.98
R5048 Vbias.n2708 Vbias.n2698 1010.98
R5049 Vbias.n4791 Vbias.n2708 1010.98
R5050 Vbias.n4791 Vbias.n2709 1010.98
R5051 Vbias.n4785 Vbias.n2709 1010.98
R5052 Vbias.n2713 Vbias.n2697 1010.98
R5053 Vbias.n4790 Vbias.n2713 1010.98
R5054 Vbias.n4790 Vbias.n2714 1010.98
R5055 Vbias.n4786 Vbias.n2714 1010.98
R5056 Vbias.n2679 Vbias.n2669 1010.98
R5057 Vbias.n4829 Vbias.n2679 1010.98
R5058 Vbias.n4829 Vbias.n2680 1010.98
R5059 Vbias.n4823 Vbias.n2680 1010.98
R5060 Vbias.n2684 Vbias.n2668 1010.98
R5061 Vbias.n4828 Vbias.n2684 1010.98
R5062 Vbias.n4828 Vbias.n2685 1010.98
R5063 Vbias.n4824 Vbias.n2685 1010.98
R5064 Vbias.n4694 Vbias.n4693 1010.98
R5065 Vbias.n4693 Vbias.n2758 1010.98
R5066 Vbias.n4700 Vbias.n2758 1010.98
R5067 Vbias.n4700 Vbias.n2771 1010.98
R5068 Vbias.n4691 Vbias.n2748 1010.98
R5069 Vbias.n4691 Vbias.n2753 1010.98
R5070 Vbias.n4699 Vbias.n2753 1010.98
R5071 Vbias.n4699 Vbias.n2770 1010.98
R5072 Vbias.n4738 Vbias.n4737 1010.98
R5073 Vbias.n4737 Vbias.n2742 1010.98
R5074 Vbias.n2740 Vbias.n2733 1010.98
R5075 Vbias.n2741 Vbias.n2740 1010.98
R5076 Vbias.n4770 Vbias.n4769 1010.98
R5077 Vbias.n4769 Vbias.n2711 1010.98
R5078 Vbias.n4776 Vbias.n2711 1010.98
R5079 Vbias.n4776 Vbias.n2724 1010.98
R5080 Vbias.n4767 Vbias.n2701 1010.98
R5081 Vbias.n4767 Vbias.n2706 1010.98
R5082 Vbias.n4775 Vbias.n2706 1010.98
R5083 Vbias.n4775 Vbias.n2723 1010.98
R5084 Vbias.n4808 Vbias.n4807 1010.98
R5085 Vbias.n4807 Vbias.n2682 1010.98
R5086 Vbias.n4814 Vbias.n2682 1010.98
R5087 Vbias.n4814 Vbias.n2695 1010.98
R5088 Vbias.n4805 Vbias.n2672 1010.98
R5089 Vbias.n4805 Vbias.n2677 1010.98
R5090 Vbias.n4813 Vbias.n2677 1010.98
R5091 Vbias.n4813 Vbias.n2694 1010.98
R5092 Vbias.n4561 Vbias.n4551 1010.98
R5093 Vbias.n4569 Vbias.n4561 1010.98
R5094 Vbias.n4570 Vbias.n4569 1010.98
R5095 Vbias.n4570 Vbias.n4560 1010.98
R5096 Vbias.n4562 Vbias.n4552 1010.98
R5097 Vbias.n4562 Vbias.n4556 1010.98
R5098 Vbias.n4571 Vbias.n4556 1010.98
R5099 Vbias.n4571 Vbias.n4558 1010.98
R5100 Vbias.n6214 Vbias.n6203 1010.98
R5101 Vbias.n6214 Vbias.n6208 1010.98
R5102 Vbias.n6223 Vbias.n6208 1010.98
R5103 Vbias.n6223 Vbias.n6210 1010.98
R5104 Vbias.n6213 Vbias.n6202 1010.98
R5105 Vbias.n6221 Vbias.n6213 1010.98
R5106 Vbias.n6222 Vbias.n6221 1010.98
R5107 Vbias.n6222 Vbias.n6212 1010.98
R5108 Vbias.n6197 Vbias.n6189 1010.98
R5109 Vbias.n6197 Vbias.n6193 1010.98
R5110 Vbias.n6196 Vbias.n6188 1010.98
R5111 Vbias.n6196 Vbias.n6195 1010.98
R5112 Vbias.n6173 Vbias.n6156 1010.98
R5113 Vbias.n6173 Vbias.n6158 1010.98
R5114 Vbias.n6176 Vbias.n6158 1010.98
R5115 Vbias.n6176 Vbias.n6160 1010.98
R5116 Vbias.n6172 Vbias.n6168 1010.98
R5117 Vbias.n6179 Vbias.n6168 1010.98
R5118 Vbias.n6179 Vbias.n6166 1010.98
R5119 Vbias.n6183 Vbias.n6166 1010.98
R5120 Vbias.n6451 Vbias.n6440 1010.98
R5121 Vbias.n6451 Vbias.n6445 1010.98
R5122 Vbias.n6460 Vbias.n6445 1010.98
R5123 Vbias.n6460 Vbias.n6447 1010.98
R5124 Vbias.n6450 Vbias.n6439 1010.98
R5125 Vbias.n6458 Vbias.n6450 1010.98
R5126 Vbias.n6459 Vbias.n6458 1010.98
R5127 Vbias.n6459 Vbias.n6449 1010.98
R5128 Vbias.n6434 Vbias.n6426 1010.98
R5129 Vbias.n6434 Vbias.n6430 1010.98
R5130 Vbias.n6433 Vbias.n6425 1010.98
R5131 Vbias.n6433 Vbias.n6432 1010.98
R5132 Vbias.n6410 Vbias.n6374 1010.98
R5133 Vbias.n6410 Vbias.n6376 1010.98
R5134 Vbias.n6413 Vbias.n6376 1010.98
R5135 Vbias.n6413 Vbias.n6378 1010.98
R5136 Vbias.n6409 Vbias.n6386 1010.98
R5137 Vbias.n6416 Vbias.n6386 1010.98
R5138 Vbias.n6416 Vbias.n6384 1010.98
R5139 Vbias.n6420 Vbias.n6384 1010.98
R5140 Vbias.n6393 Vbias.n6366 1010.98
R5141 Vbias.n6393 Vbias.n6368 1010.98
R5142 Vbias.n6396 Vbias.n6368 1010.98
R5143 Vbias.n6396 Vbias.n6370 1010.98
R5144 Vbias.n6392 Vbias.n6389 1010.98
R5145 Vbias.n6399 Vbias.n6389 1010.98
R5146 Vbias.n6399 Vbias.n6387 1010.98
R5147 Vbias.n6403 Vbias.n6387 1010.98
R5148 Vbias.n905 Vbias.n894 1010.98
R5149 Vbias.n905 Vbias.n899 1010.98
R5150 Vbias.n914 Vbias.n899 1010.98
R5151 Vbias.n914 Vbias.n901 1010.98
R5152 Vbias.n904 Vbias.n893 1010.98
R5153 Vbias.n912 Vbias.n904 1010.98
R5154 Vbias.n913 Vbias.n912 1010.98
R5155 Vbias.n913 Vbias.n903 1010.98
R5156 Vbias.n888 Vbias.n880 1010.98
R5157 Vbias.n888 Vbias.n884 1010.98
R5158 Vbias.n887 Vbias.n879 1010.98
R5159 Vbias.n887 Vbias.n886 1010.98
R5160 Vbias.n6472 Vbias.n869 1010.98
R5161 Vbias.n6472 Vbias.n871 1010.98
R5162 Vbias.n6481 Vbias.n871 1010.98
R5163 Vbias.n6481 Vbias.n873 1010.98
R5164 Vbias.n6488 Vbias.n6469 1010.98
R5165 Vbias.n6484 Vbias.n6469 1010.98
R5166 Vbias.n6484 Vbias.n6471 1010.98
R5167 Vbias.n6480 Vbias.n6471 1010.98
R5168 Vbias.n6466 Vbias.n861 1010.98
R5169 Vbias.n6466 Vbias.n863 1010.98
R5170 Vbias.n6495 Vbias.n863 1010.98
R5171 Vbias.n6495 Vbias.n865 1010.98
R5172 Vbias.n6502 Vbias.n6463 1010.98
R5173 Vbias.n6498 Vbias.n6463 1010.98
R5174 Vbias.n6498 Vbias.n6465 1010.98
R5175 Vbias.n6494 Vbias.n6465 1010.98
R5176 Vbias.n7387 Vbias.n7381 1010.98
R5177 Vbias.n7408 Vbias.n7387 1010.98
R5178 Vbias.n7408 Vbias.n7388 1010.98
R5179 Vbias.n7401 Vbias.n7388 1010.98
R5180 Vbias.n7391 Vbias.n7380 1010.98
R5181 Vbias.n7407 Vbias.n7391 1010.98
R5182 Vbias.n7407 Vbias.n7392 1010.98
R5183 Vbias.n7403 Vbias.n7392 1010.98
R5184 Vbias.n7373 Vbias.n7369 1010.98
R5185 Vbias.n7417 Vbias.n7373 1010.98
R5186 Vbias.n7379 Vbias.n7372 1010.98
R5187 Vbias.n7421 Vbias.n7372 1010.98
R5188 Vbias.n7349 Vbias.n7343 1010.98
R5189 Vbias.n7442 Vbias.n7349 1010.98
R5190 Vbias.n7442 Vbias.n7350 1010.98
R5191 Vbias.n7436 Vbias.n7350 1010.98
R5192 Vbias.n7353 Vbias.n7342 1010.98
R5193 Vbias.n7441 Vbias.n7353 1010.98
R5194 Vbias.n7441 Vbias.n7354 1010.98
R5195 Vbias.n7437 Vbias.n7354 1010.98
R5196 Vbias.n7463 Vbias.n7328 1010.98
R5197 Vbias.n7457 Vbias.n7328 1010.98
R5198 Vbias.n7457 Vbias.n7336 1010.98
R5199 Vbias.n7453 Vbias.n7336 1010.98
R5200 Vbias.n7462 Vbias.n7330 1010.98
R5201 Vbias.n7458 Vbias.n7330 1010.98
R5202 Vbias.n7458 Vbias.n7334 1010.98
R5203 Vbias.n7452 Vbias.n7334 1010.98
R5204 Vbias.n6143 Vbias.n6139 1010.98
R5205 Vbias.n6642 Vbias.n6139 1010.98
R5206 Vbias.n6642 Vbias.n6146 1010.98
R5207 Vbias.n6638 Vbias.n6146 1010.98
R5208 Vbias.n6140 Vbias.n6136 1010.98
R5209 Vbias.n6145 Vbias.n6140 1010.98
R5210 Vbias.n6152 Vbias.n6145 1010.98
R5211 Vbias.n6637 Vbias.n6152 1010.98
R5212 Vbias.n1712 Vbias.n1704 1010.98
R5213 Vbias.n2052 Vbias.n1712 1010.98
R5214 Vbias.n2052 Vbias.n1713 1010.98
R5215 Vbias.n2047 Vbias.n1713 1010.98
R5216 Vbias.n1709 Vbias.n1705 1010.98
R5217 Vbias.n2053 Vbias.n1709 1010.98
R5218 Vbias.n2053 Vbias.n1710 1010.98
R5219 Vbias.n2046 Vbias.n1710 1010.98
R5220 Vbias.n6681 Vbias.n1453 1010.98
R5221 Vbias.n6687 Vbias.n1453 1010.98
R5222 Vbias.n1457 Vbias.n1454 1010.98
R5223 Vbias.n1454 Vbias.n1451 1010.98
R5224 Vbias.n4882 Vbias.n4852 918.212
R5225 Vbias.n4888 Vbias.n4850 918.212
R5226 Vbias.n4863 Vbias.n4856 866.087
R5227 Vbias.n4867 Vbias.n4863 866.087
R5228 Vbias.n4877 Vbias.n4858 866.087
R5229 Vbias.n4873 Vbias.n4858 866.087
R5230 Vbias.n4853 Vbias.n4849 866.087
R5231 Vbias.n4884 Vbias.n4853 866.087
R5232 Vbias.n4880 Vbias.n4848 866.087
R5233 Vbias.n4883 Vbias.n4880 866.087
R5234 Vbias.n7402 Vbias.n7399 858.293
R5235 Vbias.n4885 Vbias.n4852 845.5
R5236 Vbias.n4888 Vbias.n4887 845.5
R5237 Vbias.n4881 Vbias.n4851 819.201
R5238 Vbias.n4886 Vbias.n4851 819.201
R5239 Vbias.n7887 Vbias.n447 770.634
R5240 Vbias.n7871 Vbias.n457 770.634
R5241 Vbias.n7752 Vbias.n667 770.634
R5242 Vbias.n7736 Vbias.n678 770.634
R5243 Vbias.t835 Vbias.n7 770.125
R5244 Vbias.t835 Vbias.n3701 770.125
R5245 Vbias.n3700 Vbias.t170 770.125
R5246 Vbias.n3459 Vbias.t170 770.125
R5247 Vbias.t575 Vbias.n3459 770.125
R5248 Vbias.t575 Vbias.n3461 770.125
R5249 Vbias.t389 Vbias.n3461 770.125
R5250 Vbias.t389 Vbias.n3663 770.125
R5251 Vbias.n3662 Vbias.t462 770.125
R5252 Vbias.n3488 Vbias.t462 770.125
R5253 Vbias.t624 Vbias.n3488 770.125
R5254 Vbias.t624 Vbias.n3490 770.125
R5255 Vbias.t417 Vbias.n3490 770.125
R5256 Vbias.t417 Vbias.n3625 770.125
R5257 Vbias.n3624 Vbias.t809 770.125
R5258 Vbias.n3593 Vbias.t809 770.125
R5259 Vbias.n3598 Vbias.t148 770.125
R5260 Vbias.n3612 Vbias.t148 770.125
R5261 Vbias.n3612 Vbias.t693 770.125
R5262 Vbias.t693 Vbias.n3587 770.125
R5263 Vbias.n3586 Vbias.t609 770.125
R5264 Vbias.n3535 Vbias.t609 770.125
R5265 Vbias.t684 Vbias.n3535 770.125
R5266 Vbias.t684 Vbias.n3537 770.125
R5267 Vbias.t6 Vbias.n3537 770.125
R5268 Vbias.t6 Vbias.n2773 770.125
R5269 Vbias.t877 Vbias.n8 770.125
R5270 Vbias.t877 Vbias.n3432 770.125
R5271 Vbias.n3431 Vbias.t550 770.125
R5272 Vbias.n3190 Vbias.t550 770.125
R5273 Vbias.t653 Vbias.n3190 770.125
R5274 Vbias.t653 Vbias.n3192 770.125
R5275 Vbias.t314 Vbias.n3192 770.125
R5276 Vbias.t314 Vbias.n3394 770.125
R5277 Vbias.n3393 Vbias.t374 770.125
R5278 Vbias.n3219 Vbias.t374 770.125
R5279 Vbias.t692 Vbias.n3219 770.125
R5280 Vbias.t692 Vbias.n3221 770.125
R5281 Vbias.t150 Vbias.n3221 770.125
R5282 Vbias.t150 Vbias.n3356 770.125
R5283 Vbias.n3355 Vbias.t387 770.125
R5284 Vbias.n3324 Vbias.t387 770.125
R5285 Vbias.n3329 Vbias.t583 770.125
R5286 Vbias.n3343 Vbias.t583 770.125
R5287 Vbias.n3343 Vbias.t308 770.125
R5288 Vbias.t308 Vbias.n3318 770.125
R5289 Vbias.n3317 Vbias.t881 770.125
R5290 Vbias.n3266 Vbias.t881 770.125
R5291 Vbias.t514 Vbias.n3266 770.125
R5292 Vbias.t514 Vbias.n3268 770.125
R5293 Vbias.t363 Vbias.n3268 770.125
R5294 Vbias.t363 Vbias.n2774 770.125
R5295 Vbias.t651 Vbias.n9 770.125
R5296 Vbias.t651 Vbias.n3970 770.125
R5297 Vbias.n3969 Vbias.t458 770.125
R5298 Vbias.n3728 Vbias.t458 770.125
R5299 Vbias.t310 Vbias.n3728 770.125
R5300 Vbias.t310 Vbias.n3730 770.125
R5301 Vbias.t127 Vbias.n3730 770.125
R5302 Vbias.t127 Vbias.n3932 770.125
R5303 Vbias.n3931 Vbias.t351 770.125
R5304 Vbias.n3757 Vbias.t351 770.125
R5305 Vbias.t696 Vbias.n3757 770.125
R5306 Vbias.t696 Vbias.n3759 770.125
R5307 Vbias.t435 Vbias.n3759 770.125
R5308 Vbias.t435 Vbias.n3894 770.125
R5309 Vbias.n3893 Vbias.t450 770.125
R5310 Vbias.n3862 Vbias.t450 770.125
R5311 Vbias.n3867 Vbias.t124 770.125
R5312 Vbias.n3881 Vbias.t124 770.125
R5313 Vbias.n3881 Vbias.t545 770.125
R5314 Vbias.t545 Vbias.n3856 770.125
R5315 Vbias.n3855 Vbias.t524 770.125
R5316 Vbias.n3804 Vbias.t524 770.125
R5317 Vbias.t620 Vbias.n3804 770.125
R5318 Vbias.t620 Vbias.n3806 770.125
R5319 Vbias.t438 Vbias.n3806 770.125
R5320 Vbias.t438 Vbias.n2775 770.125
R5321 Vbias.t833 Vbias.n2905 770.125
R5322 Vbias.t833 Vbias.n3162 770.125
R5323 Vbias.n3161 Vbias.t137 770.125
R5324 Vbias.n2920 Vbias.t137 770.125
R5325 Vbias.t365 Vbias.n2920 770.125
R5326 Vbias.t365 Vbias.n2922 770.125
R5327 Vbias.t639 Vbias.n2922 770.125
R5328 Vbias.t639 Vbias.n3124 770.125
R5329 Vbias.n3123 Vbias.t726 770.125
R5330 Vbias.n2949 Vbias.t726 770.125
R5331 Vbias.t147 Vbias.n2949 770.125
R5332 Vbias.t147 Vbias.n2951 770.125
R5333 Vbias.t130 Vbias.n2951 770.125
R5334 Vbias.t130 Vbias.n3086 770.125
R5335 Vbias.n3085 Vbias.t871 770.125
R5336 Vbias.n3054 Vbias.t871 770.125
R5337 Vbias.n3059 Vbias.t280 770.125
R5338 Vbias.n3073 Vbias.t280 770.125
R5339 Vbias.n3073 Vbias.t311 770.125
R5340 Vbias.t311 Vbias.n3048 770.125
R5341 Vbias.n3047 Vbias.t165 770.125
R5342 Vbias.n2996 Vbias.t165 770.125
R5343 Vbias.t362 Vbias.n2996 770.125
R5344 Vbias.t362 Vbias.n2998 770.125
R5345 Vbias.t775 Vbias.n2998 770.125
R5346 Vbias.t775 Vbias.n2776 770.125
R5347 Vbias.n4844 Vbias.t875 770.125
R5348 Vbias.n4838 Vbias.t875 770.125
R5349 Vbias.n4837 Vbias.t227 770.125
R5350 Vbias.n2681 Vbias.t227 770.125
R5351 Vbias.t400 Vbias.n2681 770.125
R5352 Vbias.t400 Vbias.n2683 770.125
R5353 Vbias.t448 Vbias.n2683 770.125
R5354 Vbias.t448 Vbias.n4800 770.125
R5355 Vbias.n4799 Vbias.t133 770.125
R5356 Vbias.n2710 Vbias.t133 770.125
R5357 Vbias.t626 Vbias.n2710 770.125
R5358 Vbias.t626 Vbias.n2712 770.125
R5359 Vbias.t282 Vbias.n2712 770.125
R5360 Vbias.t282 Vbias.n4762 770.125
R5361 Vbias.n4761 Vbias.t446 770.125
R5362 Vbias.n4730 Vbias.t446 770.125
R5363 Vbias.n4735 Vbias.t348 770.125
R5364 Vbias.n4749 Vbias.t348 770.125
R5365 Vbias.n4749 Vbias.t312 770.125
R5366 Vbias.t312 Vbias.n4724 770.125
R5367 Vbias.n4723 Vbias.t460 770.125
R5368 Vbias.n2757 Vbias.t460 770.125
R5369 Vbias.t304 Vbias.n2757 770.125
R5370 Vbias.t304 Vbias.n2759 770.125
R5371 Vbias.t297 Vbias.n2759 770.125
R5372 Vbias.t297 Vbias.n4686 770.125
R5373 Vbias.t837 Vbias.n4261 770.125
R5374 Vbias.n4262 Vbias.t837 770.125
R5375 Vbias.t84 Vbias.n2883 770.125
R5376 Vbias.t84 Vbias.n2874 770.125
R5377 Vbias.t576 Vbias.n2874 770.125
R5378 Vbias.t576 Vbias.n2866 770.125
R5379 Vbias.t502 Vbias.n2866 770.125
R5380 Vbias.t502 Vbias.n2868 770.125
R5381 Vbias.t167 Vbias.n2849 770.125
R5382 Vbias.t167 Vbias.n2840 770.125
R5383 Vbias.t596 Vbias.n2840 770.125
R5384 Vbias.t596 Vbias.n2830 770.125
R5385 Vbias.t343 Vbias.n2830 770.125
R5386 Vbias.t343 Vbias.n2834 770.125
R5387 Vbias.n2833 Vbias.t637 770.125
R5388 Vbias.n4338 Vbias.t637 770.125
R5389 Vbias.n4343 Vbias.t128 770.125
R5390 Vbias.n4352 Vbias.t128 770.125
R5391 Vbias.n4352 Vbias.t466 770.125
R5392 Vbias.n4364 Vbias.t466 770.125
R5393 Vbias.t507 Vbias.n4365 770.125
R5394 Vbias.t507 Vbias.n2786 770.125
R5395 Vbias.t372 Vbias.n2786 770.125
R5396 Vbias.t372 Vbias.n2790 770.125
R5397 Vbias.n2790 Vbias.t162 770.125
R5398 Vbias.n4406 Vbias.t162 770.125
R5399 Vbias.n7225 Vbias.n976 753.46
R5400 Vbias.n6710 Vbias.n976 751.688
R5401 Vbias.n4874 Vbias.n4861 729.976
R5402 Vbias.n4866 Vbias.n4861 729.976
R5403 Vbias.n4864 Vbias.n4859 729.976
R5404 Vbias.n4876 Vbias.n4859 729.976
R5405 Vbias.n8076 Vbias.n8075 726.005
R5406 Vbias.n6751 Vbias.n1443 696.773
R5407 Vbias.n6701 Vbias.n1305 696.773
R5408 Vbias.n5012 Vbias.n5011 696.773
R5409 Vbias.n5016 Vbias.n2228 696.773
R5410 Vbias.n5533 Vbias.n5532 696.773
R5411 Vbias.n5878 Vbias.n1673 696.773
R5412 Vbias.n6675 Vbias.t293 648.799
R5413 Vbias.n1475 Vbias.t293 648.799
R5414 Vbias.t539 Vbias.n1475 648.799
R5415 Vbias.t539 Vbias.n1476 648.799
R5416 Vbias.n1488 Vbias.t52 648.799
R5417 Vbias.t537 Vbias.n1488 648.799
R5418 Vbias.t537 Vbias.n1489 648.799
R5419 Vbias.t549 Vbias.n1489 648.799
R5420 Vbias.t549 Vbias.n6132 648.799
R5421 Vbias.n6131 Vbias.t615 648.799
R5422 Vbias.n1504 Vbias.t615 648.799
R5423 Vbias.t646 Vbias.n757 648.799
R5424 Vbias.t481 Vbias.n757 648.799
R5425 Vbias.t481 Vbias.n765 648.799
R5426 Vbias.t611 Vbias.n6303 648.799
R5427 Vbias.n6308 Vbias.t611 648.799
R5428 Vbias.n6307 Vbias.t253 648.799
R5429 Vbias.t253 Vbias.n6291 648.799
R5430 Vbias.t608 Vbias.n6291 648.799
R5431 Vbias.t608 Vbias.n6280 648.799
R5432 Vbias.t444 Vbias.n6280 648.799
R5433 Vbias.t444 Vbias.n6285 648.799
R5434 Vbias.n6284 Vbias.t18 648.799
R5435 Vbias.t18 Vbias.n6269 648.799
R5436 Vbias.t755 Vbias.n6269 648.799
R5437 Vbias.t755 Vbias.n6263 648.799
R5438 Vbias.t735 Vbias.n6263 648.799
R5439 Vbias.t464 Vbias.n6252 648.799
R5440 Vbias.t464 Vbias.n6253 648.799
R5441 Vbias.n6253 Vbias.t748 648.799
R5442 Vbias.n6352 Vbias.t748 648.799
R5443 Vbias.t78 Vbias.n6353 648.799
R5444 Vbias.t78 Vbias.n6234 648.799
R5445 Vbias.t521 Vbias.n6234 648.799
R5446 Vbias.t521 Vbias.n6235 648.799
R5447 Vbias.n6235 Vbias.t501 648.799
R5448 Vbias.n6589 Vbias.t501 648.799
R5449 Vbias.n6590 Vbias.t607 648.799
R5450 Vbias.n6598 Vbias.t607 648.799
R5451 Vbias.n6598 Vbias.t14 648.799
R5452 Vbias.n7652 Vbias.t14 648.799
R5453 Vbias.n7651 Vbias.t366 648.799
R5454 Vbias.n7645 Vbias.t366 648.799
R5455 Vbias.n7644 Vbias.t233 648.799
R5456 Vbias.n788 Vbias.t233 648.799
R5457 Vbias.t769 Vbias.n788 648.799
R5458 Vbias.t769 Vbias.n789 648.799
R5459 Vbias.t657 Vbias.n789 648.799
R5460 Vbias.t657 Vbias.n7630 648.799
R5461 Vbias.n7629 Vbias.t96 648.799
R5462 Vbias.n807 Vbias.t96 648.799
R5463 Vbias.t847 Vbias.n807 648.799
R5464 Vbias.t847 Vbias.n808 648.799
R5465 Vbias.t346 Vbias.n7615 648.799
R5466 Vbias.n7614 Vbias.t564 648.799
R5467 Vbias.n829 Vbias.t564 648.799
R5468 Vbias.t353 Vbias.n829 648.799
R5469 Vbias.t353 Vbias.n830 648.799
R5470 Vbias.t34 Vbias.n849 648.799
R5471 Vbias.t34 Vbias.n843 648.799
R5472 Vbias.t0 Vbias.n843 648.799
R5473 Vbias.t0 Vbias.n844 648.799
R5474 Vbias.t649 Vbias.n844 648.799
R5475 Vbias.t649 Vbias.n857 648.799
R5476 Vbias.n6508 Vbias.t368 648.799
R5477 Vbias.n6517 Vbias.t368 648.799
R5478 Vbias.t402 Vbias.n6519 648.799
R5479 Vbias.n6519 Vbias.t328 648.799
R5480 Vbias.n7531 Vbias.t328 648.799
R5481 Vbias.n7530 Vbias.t156 648.799
R5482 Vbias.n7524 Vbias.t156 648.799
R5483 Vbias.n7523 Vbias.t208 648.799
R5484 Vbias.n939 Vbias.t208 648.799
R5485 Vbias.t376 Vbias.n939 648.799
R5486 Vbias.t376 Vbias.n940 648.799
R5487 Vbias.t399 Vbias.n940 648.799
R5488 Vbias.t399 Vbias.n7509 648.799
R5489 Vbias.n7508 Vbias.t16 648.799
R5490 Vbias.n962 Vbias.t16 648.799
R5491 Vbias.t377 Vbias.n962 648.799
R5492 Vbias.t377 Vbias.n963 648.799
R5493 Vbias.t806 Vbias.n963 648.799
R5494 Vbias.n7492 Vbias.t571 648.799
R5495 Vbias.n984 Vbias.t571 648.799
R5496 Vbias.t390 Vbias.n984 648.799
R5497 Vbias.t390 Vbias.n985 648.799
R5498 Vbias.t48 Vbias.n1004 648.799
R5499 Vbias.t48 Vbias.n998 648.799
R5500 Vbias.t703 Vbias.n998 648.799
R5501 Vbias.t703 Vbias.n999 648.799
R5502 Vbias.t699 Vbias.n999 648.799
R5503 Vbias.t699 Vbias.n1018 648.799
R5504 Vbias.n1017 Vbias.t888 648.799
R5505 Vbias.n7544 Vbias.t888 648.799
R5506 Vbias.n7544 Vbias.t717 648.799
R5507 Vbias.n1026 Vbias.t717 648.799
R5508 Vbias.t477 Vbias.n1028 648.799
R5509 Vbias.n7317 Vbias.t477 648.799
R5510 Vbias.n7316 Vbias.t261 648.799
R5511 Vbias.n1036 Vbias.t261 648.799
R5512 Vbias.t475 Vbias.n1036 648.799
R5513 Vbias.t475 Vbias.n1037 648.799
R5514 Vbias.t819 Vbias.n1037 648.799
R5515 Vbias.t819 Vbias.n7302 648.799
R5516 Vbias.n7301 Vbias.t68 648.799
R5517 Vbias.n1057 Vbias.t68 648.799
R5518 Vbias.t619 Vbias.n1057 648.799
R5519 Vbias.t619 Vbias.n1058 648.799
R5520 Vbias.t669 Vbias.n7287 648.799
R5521 Vbias.n7286 Vbias.t143 648.799
R5522 Vbias.n7234 Vbias.t143 648.799
R5523 Vbias.t580 Vbias.n7234 648.799
R5524 Vbias.t580 Vbias.n7235 648.799
R5525 Vbias.t116 Vbias.n7254 648.799
R5526 Vbias.t116 Vbias.n7248 648.799
R5527 Vbias.t788 Vbias.n7248 648.799
R5528 Vbias.t788 Vbias.n7249 648.799
R5529 Vbias.t566 Vbias.n7249 648.799
R5530 Vbias.n6750 Vbias.n6749 641.857
R5531 Vbias.n6737 Vbias.n6736 641.857
R5532 Vbias.n5553 Vbias.n5552 641.857
R5533 Vbias.n5535 Vbias.n5534 641.857
R5534 Vbias.n5877 Vbias.n5876 641.857
R5535 Vbias.n4875 Vbias.n4860 630.966
R5536 Vbias.n4865 Vbias.n4860 630.966
R5537 Vbias.n7790 Vbias.n7789 625.822
R5538 Vbias.n7778 Vbias.n7777 625.822
R5539 Vbias.n634 Vbias.n633 625.822
R5540 Vbias.n7765 Vbias.n7764 625.822
R5541 Vbias.n7859 Vbias.n7858 625.822
R5542 Vbias.n7847 Vbias.n7846 625.822
R5543 Vbias.n520 Vbias.n519 625.822
R5544 Vbias.n7834 Vbias.n7833 625.822
R5545 Vbias.n7925 Vbias.n7924 625.822
R5546 Vbias.n7913 Vbias.n7912 625.822
R5547 Vbias.n414 Vbias.n413 625.822
R5548 Vbias.n7900 Vbias.n7899 625.822
R5549 Vbias.n268 Vbias.n223 625.822
R5550 Vbias.n287 Vbias.n286 625.822
R5551 Vbias.n299 Vbias.n298 625.822
R5552 Vbias.n307 Vbias.n190 625.822
R5553 Vbias.n1256 Vbias.n1255 625.822
R5554 Vbias.n1225 Vbias.n1224 625.822
R5555 Vbias.n7218 Vbias.n7217 625.822
R5556 Vbias.n6989 Vbias.n6988 625.822
R5557 Vbias.n6958 Vbias.n6957 625.822
R5558 Vbias.n7114 Vbias.n7113 625.822
R5559 Vbias.n1393 Vbias.n1383 625.822
R5560 Vbias.n6870 Vbias.n6869 625.822
R5561 Vbias.n6893 Vbias.n6892 625.822
R5562 Vbias.n1604 Vbias.n1594 625.822
R5563 Vbias.n6012 Vbias.n6011 625.822
R5564 Vbias.n6038 Vbias.n6037 625.822
R5565 Vbias.n5397 Vbias.n5396 625.822
R5566 Vbias.n5366 Vbias.n5365 625.822
R5567 Vbias.n5350 Vbias.n5349 625.822
R5568 Vbias.n2341 Vbias.n2331 625.822
R5569 Vbias.n5239 Vbias.n5238 625.822
R5570 Vbias.n5262 Vbias.n5261 625.822
R5571 Vbias.n2565 Vbias.n2564 625.822
R5572 Vbias.n2534 Vbias.n2533 625.822
R5573 Vbias.n2518 Vbias.n2517 625.822
R5574 Vbias.n4535 Vbias.n4534 625.822
R5575 Vbias.n4474 Vbias.n4460 625.822
R5576 Vbias.n4490 Vbias.n4482 625.822
R5577 Vbias.n7450 Vbias.n7449 625.822
R5578 Vbias.n7434 Vbias.n7433 625.822
R5579 Vbias.n7376 Vbias.n7375 625.822
R5580 Vbias.n7416 Vbias.n7415 625.822
R5581 Vbias.n6491 Vbias.n6490 625.822
R5582 Vbias.n6477 Vbias.n6476 625.822
R5583 Vbias.n7567 Vbias.n7566 625.822
R5584 Vbias.n7557 Vbias.n7556 625.822
R5585 Vbias.n6406 Vbias.n6405 625.822
R5586 Vbias.n6424 Vbias.n6422 625.822
R5587 Vbias.n6554 Vbias.n6553 625.822
R5588 Vbias.n6544 Vbias.n6543 625.822
R5589 Vbias.n6169 Vbias.n6150 625.822
R5590 Vbias.n6187 Vbias.n6185 625.822
R5591 Vbias.n6621 Vbias.n6620 625.822
R5592 Vbias.n6611 Vbias.n6610 625.822
R5593 Vbias.n706 Vbias.n698 625.822
R5594 Vbias.n725 Vbias.n716 625.822
R5595 Vbias.n7700 Vbias.n7699 625.822
R5596 Vbias.n7685 Vbias.n7684 625.822
R5597 Vbias.t511 Vbias.n7123 615.399
R5598 Vbias.t511 Vbias.n1143 615.399
R5599 Vbias.t776 Vbias.n1143 615.399
R5600 Vbias.t776 Vbias.n1144 615.399
R5601 Vbias.n1144 Vbias.t32 615.399
R5602 Vbias.n7142 Vbias.t32 615.399
R5603 Vbias.t354 Vbias.n7143 615.399
R5604 Vbias.t354 Vbias.n7144 615.399
R5605 Vbias.n7144 Vbias.t845 615.399
R5606 Vbias.n7159 Vbias.t845 615.399
R5607 Vbias.t498 Vbias.n7161 615.399
R5608 Vbias.n7162 Vbias.t498 615.399
R5609 Vbias.t493 Vbias.n1116 615.399
R5610 Vbias.t493 Vbias.n1117 615.399
R5611 Vbias.n1117 Vbias.t782 615.399
R5612 Vbias.n7178 Vbias.t782 615.399
R5613 Vbias.t62 Vbias.n7178 615.399
R5614 Vbias.n7179 Vbias.t62 615.399
R5615 Vbias.t658 Vbias.n1097 615.399
R5616 Vbias.t658 Vbias.n1098 615.399
R5617 Vbias.n1098 Vbias.t599 615.399
R5618 Vbias.n7195 Vbias.t599 615.399
R5619 Vbias.t176 Vbias.n7195 615.399
R5620 Vbias.t176 Vbias.n1071 615.399
R5621 Vbias.t230 Vbias.n7017 615.399
R5622 Vbias.t230 Vbias.n1331 615.399
R5623 Vbias.t496 Vbias.n1331 615.399
R5624 Vbias.t496 Vbias.n1332 615.399
R5625 Vbias.n1332 Vbias.t239 615.399
R5626 Vbias.n7036 Vbias.t239 615.399
R5627 Vbias.t556 Vbias.n7037 615.399
R5628 Vbias.t556 Vbias.n7038 615.399
R5629 Vbias.n7038 Vbias.t542 615.399
R5630 Vbias.n7053 Vbias.t542 615.399
R5631 Vbias.t381 Vbias.n7055 615.399
R5632 Vbias.n7056 Vbias.t381 615.399
R5633 Vbias.t715 Vbias.n1303 615.399
R5634 Vbias.n1304 Vbias.t355 615.399
R5635 Vbias.n7072 Vbias.t355 615.399
R5636 Vbias.t198 Vbias.n7072 615.399
R5637 Vbias.n7073 Vbias.t198 615.399
R5638 Vbias.t593 Vbias.n1284 615.399
R5639 Vbias.t593 Vbias.n1285 615.399
R5640 Vbias.n1285 Vbias.t636 615.399
R5641 Vbias.n7089 Vbias.t636 615.399
R5642 Vbias.t114 Vbias.n7089 615.399
R5643 Vbias.t114 Vbias.n1151 615.399
R5644 Vbias.n6074 Vbias.t731 615.399
R5645 Vbias.n6051 Vbias.t731 615.399
R5646 Vbias.t541 Vbias.n6051 615.399
R5647 Vbias.t541 Vbias.n6067 615.399
R5648 Vbias.n6067 Vbias.t267 615.399
R5649 Vbias.t267 Vbias.n6061 615.399
R5650 Vbias.n6060 Vbias.t756 615.399
R5651 Vbias.n6053 Vbias.t756 615.399
R5652 Vbias.n6053 Vbias.t490 615.399
R5653 Vbias.n6799 Vbias.t490 615.399
R5654 Vbias.n6798 Vbias.t330 615.399
R5655 Vbias.n6753 Vbias.t330 615.399
R5656 Vbias.n6760 Vbias.t781 615.399
R5657 Vbias.t799 Vbias.n6760 615.399
R5658 Vbias.t799 Vbias.n6763 615.399
R5659 Vbias.n6763 Vbias.t265 615.399
R5660 Vbias.n6770 Vbias.t265 615.399
R5661 Vbias.t340 Vbias.n6771 615.399
R5662 Vbias.t340 Vbias.n1434 615.399
R5663 Vbias.t647 Vbias.n1434 615.399
R5664 Vbias.t647 Vbias.n1435 615.399
R5665 Vbias.n1435 Vbias.t92 615.399
R5666 Vbias.n7014 Vbias.t92 615.399
R5667 Vbias.n1790 Vbias.t182 615.399
R5668 Vbias.n1789 Vbias.t500 615.399
R5669 Vbias.n1776 Vbias.t500 615.399
R5670 Vbias.n1776 Vbias.t305 615.399
R5671 Vbias.t76 Vbias.n1458 615.399
R5672 Vbias.n6076 Vbias.t76 615.399
R5673 Vbias.t155 Vbias.n5920 615.399
R5674 Vbias.t155 Vbias.n1630 615.399
R5675 Vbias.t730 Vbias.n1630 615.399
R5676 Vbias.n5929 Vbias.t730 615.399
R5677 Vbias.t212 Vbias.n5929 615.399
R5678 Vbias.t867 Vbias.n5933 615.399
R5679 Vbias.n5940 Vbias.t867 615.399
R5680 Vbias.t750 Vbias.n5940 615.399
R5681 Vbias.t750 Vbias.n1532 615.399
R5682 Vbias.n5484 Vbias.t710 615.399
R5683 Vbias.n5425 Vbias.t710 615.399
R5684 Vbias.n5425 Vbias.t479 615.399
R5685 Vbias.n5435 Vbias.t479 615.399
R5686 Vbias.t178 Vbias.n5435 615.399
R5687 Vbias.n5473 Vbias.t178 615.399
R5688 Vbias.n5472 Vbias.t736 615.399
R5689 Vbias.n5450 Vbias.t736 615.399
R5690 Vbias.t11 Vbias.n5450 615.399
R5691 Vbias.n5463 Vbias.t11 615.399
R5692 Vbias.n5462 Vbias.t395 615.399
R5693 Vbias.n5454 Vbias.t395 615.399
R5694 Vbias.t403 Vbias.n1664 615.399
R5695 Vbias.t449 Vbias.n1664 615.399
R5696 Vbias.t449 Vbias.n1665 615.399
R5697 Vbias.n1665 Vbias.t237 615.399
R5698 Vbias.n5897 Vbias.t237 615.399
R5699 Vbias.t592 Vbias.n5898 615.399
R5700 Vbias.t592 Vbias.n1648 615.399
R5701 Vbias.t757 Vbias.n1648 615.399
R5702 Vbias.t757 Vbias.n1649 615.399
R5703 Vbias.n1649 Vbias.t26 615.399
R5704 Vbias.n5917 Vbias.t26 615.399
R5705 Vbias.t605 Vbias.n5123 615.399
R5706 Vbias.n5129 Vbias.t605 615.399
R5707 Vbias.t520 Vbias.n5129 615.399
R5708 Vbias.t520 Vbias.n5132 615.399
R5709 Vbias.n5132 Vbias.t220 615.399
R5710 Vbias.n5139 Vbias.t220 615.399
R5711 Vbias.n5140 Vbias.t406 615.399
R5712 Vbias.n5148 Vbias.t406 615.399
R5713 Vbias.t686 Vbias.n5148 615.399
R5714 Vbias.n5168 Vbias.t686 615.399
R5715 Vbias.n5167 Vbias.t586 615.399
R5716 Vbias.n5158 Vbias.t586 615.399
R5717 Vbias.n5157 Vbias.t666 615.399
R5718 Vbias.n5508 Vbias.t554 615.399
R5719 Vbias.n2264 Vbias.t554 615.399
R5720 Vbias.t259 Vbias.n2264 615.399
R5721 Vbias.n5498 Vbias.t259 615.399
R5722 Vbias.n5497 Vbias.t339 615.399
R5723 Vbias.n2277 Vbias.t339 615.399
R5724 Vbias.n2277 Vbias.t894 615.399
R5725 Vbias.n2287 Vbias.t894 615.399
R5726 Vbias.t100 Vbias.n2287 615.399
R5727 Vbias.n5486 Vbias.t100 615.399
R5728 Vbias.t828 Vbias.n5038 615.399
R5729 Vbias.t828 Vbias.n2425 615.399
R5730 Vbias.t325 Vbias.n2425 615.399
R5731 Vbias.t325 Vbias.n2426 615.399
R5732 Vbias.n2426 Vbias.t241 615.399
R5733 Vbias.n5057 Vbias.t241 615.399
R5734 Vbias.n5058 Vbias.t892 615.399
R5735 Vbias.n5065 Vbias.t892 615.399
R5736 Vbias.t640 Vbias.n5065 615.399
R5737 Vbias.n5068 Vbias.t640 615.399
R5738 Vbias.n5067 Vbias.t385 615.399
R5739 Vbias.n5079 Vbias.t385 615.399
R5740 Vbias.t287 Vbias.n2396 615.399
R5741 Vbias.t722 Vbias.n2396 615.399
R5742 Vbias.t722 Vbias.n2397 615.399
R5743 Vbias.n2397 Vbias.t271 615.399
R5744 Vbias.n5100 Vbias.t271 615.399
R5745 Vbias.t411 Vbias.n5101 615.399
R5746 Vbias.t411 Vbias.n2380 615.399
R5747 Vbias.t627 Vbias.n2380 615.399
R5748 Vbias.t627 Vbias.n2381 615.399
R5749 Vbias.n2381 Vbias.t56 615.399
R5750 Vbias.n5120 Vbias.t56 615.399
R5751 Vbias.n4681 Vbias.t789 615.399
R5752 Vbias.n4563 Vbias.t789 615.399
R5753 Vbias.n4563 Vbias.t513 615.399
R5754 Vbias.n4573 Vbias.t513 615.399
R5755 Vbias.t269 Vbias.n4573 615.399
R5756 Vbias.n4671 Vbias.t269 615.399
R5757 Vbias.n4670 Vbias.t679 615.399
R5758 Vbias.n4588 Vbias.t679 615.399
R5759 Vbias.t452 Vbias.n4588 615.399
R5760 Vbias.n4661 Vbias.t452 615.399
R5761 Vbias.n4660 Vbias.t334 615.399
R5762 Vbias.n4617 Vbias.t334 615.399
R5763 Vbias.n4618 Vbias.t285 615.399
R5764 Vbias.t716 Vbias.n2592 615.399
R5765 Vbias.t716 Vbias.n4625 615.399
R5766 Vbias.n4625 Vbias.t214 615.399
R5767 Vbias.n4632 Vbias.t214 615.399
R5768 Vbias.t861 Vbias.n4633 615.399
R5769 Vbias.t861 Vbias.n4606 615.399
R5770 Vbias.t439 Vbias.n4606 615.399
R5771 Vbias.t439 Vbias.n4607 615.399
R5772 Vbias.n4607 Vbias.t42 615.399
R5773 Vbias.n5036 Vbias.t42 615.399
R5774 Vbias.t427 Vbias.n1527 600.622
R5775 Vbias.t427 Vbias.n1853 600.622
R5776 Vbias.t779 Vbias.n1853 600.622
R5777 Vbias.t779 Vbias.n1854 600.622
R5778 Vbias.t358 Vbias.n1854 600.622
R5779 Vbias.t358 Vbias.n1465 600.622
R5780 Vbias.n6677 Vbias.n1459 583.285
R5781 Vbias.n4904 Vbias.n4903 581.408
R5782 Vbias.n4956 Vbias.n4955 579.418
R5783 Vbias.n6678 Vbias.t305 571.298
R5784 Vbias.n3 Vbias.n1 541.741
R5785 Vbias.n8080 Vbias.n3 541.741
R5786 Vbias.t735 Vbias.n1444 530.452
R5787 Vbias.t806 Vbias.n7494 530.452
R5788 Vbias.n6676 Vbias.t182 527.198
R5789 Vbias.n7265 Vbias.n7261 516.5
R5790 Vbias.n7668 Vbias.n756 511.432
R5791 Vbias.n6531 Vbias.n6518 511.432
R5792 Vbias.t781 Vbias.n6751 503.144
R5793 Vbias.t403 Vbias.n5878 503.144
R5794 Vbias.t287 Vbias.n2228 503.144
R5795 Vbias.t758 Vbias.n1523 502.156
R5796 Vbias.t758 Vbias.n1887 502.156
R5797 Vbias.t883 Vbias.n1887 502.156
R5798 Vbias.t883 Vbias.n1893 502.156
R5799 Vbias.t644 Vbias.n1893 502.156
R5800 Vbias.t644 Vbias.n1460 502.156
R5801 Vbias.t662 Vbias.n1525 502.156
R5802 Vbias.t662 Vbias.n1994 502.156
R5803 Vbias.n1994 Vbias.t5 502.156
R5804 Vbias.n2010 Vbias.t5 502.156
R5805 Vbias.t853 Vbias.n2010 502.156
R5806 Vbias.t853 Vbias.n1463 502.156
R5807 Vbias.t868 Vbias.n1526 502.156
R5808 Vbias.t868 Vbias.n1921 502.156
R5809 Vbias.t870 Vbias.n1921 502.156
R5810 Vbias.t870 Vbias.n1922 502.156
R5811 Vbias.t422 Vbias.n1922 502.156
R5812 Vbias.t422 Vbias.n1464 502.156
R5813 Vbias.t140 Vbias.n6102 501.411
R5814 Vbias.t140 Vbias.n1515 501.411
R5815 Vbias.t142 Vbias.n1515 501.411
R5816 Vbias.t142 Vbias.n1516 501.411
R5817 Vbias.t594 Vbias.n1516 501.411
R5818 Vbias.t594 Vbias.n1462 501.411
R5819 Vbias.n5010 Vbias.n5009 492.76
R5820 Vbias.n4901 Vbias.n4891 482.887
R5821 Vbias.n8081 Vbias.n1 469.029
R5822 Vbias.n8081 Vbias.n8080 469.029
R5823 Vbias.n5932 Vbias.n1528 463.053
R5824 Vbias.n6132 Vbias.n6131 460.712
R5825 Vbias.n6303 Vbias.n765 460.712
R5826 Vbias.n6508 Vbias.n857 460.712
R5827 Vbias.n7531 Vbias.n7530 460.712
R5828 Vbias.t415 Vbias.n174 455.736
R5829 Vbias.n5601 Vbias.t415 455.736
R5830 Vbias.t235 Vbias.n5602 455.736
R5831 Vbias.t235 Vbias.n5579 455.736
R5832 Vbias.t2 Vbias.n5579 455.736
R5833 Vbias.t2 Vbias.n5580 455.736
R5834 Vbias.n5580 Vbias.t659 455.736
R5835 Vbias.n5619 Vbias.t659 455.736
R5836 Vbias.t90 Vbias.n5620 455.736
R5837 Vbias.t90 Vbias.n5561 455.736
R5838 Vbias.t306 Vbias.n5561 455.736
R5839 Vbias.t306 Vbias.n5562 455.736
R5840 Vbias.n5562 Vbias.t322 455.736
R5841 Vbias.t431 Vbias.n5639 455.736
R5842 Vbias.t431 Vbias.n2217 455.736
R5843 Vbias.t634 Vbias.n2217 455.736
R5844 Vbias.t634 Vbias.n2222 455.736
R5845 Vbias.n2221 Vbias.t72 455.736
R5846 Vbias.t72 Vbias.n2206 455.736
R5847 Vbias.t291 Vbias.n2206 455.736
R5848 Vbias.t291 Vbias.n2200 455.736
R5849 Vbias.t630 Vbias.n2200 455.736
R5850 Vbias.t630 Vbias.n447 455.736
R5851 Vbias.t772 Vbias.n457 455.736
R5852 Vbias.n5675 Vbias.t772 455.736
R5853 Vbias.t210 Vbias.n5676 455.736
R5854 Vbias.t210 Vbias.n2182 455.736
R5855 Vbias.t766 Vbias.n2182 455.736
R5856 Vbias.t766 Vbias.n2183 455.736
R5857 Vbias.n2183 Vbias.t379 455.736
R5858 Vbias.n5693 Vbias.t379 455.736
R5859 Vbias.t44 Vbias.n5694 455.736
R5860 Vbias.t44 Vbias.n2164 455.736
R5861 Vbias.t849 Vbias.n2164 455.736
R5862 Vbias.t849 Vbias.n2165 455.736
R5863 Vbias.n5712 Vbias.t457 455.736
R5864 Vbias.t151 Vbias.n5713 455.736
R5865 Vbias.t151 Vbias.n2146 455.736
R5866 Vbias.t697 Vbias.n2146 455.736
R5867 Vbias.t697 Vbias.n2151 455.736
R5868 Vbias.n2150 Vbias.t80 455.736
R5869 Vbias.t80 Vbias.n2135 455.736
R5870 Vbias.t568 Vbias.n2135 455.736
R5871 Vbias.t568 Vbias.n2129 455.736
R5872 Vbias.t643 Vbias.n2129 455.736
R5873 Vbias.t643 Vbias.n553 455.736
R5874 Vbias.t821 Vbias.n571 455.736
R5875 Vbias.n5751 Vbias.t821 455.736
R5876 Vbias.n5750 Vbias.t174 455.736
R5877 Vbias.t174 Vbias.n2118 455.736
R5878 Vbias.t350 Vbias.n2118 455.736
R5879 Vbias.t350 Vbias.n2107 455.736
R5880 Vbias.t585 Vbias.n2107 455.736
R5881 Vbias.t585 Vbias.n2112 455.736
R5882 Vbias.n2111 Vbias.t102 455.736
R5883 Vbias.t102 Vbias.n2094 455.736
R5884 Vbias.t805 Vbias.n2094 455.736
R5885 Vbias.t805 Vbias.n2096 455.736
R5886 Vbias.n2096 Vbias.t857 455.736
R5887 Vbias.t682 Vbias.n5802 455.736
R5888 Vbias.t682 Vbias.n5791 455.736
R5889 Vbias.t401 Vbias.n5791 455.736
R5890 Vbias.t401 Vbias.n5796 455.736
R5891 Vbias.n5795 Vbias.t106 455.736
R5892 Vbias.t106 Vbias.n2080 455.736
R5893 Vbias.t648 Vbias.n2080 455.736
R5894 Vbias.t648 Vbias.n2074 455.736
R5895 Vbias.t494 Vbias.n2074 455.736
R5896 Vbias.t494 Vbias.n667 455.736
R5897 Vbias.t784 Vbias.n678 455.736
R5898 Vbias.n5837 Vbias.t784 455.736
R5899 Vbias.t202 Vbias.n2068 455.736
R5900 Vbias.t202 Vbias.n1693 455.736
R5901 Vbias.t712 Vbias.n1694 455.736
R5902 Vbias.t392 Vbias.n1694 455.736
R5903 Vbias.t392 Vbias.n2060 455.736
R5904 Vbias.n2059 Vbias.t30 455.736
R5905 Vbias.t30 Vbias.n1530 455.736
R5906 Vbias.n8007 Vbias.t791 455.736
R5907 Vbias.n8001 Vbias.t791 455.736
R5908 Vbias.n8000 Vbias.t257 455.736
R5909 Vbias.n97 Vbias.t257 455.736
R5910 Vbias.t790 Vbias.n97 455.736
R5911 Vbias.t790 Vbias.n98 455.736
R5912 Vbias.t813 Vbias.n98 455.736
R5913 Vbias.t813 Vbias.n7986 455.736
R5914 Vbias.n7985 Vbias.t46 455.736
R5915 Vbias.t288 Vbias.n116 455.736
R5916 Vbias.t288 Vbias.n117 455.736
R5917 Vbias.t538 Vbias.n117 455.736
R5918 Vbias.t538 Vbias.n7971 455.736
R5919 Vbias.n7970 Vbias.t356 455.736
R5920 Vbias.n137 Vbias.t356 455.736
R5921 Vbias.t858 Vbias.n137 455.736
R5922 Vbias.t858 Vbias.n138 455.736
R5923 Vbias.t20 Vbias.n157 455.736
R5924 Vbias.t20 Vbias.n151 455.736
R5925 Vbias.t801 Vbias.n151 455.736
R5926 Vbias.t801 Vbias.n152 455.736
R5927 Vbias.t518 Vbias.n152 455.736
R5928 Vbias.t518 Vbias.n165 455.736
R5929 Vbias.n6750 Vbias.n1444 416.842
R5930 Vbias.n6736 Vbias.n821 416.842
R5931 Vbias.n7494 Vbias.n976 416.842
R5932 Vbias.n821 Vbias.n808 393.084
R5933 Vbias.n1305 Vbias.n1304 372.848
R5934 Vbias.n5533 Vbias.n5508 372.848
R5935 Vbias.n5011 Vbias.n2592 372.848
R5936 Vbias.t322 Vbias.n5553 372.606
R5937 Vbias.n5877 Vbias.t857 372.606
R5938 Vbias.n4902 Vbias.n4846 359
R5939 Vbias.n5858 Vbias.t712 356.276
R5940 Vbias.t573 Vbias.n6 349.135
R5941 Vbias.t573 Vbias.n4107 349.135
R5942 Vbias.t528 Vbias.n3985 349.135
R5943 Vbias.t528 Vbias.n3988 349.135
R5944 Vbias.t286 Vbias.n3988 349.135
R5945 Vbias.t286 Vbias.n3996 349.135
R5946 Vbias.t131 Vbias.n3996 349.135
R5947 Vbias.t131 Vbias.n4235 349.135
R5948 Vbias.n4234 Vbias.t82 349.135
R5949 Vbias.n4016 Vbias.t82 349.135
R5950 Vbias.t163 Vbias.n4016 349.135
R5951 Vbias.t163 Vbias.n4019 349.135
R5952 Vbias.t296 Vbias.n4019 349.135
R5953 Vbias.t296 Vbias.n4219 349.135
R5954 Vbias.n4218 Vbias.t503 349.135
R5955 Vbias.n4151 Vbias.t503 349.135
R5956 Vbias.n4155 Vbias.t289 349.135
R5957 Vbias.n4207 Vbias.t289 349.135
R5958 Vbias.n4207 Vbias.t467 349.135
R5959 Vbias.t467 Vbias.n4201 349.135
R5960 Vbias.n4200 Vbias.t36 349.135
R5961 Vbias.n4058 Vbias.t36 349.135
R5962 Vbias.t10 Vbias.n4058 349.135
R5963 Vbias.t10 Vbias.n4061 349.135
R5964 Vbias.t783 Vbias.n4061 349.135
R5965 Vbias.t783 Vbias.n2772 349.135
R5966 Vbias.t669 Vbias.n7226 348.704
R5967 Vbias.n2039 Vbias.t341 336.942
R5968 Vbias.t341 Vbias.n1467 336.942
R5969 Vbias.n3701 Vbias.n3700 326.113
R5970 Vbias.n3663 Vbias.n3662 326.113
R5971 Vbias.n3625 Vbias.n3624 326.113
R5972 Vbias.n3598 Vbias.n3593 326.113
R5973 Vbias.n3587 Vbias.n3586 326.113
R5974 Vbias.n3432 Vbias.n3431 326.113
R5975 Vbias.n3394 Vbias.n3393 326.113
R5976 Vbias.n3356 Vbias.n3355 326.113
R5977 Vbias.n3329 Vbias.n3324 326.113
R5978 Vbias.n3318 Vbias.n3317 326.113
R5979 Vbias.n3970 Vbias.n3969 326.113
R5980 Vbias.n3932 Vbias.n3931 326.113
R5981 Vbias.n3894 Vbias.n3893 326.113
R5982 Vbias.n3867 Vbias.n3862 326.113
R5983 Vbias.n3856 Vbias.n3855 326.113
R5984 Vbias.n3162 Vbias.n3161 326.113
R5985 Vbias.n3124 Vbias.n3123 326.113
R5986 Vbias.n3086 Vbias.n3085 326.113
R5987 Vbias.n3059 Vbias.n3054 326.113
R5988 Vbias.n3048 Vbias.n3047 326.113
R5989 Vbias.n4838 Vbias.n4837 326.113
R5990 Vbias.n4800 Vbias.n4799 326.113
R5991 Vbias.n4762 Vbias.n4761 326.113
R5992 Vbias.n4735 Vbias.n4730 326.113
R5993 Vbias.n4724 Vbias.n4723 326.113
R5994 Vbias.n4262 Vbias.n2883 326.113
R5995 Vbias.n2868 Vbias.n2849 326.113
R5996 Vbias.n2834 Vbias.n2833 326.113
R5997 Vbias.n4343 Vbias.n4338 326.113
R5998 Vbias.n4365 Vbias.n4364 326.113
R5999 Vbias.n5010 Vbias.n116 311.741
R6000 Vbias.n7017 Vbias.n7016 306.584
R6001 Vbias.n5920 Vbias.n5919 306.584
R6002 Vbias.n5123 Vbias.n5122 306.584
R6003 Vbias.n4682 Vbias.n4681 306.584
R6004 Vbias.n7226 Vbias.n1058 300.096
R6005 Vbias.n6679 Vbias.n6678 290.815
R6006 Vbias.n348 Vbias.t621 281.065
R6007 Vbias.n342 Vbias.t621 281.065
R6008 Vbias.n341 Vbias.t440 281.065
R6009 Vbias.n332 Vbias.t440 281.065
R6010 Vbias.n332 Vbias.t811 281.065
R6011 Vbias.n7938 Vbias.t811 281.065
R6012 Vbias.n7886 Vbias.t3 281.065
R6013 Vbias.n456 Vbias.t3 281.065
R6014 Vbias.t767 Vbias.n456 281.065
R6015 Vbias.t767 Vbias.n7872 281.065
R6016 Vbias.n7820 Vbias.t628 281.065
R6017 Vbias.n566 Vbias.t628 281.065
R6018 Vbias.t850 Vbias.n567 281.065
R6019 Vbias.n7809 Vbias.t850 281.065
R6020 Vbias.n7809 Vbias.t485 281.065
R6021 Vbias.t485 Vbias.n7803 281.065
R6022 Vbias.n7751 Vbias.t820 281.065
R6023 Vbias.n677 Vbias.t820 281.065
R6024 Vbias.t713 Vbias.n677 281.065
R6025 Vbias.t713 Vbias.n7737 281.065
R6026 Vbias.n5534 Vbias.n2165 276.113
R6027 Vbias.n8075 Vbias.t158 275.505
R6028 Vbias.n19 Vbias.t158 275.505
R6029 Vbias.t631 Vbias.n19 275.505
R6030 Vbias.t631 Vbias.n20 275.505
R6031 Vbias.t313 Vbias.n20 275.505
R6032 Vbias.t313 Vbias.n29 275.505
R6033 Vbias.t674 Vbias.n37 275.505
R6034 Vbias.n8054 Vbias.t674 275.505
R6035 Vbias.n8054 Vbias.t360 275.505
R6036 Vbias.t360 Vbias.n41 275.505
R6037 Vbias.t798 Vbias.n41 275.505
R6038 Vbias.t798 Vbias.n47 275.505
R6039 Vbias.t323 Vbias.n56 275.505
R6040 Vbias.n8040 Vbias.t323 275.505
R6041 Vbias.n8039 Vbias.t418 275.505
R6042 Vbias.n65 Vbias.t418 275.505
R6043 Vbias.t307 Vbias.n65 275.505
R6044 Vbias.t307 Vbias.n8025 275.505
R6045 Vbias.n8024 Vbias.t522 275.505
R6046 Vbias.n75 Vbias.t522 275.505
R6047 Vbias.t533 Vbias.n75 275.505
R6048 Vbias.t533 Vbias.n76 275.505
R6049 Vbias.t694 Vbias.n76 275.505
R6050 Vbias.t694 Vbias.n8009 275.505
R6051 Vbias.t795 Vbias.n1765 274.82
R6052 Vbias.t317 Vbias.n1767 274.82
R6053 Vbias.t560 Vbias.n1759 274.82
R6054 Vbias.t414 Vbias.n1760 274.82
R6055 Vbias.n1476 Vbias.n1459 274.736
R6056 Vbias.n1504 Vbias.n756 274.736
R6057 Vbias.n6308 Vbias.n6307 274.736
R6058 Vbias.n6285 Vbias.n6284 274.736
R6059 Vbias.n6353 Vbias.n6352 274.736
R6060 Vbias.n7645 Vbias.n7644 274.736
R6061 Vbias.n7630 Vbias.n7629 274.736
R6062 Vbias.n849 Vbias.n830 274.736
R6063 Vbias.n6518 Vbias.n6517 274.736
R6064 Vbias.n7524 Vbias.n7523 274.736
R6065 Vbias.n7509 Vbias.n7508 274.736
R6066 Vbias.n1004 Vbias.n985 274.736
R6067 Vbias.n7317 Vbias.n7316 274.736
R6068 Vbias.n7302 Vbias.n7301 274.736
R6069 Vbias.n7254 Vbias.n7235 274.736
R6070 Vbias.n7143 Vbias.n7142 260.592
R6071 Vbias.n7161 Vbias.n7159 260.592
R6072 Vbias.n7162 Vbias.n1116 260.592
R6073 Vbias.n7179 Vbias.n1097 260.592
R6074 Vbias.n7037 Vbias.n7036 260.592
R6075 Vbias.n7055 Vbias.n7053 260.592
R6076 Vbias.n7056 Vbias.n1303 260.592
R6077 Vbias.n7073 Vbias.n1284 260.592
R6078 Vbias.n6061 Vbias.n6060 260.592
R6079 Vbias.n6799 Vbias.n6798 260.592
R6080 Vbias.n6754 Vbias.n6753 260.592
R6081 Vbias.n6771 Vbias.n6770 260.592
R6082 Vbias.n1790 Vbias.n1789 260.592
R6083 Vbias.n5933 Vbias.n5932 260.592
R6084 Vbias.n6100 Vbias.n1532 260.592
R6085 Vbias.n5473 Vbias.n5472 260.592
R6086 Vbias.n5463 Vbias.n5462 260.592
R6087 Vbias.n5454 Vbias.n1672 260.592
R6088 Vbias.n5898 Vbias.n5897 260.592
R6089 Vbias.n5140 Vbias.n5139 260.592
R6090 Vbias.n5168 Vbias.n5167 260.592
R6091 Vbias.n5158 Vbias.n5157 260.592
R6092 Vbias.n5498 Vbias.n5497 260.592
R6093 Vbias.n5058 Vbias.n5057 260.592
R6094 Vbias.n5068 Vbias.n5067 260.592
R6095 Vbias.n5080 Vbias.n5079 260.592
R6096 Vbias.n5101 Vbias.n5100 260.592
R6097 Vbias.n4671 Vbias.n4670 260.592
R6098 Vbias.n4661 Vbias.n4660 260.592
R6099 Vbias.n4618 Vbias.n4617 260.592
R6100 Vbias.n4633 Vbias.n4632 260.592
R6101 Vbias.n6101 Vbias.n1528 260.257
R6102 Vbias.t346 Vbias.n821 255.716
R6103 Vbias.n6677 Vbias.n6676 246.612
R6104 Vbias.t715 Vbias.n1305 242.552
R6105 Vbias.n5533 Vbias.t666 242.552
R6106 Vbias.n5011 Vbias.t285 242.552
R6107 Vbias.n5859 Vbias.n5858 242.542
R6108 Vbias.n8013 Vbias.n84 236.048
R6109 Vbias.n8022 Vbias.n68 236.048
R6110 Vbias.n8030 Vbias.n62 236.048
R6111 Vbias.n8037 Vbias.n59 236.048
R6112 Vbias.n8042 Vbias.n53 236.048
R6113 Vbias.n53 Vbias.n51 236.048
R6114 Vbias.n8050 Vbias.n45 236.048
R6115 Vbias.n39 Vbias.n31 236.048
R6116 Vbias.n4371 Vbias.n2800 236.048
R6117 Vbias.n4404 Vbias.n2780 236.048
R6118 Vbias.n4402 Vbias.n4401 236.048
R6119 Vbias.n4368 Vbias.n4367 236.048
R6120 Vbias.n4362 Vbias.n2805 236.048
R6121 Vbias.n4346 Vbias.n2819 236.048
R6122 Vbias.n4348 Vbias.n2806 236.048
R6123 Vbias.n4341 Vbias.n4340 236.048
R6124 Vbias.n4336 Vbias.n2822 236.048
R6125 Vbias.n2823 Vbias.n2822 236.048
R6126 Vbias.n4308 Vbias.n2846 236.048
R6127 Vbias.n4328 Vbias.n4327 236.048
R6128 Vbias.n4313 Vbias.n4312 236.048
R6129 Vbias.n4305 Vbias.n4304 236.048
R6130 Vbias.n4275 Vbias.n2880 236.048
R6131 Vbias.n4295 Vbias.n4294 236.048
R6132 Vbias.n4280 Vbias.n4279 236.048
R6133 Vbias.n4272 Vbias.n4271 236.048
R6134 Vbias.n4264 Vbias.n4258 236.048
R6135 Vbias.n4258 Vbias.n4256 236.048
R6136 Vbias.n5007 Vbias.n2595 236.048
R6137 Vbias.n4999 Vbias.n2597 236.048
R6138 Vbias.n4990 Vbias.n2602 236.048
R6139 Vbias.n2603 Vbias.n2602 236.048
R6140 Vbias.n6712 Vbias.n6699 236.048
R6141 Vbias.n6704 Vbias.n6695 236.048
R6142 Vbias.n6739 Vbias.n6723 236.048
R6143 Vbias.n6730 Vbias.n6719 236.048
R6144 Vbias.n1448 Vbias.n1447 236.048
R6145 Vbias.n6747 Vbias.n1447 236.048
R6146 Vbias.n7742 Vbias.n674 236.048
R6147 Vbias.n7749 Vbias.n670 236.048
R6148 Vbias.n7807 Vbias.n7806 236.048
R6149 Vbias.n569 Vbias.n559 236.048
R6150 Vbias.n557 Vbias.n556 236.048
R6151 Vbias.n7818 Vbias.n556 236.048
R6152 Vbias.n7877 Vbias.n453 236.048
R6153 Vbias.n7884 Vbias.n450 236.048
R6154 Vbias.n7940 Vbias.n172 236.048
R6155 Vbias.n339 Vbias.n336 236.048
R6156 Vbias.n1023 Vbias.n923 236.048
R6157 Vbias.n1015 Vbias.n1014 236.048
R6158 Vbias.n7533 Vbias.n927 236.048
R6159 Vbias.n6529 Vbias.n6524 236.048
R6160 Vbias.n6515 Vbias.n6507 236.048
R6161 Vbias.n6510 Vbias.n6507 236.048
R6162 Vbias.n7654 Vbias.n776 236.048
R6163 Vbias.n6593 Vbias.n772 236.048
R6164 Vbias.n7664 Vbias.n763 236.048
R6165 Vbias.n7666 Vbias.n761 236.048
R6166 Vbias.n7673 Vbias.n753 236.048
R6167 Vbias.n7682 Vbias.n737 236.048
R6168 Vbias.n7690 Vbias.n731 236.048
R6169 Vbias.n7697 Vbias.n728 236.048
R6170 Vbias.n7702 Vbias.n722 236.048
R6171 Vbias.n722 Vbias.n720 236.048
R6172 Vbias.n7710 Vbias.n714 236.048
R6173 Vbias.n708 Vbias.n700 236.048
R6174 Vbias.n7755 Vbias.n652 236.048
R6175 Vbias.n7762 Vbias.n645 236.048
R6176 Vbias.n7767 Vbias.n630 236.048
R6177 Vbias.n637 Vbias.n626 236.048
R6178 Vbias.n623 Vbias.n622 236.048
R6179 Vbias.n7775 Vbias.n622 236.048
R6180 Vbias.n7780 Vbias.n605 236.048
R6181 Vbias.n7787 Vbias.n598 236.048
R6182 Vbias.n7792 Vbias.n581 236.048
R6183 Vbias.n7799 Vbias.n574 236.048
R6184 Vbias.n7824 Vbias.n538 236.048
R6185 Vbias.n7831 Vbias.n531 236.048
R6186 Vbias.n7836 Vbias.n516 236.048
R6187 Vbias.n523 Vbias.n512 236.048
R6188 Vbias.n509 Vbias.n508 236.048
R6189 Vbias.n7844 Vbias.n508 236.048
R6190 Vbias.n7849 Vbias.n491 236.048
R6191 Vbias.n7856 Vbias.n484 236.048
R6192 Vbias.n7861 Vbias.n467 236.048
R6193 Vbias.n7868 Vbias.n460 236.048
R6194 Vbias.n7890 Vbias.n432 236.048
R6195 Vbias.n7897 Vbias.n425 236.048
R6196 Vbias.n7902 Vbias.n410 236.048
R6197 Vbias.n417 Vbias.n406 236.048
R6198 Vbias.n403 Vbias.n402 236.048
R6199 Vbias.n7910 Vbias.n402 236.048
R6200 Vbias.n7915 Vbias.n385 236.048
R6201 Vbias.n7922 Vbias.n378 236.048
R6202 Vbias.n7927 Vbias.n361 236.048
R6203 Vbias.n7934 Vbias.n177 236.048
R6204 Vbias.n352 Vbias.n182 236.048
R6205 Vbias.n193 Vbias.n189 236.048
R6206 Vbias.n309 Vbias.n201 236.048
R6207 Vbias.n302 Vbias.n205 236.048
R6208 Vbias.n296 Vbias.n210 236.048
R6209 Vbias.n211 Vbias.n210 236.048
R6210 Vbias.n289 Vbias.n215 236.048
R6211 Vbias.n226 Vbias.n222 236.048
R6212 Vbias.n270 Vbias.n234 236.048
R6213 Vbias.n244 Vbias.n241 236.048
R6214 Vbias.n7951 Vbias.n163 236.048
R6215 Vbias.n159 Vbias.n145 236.048
R6216 Vbias.n7965 Vbias.n134 236.048
R6217 Vbias.n7968 Vbias.n7967 236.048
R6218 Vbias.n7972 Vbias.n128 236.048
R6219 Vbias.n7983 Vbias.n7982 236.048
R6220 Vbias.n7987 Vbias.n107 236.048
R6221 Vbias.n7998 Vbias.n7997 236.048
R6222 Vbias.n8004 Vbias.n8003 236.048
R6223 Vbias.n8005 Vbias.n8004 236.048
R6224 Vbias.n5034 Vbias.n2436 236.048
R6225 Vbias.n4635 Vbias.n4601 236.048
R6226 Vbias.n4629 Vbias.n4600 236.048
R6227 Vbias.n4620 Vbias.n4594 236.048
R6228 Vbias.n4592 Vbias.n4591 236.048
R6229 Vbias.n4658 Vbias.n4591 236.048
R6230 Vbias.n4663 Vbias.n4581 236.048
R6231 Vbias.n4668 Vbias.n4576 236.048
R6232 Vbias.n4493 Vbias.n4487 236.048
R6233 Vbias.n4487 Vbias.n4485 236.048
R6234 Vbias.n4501 Vbias.n4480 236.048
R6235 Vbias.n4476 Vbias.n4462 236.048
R6236 Vbias.n4515 Vbias.n4458 236.048
R6237 Vbias.n4454 Vbias.n4440 236.048
R6238 Vbias.n4529 Vbias.n4430 236.048
R6239 Vbias.n4532 Vbias.n4531 236.048
R6240 Vbias.n5118 Vbias.n2374 236.048
R6241 Vbias.n5105 Vbias.n2386 236.048
R6242 Vbias.n5098 Vbias.n2390 236.048
R6243 Vbias.n5085 Vbias.n2402 236.048
R6244 Vbias.n5077 Vbias.n2405 236.048
R6245 Vbias.n2406 Vbias.n2405 236.048
R6246 Vbias.n5070 Vbias.n2410 236.048
R6247 Vbias.n5061 Vbias.n2414 236.048
R6248 Vbias.n5488 Vbias.n2273 236.048
R6249 Vbias.n5495 Vbias.n2267 236.048
R6250 Vbias.n5500 Vbias.n2255 236.048
R6251 Vbias.n5155 Vbias.n5154 236.048
R6252 Vbias.n5160 Vbias.n5151 236.048
R6253 Vbias.n5165 Vbias.n5151 236.048
R6254 Vbias.n5170 Vbias.n2362 236.048
R6255 Vbias.n5143 Vbias.n2358 236.048
R6256 Vbias.n5136 Vbias.n2356 236.048
R6257 Vbias.n5125 Vbias.n2350 236.048
R6258 Vbias.n5915 Vbias.n1642 236.048
R6259 Vbias.n5902 Vbias.n1654 236.048
R6260 Vbias.n5895 Vbias.n1658 236.048
R6261 Vbias.n5882 Vbias.n1670 236.048
R6262 Vbias.n5456 Vbias.n5453 236.048
R6263 Vbias.n5460 Vbias.n5453 236.048
R6264 Vbias.n5465 Vbias.n5443 236.048
R6265 Vbias.n5470 Vbias.n5438 236.048
R6266 Vbias.n5475 Vbias.n5421 236.048
R6267 Vbias.n5482 Vbias.n2291 236.048
R6268 Vbias.n5943 Vbias.n1626 236.048
R6269 Vbias.n5936 Vbias.n1622 236.048
R6270 Vbias.n1629 Vbias.n1619 236.048
R6271 Vbias.n5922 Vbias.n1613 236.048
R6272 Vbias.n1536 Vbias.n1535 236.048
R6273 Vbias.n6098 Vbias.n1535 236.048
R6274 Vbias.n6105 Vbias.n1521 236.048
R6275 Vbias.n6114 Vbias.n6107 236.048
R6276 Vbias.n1996 Vbias.n1993 236.048
R6277 Vbias.n2013 Vbias.n1987 236.048
R6278 Vbias.n1965 Vbias.n1961 236.048
R6279 Vbias.n1974 Vbias.n1967 236.048
R6280 Vbias.n1931 Vbias.n1927 236.048
R6281 Vbias.n1940 Vbias.n1933 236.048
R6282 Vbias.n1816 Vbias.n1756 236.048
R6283 Vbias.n1808 Vbias.n1807 236.048
R6284 Vbias.n1874 Vbias.n1867 236.048
R6285 Vbias.n1863 Vbias.n1859 236.048
R6286 Vbias.n2036 Vbias.n1730 236.048
R6287 Vbias.n1737 Vbias.n1736 236.048
R6288 Vbias.n1910 Vbias.n1883 236.048
R6289 Vbias.n1902 Vbias.n1901 236.048
R6290 Vbias.n6078 Vbias.n1552 236.048
R6291 Vbias.n1786 Vbias.n1546 236.048
R6292 Vbias.n1792 Vbias.n1544 236.048
R6293 Vbias.n1798 Vbias.n1538 236.048
R6294 Vbias.n7012 Vbias.n1343 236.048
R6295 Vbias.n6773 Vbias.n1429 236.048
R6296 Vbias.n6767 Vbias.n1428 236.048
R6297 Vbias.n6756 Vbias.n1422 236.048
R6298 Vbias.n1419 Vbias.n1418 236.048
R6299 Vbias.n6796 Vbias.n1418 236.048
R6300 Vbias.n6801 Vbias.n1414 236.048
R6301 Vbias.n6057 Vbias.n1410 236.048
R6302 Vbias.n6063 Vbias.n1408 236.048
R6303 Vbias.n6071 Vbias.n1402 236.048
R6304 Vbias.n7092 Vbias.n1277 236.048
R6305 Vbias.n1287 Vbias.n1283 236.048
R6306 Vbias.n7075 Vbias.n1295 236.048
R6307 Vbias.n1307 Vbias.n1302 236.048
R6308 Vbias.n7058 Vbias.n1314 236.048
R6309 Vbias.n1314 Vbias.n1312 236.048
R6310 Vbias.n7051 Vbias.n1318 236.048
R6311 Vbias.n7043 Vbias.n1320 236.048
R6312 Vbias.n7034 Vbias.n1325 236.048
R6313 Vbias.n7021 Vbias.n1337 236.048
R6314 Vbias.n7198 Vbias.n1090 236.048
R6315 Vbias.n1100 Vbias.n1096 236.048
R6316 Vbias.n7181 Vbias.n1108 236.048
R6317 Vbias.n1119 Vbias.n1115 236.048
R6318 Vbias.n7164 Vbias.n1126 236.048
R6319 Vbias.n1126 Vbias.n1124 236.048
R6320 Vbias.n7157 Vbias.n1130 236.048
R6321 Vbias.n7149 Vbias.n1132 236.048
R6322 Vbias.n7140 Vbias.n1137 236.048
R6323 Vbias.n7127 Vbias.n1149 236.048
R6324 Vbias.n7222 Vbias.n7221 236.048
R6325 Vbias.n7221 Vbias.n7220 236.048
R6326 Vbias.n1222 Vbias.n1221 236.048
R6327 Vbias.n7215 Vbias.n7214 236.048
R6328 Vbias.n1205 Vbias.n1197 236.048
R6329 Vbias.n1232 Vbias.n1231 236.048
R6330 Vbias.n1253 Vbias.n1252 236.048
R6331 Vbias.n1245 Vbias.n1186 236.048
R6332 Vbias.n1176 Vbias.n1169 236.048
R6333 Vbias.n1263 Vbias.n1262 236.048
R6334 Vbias.n7118 Vbias.n7117 236.048
R6335 Vbias.n7117 Vbias.n7116 236.048
R6336 Vbias.n6955 Vbias.n6954 236.048
R6337 Vbias.n7111 Vbias.n7110 236.048
R6338 Vbias.n6938 Vbias.n6930 236.048
R6339 Vbias.n6965 Vbias.n6964 236.048
R6340 Vbias.n6986 Vbias.n6985 236.048
R6341 Vbias.n6978 Vbias.n6919 236.048
R6342 Vbias.n6909 Vbias.n6902 236.048
R6343 Vbias.n6996 Vbias.n6995 236.048
R6344 Vbias.n6894 Vbias.n1347 236.048
R6345 Vbias.n6894 Vbias.n1346 236.048
R6346 Vbias.n6875 Vbias.n1361 236.048
R6347 Vbias.n6890 Vbias.n6889 236.048
R6348 Vbias.n6852 Vbias.n1374 236.048
R6349 Vbias.n6867 Vbias.n6866 236.048
R6350 Vbias.n1386 Vbias.n1379 236.048
R6351 Vbias.n6844 Vbias.n6843 236.048
R6352 Vbias.n1554 Vbias.n1399 236.048
R6353 Vbias.n6828 Vbias.n1389 236.048
R6354 Vbias.n6042 Vbias.n6041 236.048
R6355 Vbias.n6041 Vbias.n6040 236.048
R6356 Vbias.n6017 Vbias.n1572 236.048
R6357 Vbias.n6035 Vbias.n6034 236.048
R6358 Vbias.n5994 Vbias.n1585 236.048
R6359 Vbias.n6009 Vbias.n6008 236.048
R6360 Vbias.n1597 Vbias.n1590 236.048
R6361 Vbias.n5986 Vbias.n5985 236.048
R6362 Vbias.n1635 Vbias.n1610 236.048
R6363 Vbias.n5970 Vbias.n1600 236.048
R6364 Vbias.n5346 Vbias.n5345 236.048
R6365 Vbias.n5347 Vbias.n5346 236.048
R6366 Vbias.n5363 Vbias.n5362 236.048
R6367 Vbias.n5351 Vbias.n5336 236.048
R6368 Vbias.n5309 Vbias.n5301 236.048
R6369 Vbias.n5373 Vbias.n5372 236.048
R6370 Vbias.n5394 Vbias.n5393 236.048
R6371 Vbias.n5386 Vbias.n5290 236.048
R6372 Vbias.n5280 Vbias.n5272 236.048
R6373 Vbias.n5404 Vbias.n5403 236.048
R6374 Vbias.n5264 Vbias.n2295 236.048
R6375 Vbias.n5264 Vbias.n2294 236.048
R6376 Vbias.n5244 Vbias.n2309 236.048
R6377 Vbias.n5259 Vbias.n5258 236.048
R6378 Vbias.n5221 Vbias.n2322 236.048
R6379 Vbias.n5236 Vbias.n5235 236.048
R6380 Vbias.n2334 Vbias.n2327 236.048
R6381 Vbias.n5213 Vbias.n5212 236.048
R6382 Vbias.n2367 Vbias.n2347 236.048
R6383 Vbias.n5197 Vbias.n2337 236.048
R6384 Vbias.n2514 Vbias.n2513 236.048
R6385 Vbias.n2515 Vbias.n2514 236.048
R6386 Vbias.n2531 Vbias.n2530 236.048
R6387 Vbias.n2519 Vbias.n2504 236.048
R6388 Vbias.n2477 Vbias.n2469 236.048
R6389 Vbias.n2541 Vbias.n2540 236.048
R6390 Vbias.n2562 Vbias.n2561 236.048
R6391 Vbias.n2554 Vbias.n2458 236.048
R6392 Vbias.n2448 Vbias.n2440 236.048
R6393 Vbias.n2572 Vbias.n2571 236.048
R6394 Vbias.n5055 Vbias.n2419 236.048
R6395 Vbias.n5042 Vbias.n2431 236.048
R6396 Vbias.n4548 Vbias.n4547 236.048
R6397 Vbias.n4536 Vbias.n4424 236.048
R6398 Vbias.n3827 Vbias.n3794 236.048
R6399 Vbias.n3843 Vbias.n3815 236.048
R6400 Vbias.n3838 Vbias.n3836 236.048
R6401 Vbias.n3853 Vbias.n3793 236.048
R6402 Vbias.n3879 Vbias.n3878 236.048
R6403 Vbias.n3871 Vbias.n3860 236.048
R6404 Vbias.n3875 Vbias.n3873 236.048
R6405 Vbias.n3865 Vbias.n3864 236.048
R6406 Vbias.n3775 Vbias.n3774 236.048
R6407 Vbias.n3891 Vbias.n3774 236.048
R6408 Vbias.n3903 Vbias.n3747 236.048
R6409 Vbias.n3919 Vbias.n3768 236.048
R6410 Vbias.n3914 Vbias.n3912 236.048
R6411 Vbias.n3929 Vbias.n3746 236.048
R6412 Vbias.n3941 Vbias.n3718 236.048
R6413 Vbias.n3957 Vbias.n3739 236.048
R6414 Vbias.n3952 Vbias.n3950 236.048
R6415 Vbias.n3967 Vbias.n3717 236.048
R6416 Vbias.n3971 Vbias.n3711 236.048
R6417 Vbias.n3971 Vbias.n3710 236.048
R6418 Vbias.n3289 Vbias.n3256 236.048
R6419 Vbias.n3305 Vbias.n3277 236.048
R6420 Vbias.n3300 Vbias.n3298 236.048
R6421 Vbias.n3315 Vbias.n3255 236.048
R6422 Vbias.n3341 Vbias.n3340 236.048
R6423 Vbias.n3333 Vbias.n3322 236.048
R6424 Vbias.n3337 Vbias.n3335 236.048
R6425 Vbias.n3327 Vbias.n3326 236.048
R6426 Vbias.n3237 Vbias.n3236 236.048
R6427 Vbias.n3353 Vbias.n3236 236.048
R6428 Vbias.n3365 Vbias.n3209 236.048
R6429 Vbias.n3381 Vbias.n3230 236.048
R6430 Vbias.n3376 Vbias.n3374 236.048
R6431 Vbias.n3391 Vbias.n3208 236.048
R6432 Vbias.n3403 Vbias.n3180 236.048
R6433 Vbias.n3419 Vbias.n3201 236.048
R6434 Vbias.n3414 Vbias.n3412 236.048
R6435 Vbias.n3429 Vbias.n3179 236.048
R6436 Vbias.n3433 Vbias.n3173 236.048
R6437 Vbias.n3433 Vbias.n3172 236.048
R6438 Vbias.n3558 Vbias.n3525 236.048
R6439 Vbias.n3574 Vbias.n3546 236.048
R6440 Vbias.n3569 Vbias.n3567 236.048
R6441 Vbias.n3584 Vbias.n3524 236.048
R6442 Vbias.n3610 Vbias.n3609 236.048
R6443 Vbias.n3602 Vbias.n3591 236.048
R6444 Vbias.n3606 Vbias.n3604 236.048
R6445 Vbias.n3596 Vbias.n3595 236.048
R6446 Vbias.n3506 Vbias.n3505 236.048
R6447 Vbias.n3622 Vbias.n3505 236.048
R6448 Vbias.n3634 Vbias.n3478 236.048
R6449 Vbias.n3650 Vbias.n3499 236.048
R6450 Vbias.n3645 Vbias.n3643 236.048
R6451 Vbias.n3660 Vbias.n3477 236.048
R6452 Vbias.n3672 Vbias.n3449 236.048
R6453 Vbias.n3688 Vbias.n3470 236.048
R6454 Vbias.n3683 Vbias.n3681 236.048
R6455 Vbias.n3698 Vbias.n3448 236.048
R6456 Vbias.n3702 Vbias.n3442 236.048
R6457 Vbias.n3702 Vbias.n3441 236.048
R6458 Vbias.n4189 Vbias.n4069 236.048
R6459 Vbias.n4198 Vbias.n4051 236.048
R6460 Vbias.n4205 Vbias.n4204 236.048
R6461 Vbias.n4152 Vbias.n4038 236.048
R6462 Vbias.n4035 Vbias.n4034 236.048
R6463 Vbias.n4216 Vbias.n4034 236.048
R6464 Vbias.n4223 Vbias.n4027 236.048
R6465 Vbias.n4232 Vbias.n4009 236.048
R6466 Vbias.n4236 Vbias.n4001 236.048
R6467 Vbias.n4246 Vbias.n3981 236.048
R6468 Vbias.n4184 Vbias.n4183 236.048
R6469 Vbias.n4171 Vbias.n4168 236.048
R6470 Vbias.n4162 Vbias.n4161 236.048
R6471 Vbias.n4159 Vbias.n4146 236.048
R6472 Vbias.n4139 Vbias.n4138 236.048
R6473 Vbias.n4134 Vbias.n4086 236.048
R6474 Vbias.n4123 Vbias.n4122 236.048
R6475 Vbias.n4118 Vbias.n4117 236.048
R6476 Vbias.n4108 Vbias.n4104 236.048
R6477 Vbias.n4108 Vbias.n4103 236.048
R6478 Vbias.n2624 Vbias.n2616 236.048
R6479 Vbias.n4982 Vbias.n2606 236.048
R6480 Vbias.n4960 Vbias.n2630 236.048
R6481 Vbias.n4964 Vbias.n2620 236.048
R6482 Vbias.n4938 Vbias.n2644 236.048
R6483 Vbias.n4953 Vbias.n4952 236.048
R6484 Vbias.n4916 Vbias.n2658 236.048
R6485 Vbias.n4930 Vbias.n4929 236.048
R6486 Vbias.n4908 Vbias.n4907 236.048
R6487 Vbias.n4907 Vbias.n4906 236.048
R6488 Vbias.n3019 Vbias.n2986 236.048
R6489 Vbias.n3035 Vbias.n3007 236.048
R6490 Vbias.n3030 Vbias.n3028 236.048
R6491 Vbias.n3045 Vbias.n2985 236.048
R6492 Vbias.n3071 Vbias.n3070 236.048
R6493 Vbias.n3063 Vbias.n3052 236.048
R6494 Vbias.n3067 Vbias.n3065 236.048
R6495 Vbias.n3057 Vbias.n3056 236.048
R6496 Vbias.n2967 Vbias.n2966 236.048
R6497 Vbias.n3083 Vbias.n2966 236.048
R6498 Vbias.n3095 Vbias.n2939 236.048
R6499 Vbias.n3111 Vbias.n2960 236.048
R6500 Vbias.n3106 Vbias.n3104 236.048
R6501 Vbias.n3121 Vbias.n2938 236.048
R6502 Vbias.n3133 Vbias.n2910 236.048
R6503 Vbias.n3149 Vbias.n2931 236.048
R6504 Vbias.n3144 Vbias.n3142 236.048
R6505 Vbias.n3159 Vbias.n2909 236.048
R6506 Vbias.n3163 Vbias.n2902 236.048
R6507 Vbias.n3163 Vbias.n2901 236.048
R6508 Vbias.n4695 Vbias.n2747 236.048
R6509 Vbias.n4711 Vbias.n2768 236.048
R6510 Vbias.n4706 Vbias.n4704 236.048
R6511 Vbias.n4721 Vbias.n2746 236.048
R6512 Vbias.n4747 Vbias.n4746 236.048
R6513 Vbias.n4739 Vbias.n4728 236.048
R6514 Vbias.n4743 Vbias.n4741 236.048
R6515 Vbias.n4733 Vbias.n4732 236.048
R6516 Vbias.n2728 Vbias.n2727 236.048
R6517 Vbias.n4759 Vbias.n2727 236.048
R6518 Vbias.n4771 Vbias.n2700 236.048
R6519 Vbias.n4787 Vbias.n2721 236.048
R6520 Vbias.n4782 Vbias.n4780 236.048
R6521 Vbias.n4797 Vbias.n2699 236.048
R6522 Vbias.n4809 Vbias.n2671 236.048
R6523 Vbias.n4825 Vbias.n2692 236.048
R6524 Vbias.n4820 Vbias.n4818 236.048
R6525 Vbias.n4835 Vbias.n2670 236.048
R6526 Vbias.n4841 Vbias.n4840 236.048
R6527 Vbias.n4842 Vbias.n4841 236.048
R6528 Vbias.n4673 Vbias.n4559 236.048
R6529 Vbias.n4679 Vbias.n4553 236.048
R6530 Vbias.n5659 Vbias.n2197 236.048
R6531 Vbias.n2218 Vbias.n2210 236.048
R6532 Vbias.n5645 Vbias.n2214 236.048
R6533 Vbias.n5643 Vbias.n2226 236.048
R6534 Vbias.n5636 Vbias.n5635 236.048
R6535 Vbias.n5621 Vbias.n5570 236.048
R6536 Vbias.n5617 Vbias.n5616 236.048
R6537 Vbias.n5603 Vbias.n5588 236.048
R6538 Vbias.n5599 Vbias.n5598 236.048
R6539 Vbias.n5598 Vbias.n5597 236.048
R6540 Vbias.n5733 Vbias.n2126 236.048
R6541 Vbias.n2147 Vbias.n2139 236.048
R6542 Vbias.n5719 Vbias.n2143 236.048
R6543 Vbias.n5717 Vbias.n2155 236.048
R6544 Vbias.n5710 Vbias.n5709 236.048
R6545 Vbias.n5695 Vbias.n2173 236.048
R6546 Vbias.n5691 Vbias.n5690 236.048
R6547 Vbias.n5677 Vbias.n2191 236.048
R6548 Vbias.n5673 Vbias.n5672 236.048
R6549 Vbias.n5672 Vbias.n5671 236.048
R6550 Vbias.n5822 Vbias.n2071 236.048
R6551 Vbias.n5792 Vbias.n2084 236.048
R6552 Vbias.n5808 Vbias.n5788 236.048
R6553 Vbias.n5806 Vbias.n5800 236.048
R6554 Vbias.n5779 Vbias.n2088 236.048
R6555 Vbias.n2108 Vbias.n2100 236.048
R6556 Vbias.n5765 Vbias.n2104 236.048
R6557 Vbias.n5747 Vbias.n2122 236.048
R6558 Vbias.n5753 Vbias.n5744 236.048
R6559 Vbias.n5744 Vbias.n5742 236.048
R6560 Vbias.n6656 Vbias.n1499 236.048
R6561 Vbias.n1495 Vbias.n1482 236.048
R6562 Vbias.n6670 Vbias.n1472 236.048
R6563 Vbias.n6673 Vbias.n6672 236.048
R6564 Vbias.n5851 Vbias.n1702 236.048
R6565 Vbias.n5847 Vbias.n2064 236.048
R6566 Vbias.n5839 Vbias.n5834 236.048
R6567 Vbias.n5834 Vbias.n5832 236.048
R6568 Vbias.n6587 Vbias.n6586 236.048
R6569 Vbias.n6354 Vbias.n6243 236.048
R6570 Vbias.n6350 Vbias.n6349 236.048
R6571 Vbias.n6347 Vbias.n6249 236.048
R6572 Vbias.n6336 Vbias.n6259 236.048
R6573 Vbias.n6281 Vbias.n6273 236.048
R6574 Vbias.n6322 Vbias.n6277 236.048
R6575 Vbias.n6304 Vbias.n6295 236.048
R6576 Vbias.n6310 Vbias.n6300 236.048
R6577 Vbias.n6300 Vbias.n6298 236.048
R6578 Vbias.n7595 Vbias.n855 236.048
R6579 Vbias.n851 Vbias.n837 236.048
R6580 Vbias.n7609 Vbias.n826 236.048
R6581 Vbias.n7612 Vbias.n7611 236.048
R6582 Vbias.n7616 Vbias.n819 236.048
R6583 Vbias.n7627 Vbias.n7626 236.048
R6584 Vbias.n7631 Vbias.n798 236.048
R6585 Vbias.n7642 Vbias.n7641 236.048
R6586 Vbias.n7648 Vbias.n7647 236.048
R6587 Vbias.n7649 Vbias.n7648 236.048
R6588 Vbias.n7473 Vbias.n1010 236.048
R6589 Vbias.n1006 Vbias.n992 236.048
R6590 Vbias.n7487 Vbias.n981 236.048
R6591 Vbias.n7490 Vbias.n7489 236.048
R6592 Vbias.n7495 Vbias.n974 236.048
R6593 Vbias.n7506 Vbias.n7505 236.048
R6594 Vbias.n7510 Vbias.n953 236.048
R6595 Vbias.n7521 Vbias.n7520 236.048
R6596 Vbias.n7527 Vbias.n7526 236.048
R6597 Vbias.n7528 Vbias.n7527 236.048
R6598 Vbias.n6601 Vbias.n6211 236.048
R6599 Vbias.n6608 Vbias.n6204 236.048
R6600 Vbias.n6613 Vbias.n6194 236.048
R6601 Vbias.n6618 Vbias.n6190 236.048
R6602 Vbias.n6623 Vbias.n6164 236.048
R6603 Vbias.n6164 Vbias.n6162 236.048
R6604 Vbias.n6182 Vbias.n6161 236.048
R6605 Vbias.n6171 Vbias.n6155 236.048
R6606 Vbias.n6534 Vbias.n6448 236.048
R6607 Vbias.n6541 Vbias.n6441 236.048
R6608 Vbias.n6546 Vbias.n6431 236.048
R6609 Vbias.n6551 Vbias.n6427 236.048
R6610 Vbias.n6556 Vbias.n6382 236.048
R6611 Vbias.n6382 Vbias.n6380 236.048
R6612 Vbias.n6419 Vbias.n6379 236.048
R6613 Vbias.n6408 Vbias.n6373 236.048
R6614 Vbias.n6402 Vbias.n6371 236.048
R6615 Vbias.n6391 Vbias.n6365 236.048
R6616 Vbias.n7547 Vbias.n902 236.048
R6617 Vbias.n7554 Vbias.n895 236.048
R6618 Vbias.n7559 Vbias.n885 236.048
R6619 Vbias.n7564 Vbias.n881 236.048
R6620 Vbias.n7569 Vbias.n877 236.048
R6621 Vbias.n877 Vbias.n875 236.048
R6622 Vbias.n6479 Vbias.n874 236.048
R6623 Vbias.n6487 Vbias.n868 236.048
R6624 Vbias.n6493 Vbias.n866 236.048
R6625 Vbias.n6501 Vbias.n860 236.048
R6626 Vbias.n7404 Vbias.n7398 236.048
R6627 Vbias.n7413 Vbias.n7382 236.048
R6628 Vbias.n7420 Vbias.n7419 236.048
R6629 Vbias.n7378 Vbias.n7368 236.048
R6630 Vbias.n7365 Vbias.n7364 236.048
R6631 Vbias.n7431 Vbias.n7364 236.048
R6632 Vbias.n7438 Vbias.n7360 236.048
R6633 Vbias.n7447 Vbias.n7344 236.048
R6634 Vbias.n7451 Vbias.n7340 236.048
R6635 Vbias.n7461 Vbias.n7325 236.048
R6636 Vbias.n6639 Vbias.n6148 236.048
R6637 Vbias.n6142 Vbias.n6135 236.048
R6638 Vbias.n7267 Vbias.n7260 236.048
R6639 Vbias.n7256 Vbias.n7242 236.048
R6640 Vbias.n7281 Vbias.n7231 236.048
R6641 Vbias.n7284 Vbias.n7283 236.048
R6642 Vbias.n7288 Vbias.n1069 236.048
R6643 Vbias.n7299 Vbias.n7298 236.048
R6644 Vbias.n7303 Vbias.n1048 236.048
R6645 Vbias.n7314 Vbias.n7313 236.048
R6646 Vbias.n7319 Vbias.n1021 236.048
R6647 Vbias.n1021 Vbias.n1019 236.048
R6648 Vbias.n7725 Vbias.n696 236.048
R6649 Vbias.n7733 Vbias.n681 236.048
R6650 Vbias.n1506 Vbias.n1503 236.048
R6651 Vbias.n6129 Vbias.n1503 236.048
R6652 Vbias.n344 Vbias.n326 236.048
R6653 Vbias.n346 Vbias.n326 236.048
R6654 Vbias.n2057 Vbias.n2056 236.048
R6655 Vbias.n2045 Vbias.n1719 236.048
R6656 Vbias.n6689 Vbias.n1452 236.048
R6657 Vbias.n6682 Vbias.n1455 236.048
R6658 Vbias.n5863 Vbias.n5862 236.048
R6659 Vbias.n1691 Vbias.n1681 236.048
R6660 Vbias.n1678 Vbias.n1677 236.048
R6661 Vbias.n5874 Vbias.n1677 236.048
R6662 Vbias.n5523 Vbias.n5515 236.048
R6663 Vbias.n5530 Vbias.n5511 236.048
R6664 Vbias.n5539 Vbias.n5538 236.048
R6665 Vbias.n2244 Vbias.n2234 236.048
R6666 Vbias.n2232 Vbias.n2231 236.048
R6667 Vbias.n5550 Vbias.n2231 236.048
R6668 Vbias.n5020 Vbias.n5019 236.048
R6669 Vbias.n5014 Vbias.n2586 236.048
R6670 Vbias.n8065 Vbias.n27 236.048
R6671 Vbias.n8073 Vbias.n12 236.048
R6672 Vbias.n7937 Vbias.n174 227.064
R6673 Vbias.n7821 Vbias.n553 227.064
R6674 Vbias.n7802 Vbias.n571 227.064
R6675 Vbias.n349 Vbias.n165 227.064
R6676 Vbias.t777 Vbias.n1529 217.311
R6677 Vbias.n1723 Vbias.t557 217.311
R6678 Vbias.t670 Vbias.n1724 217.311
R6679 Vbias.t559 Vbias.n1725 217.311
R6680 Vbias.t746 Vbias.n1524 215.714
R6681 Vbias.t746 Vbias.n1955 215.714
R6682 Vbias.t436 Vbias.n1955 215.714
R6683 Vbias.t436 Vbias.n1956 215.714
R6684 Vbias.t763 Vbias.n1956 215.714
R6685 Vbias.t763 Vbias.n1461 215.714
R6686 Vbias.n5011 Vbias.n5010 204.013
R6687 Vbias.n4904 Vbias.t839 203.526
R6688 Vbias.n4910 Vbias.t839 203.526
R6689 Vbias.t526 Vbias.n4911 203.526
R6690 Vbias.t526 Vbias.n2653 203.526
R6691 Vbias.t577 Vbias.n2653 203.526
R6692 Vbias.n4925 Vbias.t577 203.526
R6693 Vbias.n4925 Vbias.t445 203.526
R6694 Vbias.n4932 Vbias.t445 203.526
R6695 Vbias.t831 Vbias.n4933 203.526
R6696 Vbias.t831 Vbias.n2639 203.526
R6697 Vbias.t632 Vbias.n2639 203.526
R6698 Vbias.n4948 Vbias.t632 203.526
R6699 Vbias.n4948 Vbias.t517 203.526
R6700 Vbias.n4955 Vbias.t517 203.526
R6701 Vbias.t424 Vbias.n4956 203.526
R6702 Vbias.t424 Vbias.n2623 203.526
R6703 Vbias.t650 Vbias.n2623 203.526
R6704 Vbias.t650 Vbias.n2628 203.526
R6705 Vbias.n2627 Vbias.t826 203.526
R6706 Vbias.t826 Vbias.n2614 203.526
R6707 Vbias.t164 Vbias.n2614 203.526
R6708 Vbias.t164 Vbias.n2609 203.526
R6709 Vbias.t283 Vbias.n2609 203.526
R6710 Vbias.t283 Vbias.n2610 203.526
R6711 Vbias.n5602 Vbias.n5601 192.982
R6712 Vbias.n5620 Vbias.n5619 192.982
R6713 Vbias.n2222 Vbias.n2221 192.982
R6714 Vbias.n5676 Vbias.n5675 192.982
R6715 Vbias.n5694 Vbias.n5693 192.982
R6716 Vbias.n2151 Vbias.n2150 192.982
R6717 Vbias.n5751 Vbias.n5750 192.982
R6718 Vbias.n2112 Vbias.n2111 192.982
R6719 Vbias.n5796 Vbias.n5795 192.982
R6720 Vbias.n5837 Vbias.n2068 192.982
R6721 Vbias.n2060 Vbias.n2059 192.982
R6722 Vbias.n8001 Vbias.n8000 192.982
R6723 Vbias.n7986 Vbias.n7985 192.982
R6724 Vbias.n157 Vbias.n138 192.982
R6725 Vbias.t815 Vbias.n1531 190.261
R6726 Vbias.t793 Vbias.n1806 190.261
R6727 Vbias.n6676 Vbias.n6675 181.749
R6728 Vbias.n5534 Vbias.t457 179.623
R6729 Vbias.n2028 Vbias.t695 176.65
R6730 Vbias.n2027 Vbias.t364 176.65
R6731 Vbias.n2022 Vbias.t661 176.65
R6732 Vbias.n1748 Vbias.t437 176.65
R6733 Vbias.n1826 Vbias.t284 176.65
R6734 Vbias.n1831 Vbias.t884 176.65
R6735 Vbias.n1836 Vbias.t426 176.65
R6736 Vbias.n1841 Vbias.t279 176.65
R6737 Vbias.n8010 Vbias.n84 173.012
R6738 Vbias.n8022 Vbias.n8021 173.012
R6739 Vbias.n8033 Vbias.n62 173.012
R6740 Vbias.n8037 Vbias.n8036 173.012
R6741 Vbias.n8043 Vbias.n8042 173.012
R6742 Vbias.n8043 Vbias.n51 173.012
R6743 Vbias.n8047 Vbias.n45 173.012
R6744 Vbias.n8058 Vbias.n31 173.012
R6745 Vbias.n4336 Vbias.n4335 173.012
R6746 Vbias.n4335 Vbias.n2823 173.012
R6747 Vbias.n4265 Vbias.n4264 173.012
R6748 Vbias.n4265 Vbias.n4256 173.012
R6749 Vbias.n5007 Vbias.n5006 173.012
R6750 Vbias.n5002 Vbias.n2597 173.012
R6751 Vbias.n4990 Vbias.n4989 173.012
R6752 Vbias.n4989 Vbias.n2603 173.012
R6753 Vbias.n6713 Vbias.n6712 173.012
R6754 Vbias.n6715 Vbias.n6695 173.012
R6755 Vbias.n6740 Vbias.n6739 173.012
R6756 Vbias.n6742 Vbias.n6719 173.012
R6757 Vbias.n6746 Vbias.n1448 173.012
R6758 Vbias.n6747 Vbias.n6746 173.012
R6759 Vbias.n7745 Vbias.n674 173.012
R6760 Vbias.n7749 Vbias.n7748 173.012
R6761 Vbias.n7806 Vbias.n561 173.012
R6762 Vbias.n7813 Vbias.n559 173.012
R6763 Vbias.n7817 Vbias.n557 173.012
R6764 Vbias.n7818 Vbias.n7817 173.012
R6765 Vbias.n7880 Vbias.n453 173.012
R6766 Vbias.n7884 Vbias.n7883 173.012
R6767 Vbias.n7941 Vbias.n7940 173.012
R6768 Vbias.n339 Vbias.n338 173.012
R6769 Vbias.n7540 Vbias.n923 173.012
R6770 Vbias.n1015 Vbias.n921 173.012
R6771 Vbias.n7534 Vbias.n7533 173.012
R6772 Vbias.n6524 Vbias.n6523 173.012
R6773 Vbias.n6515 Vbias.n6514 173.012
R6774 Vbias.n6514 Vbias.n6510 173.012
R6775 Vbias.n7655 Vbias.n7654 173.012
R6776 Vbias.n7657 Vbias.n772 173.012
R6777 Vbias.n7661 Vbias.n763 173.012
R6778 Vbias.n769 Vbias.n761 173.012
R6779 Vbias.n7670 Vbias.n753 173.012
R6780 Vbias.n7682 Vbias.n7681 173.012
R6781 Vbias.n7693 Vbias.n731 173.012
R6782 Vbias.n7697 Vbias.n7696 173.012
R6783 Vbias.n7703 Vbias.n7702 173.012
R6784 Vbias.n7703 Vbias.n720 173.012
R6785 Vbias.n7707 Vbias.n714 173.012
R6786 Vbias.n7718 Vbias.n700 173.012
R6787 Vbias.n7756 Vbias.n7755 173.012
R6788 Vbias.n7762 Vbias.n7761 173.012
R6789 Vbias.n7768 Vbias.n7767 173.012
R6790 Vbias.n7770 Vbias.n626 173.012
R6791 Vbias.n7774 Vbias.n623 173.012
R6792 Vbias.n7775 Vbias.n7774 173.012
R6793 Vbias.n7781 Vbias.n7780 173.012
R6794 Vbias.n7787 Vbias.n7786 173.012
R6795 Vbias.n7793 Vbias.n7792 173.012
R6796 Vbias.n7799 Vbias.n7798 173.012
R6797 Vbias.n7825 Vbias.n7824 173.012
R6798 Vbias.n7831 Vbias.n7830 173.012
R6799 Vbias.n7837 Vbias.n7836 173.012
R6800 Vbias.n7839 Vbias.n512 173.012
R6801 Vbias.n7843 Vbias.n509 173.012
R6802 Vbias.n7844 Vbias.n7843 173.012
R6803 Vbias.n7850 Vbias.n7849 173.012
R6804 Vbias.n7856 Vbias.n7855 173.012
R6805 Vbias.n7862 Vbias.n7861 173.012
R6806 Vbias.n7868 Vbias.n7867 173.012
R6807 Vbias.n7891 Vbias.n7890 173.012
R6808 Vbias.n7897 Vbias.n7896 173.012
R6809 Vbias.n7903 Vbias.n7902 173.012
R6810 Vbias.n7905 Vbias.n406 173.012
R6811 Vbias.n7909 Vbias.n403 173.012
R6812 Vbias.n7910 Vbias.n7909 173.012
R6813 Vbias.n7916 Vbias.n7915 173.012
R6814 Vbias.n7922 Vbias.n7921 173.012
R6815 Vbias.n7928 Vbias.n7927 173.012
R6816 Vbias.n7934 Vbias.n7933 173.012
R6817 Vbias.n353 Vbias.n352 173.012
R6818 Vbias.n314 Vbias.n193 173.012
R6819 Vbias.n310 Vbias.n309 173.012
R6820 Vbias.n206 Vbias.n205 173.012
R6821 Vbias.n296 Vbias.n295 173.012
R6822 Vbias.n295 Vbias.n211 173.012
R6823 Vbias.n290 Vbias.n289 173.012
R6824 Vbias.n275 Vbias.n226 173.012
R6825 Vbias.n271 Vbias.n270 173.012
R6826 Vbias.n258 Vbias.n244 173.012
R6827 Vbias.n7948 Vbias.n163 173.012
R6828 Vbias.n7958 Vbias.n145 173.012
R6829 Vbias.n7962 Vbias.n134 173.012
R6830 Vbias.n7968 Vbias.n132 173.012
R6831 Vbias.n7975 Vbias.n128 173.012
R6832 Vbias.n7983 Vbias.n111 173.012
R6833 Vbias.n7990 Vbias.n107 173.012
R6834 Vbias.n7998 Vbias.n92 173.012
R6835 Vbias.n8003 Vbias.n89 173.012
R6836 Vbias.n8005 Vbias.n89 173.012
R6837 Vbias.n5034 Vbias.n5033 173.012
R6838 Vbias.n4645 Vbias.n4601 173.012
R6839 Vbias.n4649 Vbias.n4600 173.012
R6840 Vbias.n4653 Vbias.n4594 173.012
R6841 Vbias.n4657 Vbias.n4592 173.012
R6842 Vbias.n4658 Vbias.n4657 173.012
R6843 Vbias.n4664 Vbias.n4663 173.012
R6844 Vbias.n4668 Vbias.n4667 173.012
R6845 Vbias.n4494 Vbias.n4493 173.012
R6846 Vbias.n4494 Vbias.n4485 173.012
R6847 Vbias.n4498 Vbias.n4480 173.012
R6848 Vbias.n4508 Vbias.n4462 173.012
R6849 Vbias.n4512 Vbias.n4458 173.012
R6850 Vbias.n4522 Vbias.n4440 173.012
R6851 Vbias.n4526 Vbias.n4430 173.012
R6852 Vbias.n4532 Vbias.n4428 173.012
R6853 Vbias.n5118 Vbias.n5117 173.012
R6854 Vbias.n5102 Vbias.n2386 173.012
R6855 Vbias.n5098 Vbias.n5097 173.012
R6856 Vbias.n5082 Vbias.n2402 173.012
R6857 Vbias.n5077 Vbias.n5076 173.012
R6858 Vbias.n5076 Vbias.n2406 173.012
R6859 Vbias.n5071 Vbias.n5070 173.012
R6860 Vbias.n2415 Vbias.n2414 173.012
R6861 Vbias.n5489 Vbias.n5488 173.012
R6862 Vbias.n5495 Vbias.n5494 173.012
R6863 Vbias.n5501 Vbias.n5500 173.012
R6864 Vbias.n5155 Vbias.n2249 173.012
R6865 Vbias.n5164 Vbias.n5160 173.012
R6866 Vbias.n5165 Vbias.n5164 173.012
R6867 Vbias.n5171 Vbias.n5170 173.012
R6868 Vbias.n5173 Vbias.n2358 173.012
R6869 Vbias.n5177 Vbias.n2356 173.012
R6870 Vbias.n5181 Vbias.n2350 173.012
R6871 Vbias.n5915 Vbias.n5914 173.012
R6872 Vbias.n5899 Vbias.n1654 173.012
R6873 Vbias.n5895 Vbias.n5894 173.012
R6874 Vbias.n5879 Vbias.n1670 173.012
R6875 Vbias.n5459 Vbias.n5456 173.012
R6876 Vbias.n5460 Vbias.n5459 173.012
R6877 Vbias.n5466 Vbias.n5465 173.012
R6878 Vbias.n5470 Vbias.n5469 173.012
R6879 Vbias.n5476 Vbias.n5475 173.012
R6880 Vbias.n5482 Vbias.n5481 173.012
R6881 Vbias.n5944 Vbias.n5943 173.012
R6882 Vbias.n5946 Vbias.n1622 173.012
R6883 Vbias.n5950 Vbias.n1619 173.012
R6884 Vbias.n5954 Vbias.n1613 173.012
R6885 Vbias.n6097 Vbias.n1536 173.012
R6886 Vbias.n6098 Vbias.n6097 173.012
R6887 Vbias.n1521 Vbias.n1510 173.012
R6888 Vbias.n6111 Vbias.n6107 173.012
R6889 Vbias.n2001 Vbias.n1996 173.012
R6890 Vbias.n2014 Vbias.n2013 173.012
R6891 Vbias.n1961 Vbias.n1950 173.012
R6892 Vbias.n1971 Vbias.n1967 173.012
R6893 Vbias.n1927 Vbias.n1916 173.012
R6894 Vbias.n1937 Vbias.n1933 173.012
R6895 Vbias.n1819 Vbias.n1756 173.012
R6896 Vbias.n1807 Vbias.n1754 173.012
R6897 Vbias.n1871 Vbias.n1867 173.012
R6898 Vbias.n1859 Vbias.n1848 173.012
R6899 Vbias.n2036 Vbias.n2035 173.012
R6900 Vbias.n1743 Vbias.n1736 173.012
R6901 Vbias.n1913 Vbias.n1883 173.012
R6902 Vbias.n1901 Vbias.n1900 173.012
R6903 Vbias.n6081 Vbias.n6078 173.012
R6904 Vbias.n6085 Vbias.n1546 173.012
R6905 Vbias.n6089 Vbias.n1544 173.012
R6906 Vbias.n6093 Vbias.n1538 173.012
R6907 Vbias.n7012 Vbias.n7011 173.012
R6908 Vbias.n6783 Vbias.n1429 173.012
R6909 Vbias.n6787 Vbias.n1428 173.012
R6910 Vbias.n6791 Vbias.n1422 173.012
R6911 Vbias.n6795 Vbias.n1419 173.012
R6912 Vbias.n6796 Vbias.n6795 173.012
R6913 Vbias.n6802 Vbias.n6801 173.012
R6914 Vbias.n6804 Vbias.n1410 173.012
R6915 Vbias.n6808 Vbias.n1408 173.012
R6916 Vbias.n6812 Vbias.n1402 173.012
R6917 Vbias.n7093 Vbias.n7092 173.012
R6918 Vbias.n7080 Vbias.n1287 173.012
R6919 Vbias.n7076 Vbias.n7075 173.012
R6920 Vbias.n7063 Vbias.n1307 173.012
R6921 Vbias.n7059 Vbias.n7058 173.012
R6922 Vbias.n7059 Vbias.n1312 173.012
R6923 Vbias.n7051 Vbias.n7050 173.012
R6924 Vbias.n7046 Vbias.n1320 173.012
R6925 Vbias.n7034 Vbias.n7033 173.012
R6926 Vbias.n7018 Vbias.n1337 173.012
R6927 Vbias.n7199 Vbias.n7198 173.012
R6928 Vbias.n7186 Vbias.n1100 173.012
R6929 Vbias.n7182 Vbias.n7181 173.012
R6930 Vbias.n7169 Vbias.n1119 173.012
R6931 Vbias.n7165 Vbias.n7164 173.012
R6932 Vbias.n7165 Vbias.n1124 173.012
R6933 Vbias.n7157 Vbias.n7156 173.012
R6934 Vbias.n7152 Vbias.n1132 173.012
R6935 Vbias.n7140 Vbias.n7139 173.012
R6936 Vbias.n7124 Vbias.n1149 173.012
R6937 Vbias.n7220 Vbias.n1074 173.012
R6938 Vbias.n7222 Vbias.n1074 173.012
R6939 Vbias.n1222 Vbias.n1216 173.012
R6940 Vbias.n7215 Vbias.n1077 173.012
R6941 Vbias.n1241 Vbias.n1197 173.012
R6942 Vbias.n1231 Vbias.n1213 173.012
R6943 Vbias.n1253 Vbias.n1185 173.012
R6944 Vbias.n1246 Vbias.n1245 173.012
R6945 Vbias.n1272 Vbias.n1169 173.012
R6946 Vbias.n1262 Vbias.n1182 173.012
R6947 Vbias.n7118 Vbias.n1155 173.012
R6948 Vbias.n7116 Vbias.n1155 173.012
R6949 Vbias.n6955 Vbias.n6949 173.012
R6950 Vbias.n7111 Vbias.n1158 173.012
R6951 Vbias.n6974 Vbias.n6930 173.012
R6952 Vbias.n6964 Vbias.n6946 173.012
R6953 Vbias.n6986 Vbias.n6918 173.012
R6954 Vbias.n6979 Vbias.n6978 173.012
R6955 Vbias.n7005 Vbias.n6902 173.012
R6956 Vbias.n6995 Vbias.n6915 173.012
R6957 Vbias.n6897 Vbias.n1347 173.012
R6958 Vbias.n6897 Vbias.n1346 173.012
R6959 Vbias.n6878 Vbias.n1361 173.012
R6960 Vbias.n6890 Vbias.n1352 173.012
R6961 Vbias.n6855 Vbias.n1374 173.012
R6962 Vbias.n6867 Vbias.n1365 173.012
R6963 Vbias.n6837 Vbias.n1386 173.012
R6964 Vbias.n6844 Vbias.n1378 173.012
R6965 Vbias.n6817 Vbias.n1399 173.012
R6966 Vbias.n6831 Vbias.n1389 173.012
R6967 Vbias.n6042 Vbias.n1560 173.012
R6968 Vbias.n6040 Vbias.n1560 173.012
R6969 Vbias.n6020 Vbias.n1572 173.012
R6970 Vbias.n6035 Vbias.n1563 173.012
R6971 Vbias.n5997 Vbias.n1585 173.012
R6972 Vbias.n6009 Vbias.n1576 173.012
R6973 Vbias.n5979 Vbias.n1597 173.012
R6974 Vbias.n5986 Vbias.n1589 173.012
R6975 Vbias.n5959 Vbias.n1610 173.012
R6976 Vbias.n5973 Vbias.n1600 173.012
R6977 Vbias.n5345 Vbias.n5343 173.012
R6978 Vbias.n5347 Vbias.n5343 173.012
R6979 Vbias.n5363 Vbias.n5318 173.012
R6980 Vbias.n5354 Vbias.n5336 173.012
R6981 Vbias.n5382 Vbias.n5301 173.012
R6982 Vbias.n5372 Vbias.n5315 173.012
R6983 Vbias.n5394 Vbias.n5289 173.012
R6984 Vbias.n5387 Vbias.n5386 173.012
R6985 Vbias.n5413 Vbias.n5272 173.012
R6986 Vbias.n5403 Vbias.n5286 173.012
R6987 Vbias.n5267 Vbias.n2295 173.012
R6988 Vbias.n5267 Vbias.n2294 173.012
R6989 Vbias.n5247 Vbias.n2309 173.012
R6990 Vbias.n5259 Vbias.n2300 173.012
R6991 Vbias.n5224 Vbias.n2322 173.012
R6992 Vbias.n5236 Vbias.n2313 173.012
R6993 Vbias.n5206 Vbias.n2334 173.012
R6994 Vbias.n5213 Vbias.n2326 173.012
R6995 Vbias.n5186 Vbias.n2347 173.012
R6996 Vbias.n5200 Vbias.n2337 173.012
R6997 Vbias.n2513 Vbias.n2511 173.012
R6998 Vbias.n2515 Vbias.n2511 173.012
R6999 Vbias.n2531 Vbias.n2486 173.012
R7000 Vbias.n2522 Vbias.n2504 173.012
R7001 Vbias.n2550 Vbias.n2469 173.012
R7002 Vbias.n2540 Vbias.n2483 173.012
R7003 Vbias.n2562 Vbias.n2457 173.012
R7004 Vbias.n2555 Vbias.n2554 173.012
R7005 Vbias.n2581 Vbias.n2440 173.012
R7006 Vbias.n2571 Vbias.n2454 173.012
R7007 Vbias.n5055 Vbias.n5054 173.012
R7008 Vbias.n5039 Vbias.n2431 173.012
R7009 Vbias.n4548 Vbias.n4409 173.012
R7010 Vbias.n4539 Vbias.n4424 173.012
R7011 Vbias.n3890 Vbias.n3775 173.012
R7012 Vbias.n3891 Vbias.n3890 173.012
R7013 Vbias.n3974 Vbias.n3711 173.012
R7014 Vbias.n3974 Vbias.n3710 173.012
R7015 Vbias.n3352 Vbias.n3237 173.012
R7016 Vbias.n3353 Vbias.n3352 173.012
R7017 Vbias.n3436 Vbias.n3173 173.012
R7018 Vbias.n3436 Vbias.n3172 173.012
R7019 Vbias.n3621 Vbias.n3506 173.012
R7020 Vbias.n3622 Vbias.n3621 173.012
R7021 Vbias.n3705 Vbias.n3442 173.012
R7022 Vbias.n3705 Vbias.n3441 173.012
R7023 Vbias.n4186 Vbias.n4069 173.012
R7024 Vbias.n4198 Vbias.n4197 173.012
R7025 Vbias.n4204 Vbias.n4040 173.012
R7026 Vbias.n4211 Vbias.n4038 173.012
R7027 Vbias.n4215 Vbias.n4035 173.012
R7028 Vbias.n4216 Vbias.n4215 173.012
R7029 Vbias.n4220 Vbias.n4027 173.012
R7030 Vbias.n4232 Vbias.n4231 173.012
R7031 Vbias.n4239 Vbias.n4001 173.012
R7032 Vbias.n4249 Vbias.n3981 173.012
R7033 Vbias.n4183 Vbias.n4182 173.012
R7034 Vbias.n4177 Vbias.n4168 173.012
R7035 Vbias.n4163 Vbias.n4162 173.012
R7036 Vbias.n4148 Vbias.n4146 173.012
R7037 Vbias.n4140 Vbias.n4139 173.012
R7038 Vbias.n4128 Vbias.n4086 173.012
R7039 Vbias.n4124 Vbias.n4123 173.012
R7040 Vbias.n4117 Vbias.n4115 173.012
R7041 Vbias.n4111 Vbias.n4104 173.012
R7042 Vbias.n4111 Vbias.n4103 173.012
R7043 Vbias.n4971 Vbias.n2616 173.012
R7044 Vbias.n4985 Vbias.n2606 173.012
R7045 Vbias.n4957 Vbias.n2630 173.012
R7046 Vbias.n4967 Vbias.n2620 173.012
R7047 Vbias.n4941 Vbias.n2644 173.012
R7048 Vbias.n4953 Vbias.n2634 173.012
R7049 Vbias.n4919 Vbias.n2658 173.012
R7050 Vbias.n4930 Vbias.n2648 173.012
R7051 Vbias.n4908 Vbias.n2662 173.012
R7052 Vbias.n4906 Vbias.n2662 173.012
R7053 Vbias.n3082 Vbias.n2967 173.012
R7054 Vbias.n3083 Vbias.n3082 173.012
R7055 Vbias.n3166 Vbias.n2902 173.012
R7056 Vbias.n3166 Vbias.n2901 173.012
R7057 Vbias.n4758 Vbias.n2728 173.012
R7058 Vbias.n4759 Vbias.n4758 173.012
R7059 Vbias.n4840 Vbias.n2666 173.012
R7060 Vbias.n4842 Vbias.n2666 173.012
R7061 Vbias.n4674 Vbias.n4673 173.012
R7062 Vbias.n4679 Vbias.n4678 173.012
R7063 Vbias.n5662 Vbias.n2197 173.012
R7064 Vbias.n5652 Vbias.n2210 173.012
R7065 Vbias.n5648 Vbias.n2214 173.012
R7066 Vbias.n5640 Vbias.n2226 173.012
R7067 Vbias.n5636 Vbias.n5556 173.012
R7068 Vbias.n5624 Vbias.n5570 173.012
R7069 Vbias.n5617 Vbias.n5574 173.012
R7070 Vbias.n5606 Vbias.n5588 173.012
R7071 Vbias.n5599 Vbias.n5595 173.012
R7072 Vbias.n5597 Vbias.n5595 173.012
R7073 Vbias.n5736 Vbias.n2126 173.012
R7074 Vbias.n5726 Vbias.n2139 173.012
R7075 Vbias.n5722 Vbias.n2143 173.012
R7076 Vbias.n5714 Vbias.n2155 173.012
R7077 Vbias.n5710 Vbias.n2159 173.012
R7078 Vbias.n5698 Vbias.n2173 173.012
R7079 Vbias.n5691 Vbias.n2177 173.012
R7080 Vbias.n5680 Vbias.n2191 173.012
R7081 Vbias.n5673 Vbias.n5669 173.012
R7082 Vbias.n5671 Vbias.n5669 173.012
R7083 Vbias.n5825 Vbias.n2071 173.012
R7084 Vbias.n5815 Vbias.n2084 173.012
R7085 Vbias.n5811 Vbias.n5788 173.012
R7086 Vbias.n5803 Vbias.n5800 173.012
R7087 Vbias.n5783 Vbias.n2088 173.012
R7088 Vbias.n5772 Vbias.n2100 173.012
R7089 Vbias.n5768 Vbias.n2104 173.012
R7090 Vbias.n5758 Vbias.n2122 173.012
R7091 Vbias.n5754 Vbias.n5753 173.012
R7092 Vbias.n5754 Vbias.n5742 173.012
R7093 Vbias.n6653 Vbias.n1499 173.012
R7094 Vbias.n6663 Vbias.n1482 173.012
R7095 Vbias.n6667 Vbias.n1472 173.012
R7096 Vbias.n6673 Vbias.n1470 173.012
R7097 Vbias.n5854 Vbias.n1702 173.012
R7098 Vbias.n5844 Vbias.n2064 173.012
R7099 Vbias.n5840 Vbias.n5839 173.012
R7100 Vbias.n5840 Vbias.n5832 173.012
R7101 Vbias.n6587 Vbias.n6229 173.012
R7102 Vbias.n6357 Vbias.n6243 173.012
R7103 Vbias.n6350 Vbias.n6247 173.012
R7104 Vbias.n6344 Vbias.n6249 173.012
R7105 Vbias.n6339 Vbias.n6259 173.012
R7106 Vbias.n6329 Vbias.n6273 173.012
R7107 Vbias.n6325 Vbias.n6277 173.012
R7108 Vbias.n6315 Vbias.n6295 173.012
R7109 Vbias.n6311 Vbias.n6310 173.012
R7110 Vbias.n6311 Vbias.n6298 173.012
R7111 Vbias.n7592 Vbias.n855 173.012
R7112 Vbias.n7602 Vbias.n837 173.012
R7113 Vbias.n7606 Vbias.n826 173.012
R7114 Vbias.n7612 Vbias.n824 173.012
R7115 Vbias.n7619 Vbias.n819 173.012
R7116 Vbias.n7627 Vbias.n802 173.012
R7117 Vbias.n7634 Vbias.n798 173.012
R7118 Vbias.n7642 Vbias.n783 173.012
R7119 Vbias.n7647 Vbias.n780 173.012
R7120 Vbias.n7649 Vbias.n780 173.012
R7121 Vbias.n7470 Vbias.n1010 173.012
R7122 Vbias.n7480 Vbias.n992 173.012
R7123 Vbias.n7484 Vbias.n981 173.012
R7124 Vbias.n7490 Vbias.n979 173.012
R7125 Vbias.n7498 Vbias.n974 173.012
R7126 Vbias.n7506 Vbias.n957 173.012
R7127 Vbias.n7513 Vbias.n953 173.012
R7128 Vbias.n7521 Vbias.n934 173.012
R7129 Vbias.n7526 Vbias.n931 173.012
R7130 Vbias.n7528 Vbias.n931 173.012
R7131 Vbias.n6602 Vbias.n6601 173.012
R7132 Vbias.n6608 Vbias.n6607 173.012
R7133 Vbias.n6614 Vbias.n6613 173.012
R7134 Vbias.n6618 Vbias.n6617 173.012
R7135 Vbias.n6624 Vbias.n6623 173.012
R7136 Vbias.n6624 Vbias.n6162 173.012
R7137 Vbias.n6628 Vbias.n6161 173.012
R7138 Vbias.n6632 Vbias.n6155 173.012
R7139 Vbias.n6535 Vbias.n6534 173.012
R7140 Vbias.n6541 Vbias.n6540 173.012
R7141 Vbias.n6547 Vbias.n6546 173.012
R7142 Vbias.n6551 Vbias.n6550 173.012
R7143 Vbias.n6557 Vbias.n6556 173.012
R7144 Vbias.n6557 Vbias.n6380 173.012
R7145 Vbias.n6561 Vbias.n6379 173.012
R7146 Vbias.n6565 Vbias.n6373 173.012
R7147 Vbias.n6569 Vbias.n6371 173.012
R7148 Vbias.n6573 Vbias.n6365 173.012
R7149 Vbias.n7548 Vbias.n7547 173.012
R7150 Vbias.n7554 Vbias.n7553 173.012
R7151 Vbias.n7560 Vbias.n7559 173.012
R7152 Vbias.n7564 Vbias.n7563 173.012
R7153 Vbias.n7570 Vbias.n7569 173.012
R7154 Vbias.n7570 Vbias.n875 173.012
R7155 Vbias.n7574 Vbias.n874 173.012
R7156 Vbias.n7578 Vbias.n868 173.012
R7157 Vbias.n7582 Vbias.n866 173.012
R7158 Vbias.n7586 Vbias.n860 173.012
R7159 Vbias.n7400 Vbias.n7398 173.012
R7160 Vbias.n7413 Vbias.n7412 173.012
R7161 Vbias.n7419 Vbias.n7370 173.012
R7162 Vbias.n7426 Vbias.n7368 173.012
R7163 Vbias.n7430 Vbias.n7365 173.012
R7164 Vbias.n7431 Vbias.n7430 173.012
R7165 Vbias.n7435 Vbias.n7360 173.012
R7166 Vbias.n7447 Vbias.n7446 173.012
R7167 Vbias.n7454 Vbias.n7340 173.012
R7168 Vbias.n7464 Vbias.n7325 173.012
R7169 Vbias.n6636 Vbias.n6148 173.012
R7170 Vbias.n6647 Vbias.n6135 173.012
R7171 Vbias.n7263 Vbias.n7260 173.012
R7172 Vbias.n7274 Vbias.n7242 173.012
R7173 Vbias.n7278 Vbias.n7231 173.012
R7174 Vbias.n7284 Vbias.n7229 173.012
R7175 Vbias.n7291 Vbias.n1069 173.012
R7176 Vbias.n7299 Vbias.n1052 173.012
R7177 Vbias.n7306 Vbias.n1048 173.012
R7178 Vbias.n7314 Vbias.n1031 173.012
R7179 Vbias.n7320 Vbias.n7319 173.012
R7180 Vbias.n7320 Vbias.n1019 173.012
R7181 Vbias.n7722 Vbias.n696 173.012
R7182 Vbias.n7733 Vbias.n7732 173.012
R7183 Vbias.n6128 Vbias.n1506 173.012
R7184 Vbias.n6129 Vbias.n6128 173.012
R7185 Vbias.n345 Vbias.n344 173.012
R7186 Vbias.n346 Vbias.n345 173.012
R7187 Vbias.n2057 Vbias.n1706 173.012
R7188 Vbias.n2048 Vbias.n1719 173.012
R7189 Vbias.n6690 Vbias.n6689 173.012
R7190 Vbias.n1456 Vbias.n1455 173.012
R7191 Vbias.n5862 Vbias.n1683 173.012
R7192 Vbias.n5869 Vbias.n1681 173.012
R7193 Vbias.n5873 Vbias.n1678 173.012
R7194 Vbias.n5874 Vbias.n5873 173.012
R7195 Vbias.n5526 Vbias.n5515 173.012
R7196 Vbias.n5530 Vbias.n5529 173.012
R7197 Vbias.n5538 Vbias.n2236 173.012
R7198 Vbias.n5545 Vbias.n2234 173.012
R7199 Vbias.n5549 Vbias.n2232 173.012
R7200 Vbias.n5550 Vbias.n5549 173.012
R7201 Vbias.n5019 Vbias.n2588 173.012
R7202 Vbias.n5026 Vbias.n2586 173.012
R7203 Vbias.n8062 Vbias.n27 173.012
R7204 Vbias.n8073 Vbias.n8072 173.012
R7205 Vbias.n8078 Vbias.n8077 168.537
R7206 Vbias.n8076 Vbias.n7 163.056
R7207 Vbias.n4685 Vbias.n2773 163.056
R7208 Vbias.n8076 Vbias.n8 163.056
R7209 Vbias.n4685 Vbias.n2774 163.056
R7210 Vbias.n8076 Vbias.n9 163.056
R7211 Vbias.n4685 Vbias.n2775 163.056
R7212 Vbias.n4685 Vbias.n2776 163.056
R7213 Vbias.n4686 Vbias.n4685 163.056
R7214 Vbias.n4685 Vbias.n4406 163.056
R7215 Vbias.n8077 Vbias.n8076 159.131
R7216 Vbias.t212 Vbias.n1528 152.346
R7217 Vbias.n2800 Vbias.n2797 150.213
R7218 Vbias.n4404 Vbias.n4403 150.213
R7219 Vbias.n4403 Vbias.n4402 150.213
R7220 Vbias.n4367 Vbias.n2797 150.213
R7221 Vbias.n4362 Vbias.n4361 150.213
R7222 Vbias.n2819 Vbias.n2810 150.213
R7223 Vbias.n4361 Vbias.n2806 150.213
R7224 Vbias.n4341 Vbias.n2810 150.213
R7225 Vbias.n4303 Vbias.n2846 150.213
R7226 Vbias.n4327 Vbias.n2827 150.213
R7227 Vbias.n4312 Vbias.n2827 150.213
R7228 Vbias.n4304 Vbias.n4303 150.213
R7229 Vbias.n4270 Vbias.n2880 150.213
R7230 Vbias.n4294 Vbias.n2863 150.213
R7231 Vbias.n4279 Vbias.n2863 150.213
R7232 Vbias.n4271 Vbias.n4270 150.213
R7233 Vbias.n3852 Vbias.n3794 150.213
R7234 Vbias.n3839 Vbias.n3815 150.213
R7235 Vbias.n3839 Vbias.n3838 150.213
R7236 Vbias.n3853 Vbias.n3852 150.213
R7237 Vbias.n3878 Vbias.n3877 150.213
R7238 Vbias.n3860 Vbias.n3778 150.213
R7239 Vbias.n3877 Vbias.n3875 150.213
R7240 Vbias.n3865 Vbias.n3778 150.213
R7241 Vbias.n3928 Vbias.n3747 150.213
R7242 Vbias.n3915 Vbias.n3768 150.213
R7243 Vbias.n3915 Vbias.n3914 150.213
R7244 Vbias.n3929 Vbias.n3928 150.213
R7245 Vbias.n3966 Vbias.n3718 150.213
R7246 Vbias.n3953 Vbias.n3739 150.213
R7247 Vbias.n3953 Vbias.n3952 150.213
R7248 Vbias.n3967 Vbias.n3966 150.213
R7249 Vbias.n3314 Vbias.n3256 150.213
R7250 Vbias.n3301 Vbias.n3277 150.213
R7251 Vbias.n3301 Vbias.n3300 150.213
R7252 Vbias.n3315 Vbias.n3314 150.213
R7253 Vbias.n3340 Vbias.n3339 150.213
R7254 Vbias.n3322 Vbias.n3240 150.213
R7255 Vbias.n3339 Vbias.n3337 150.213
R7256 Vbias.n3327 Vbias.n3240 150.213
R7257 Vbias.n3390 Vbias.n3209 150.213
R7258 Vbias.n3377 Vbias.n3230 150.213
R7259 Vbias.n3377 Vbias.n3376 150.213
R7260 Vbias.n3391 Vbias.n3390 150.213
R7261 Vbias.n3428 Vbias.n3180 150.213
R7262 Vbias.n3415 Vbias.n3201 150.213
R7263 Vbias.n3415 Vbias.n3414 150.213
R7264 Vbias.n3429 Vbias.n3428 150.213
R7265 Vbias.n3583 Vbias.n3525 150.213
R7266 Vbias.n3570 Vbias.n3546 150.213
R7267 Vbias.n3570 Vbias.n3569 150.213
R7268 Vbias.n3584 Vbias.n3583 150.213
R7269 Vbias.n3609 Vbias.n3608 150.213
R7270 Vbias.n3591 Vbias.n3509 150.213
R7271 Vbias.n3608 Vbias.n3606 150.213
R7272 Vbias.n3596 Vbias.n3509 150.213
R7273 Vbias.n3659 Vbias.n3478 150.213
R7274 Vbias.n3646 Vbias.n3499 150.213
R7275 Vbias.n3646 Vbias.n3645 150.213
R7276 Vbias.n3660 Vbias.n3659 150.213
R7277 Vbias.n3697 Vbias.n3449 150.213
R7278 Vbias.n3684 Vbias.n3470 150.213
R7279 Vbias.n3684 Vbias.n3683 150.213
R7280 Vbias.n3698 Vbias.n3697 150.213
R7281 Vbias.n3044 Vbias.n2986 150.213
R7282 Vbias.n3031 Vbias.n3007 150.213
R7283 Vbias.n3031 Vbias.n3030 150.213
R7284 Vbias.n3045 Vbias.n3044 150.213
R7285 Vbias.n3070 Vbias.n3069 150.213
R7286 Vbias.n3052 Vbias.n2970 150.213
R7287 Vbias.n3069 Vbias.n3067 150.213
R7288 Vbias.n3057 Vbias.n2970 150.213
R7289 Vbias.n3120 Vbias.n2939 150.213
R7290 Vbias.n3107 Vbias.n2960 150.213
R7291 Vbias.n3107 Vbias.n3106 150.213
R7292 Vbias.n3121 Vbias.n3120 150.213
R7293 Vbias.n3158 Vbias.n2910 150.213
R7294 Vbias.n3145 Vbias.n2931 150.213
R7295 Vbias.n3145 Vbias.n3144 150.213
R7296 Vbias.n3159 Vbias.n3158 150.213
R7297 Vbias.n4720 Vbias.n2747 150.213
R7298 Vbias.n4707 Vbias.n2768 150.213
R7299 Vbias.n4707 Vbias.n4706 150.213
R7300 Vbias.n4721 Vbias.n4720 150.213
R7301 Vbias.n4746 Vbias.n4745 150.213
R7302 Vbias.n4728 Vbias.n2731 150.213
R7303 Vbias.n4745 Vbias.n4743 150.213
R7304 Vbias.n4733 Vbias.n2731 150.213
R7305 Vbias.n4796 Vbias.n2700 150.213
R7306 Vbias.n4783 Vbias.n2721 150.213
R7307 Vbias.n4783 Vbias.n4782 150.213
R7308 Vbias.n4797 Vbias.n4796 150.213
R7309 Vbias.n4834 Vbias.n2671 150.213
R7310 Vbias.n4821 Vbias.n2692 150.213
R7311 Vbias.n4821 Vbias.n4820 150.213
R7312 Vbias.n4835 Vbias.n4834 150.213
R7313 Vbias.n4107 Vbias.n3985 147.843
R7314 Vbias.n4235 Vbias.n4234 147.843
R7315 Vbias.n4219 Vbias.n4218 147.843
R7316 Vbias.n4155 Vbias.n4151 147.843
R7317 Vbias.n4201 Vbias.n4200 147.843
R7318 Vbias.n5010 Vbias.t46 143.995
R7319 Vbias.n7668 Vbias.t646 137.369
R7320 Vbias.n6531 Vbias.t402 137.369
R7321 Vbias.n4895 Vbias.n4892 135.484
R7322 Vbias.t702 Vbias.n4900 134.439
R7323 Vbias.n4871 Vbias.n4870 127.775
R7324 Vbias.n6101 Vbias.n1527 127.168
R7325 Vbias.n6676 Vbias.n1465 127.168
R7326 Vbias.n8014 Vbias.n83 120.472
R7327 Vbias.n83 Vbias.n72 120.472
R7328 Vbias.n81 Vbias.n80 120.472
R7329 Vbias.n80 Vbias.n69 120.472
R7330 Vbias.n8029 Vbias.n8028 120.472
R7331 Vbias.n8028 Vbias.n60 120.472
R7332 Vbias.n8051 Vbias.n44 120.472
R7333 Vbias.n50 Vbias.n44 120.472
R7334 Vbias.n8056 Vbias.n34 120.472
R7335 Vbias.n8057 Vbias.n8056 120.472
R7336 Vbias.n4395 Vbias.n4394 120.472
R7337 Vbias.n4394 Vbias.n4391 120.472
R7338 Vbias.n4376 Vbias.n4375 120.472
R7339 Vbias.n4375 Vbias.n4372 120.472
R7340 Vbias.n4389 Vbias.n4388 120.472
R7341 Vbias.n4388 Vbias.n2782 120.472
R7342 Vbias.n4379 Vbias.n2794 120.472
R7343 Vbias.n4380 Vbias.n4379 120.472
R7344 Vbias.n4350 Vbias.n2813 120.472
R7345 Vbias.n4350 Vbias.n4349 120.472
R7346 Vbias.n4354 Vbias.n2814 120.472
R7347 Vbias.n4355 Vbias.n4354 120.472
R7348 Vbias.n4326 Vbias.n2837 120.472
R7349 Vbias.n4320 Vbias.n2837 120.472
R7350 Vbias.n2855 Vbias.n2845 120.472
R7351 Vbias.n4309 Vbias.n2845 120.472
R7352 Vbias.n4319 Vbias.n4318 120.472
R7353 Vbias.n4318 Vbias.n4314 120.472
R7354 Vbias.n2857 Vbias.n2838 120.472
R7355 Vbias.n2858 Vbias.n2857 120.472
R7356 Vbias.n4293 Vbias.n2871 120.472
R7357 Vbias.n4287 Vbias.n2871 120.472
R7358 Vbias.n2889 Vbias.n2879 120.472
R7359 Vbias.n4276 Vbias.n2879 120.472
R7360 Vbias.n4286 Vbias.n4285 120.472
R7361 Vbias.n4285 Vbias.n4281 120.472
R7362 Vbias.n2891 Vbias.n2872 120.472
R7363 Vbias.n2892 Vbias.n2891 120.472
R7364 Vbias.n4998 Vbias.n4997 120.472
R7365 Vbias.n4997 Vbias.n2596 120.472
R7366 Vbias.n6703 Vbias.n6697 120.472
R7367 Vbias.n6714 Vbias.n6697 120.472
R7368 Vbias.n6729 Vbias.n6721 120.472
R7369 Vbias.n6741 Vbias.n6721 120.472
R7370 Vbias.n7741 Vbias.n7740 120.472
R7371 Vbias.n7740 Vbias.n671 120.472
R7372 Vbias.n7811 Vbias.n562 120.472
R7373 Vbias.n7812 Vbias.n7811 120.472
R7374 Vbias.n7876 Vbias.n7875 120.472
R7375 Vbias.n7875 Vbias.n451 120.472
R7376 Vbias.n335 Vbias.n334 120.472
R7377 Vbias.n334 Vbias.n170 120.472
R7378 Vbias.n7542 Vbias.n920 120.472
R7379 Vbias.n7542 Vbias.n7541 120.472
R7380 Vbias.n6528 Vbias.n6527 120.472
R7381 Vbias.n6527 Vbias.n925 120.472
R7382 Vbias.n6592 Vbias.n774 120.472
R7383 Vbias.n7656 Vbias.n774 120.472
R7384 Vbias.n7665 Vbias.n762 120.472
R7385 Vbias.n768 Vbias.n762 120.472
R7386 Vbias.n7674 Vbias.n752 120.472
R7387 Vbias.n752 Vbias.n741 120.472
R7388 Vbias.n750 Vbias.n749 120.472
R7389 Vbias.n749 Vbias.n738 120.472
R7390 Vbias.n7689 Vbias.n7688 120.472
R7391 Vbias.n7688 Vbias.n729 120.472
R7392 Vbias.n7711 Vbias.n713 120.472
R7393 Vbias.n719 Vbias.n713 120.472
R7394 Vbias.n7716 Vbias.n703 120.472
R7395 Vbias.n7717 Vbias.n7716 120.472
R7396 Vbias.n660 Vbias.n650 120.472
R7397 Vbias.n7757 Vbias.n650 120.472
R7398 Vbias.n659 Vbias.n658 120.472
R7399 Vbias.n658 Vbias.n646 120.472
R7400 Vbias.n636 Vbias.n628 120.472
R7401 Vbias.n7769 Vbias.n628 120.472
R7402 Vbias.n613 Vbias.n603 120.472
R7403 Vbias.n7782 Vbias.n603 120.472
R7404 Vbias.n612 Vbias.n611 120.472
R7405 Vbias.n611 Vbias.n599 120.472
R7406 Vbias.n589 Vbias.n579 120.472
R7407 Vbias.n7794 Vbias.n579 120.472
R7408 Vbias.n588 Vbias.n587 120.472
R7409 Vbias.n587 Vbias.n575 120.472
R7410 Vbias.n546 Vbias.n536 120.472
R7411 Vbias.n7826 Vbias.n536 120.472
R7412 Vbias.n545 Vbias.n544 120.472
R7413 Vbias.n544 Vbias.n532 120.472
R7414 Vbias.n522 Vbias.n514 120.472
R7415 Vbias.n7838 Vbias.n514 120.472
R7416 Vbias.n499 Vbias.n489 120.472
R7417 Vbias.n7851 Vbias.n489 120.472
R7418 Vbias.n498 Vbias.n497 120.472
R7419 Vbias.n497 Vbias.n485 120.472
R7420 Vbias.n475 Vbias.n465 120.472
R7421 Vbias.n7863 Vbias.n465 120.472
R7422 Vbias.n474 Vbias.n473 120.472
R7423 Vbias.n473 Vbias.n461 120.472
R7424 Vbias.n440 Vbias.n430 120.472
R7425 Vbias.n7892 Vbias.n430 120.472
R7426 Vbias.n439 Vbias.n438 120.472
R7427 Vbias.n438 Vbias.n426 120.472
R7428 Vbias.n416 Vbias.n408 120.472
R7429 Vbias.n7904 Vbias.n408 120.472
R7430 Vbias.n393 Vbias.n383 120.472
R7431 Vbias.n7917 Vbias.n383 120.472
R7432 Vbias.n392 Vbias.n391 120.472
R7433 Vbias.n391 Vbias.n379 120.472
R7434 Vbias.n369 Vbias.n359 120.472
R7435 Vbias.n7929 Vbias.n359 120.472
R7436 Vbias.n368 Vbias.n367 120.472
R7437 Vbias.n367 Vbias.n178 120.472
R7438 Vbias.n321 Vbias.n320 120.472
R7439 Vbias.n321 Vbias.n180 120.472
R7440 Vbias.n194 Vbias.n186 120.472
R7441 Vbias.n197 Vbias.n194 120.472
R7442 Vbias.n304 Vbias.n303 120.472
R7443 Vbias.n304 Vbias.n199 120.472
R7444 Vbias.n282 Vbias.n281 120.472
R7445 Vbias.n282 Vbias.n213 120.472
R7446 Vbias.n227 Vbias.n219 120.472
R7447 Vbias.n230 Vbias.n227 120.472
R7448 Vbias.n265 Vbias.n264 120.472
R7449 Vbias.n265 Vbias.n232 120.472
R7450 Vbias.n247 Vbias.n238 120.472
R7451 Vbias.n248 Vbias.n247 120.472
R7452 Vbias.n7957 Vbias.n147 120.472
R7453 Vbias.n160 Vbias.n147 120.472
R7454 Vbias.n162 Vbias.n148 120.472
R7455 Vbias.n7952 Vbias.n162 120.472
R7456 Vbias.n141 Vbias.n133 120.472
R7457 Vbias.n7966 Vbias.n133 120.472
R7458 Vbias.n121 Vbias.n112 120.472
R7459 Vbias.n7981 Vbias.n112 120.472
R7460 Vbias.n7976 Vbias.n126 120.472
R7461 Vbias.n126 Vbias.n113 120.472
R7462 Vbias.n102 Vbias.n93 120.472
R7463 Vbias.n7996 Vbias.n93 120.472
R7464 Vbias.n7991 Vbias.n105 120.472
R7465 Vbias.n105 Vbias.n94 120.472
R7466 Vbias.n4639 Vbias.n4638 120.472
R7467 Vbias.n4638 Vbias.n2437 120.472
R7468 Vbias.n4636 Vbias.n4603 120.472
R7469 Vbias.n4644 Vbias.n4603 120.472
R7470 Vbias.n4628 Vbias.n4598 120.472
R7471 Vbias.n4650 Vbias.n4598 120.472
R7472 Vbias.n4613 Vbias.n4596 120.472
R7473 Vbias.n4652 Vbias.n4596 120.472
R7474 Vbias.n4586 Vbias.n4585 120.472
R7475 Vbias.n4586 Vbias.n4577 120.472
R7476 Vbias.n4507 Vbias.n4464 120.472
R7477 Vbias.n4477 Vbias.n4464 120.472
R7478 Vbias.n4479 Vbias.n4465 120.472
R7479 Vbias.n4502 Vbias.n4479 120.472
R7480 Vbias.n4521 Vbias.n4442 120.472
R7481 Vbias.n4455 Vbias.n4442 120.472
R7482 Vbias.n4457 Vbias.n4443 120.472
R7483 Vbias.n4516 Vbias.n4457 120.472
R7484 Vbias.n4437 Vbias.n4429 120.472
R7485 Vbias.n4530 Vbias.n4429 120.472
R7486 Vbias.n5109 Vbias.n5108 120.472
R7487 Vbias.n5108 Vbias.n2375 120.472
R7488 Vbias.n5106 Vbias.n2385 120.472
R7489 Vbias.n2385 Vbias.n2377 120.472
R7490 Vbias.n5089 Vbias.n5088 120.472
R7491 Vbias.n5088 Vbias.n2391 120.472
R7492 Vbias.n5086 Vbias.n2401 120.472
R7493 Vbias.n2401 Vbias.n2393 120.472
R7494 Vbias.n5063 Vbias.n5062 120.472
R7495 Vbias.n5063 Vbias.n2408 120.472
R7496 Vbias.n2281 Vbias.n2271 120.472
R7497 Vbias.n5490 Vbias.n2271 120.472
R7498 Vbias.n2280 Vbias.n2279 120.472
R7499 Vbias.n2279 Vbias.n2268 120.472
R7500 Vbias.n2262 Vbias.n2261 120.472
R7501 Vbias.n2262 Vbias.n2251 120.472
R7502 Vbias.n5506 Vbias.n2248 120.472
R7503 Vbias.n5506 Vbias.n5505 120.472
R7504 Vbias.n5142 Vbias.n2360 120.472
R7505 Vbias.n5172 Vbias.n2360 120.472
R7506 Vbias.n5135 Vbias.n2354 120.472
R7507 Vbias.n5178 Vbias.n2354 120.472
R7508 Vbias.n2365 Vbias.n2352 120.472
R7509 Vbias.n5180 Vbias.n2352 120.472
R7510 Vbias.n5906 Vbias.n5905 120.472
R7511 Vbias.n5905 Vbias.n1643 120.472
R7512 Vbias.n5903 Vbias.n1653 120.472
R7513 Vbias.n1653 Vbias.n1645 120.472
R7514 Vbias.n5886 Vbias.n5885 120.472
R7515 Vbias.n5885 Vbias.n1659 120.472
R7516 Vbias.n5883 Vbias.n1669 120.472
R7517 Vbias.n1669 Vbias.n1661 120.472
R7518 Vbias.n5448 Vbias.n5447 120.472
R7519 Vbias.n5448 Vbias.n5439 120.472
R7520 Vbias.n5429 Vbias.n5419 120.472
R7521 Vbias.n5477 Vbias.n5419 120.472
R7522 Vbias.n5428 Vbias.n5427 120.472
R7523 Vbias.n5427 Vbias.n2292 120.472
R7524 Vbias.n5935 Vbias.n1624 120.472
R7525 Vbias.n5945 Vbias.n1624 120.472
R7526 Vbias.n5924 Vbias.n1617 120.472
R7527 Vbias.n5951 Vbias.n1617 120.472
R7528 Vbias.n5923 Vbias.n1615 120.472
R7529 Vbias.n5953 Vbias.n1615 120.472
R7530 Vbias.n1520 Vbias.n1511 120.472
R7531 Vbias.n6106 Vbias.n1520 120.472
R7532 Vbias.n6116 Vbias.n1512 120.472
R7533 Vbias.n6117 Vbias.n6116 120.472
R7534 Vbias.n2000 Vbias.n1999 120.472
R7535 Vbias.n1999 Vbias.n1990 120.472
R7536 Vbias.n2008 Vbias.n1985 120.472
R7537 Vbias.n2008 Vbias.n2007 120.472
R7538 Vbias.n1960 Vbias.n1951 120.472
R7539 Vbias.n1966 Vbias.n1960 120.472
R7540 Vbias.n1976 Vbias.n1952 120.472
R7541 Vbias.n1977 Vbias.n1976 120.472
R7542 Vbias.n1926 Vbias.n1917 120.472
R7543 Vbias.n1932 Vbias.n1926 120.472
R7544 Vbias.n1942 Vbias.n1918 120.472
R7545 Vbias.n1943 Vbias.n1942 120.472
R7546 Vbias.n1801 Vbias.n1800 120.472
R7547 Vbias.n1801 Vbias.n1763 120.472
R7548 Vbias.n1762 Vbias.n1755 120.472
R7549 Vbias.n1815 Vbias.n1762 120.472
R7550 Vbias.n1858 Vbias.n1849 120.472
R7551 Vbias.n1864 Vbias.n1858 120.472
R7552 Vbias.n1866 Vbias.n1850 120.472
R7553 Vbias.n1875 Vbias.n1866 120.472
R7554 Vbias.n1735 Vbias.n1729 120.472
R7555 Vbias.n1744 Vbias.n1735 120.472
R7556 Vbias.n2042 Vbias.n2041 120.472
R7557 Vbias.n2041 Vbias.n1731 120.472
R7558 Vbias.n1890 Vbias.n1884 120.472
R7559 Vbias.n1909 Vbias.n1890 120.472
R7560 Vbias.n1897 Vbias.n1896 120.472
R7561 Vbias.n1896 Vbias.n1891 120.472
R7562 Vbias.n1779 Vbias.n1550 120.472
R7563 Vbias.n6082 Vbias.n1550 120.472
R7564 Vbias.n1785 Vbias.n1548 120.472
R7565 Vbias.n6084 Vbias.n1548 120.472
R7566 Vbias.n1772 Vbias.n1542 120.472
R7567 Vbias.n6090 Vbias.n1542 120.472
R7568 Vbias.n1797 Vbias.n1540 120.472
R7569 Vbias.n6092 Vbias.n1540 120.472
R7570 Vbias.n6777 Vbias.n6776 120.472
R7571 Vbias.n6776 Vbias.n1344 120.472
R7572 Vbias.n6774 Vbias.n1431 120.472
R7573 Vbias.n6782 Vbias.n1431 120.472
R7574 Vbias.n6766 Vbias.n1426 120.472
R7575 Vbias.n6788 Vbias.n1426 120.472
R7576 Vbias.n1441 Vbias.n1424 120.472
R7577 Vbias.n6790 Vbias.n1424 120.472
R7578 Vbias.n6056 Vbias.n1412 120.472
R7579 Vbias.n6803 Vbias.n1412 120.472
R7580 Vbias.n6047 Vbias.n1406 120.472
R7581 Vbias.n6809 Vbias.n1406 120.472
R7582 Vbias.n6070 Vbias.n1404 120.472
R7583 Vbias.n6811 Vbias.n1404 120.472
R7584 Vbias.n7087 Vbias.n7086 120.472
R7585 Vbias.n7087 Vbias.n1275 120.472
R7586 Vbias.n1288 Vbias.n1280 120.472
R7587 Vbias.n1291 Vbias.n1288 120.472
R7588 Vbias.n7070 Vbias.n7069 120.472
R7589 Vbias.n7070 Vbias.n1293 120.472
R7590 Vbias.n1308 Vbias.n1299 120.472
R7591 Vbias.n1311 Vbias.n1308 120.472
R7592 Vbias.n7042 Vbias.n7041 120.472
R7593 Vbias.n7041 Vbias.n1319 120.472
R7594 Vbias.n7025 Vbias.n7024 120.472
R7595 Vbias.n7024 Vbias.n1326 120.472
R7596 Vbias.n7022 Vbias.n1336 120.472
R7597 Vbias.n1336 Vbias.n1328 120.472
R7598 Vbias.n7193 Vbias.n7192 120.472
R7599 Vbias.n7193 Vbias.n1088 120.472
R7600 Vbias.n1101 Vbias.n1093 120.472
R7601 Vbias.n1104 Vbias.n1101 120.472
R7602 Vbias.n7176 Vbias.n7175 120.472
R7603 Vbias.n7176 Vbias.n1106 120.472
R7604 Vbias.n1120 Vbias.n1112 120.472
R7605 Vbias.n1123 Vbias.n1120 120.472
R7606 Vbias.n7148 Vbias.n7147 120.472
R7607 Vbias.n7147 Vbias.n1131 120.472
R7608 Vbias.n7131 Vbias.n7130 120.472
R7609 Vbias.n7130 Vbias.n1138 120.472
R7610 Vbias.n7128 Vbias.n1148 120.472
R7611 Vbias.n1148 Vbias.n1140 120.472
R7612 Vbias.n1219 Vbias.n1085 120.472
R7613 Vbias.n1220 Vbias.n1219 120.472
R7614 Vbias.n7212 Vbias.n1079 120.472
R7615 Vbias.n7213 Vbias.n7212 120.472
R7616 Vbias.n1240 Vbias.n1239 120.472
R7617 Vbias.n1239 Vbias.n1200 120.472
R7618 Vbias.n1229 Vbias.n1228 120.472
R7619 Vbias.n1230 Vbias.n1229 120.472
R7620 Vbias.n1250 Vbias.n1187 120.472
R7621 Vbias.n1251 Vbias.n1250 120.472
R7622 Vbias.n1271 Vbias.n1270 120.472
R7623 Vbias.n1270 Vbias.n1172 120.472
R7624 Vbias.n1260 Vbias.n1259 120.472
R7625 Vbias.n1261 Vbias.n1260 120.472
R7626 Vbias.n6952 Vbias.n1166 120.472
R7627 Vbias.n6953 Vbias.n6952 120.472
R7628 Vbias.n7108 Vbias.n1160 120.472
R7629 Vbias.n7109 Vbias.n7108 120.472
R7630 Vbias.n6973 Vbias.n6972 120.472
R7631 Vbias.n6972 Vbias.n6933 120.472
R7632 Vbias.n6962 Vbias.n6961 120.472
R7633 Vbias.n6963 Vbias.n6962 120.472
R7634 Vbias.n6983 Vbias.n6920 120.472
R7635 Vbias.n6984 Vbias.n6983 120.472
R7636 Vbias.n7004 Vbias.n7003 120.472
R7637 Vbias.n7003 Vbias.n6905 120.472
R7638 Vbias.n6993 Vbias.n6992 120.472
R7639 Vbias.n6994 Vbias.n6993 120.472
R7640 Vbias.n6873 Vbias.n1360 120.472
R7641 Vbias.n6874 Vbias.n6873 120.472
R7642 Vbias.n6887 Vbias.n1354 120.472
R7643 Vbias.n6888 Vbias.n6887 120.472
R7644 Vbias.n6850 Vbias.n1373 120.472
R7645 Vbias.n6851 Vbias.n6850 120.472
R7646 Vbias.n6864 Vbias.n1367 120.472
R7647 Vbias.n6865 Vbias.n6864 120.472
R7648 Vbias.n6841 Vbias.n1380 120.472
R7649 Vbias.n6842 Vbias.n6841 120.472
R7650 Vbias.n6820 Vbias.n6819 120.472
R7651 Vbias.n6819 Vbias.n1395 120.472
R7652 Vbias.n6826 Vbias.n1388 120.472
R7653 Vbias.n6827 Vbias.n6826 120.472
R7654 Vbias.n6015 Vbias.n1571 120.472
R7655 Vbias.n6016 Vbias.n6015 120.472
R7656 Vbias.n6032 Vbias.n1565 120.472
R7657 Vbias.n6033 Vbias.n6032 120.472
R7658 Vbias.n5992 Vbias.n1584 120.472
R7659 Vbias.n5993 Vbias.n5992 120.472
R7660 Vbias.n6006 Vbias.n1578 120.472
R7661 Vbias.n6007 Vbias.n6006 120.472
R7662 Vbias.n5983 Vbias.n1591 120.472
R7663 Vbias.n5984 Vbias.n5983 120.472
R7664 Vbias.n5962 Vbias.n5961 120.472
R7665 Vbias.n5961 Vbias.n1606 120.472
R7666 Vbias.n5968 Vbias.n1599 120.472
R7667 Vbias.n5969 Vbias.n5968 120.472
R7668 Vbias.n5328 Vbias.n5319 120.472
R7669 Vbias.n5361 Vbias.n5319 120.472
R7670 Vbias.n5331 Vbias.n5330 120.472
R7671 Vbias.n5330 Vbias.n5320 120.472
R7672 Vbias.n5381 Vbias.n5380 120.472
R7673 Vbias.n5380 Vbias.n5304 120.472
R7674 Vbias.n5370 Vbias.n5369 120.472
R7675 Vbias.n5371 Vbias.n5370 120.472
R7676 Vbias.n5391 Vbias.n5291 120.472
R7677 Vbias.n5392 Vbias.n5391 120.472
R7678 Vbias.n5412 Vbias.n5411 120.472
R7679 Vbias.n5411 Vbias.n5275 120.472
R7680 Vbias.n5401 Vbias.n5400 120.472
R7681 Vbias.n5402 Vbias.n5401 120.472
R7682 Vbias.n5242 Vbias.n2308 120.472
R7683 Vbias.n5243 Vbias.n5242 120.472
R7684 Vbias.n5256 Vbias.n2302 120.472
R7685 Vbias.n5257 Vbias.n5256 120.472
R7686 Vbias.n5219 Vbias.n2321 120.472
R7687 Vbias.n5220 Vbias.n5219 120.472
R7688 Vbias.n5233 Vbias.n2315 120.472
R7689 Vbias.n5234 Vbias.n5233 120.472
R7690 Vbias.n5210 Vbias.n2328 120.472
R7691 Vbias.n5211 Vbias.n5210 120.472
R7692 Vbias.n5189 Vbias.n5188 120.472
R7693 Vbias.n5188 Vbias.n2343 120.472
R7694 Vbias.n5195 Vbias.n2336 120.472
R7695 Vbias.n5196 Vbias.n5195 120.472
R7696 Vbias.n2496 Vbias.n2487 120.472
R7697 Vbias.n2529 Vbias.n2487 120.472
R7698 Vbias.n2499 Vbias.n2498 120.472
R7699 Vbias.n2498 Vbias.n2488 120.472
R7700 Vbias.n2549 Vbias.n2548 120.472
R7701 Vbias.n2548 Vbias.n2472 120.472
R7702 Vbias.n2538 Vbias.n2537 120.472
R7703 Vbias.n2539 Vbias.n2538 120.472
R7704 Vbias.n2559 Vbias.n2459 120.472
R7705 Vbias.n2560 Vbias.n2559 120.472
R7706 Vbias.n2580 Vbias.n2579 120.472
R7707 Vbias.n2579 Vbias.n2443 120.472
R7708 Vbias.n2569 Vbias.n2568 120.472
R7709 Vbias.n2570 Vbias.n2569 120.472
R7710 Vbias.n5046 Vbias.n5045 120.472
R7711 Vbias.n5045 Vbias.n2420 120.472
R7712 Vbias.n5043 Vbias.n2430 120.472
R7713 Vbias.n2430 Vbias.n2422 120.472
R7714 Vbias.n4419 Vbias.n4410 120.472
R7715 Vbias.n4546 Vbias.n4410 120.472
R7716 Vbias.n4422 Vbias.n4421 120.472
R7717 Vbias.n4421 Vbias.n4411 120.472
R7718 Vbias.n3844 Vbias.n3814 120.472
R7719 Vbias.n3819 Vbias.n3814 120.472
R7720 Vbias.n3822 Vbias.n3821 120.472
R7721 Vbias.n3828 Vbias.n3822 120.472
R7722 Vbias.n3834 Vbias.n3830 120.472
R7723 Vbias.n3835 Vbias.n3834 120.472
R7724 Vbias.n3812 Vbias.n3811 120.472
R7725 Vbias.n3811 Vbias.n3809 120.472
R7726 Vbias.n3859 Vbias.n3781 120.472
R7727 Vbias.n3872 Vbias.n3859 120.472
R7728 Vbias.n3883 Vbias.n3783 120.472
R7729 Vbias.n3884 Vbias.n3883 120.472
R7730 Vbias.n3920 Vbias.n3767 120.472
R7731 Vbias.n3895 Vbias.n3767 120.472
R7732 Vbias.n3898 Vbias.n3897 120.472
R7733 Vbias.n3904 Vbias.n3898 120.472
R7734 Vbias.n3910 Vbias.n3906 120.472
R7735 Vbias.n3911 Vbias.n3910 120.472
R7736 Vbias.n3765 Vbias.n3764 120.472
R7737 Vbias.n3764 Vbias.n3762 120.472
R7738 Vbias.n3958 Vbias.n3738 120.472
R7739 Vbias.n3933 Vbias.n3738 120.472
R7740 Vbias.n3936 Vbias.n3935 120.472
R7741 Vbias.n3942 Vbias.n3936 120.472
R7742 Vbias.n3948 Vbias.n3944 120.472
R7743 Vbias.n3949 Vbias.n3948 120.472
R7744 Vbias.n3736 Vbias.n3735 120.472
R7745 Vbias.n3735 Vbias.n3733 120.472
R7746 Vbias.n3306 Vbias.n3276 120.472
R7747 Vbias.n3281 Vbias.n3276 120.472
R7748 Vbias.n3284 Vbias.n3283 120.472
R7749 Vbias.n3290 Vbias.n3284 120.472
R7750 Vbias.n3296 Vbias.n3292 120.472
R7751 Vbias.n3297 Vbias.n3296 120.472
R7752 Vbias.n3274 Vbias.n3273 120.472
R7753 Vbias.n3273 Vbias.n3271 120.472
R7754 Vbias.n3321 Vbias.n3243 120.472
R7755 Vbias.n3334 Vbias.n3321 120.472
R7756 Vbias.n3345 Vbias.n3245 120.472
R7757 Vbias.n3346 Vbias.n3345 120.472
R7758 Vbias.n3382 Vbias.n3229 120.472
R7759 Vbias.n3357 Vbias.n3229 120.472
R7760 Vbias.n3360 Vbias.n3359 120.472
R7761 Vbias.n3366 Vbias.n3360 120.472
R7762 Vbias.n3372 Vbias.n3368 120.472
R7763 Vbias.n3373 Vbias.n3372 120.472
R7764 Vbias.n3227 Vbias.n3226 120.472
R7765 Vbias.n3226 Vbias.n3224 120.472
R7766 Vbias.n3420 Vbias.n3200 120.472
R7767 Vbias.n3395 Vbias.n3200 120.472
R7768 Vbias.n3398 Vbias.n3397 120.472
R7769 Vbias.n3404 Vbias.n3398 120.472
R7770 Vbias.n3410 Vbias.n3406 120.472
R7771 Vbias.n3411 Vbias.n3410 120.472
R7772 Vbias.n3198 Vbias.n3197 120.472
R7773 Vbias.n3197 Vbias.n3195 120.472
R7774 Vbias.n3575 Vbias.n3545 120.472
R7775 Vbias.n3550 Vbias.n3545 120.472
R7776 Vbias.n3553 Vbias.n3552 120.472
R7777 Vbias.n3559 Vbias.n3553 120.472
R7778 Vbias.n3565 Vbias.n3561 120.472
R7779 Vbias.n3566 Vbias.n3565 120.472
R7780 Vbias.n3543 Vbias.n3542 120.472
R7781 Vbias.n3542 Vbias.n3540 120.472
R7782 Vbias.n3590 Vbias.n3512 120.472
R7783 Vbias.n3603 Vbias.n3590 120.472
R7784 Vbias.n3614 Vbias.n3514 120.472
R7785 Vbias.n3615 Vbias.n3614 120.472
R7786 Vbias.n3651 Vbias.n3498 120.472
R7787 Vbias.n3626 Vbias.n3498 120.472
R7788 Vbias.n3629 Vbias.n3628 120.472
R7789 Vbias.n3635 Vbias.n3629 120.472
R7790 Vbias.n3641 Vbias.n3637 120.472
R7791 Vbias.n3642 Vbias.n3641 120.472
R7792 Vbias.n3496 Vbias.n3495 120.472
R7793 Vbias.n3495 Vbias.n3493 120.472
R7794 Vbias.n3689 Vbias.n3469 120.472
R7795 Vbias.n3664 Vbias.n3469 120.472
R7796 Vbias.n3667 Vbias.n3666 120.472
R7797 Vbias.n3673 Vbias.n3667 120.472
R7798 Vbias.n3679 Vbias.n3675 120.472
R7799 Vbias.n3680 Vbias.n3679 120.472
R7800 Vbias.n3467 Vbias.n3466 120.472
R7801 Vbias.n3466 Vbias.n3464 120.472
R7802 Vbias.n4190 Vbias.n4068 120.472
R7803 Vbias.n4068 Vbias.n4055 120.472
R7804 Vbias.n4066 Vbias.n4065 120.472
R7805 Vbias.n4065 Vbias.n4052 120.472
R7806 Vbias.n4209 Vbias.n4041 120.472
R7807 Vbias.n4210 Vbias.n4209 120.472
R7808 Vbias.n4224 Vbias.n4026 120.472
R7809 Vbias.n4026 Vbias.n4013 120.472
R7810 Vbias.n4024 Vbias.n4023 120.472
R7811 Vbias.n4023 Vbias.n4010 120.472
R7812 Vbias.n3999 Vbias.n3992 120.472
R7813 Vbias.n4240 Vbias.n3999 120.472
R7814 Vbias.n4245 Vbias.n3991 120.472
R7815 Vbias.n3991 Vbias.n3982 120.472
R7816 Vbias.n4178 Vbias.n4167 120.472
R7817 Vbias.n4170 Vbias.n4167 120.472
R7818 Vbias.n4078 Vbias.n4077 120.472
R7819 Vbias.n4077 Vbias.n4074 120.472
R7820 Vbias.n4145 Vbias.n4144 120.472
R7821 Vbias.n4160 Vbias.n4145 120.472
R7822 Vbias.n4088 Vbias.n4085 120.472
R7823 Vbias.n4135 Vbias.n4085 120.472
R7824 Vbias.n4084 Vbias.n4080 120.472
R7825 Vbias.n4137 Vbias.n4084 120.472
R7826 Vbias.n4100 Vbias.n4098 120.472
R7827 Vbias.n4119 Vbias.n4098 120.472
R7828 Vbias.n4094 Vbias.n4090 120.472
R7829 Vbias.n4121 Vbias.n4094 120.472
R7830 Vbias.n4974 Vbias.n4973 120.472
R7831 Vbias.n4973 Vbias.n2612 120.472
R7832 Vbias.n4980 Vbias.n2605 120.472
R7833 Vbias.n4981 Vbias.n4980 120.472
R7834 Vbias.n4962 Vbias.n2619 120.472
R7835 Vbias.n4963 Vbias.n4962 120.472
R7836 Vbias.n4936 Vbias.n2642 120.472
R7837 Vbias.n4937 Vbias.n4936 120.472
R7838 Vbias.n4950 Vbias.n2636 120.472
R7839 Vbias.n4951 Vbias.n4950 120.472
R7840 Vbias.n4914 Vbias.n2656 120.472
R7841 Vbias.n4915 Vbias.n4914 120.472
R7842 Vbias.n4927 Vbias.n2650 120.472
R7843 Vbias.n4928 Vbias.n4927 120.472
R7844 Vbias.n3036 Vbias.n3006 120.472
R7845 Vbias.n3011 Vbias.n3006 120.472
R7846 Vbias.n3014 Vbias.n3013 120.472
R7847 Vbias.n3020 Vbias.n3014 120.472
R7848 Vbias.n3026 Vbias.n3022 120.472
R7849 Vbias.n3027 Vbias.n3026 120.472
R7850 Vbias.n3004 Vbias.n3003 120.472
R7851 Vbias.n3003 Vbias.n3001 120.472
R7852 Vbias.n3051 Vbias.n2973 120.472
R7853 Vbias.n3064 Vbias.n3051 120.472
R7854 Vbias.n3075 Vbias.n2975 120.472
R7855 Vbias.n3076 Vbias.n3075 120.472
R7856 Vbias.n3112 Vbias.n2959 120.472
R7857 Vbias.n3087 Vbias.n2959 120.472
R7858 Vbias.n3090 Vbias.n3089 120.472
R7859 Vbias.n3096 Vbias.n3090 120.472
R7860 Vbias.n3102 Vbias.n3098 120.472
R7861 Vbias.n3103 Vbias.n3102 120.472
R7862 Vbias.n2957 Vbias.n2956 120.472
R7863 Vbias.n2956 Vbias.n2954 120.472
R7864 Vbias.n3150 Vbias.n2930 120.472
R7865 Vbias.n3125 Vbias.n2930 120.472
R7866 Vbias.n3128 Vbias.n3127 120.472
R7867 Vbias.n3134 Vbias.n3128 120.472
R7868 Vbias.n3140 Vbias.n3136 120.472
R7869 Vbias.n3141 Vbias.n3140 120.472
R7870 Vbias.n2928 Vbias.n2927 120.472
R7871 Vbias.n2927 Vbias.n2925 120.472
R7872 Vbias.n4712 Vbias.n2767 120.472
R7873 Vbias.n4687 Vbias.n2767 120.472
R7874 Vbias.n4690 Vbias.n4689 120.472
R7875 Vbias.n4696 Vbias.n4690 120.472
R7876 Vbias.n4702 Vbias.n4698 120.472
R7877 Vbias.n4703 Vbias.n4702 120.472
R7878 Vbias.n2765 Vbias.n2764 120.472
R7879 Vbias.n2764 Vbias.n2762 120.472
R7880 Vbias.n4727 Vbias.n2734 120.472
R7881 Vbias.n4740 Vbias.n4727 120.472
R7882 Vbias.n4751 Vbias.n2736 120.472
R7883 Vbias.n4752 Vbias.n4751 120.472
R7884 Vbias.n4788 Vbias.n2720 120.472
R7885 Vbias.n4763 Vbias.n2720 120.472
R7886 Vbias.n4766 Vbias.n4765 120.472
R7887 Vbias.n4772 Vbias.n4766 120.472
R7888 Vbias.n4778 Vbias.n4774 120.472
R7889 Vbias.n4779 Vbias.n4778 120.472
R7890 Vbias.n2718 Vbias.n2717 120.472
R7891 Vbias.n2717 Vbias.n2715 120.472
R7892 Vbias.n4826 Vbias.n2691 120.472
R7893 Vbias.n4801 Vbias.n2691 120.472
R7894 Vbias.n4804 Vbias.n4803 120.472
R7895 Vbias.n4810 Vbias.n4804 120.472
R7896 Vbias.n4816 Vbias.n4812 120.472
R7897 Vbias.n4817 Vbias.n4816 120.472
R7898 Vbias.n2689 Vbias.n2688 120.472
R7899 Vbias.n2688 Vbias.n2686 120.472
R7900 Vbias.n4567 Vbias.n4557 120.472
R7901 Vbias.n4675 Vbias.n4557 120.472
R7902 Vbias.n4566 Vbias.n4565 120.472
R7903 Vbias.n4565 Vbias.n4554 120.472
R7904 Vbias.n5653 Vbias.n2209 120.472
R7905 Vbias.n2209 Vbias.n2204 120.472
R7906 Vbias.n2203 Vbias.n2196 120.472
R7907 Vbias.n5658 Vbias.n2203 120.472
R7908 Vbias.n2225 Vbias.n2213 120.472
R7909 Vbias.n5644 Vbias.n2225 120.472
R7910 Vbias.n5568 Vbias.n5567 120.472
R7911 Vbias.n5567 Vbias.n5558 120.472
R7912 Vbias.n5629 Vbias.n5557 120.472
R7913 Vbias.n5634 Vbias.n5557 120.472
R7914 Vbias.n5586 Vbias.n5585 120.472
R7915 Vbias.n5585 Vbias.n5576 120.472
R7916 Vbias.n5610 Vbias.n5575 120.472
R7917 Vbias.n5615 Vbias.n5575 120.472
R7918 Vbias.n5727 Vbias.n2138 120.472
R7919 Vbias.n2138 Vbias.n2133 120.472
R7920 Vbias.n2132 Vbias.n2125 120.472
R7921 Vbias.n5732 Vbias.n2132 120.472
R7922 Vbias.n2154 Vbias.n2142 120.472
R7923 Vbias.n5718 Vbias.n2154 120.472
R7924 Vbias.n2171 Vbias.n2170 120.472
R7925 Vbias.n2170 Vbias.n2161 120.472
R7926 Vbias.n5703 Vbias.n2160 120.472
R7927 Vbias.n5708 Vbias.n2160 120.472
R7928 Vbias.n2189 Vbias.n2188 120.472
R7929 Vbias.n2188 Vbias.n2179 120.472
R7930 Vbias.n5684 Vbias.n2178 120.472
R7931 Vbias.n5689 Vbias.n2178 120.472
R7932 Vbias.n5816 Vbias.n2083 120.472
R7933 Vbias.n2083 Vbias.n2078 120.472
R7934 Vbias.n2077 Vbias.n2070 120.472
R7935 Vbias.n5821 Vbias.n2077 120.472
R7936 Vbias.n5799 Vbias.n5787 120.472
R7937 Vbias.n5807 Vbias.n5799 120.472
R7938 Vbias.n5773 Vbias.n2099 120.472
R7939 Vbias.n2099 Vbias.n2092 120.472
R7940 Vbias.n2091 Vbias.n2087 120.472
R7941 Vbias.n5778 Vbias.n2091 120.472
R7942 Vbias.n5759 Vbias.n2121 120.472
R7943 Vbias.n2121 Vbias.n2116 120.472
R7944 Vbias.n2115 Vbias.n2103 120.472
R7945 Vbias.n5764 Vbias.n2115 120.472
R7946 Vbias.n6662 Vbias.n1484 120.472
R7947 Vbias.n1496 Vbias.n1484 120.472
R7948 Vbias.n1498 Vbias.n1485 120.472
R7949 Vbias.n6657 Vbias.n1498 120.472
R7950 Vbias.n1479 Vbias.n1471 120.472
R7951 Vbias.n6671 Vbias.n1471 120.472
R7952 Vbias.n2063 Vbias.n1698 120.472
R7953 Vbias.n5848 Vbias.n2063 120.472
R7954 Vbias.n5855 Vbias.n1700 120.472
R7955 Vbias.n5850 Vbias.n1700 120.472
R7956 Vbias.n6241 Vbias.n6240 120.472
R7957 Vbias.n6240 Vbias.n6231 120.472
R7958 Vbias.n6580 Vbias.n6230 120.472
R7959 Vbias.n6585 Vbias.n6230 120.472
R7960 Vbias.n6256 Vbias.n6248 120.472
R7961 Vbias.n6348 Vbias.n6248 120.472
R7962 Vbias.n6330 Vbias.n6272 120.472
R7963 Vbias.n6272 Vbias.n6267 120.472
R7964 Vbias.n6266 Vbias.n6258 120.472
R7965 Vbias.n6335 Vbias.n6266 120.472
R7966 Vbias.n6316 Vbias.n6294 120.472
R7967 Vbias.n6294 Vbias.n6289 120.472
R7968 Vbias.n6288 Vbias.n6276 120.472
R7969 Vbias.n6321 Vbias.n6288 120.472
R7970 Vbias.n7601 Vbias.n839 120.472
R7971 Vbias.n852 Vbias.n839 120.472
R7972 Vbias.n854 Vbias.n840 120.472
R7973 Vbias.n7596 Vbias.n854 120.472
R7974 Vbias.n833 Vbias.n825 120.472
R7975 Vbias.n7610 Vbias.n825 120.472
R7976 Vbias.n812 Vbias.n803 120.472
R7977 Vbias.n7625 Vbias.n803 120.472
R7978 Vbias.n7620 Vbias.n817 120.472
R7979 Vbias.n817 Vbias.n804 120.472
R7980 Vbias.n793 Vbias.n784 120.472
R7981 Vbias.n7640 Vbias.n784 120.472
R7982 Vbias.n7635 Vbias.n796 120.472
R7983 Vbias.n796 Vbias.n785 120.472
R7984 Vbias.n7479 Vbias.n994 120.472
R7985 Vbias.n1007 Vbias.n994 120.472
R7986 Vbias.n1009 Vbias.n995 120.472
R7987 Vbias.n7474 Vbias.n1009 120.472
R7988 Vbias.n988 Vbias.n980 120.472
R7989 Vbias.n7488 Vbias.n980 120.472
R7990 Vbias.n967 Vbias.n958 120.472
R7991 Vbias.n7504 Vbias.n958 120.472
R7992 Vbias.n7499 Vbias.n972 120.472
R7993 Vbias.n972 Vbias.n959 120.472
R7994 Vbias.n944 Vbias.n935 120.472
R7995 Vbias.n7519 Vbias.n935 120.472
R7996 Vbias.n7514 Vbias.n951 120.472
R7997 Vbias.n951 Vbias.n936 120.472
R7998 Vbias.n6219 Vbias.n6209 120.472
R7999 Vbias.n6603 Vbias.n6209 120.472
R8000 Vbias.n6218 Vbias.n6217 120.472
R8001 Vbias.n6217 Vbias.n6205 120.472
R8002 Vbias.n6199 Vbias.n6198 120.472
R8003 Vbias.n6199 Vbias.n6191 120.472
R8004 Vbias.n6181 Vbias.n6159 120.472
R8005 Vbias.n6629 Vbias.n6159 120.472
R8006 Vbias.n6167 Vbias.n6157 120.472
R8007 Vbias.n6631 Vbias.n6157 120.472
R8008 Vbias.n6456 Vbias.n6446 120.472
R8009 Vbias.n6536 Vbias.n6446 120.472
R8010 Vbias.n6455 Vbias.n6454 120.472
R8011 Vbias.n6454 Vbias.n6442 120.472
R8012 Vbias.n6436 Vbias.n6435 120.472
R8013 Vbias.n6436 Vbias.n6428 120.472
R8014 Vbias.n6418 Vbias.n6377 120.472
R8015 Vbias.n6562 Vbias.n6377 120.472
R8016 Vbias.n6385 Vbias.n6375 120.472
R8017 Vbias.n6564 Vbias.n6375 120.472
R8018 Vbias.n6401 Vbias.n6369 120.472
R8019 Vbias.n6570 Vbias.n6369 120.472
R8020 Vbias.n6388 Vbias.n6367 120.472
R8021 Vbias.n6572 Vbias.n6367 120.472
R8022 Vbias.n910 Vbias.n900 120.472
R8023 Vbias.n7549 Vbias.n900 120.472
R8024 Vbias.n909 Vbias.n908 120.472
R8025 Vbias.n908 Vbias.n896 120.472
R8026 Vbias.n890 Vbias.n889 120.472
R8027 Vbias.n890 Vbias.n882 120.472
R8028 Vbias.n6470 Vbias.n872 120.472
R8029 Vbias.n7575 Vbias.n872 120.472
R8030 Vbias.n6486 Vbias.n870 120.472
R8031 Vbias.n7577 Vbias.n870 120.472
R8032 Vbias.n6464 Vbias.n864 120.472
R8033 Vbias.n7583 Vbias.n864 120.472
R8034 Vbias.n6500 Vbias.n862 120.472
R8035 Vbias.n7585 Vbias.n862 120.472
R8036 Vbias.n7405 Vbias.n7397 120.472
R8037 Vbias.n7397 Vbias.n7386 120.472
R8038 Vbias.n7395 Vbias.n7394 120.472
R8039 Vbias.n7394 Vbias.n7383 120.472
R8040 Vbias.n7424 Vbias.n7371 120.472
R8041 Vbias.n7425 Vbias.n7424 120.472
R8042 Vbias.n7439 Vbias.n7359 120.472
R8043 Vbias.n7359 Vbias.n7348 120.472
R8044 Vbias.n7357 Vbias.n7356 120.472
R8045 Vbias.n7356 Vbias.n7345 120.472
R8046 Vbias.n7338 Vbias.n7333 120.472
R8047 Vbias.n7455 Vbias.n7338 120.472
R8048 Vbias.n7460 Vbias.n7332 120.472
R8049 Vbias.n7332 Vbias.n7326 120.472
R8050 Vbias.n6640 Vbias.n6147 120.472
R8051 Vbias.n6153 Vbias.n6147 120.472
R8052 Vbias.n6645 Vbias.n6138 120.472
R8053 Vbias.n6646 Vbias.n6645 120.472
R8054 Vbias.n7273 Vbias.n7244 120.472
R8055 Vbias.n7257 Vbias.n7244 120.472
R8056 Vbias.n7259 Vbias.n7245 120.472
R8057 Vbias.n7268 Vbias.n7259 120.472
R8058 Vbias.n7238 Vbias.n7230 120.472
R8059 Vbias.n7282 Vbias.n7230 120.472
R8060 Vbias.n1062 Vbias.n1053 120.472
R8061 Vbias.n7297 Vbias.n1053 120.472
R8062 Vbias.n7292 Vbias.n1067 120.472
R8063 Vbias.n1067 Vbias.n1054 120.472
R8064 Vbias.n1041 Vbias.n1032 120.472
R8065 Vbias.n7312 Vbias.n1032 120.472
R8066 Vbias.n7307 Vbias.n1046 120.472
R8067 Vbias.n1046 Vbias.n1033 120.472
R8068 Vbias.n7726 Vbias.n695 120.472
R8069 Vbias.n695 Vbias.n685 120.472
R8070 Vbias.n693 Vbias.n683 120.472
R8071 Vbias.n7731 Vbias.n683 120.472
R8072 Vbias.n1714 Vbias.n1707 120.472
R8073 Vbias.n2055 Vbias.n1707 120.472
R8074 Vbias.n1721 Vbias.n1715 120.472
R8075 Vbias.n1721 Vbias.n1708 120.472
R8076 Vbias.n6684 Vbias.n6683 120.472
R8077 Vbias.n6684 Vbias.n1450 120.472
R8078 Vbias.n5867 Vbias.n1684 120.472
R8079 Vbias.n5868 Vbias.n5867 120.472
R8080 Vbias.n5522 Vbias.n5521 120.472
R8081 Vbias.n5521 Vbias.n5512 120.472
R8082 Vbias.n5543 Vbias.n2237 120.472
R8083 Vbias.n5544 Vbias.n5543 120.472
R8084 Vbias.n5024 Vbias.n2589 120.472
R8085 Vbias.n5025 Vbias.n5024 120.472
R8086 Vbias.n8066 Vbias.n26 120.472
R8087 Vbias.n26 Vbias.n16 120.472
R8088 Vbias.n24 Vbias.n14 120.472
R8089 Vbias.n8071 Vbias.n14 120.472
R8090 Vbias.t777 Vbias.t557 119.632
R8091 Vbias.n1724 Vbias.n1723 119.632
R8092 Vbias.t670 Vbias.t559 119.632
R8093 Vbias.n2039 Vbias.n1725 119.632
R8094 Vbias.n342 Vbias.n341 119.019
R8095 Vbias.n567 Vbias.n566 119.019
R8096 Vbias.n4900 Vbias.n4891 118.564
R8097 Vbias.n6261 Vbias.n1444 118.349
R8098 Vbias.n7494 Vbias.n7493 118.349
R8099 Vbias.n4883 Vbias.n4882 117.001
R8100 Vbias.t470 Vbias.n4883 117.001
R8101 Vbias.n4850 Vbias.n4848 117.001
R8102 Vbias.t472 Vbias.n4848 117.001
R8103 Vbias.n4885 Vbias.n4884 117.001
R8104 Vbias.n4884 Vbias.t470 117.001
R8105 Vbias.n4887 Vbias.n4849 117.001
R8106 Vbias.t472 Vbias.n4849 117.001
R8107 Vbias.n4874 Vbias.n4873 117.001
R8108 Vbias.n4873 Vbias.t548 117.001
R8109 Vbias.n4877 Vbias.n4876 117.001
R8110 Vbias.t893 Vbias.n4877 117.001
R8111 Vbias.n4867 Vbias.n4866 117.001
R8112 Vbias.n4867 Vbias.t548 117.001
R8113 Vbias.n4864 Vbias.n4856 117.001
R8114 Vbias.t893 Vbias.n4856 117.001
R8115 Vbias.n4 Vbias.n3 117.001
R8116 Vbias.t468 Vbias.n4 117.001
R8117 Vbias.n8081 Vbias.n2 117.001
R8118 Vbias.t468 Vbias.n2 117.001
R8119 Vbias.n37 Vbias.n29 116.663
R8120 Vbias.n56 Vbias.n47 116.663
R8121 Vbias.n8040 Vbias.n8039 116.663
R8122 Vbias.n8025 Vbias.n8024 116.663
R8123 Vbias.n81 Vbias.n68 115.576
R8124 Vbias.n8015 Vbias.n81 115.576
R8125 Vbias.n8015 Vbias.n8014 115.576
R8126 Vbias.n8014 Vbias.n8013 115.576
R8127 Vbias.n8029 Vbias.n59 115.576
R8128 Vbias.n8030 Vbias.n8029 115.576
R8129 Vbias.n39 Vbias.n34 115.576
R8130 Vbias.n8052 Vbias.n34 115.576
R8131 Vbias.n8052 Vbias.n8051 115.576
R8132 Vbias.n8051 Vbias.n8050 115.576
R8133 Vbias.n4372 Vbias.n4371 115.576
R8134 Vbias.n4372 Vbias.n2785 115.576
R8135 Vbias.n2785 Vbias.n2782 115.576
R8136 Vbias.n4401 Vbias.n2782 115.576
R8137 Vbias.n4368 Vbias.n2794 115.576
R8138 Vbias.n4396 Vbias.n2794 115.576
R8139 Vbias.n4396 Vbias.n4395 115.576
R8140 Vbias.n4395 Vbias.n2780 115.576
R8141 Vbias.n4349 Vbias.n4346 115.576
R8142 Vbias.n4349 Vbias.n4348 115.576
R8143 Vbias.n4340 Vbias.n2814 115.576
R8144 Vbias.n2814 Vbias.n2805 115.576
R8145 Vbias.n4309 Vbias.n4308 115.576
R8146 Vbias.n4310 Vbias.n4309 115.576
R8147 Vbias.n4314 Vbias.n4310 115.576
R8148 Vbias.n4314 Vbias.n4313 115.576
R8149 Vbias.n4305 Vbias.n2838 115.576
R8150 Vbias.n4325 Vbias.n2838 115.576
R8151 Vbias.n4326 Vbias.n4325 115.576
R8152 Vbias.n4328 Vbias.n4326 115.576
R8153 Vbias.n4276 Vbias.n4275 115.576
R8154 Vbias.n4277 Vbias.n4276 115.576
R8155 Vbias.n4281 Vbias.n4277 115.576
R8156 Vbias.n4281 Vbias.n4280 115.576
R8157 Vbias.n4272 Vbias.n2872 115.576
R8158 Vbias.n4292 Vbias.n2872 115.576
R8159 Vbias.n4293 Vbias.n4292 115.576
R8160 Vbias.n4295 Vbias.n4293 115.576
R8161 Vbias.n4999 Vbias.n4998 115.576
R8162 Vbias.n4998 Vbias.n2595 115.576
R8163 Vbias.n6704 Vbias.n6703 115.576
R8164 Vbias.n6703 Vbias.n6699 115.576
R8165 Vbias.n6730 Vbias.n6729 115.576
R8166 Vbias.n6729 Vbias.n6723 115.576
R8167 Vbias.n7741 Vbias.n670 115.576
R8168 Vbias.n7742 Vbias.n7741 115.576
R8169 Vbias.n569 Vbias.n562 115.576
R8170 Vbias.n7807 Vbias.n562 115.576
R8171 Vbias.n7876 Vbias.n450 115.576
R8172 Vbias.n7877 Vbias.n7876 115.576
R8173 Vbias.n336 Vbias.n335 115.576
R8174 Vbias.n335 Vbias.n172 115.576
R8175 Vbias.n1014 Vbias.n920 115.576
R8176 Vbias.n1023 Vbias.n920 115.576
R8177 Vbias.n6529 Vbias.n6528 115.576
R8178 Vbias.n6528 Vbias.n927 115.576
R8179 Vbias.n6593 Vbias.n6592 115.576
R8180 Vbias.n6592 Vbias.n776 115.576
R8181 Vbias.n7666 Vbias.n7665 115.576
R8182 Vbias.n7665 Vbias.n7664 115.576
R8183 Vbias.n750 Vbias.n737 115.576
R8184 Vbias.n7675 Vbias.n750 115.576
R8185 Vbias.n7675 Vbias.n7674 115.576
R8186 Vbias.n7674 Vbias.n7673 115.576
R8187 Vbias.n7689 Vbias.n728 115.576
R8188 Vbias.n7690 Vbias.n7689 115.576
R8189 Vbias.n708 Vbias.n703 115.576
R8190 Vbias.n7712 Vbias.n703 115.576
R8191 Vbias.n7712 Vbias.n7711 115.576
R8192 Vbias.n7711 Vbias.n7710 115.576
R8193 Vbias.n659 Vbias.n645 115.576
R8194 Vbias.n661 Vbias.n659 115.576
R8195 Vbias.n661 Vbias.n660 115.576
R8196 Vbias.n660 Vbias.n652 115.576
R8197 Vbias.n637 Vbias.n636 115.576
R8198 Vbias.n636 Vbias.n630 115.576
R8199 Vbias.n612 Vbias.n598 115.576
R8200 Vbias.n614 Vbias.n612 115.576
R8201 Vbias.n614 Vbias.n613 115.576
R8202 Vbias.n613 Vbias.n605 115.576
R8203 Vbias.n588 Vbias.n574 115.576
R8204 Vbias.n590 Vbias.n588 115.576
R8205 Vbias.n590 Vbias.n589 115.576
R8206 Vbias.n589 Vbias.n581 115.576
R8207 Vbias.n545 Vbias.n531 115.576
R8208 Vbias.n547 Vbias.n545 115.576
R8209 Vbias.n547 Vbias.n546 115.576
R8210 Vbias.n546 Vbias.n538 115.576
R8211 Vbias.n523 Vbias.n522 115.576
R8212 Vbias.n522 Vbias.n516 115.576
R8213 Vbias.n498 Vbias.n484 115.576
R8214 Vbias.n500 Vbias.n498 115.576
R8215 Vbias.n500 Vbias.n499 115.576
R8216 Vbias.n499 Vbias.n491 115.576
R8217 Vbias.n474 Vbias.n460 115.576
R8218 Vbias.n476 Vbias.n474 115.576
R8219 Vbias.n476 Vbias.n475 115.576
R8220 Vbias.n475 Vbias.n467 115.576
R8221 Vbias.n439 Vbias.n425 115.576
R8222 Vbias.n441 Vbias.n439 115.576
R8223 Vbias.n441 Vbias.n440 115.576
R8224 Vbias.n440 Vbias.n432 115.576
R8225 Vbias.n417 Vbias.n416 115.576
R8226 Vbias.n416 Vbias.n410 115.576
R8227 Vbias.n392 Vbias.n378 115.576
R8228 Vbias.n394 Vbias.n392 115.576
R8229 Vbias.n394 Vbias.n393 115.576
R8230 Vbias.n393 Vbias.n385 115.576
R8231 Vbias.n368 Vbias.n177 115.576
R8232 Vbias.n370 Vbias.n368 115.576
R8233 Vbias.n370 Vbias.n369 115.576
R8234 Vbias.n369 Vbias.n361 115.576
R8235 Vbias.n189 Vbias.n186 115.576
R8236 Vbias.n319 Vbias.n186 115.576
R8237 Vbias.n320 Vbias.n319 115.576
R8238 Vbias.n320 Vbias.n182 115.576
R8239 Vbias.n303 Vbias.n302 115.576
R8240 Vbias.n303 Vbias.n201 115.576
R8241 Vbias.n222 Vbias.n219 115.576
R8242 Vbias.n280 Vbias.n219 115.576
R8243 Vbias.n281 Vbias.n280 115.576
R8244 Vbias.n281 Vbias.n215 115.576
R8245 Vbias.n241 Vbias.n238 115.576
R8246 Vbias.n263 Vbias.n238 115.576
R8247 Vbias.n264 Vbias.n263 115.576
R8248 Vbias.n264 Vbias.n234 115.576
R8249 Vbias.n160 Vbias.n159 115.576
R8250 Vbias.n7953 Vbias.n160 115.576
R8251 Vbias.n7953 Vbias.n7952 115.576
R8252 Vbias.n7952 Vbias.n7951 115.576
R8253 Vbias.n7967 Vbias.n7966 115.576
R8254 Vbias.n7966 Vbias.n7965 115.576
R8255 Vbias.n7982 Vbias.n7981 115.576
R8256 Vbias.n7981 Vbias.n7980 115.576
R8257 Vbias.n7980 Vbias.n113 115.576
R8258 Vbias.n7972 Vbias.n113 115.576
R8259 Vbias.n7997 Vbias.n7996 115.576
R8260 Vbias.n7996 Vbias.n7995 115.576
R8261 Vbias.n7995 Vbias.n94 115.576
R8262 Vbias.n7987 Vbias.n94 115.576
R8263 Vbias.n4636 Vbias.n4635 115.576
R8264 Vbias.n4640 Vbias.n4636 115.576
R8265 Vbias.n4640 Vbias.n4639 115.576
R8266 Vbias.n4639 Vbias.n2436 115.576
R8267 Vbias.n4620 Vbias.n4613 115.576
R8268 Vbias.n4627 Vbias.n4613 115.576
R8269 Vbias.n4628 Vbias.n4627 115.576
R8270 Vbias.n4629 Vbias.n4628 115.576
R8271 Vbias.n4585 Vbias.n4576 115.576
R8272 Vbias.n4585 Vbias.n4581 115.576
R8273 Vbias.n4477 Vbias.n4476 115.576
R8274 Vbias.n4503 Vbias.n4477 115.576
R8275 Vbias.n4503 Vbias.n4502 115.576
R8276 Vbias.n4502 Vbias.n4501 115.576
R8277 Vbias.n4455 Vbias.n4454 115.576
R8278 Vbias.n4517 Vbias.n4455 115.576
R8279 Vbias.n4517 Vbias.n4516 115.576
R8280 Vbias.n4516 Vbias.n4515 115.576
R8281 Vbias.n4531 Vbias.n4530 115.576
R8282 Vbias.n4530 Vbias.n4529 115.576
R8283 Vbias.n5106 Vbias.n5105 115.576
R8284 Vbias.n5110 Vbias.n5106 115.576
R8285 Vbias.n5110 Vbias.n5109 115.576
R8286 Vbias.n5109 Vbias.n2374 115.576
R8287 Vbias.n5086 Vbias.n5085 115.576
R8288 Vbias.n5090 Vbias.n5086 115.576
R8289 Vbias.n5090 Vbias.n5089 115.576
R8290 Vbias.n5089 Vbias.n2390 115.576
R8291 Vbias.n5062 Vbias.n5061 115.576
R8292 Vbias.n5062 Vbias.n2410 115.576
R8293 Vbias.n2280 Vbias.n2267 115.576
R8294 Vbias.n2282 Vbias.n2280 115.576
R8295 Vbias.n2282 Vbias.n2281 115.576
R8296 Vbias.n2281 Vbias.n2273 115.576
R8297 Vbias.n5154 Vbias.n2248 115.576
R8298 Vbias.n2260 Vbias.n2248 115.576
R8299 Vbias.n2261 Vbias.n2260 115.576
R8300 Vbias.n2261 Vbias.n2255 115.576
R8301 Vbias.n5143 Vbias.n5142 115.576
R8302 Vbias.n5142 Vbias.n2362 115.576
R8303 Vbias.n5125 Vbias.n2365 115.576
R8304 Vbias.n5134 Vbias.n2365 115.576
R8305 Vbias.n5135 Vbias.n5134 115.576
R8306 Vbias.n5136 Vbias.n5135 115.576
R8307 Vbias.n5903 Vbias.n5902 115.576
R8308 Vbias.n5907 Vbias.n5903 115.576
R8309 Vbias.n5907 Vbias.n5906 115.576
R8310 Vbias.n5906 Vbias.n1642 115.576
R8311 Vbias.n5883 Vbias.n5882 115.576
R8312 Vbias.n5887 Vbias.n5883 115.576
R8313 Vbias.n5887 Vbias.n5886 115.576
R8314 Vbias.n5886 Vbias.n1658 115.576
R8315 Vbias.n5447 Vbias.n5438 115.576
R8316 Vbias.n5447 Vbias.n5443 115.576
R8317 Vbias.n5428 Vbias.n2291 115.576
R8318 Vbias.n5430 Vbias.n5428 115.576
R8319 Vbias.n5430 Vbias.n5429 115.576
R8320 Vbias.n5429 Vbias.n5421 115.576
R8321 Vbias.n5936 Vbias.n5935 115.576
R8322 Vbias.n5935 Vbias.n1626 115.576
R8323 Vbias.n5923 Vbias.n5922 115.576
R8324 Vbias.n5925 Vbias.n5923 115.576
R8325 Vbias.n5925 Vbias.n5924 115.576
R8326 Vbias.n5924 Vbias.n1629 115.576
R8327 Vbias.n6106 Vbias.n6105 115.576
R8328 Vbias.n6118 Vbias.n6106 115.576
R8329 Vbias.n6118 Vbias.n6117 115.576
R8330 Vbias.n6117 Vbias.n6114 115.576
R8331 Vbias.n1993 Vbias.n1990 115.576
R8332 Vbias.n2006 Vbias.n1990 115.576
R8333 Vbias.n2007 Vbias.n2006 115.576
R8334 Vbias.n2007 Vbias.n1987 115.576
R8335 Vbias.n1966 Vbias.n1965 115.576
R8336 Vbias.n1978 Vbias.n1966 115.576
R8337 Vbias.n1978 Vbias.n1977 115.576
R8338 Vbias.n1977 Vbias.n1974 115.576
R8339 Vbias.n1932 Vbias.n1931 115.576
R8340 Vbias.n1944 Vbias.n1932 115.576
R8341 Vbias.n1944 Vbias.n1943 115.576
R8342 Vbias.n1943 Vbias.n1940 115.576
R8343 Vbias.n1808 Vbias.n1763 115.576
R8344 Vbias.n1814 Vbias.n1763 115.576
R8345 Vbias.n1815 Vbias.n1814 115.576
R8346 Vbias.n1816 Vbias.n1815 115.576
R8347 Vbias.n1864 Vbias.n1863 115.576
R8348 Vbias.n1876 Vbias.n1864 115.576
R8349 Vbias.n1876 Vbias.n1875 115.576
R8350 Vbias.n1875 Vbias.n1874 115.576
R8351 Vbias.n1737 Vbias.n1729 115.576
R8352 Vbias.n2043 Vbias.n1729 115.576
R8353 Vbias.n2043 Vbias.n2042 115.576
R8354 Vbias.n2042 Vbias.n1730 115.576
R8355 Vbias.n1910 Vbias.n1909 115.576
R8356 Vbias.n1909 Vbias.n1908 115.576
R8357 Vbias.n1908 Vbias.n1891 115.576
R8358 Vbias.n1902 Vbias.n1891 115.576
R8359 Vbias.n1786 Vbias.n1785 115.576
R8360 Vbias.n1785 Vbias.n1784 115.576
R8361 Vbias.n1784 Vbias.n1779 115.576
R8362 Vbias.n1779 Vbias.n1552 115.576
R8363 Vbias.n1798 Vbias.n1797 115.576
R8364 Vbias.n1797 Vbias.n1796 115.576
R8365 Vbias.n1796 Vbias.n1772 115.576
R8366 Vbias.n1792 Vbias.n1772 115.576
R8367 Vbias.n6774 Vbias.n6773 115.576
R8368 Vbias.n6778 Vbias.n6774 115.576
R8369 Vbias.n6778 Vbias.n6777 115.576
R8370 Vbias.n6777 Vbias.n1343 115.576
R8371 Vbias.n6756 Vbias.n1441 115.576
R8372 Vbias.n6765 Vbias.n1441 115.576
R8373 Vbias.n6766 Vbias.n6765 115.576
R8374 Vbias.n6767 Vbias.n6766 115.576
R8375 Vbias.n6057 Vbias.n6056 115.576
R8376 Vbias.n6056 Vbias.n1414 115.576
R8377 Vbias.n6071 Vbias.n6070 115.576
R8378 Vbias.n6070 Vbias.n6069 115.576
R8379 Vbias.n6069 Vbias.n6047 115.576
R8380 Vbias.n6063 Vbias.n6047 115.576
R8381 Vbias.n1283 Vbias.n1280 115.576
R8382 Vbias.n7085 Vbias.n1280 115.576
R8383 Vbias.n7086 Vbias.n7085 115.576
R8384 Vbias.n7086 Vbias.n1277 115.576
R8385 Vbias.n1302 Vbias.n1299 115.576
R8386 Vbias.n7068 Vbias.n1299 115.576
R8387 Vbias.n7069 Vbias.n7068 115.576
R8388 Vbias.n7069 Vbias.n1295 115.576
R8389 Vbias.n7043 Vbias.n7042 115.576
R8390 Vbias.n7042 Vbias.n1318 115.576
R8391 Vbias.n7022 Vbias.n7021 115.576
R8392 Vbias.n7026 Vbias.n7022 115.576
R8393 Vbias.n7026 Vbias.n7025 115.576
R8394 Vbias.n7025 Vbias.n1325 115.576
R8395 Vbias.n1096 Vbias.n1093 115.576
R8396 Vbias.n7191 Vbias.n1093 115.576
R8397 Vbias.n7192 Vbias.n7191 115.576
R8398 Vbias.n7192 Vbias.n1090 115.576
R8399 Vbias.n1115 Vbias.n1112 115.576
R8400 Vbias.n7174 Vbias.n1112 115.576
R8401 Vbias.n7175 Vbias.n7174 115.576
R8402 Vbias.n7175 Vbias.n1108 115.576
R8403 Vbias.n7149 Vbias.n7148 115.576
R8404 Vbias.n7148 Vbias.n1130 115.576
R8405 Vbias.n7128 Vbias.n7127 115.576
R8406 Vbias.n7132 Vbias.n7128 115.576
R8407 Vbias.n7132 Vbias.n7131 115.576
R8408 Vbias.n7131 Vbias.n1137 115.576
R8409 Vbias.n1221 Vbias.n1220 115.576
R8410 Vbias.n1220 Vbias.n1078 115.576
R8411 Vbias.n7213 Vbias.n1078 115.576
R8412 Vbias.n7214 Vbias.n7213 115.576
R8413 Vbias.n1205 Vbias.n1200 115.576
R8414 Vbias.n1227 Vbias.n1200 115.576
R8415 Vbias.n1230 Vbias.n1227 115.576
R8416 Vbias.n1232 Vbias.n1230 115.576
R8417 Vbias.n1252 Vbias.n1251 115.576
R8418 Vbias.n1251 Vbias.n1186 115.576
R8419 Vbias.n1176 Vbias.n1172 115.576
R8420 Vbias.n1258 Vbias.n1172 115.576
R8421 Vbias.n1261 Vbias.n1258 115.576
R8422 Vbias.n1263 Vbias.n1261 115.576
R8423 Vbias.n6954 Vbias.n6953 115.576
R8424 Vbias.n6953 Vbias.n1159 115.576
R8425 Vbias.n7109 Vbias.n1159 115.576
R8426 Vbias.n7110 Vbias.n7109 115.576
R8427 Vbias.n6938 Vbias.n6933 115.576
R8428 Vbias.n6960 Vbias.n6933 115.576
R8429 Vbias.n6963 Vbias.n6960 115.576
R8430 Vbias.n6965 Vbias.n6963 115.576
R8431 Vbias.n6985 Vbias.n6984 115.576
R8432 Vbias.n6984 Vbias.n6919 115.576
R8433 Vbias.n6909 Vbias.n6905 115.576
R8434 Vbias.n6991 Vbias.n6905 115.576
R8435 Vbias.n6994 Vbias.n6991 115.576
R8436 Vbias.n6996 Vbias.n6994 115.576
R8437 Vbias.n6875 Vbias.n6874 115.576
R8438 Vbias.n6874 Vbias.n1353 115.576
R8439 Vbias.n6888 Vbias.n1353 115.576
R8440 Vbias.n6889 Vbias.n6888 115.576
R8441 Vbias.n6852 Vbias.n6851 115.576
R8442 Vbias.n6851 Vbias.n1366 115.576
R8443 Vbias.n6865 Vbias.n1366 115.576
R8444 Vbias.n6866 Vbias.n6865 115.576
R8445 Vbias.n6842 Vbias.n1379 115.576
R8446 Vbias.n6843 Vbias.n6842 115.576
R8447 Vbias.n1554 Vbias.n1395 115.576
R8448 Vbias.n6824 Vbias.n1395 115.576
R8449 Vbias.n6827 Vbias.n6824 115.576
R8450 Vbias.n6828 Vbias.n6827 115.576
R8451 Vbias.n6017 Vbias.n6016 115.576
R8452 Vbias.n6016 Vbias.n1564 115.576
R8453 Vbias.n6033 Vbias.n1564 115.576
R8454 Vbias.n6034 Vbias.n6033 115.576
R8455 Vbias.n5994 Vbias.n5993 115.576
R8456 Vbias.n5993 Vbias.n1577 115.576
R8457 Vbias.n6007 Vbias.n1577 115.576
R8458 Vbias.n6008 Vbias.n6007 115.576
R8459 Vbias.n5984 Vbias.n1590 115.576
R8460 Vbias.n5985 Vbias.n5984 115.576
R8461 Vbias.n1635 Vbias.n1606 115.576
R8462 Vbias.n5966 Vbias.n1606 115.576
R8463 Vbias.n5969 Vbias.n5966 115.576
R8464 Vbias.n5970 Vbias.n5969 115.576
R8465 Vbias.n5362 Vbias.n5361 115.576
R8466 Vbias.n5361 Vbias.n5360 115.576
R8467 Vbias.n5360 Vbias.n5320 115.576
R8468 Vbias.n5351 Vbias.n5320 115.576
R8469 Vbias.n5309 Vbias.n5304 115.576
R8470 Vbias.n5368 Vbias.n5304 115.576
R8471 Vbias.n5371 Vbias.n5368 115.576
R8472 Vbias.n5373 Vbias.n5371 115.576
R8473 Vbias.n5393 Vbias.n5392 115.576
R8474 Vbias.n5392 Vbias.n5290 115.576
R8475 Vbias.n5280 Vbias.n5275 115.576
R8476 Vbias.n5399 Vbias.n5275 115.576
R8477 Vbias.n5402 Vbias.n5399 115.576
R8478 Vbias.n5404 Vbias.n5402 115.576
R8479 Vbias.n5244 Vbias.n5243 115.576
R8480 Vbias.n5243 Vbias.n2301 115.576
R8481 Vbias.n5257 Vbias.n2301 115.576
R8482 Vbias.n5258 Vbias.n5257 115.576
R8483 Vbias.n5221 Vbias.n5220 115.576
R8484 Vbias.n5220 Vbias.n2314 115.576
R8485 Vbias.n5234 Vbias.n2314 115.576
R8486 Vbias.n5235 Vbias.n5234 115.576
R8487 Vbias.n5211 Vbias.n2327 115.576
R8488 Vbias.n5212 Vbias.n5211 115.576
R8489 Vbias.n2367 Vbias.n2343 115.576
R8490 Vbias.n5193 Vbias.n2343 115.576
R8491 Vbias.n5196 Vbias.n5193 115.576
R8492 Vbias.n5197 Vbias.n5196 115.576
R8493 Vbias.n2530 Vbias.n2529 115.576
R8494 Vbias.n2529 Vbias.n2528 115.576
R8495 Vbias.n2528 Vbias.n2488 115.576
R8496 Vbias.n2519 Vbias.n2488 115.576
R8497 Vbias.n2477 Vbias.n2472 115.576
R8498 Vbias.n2536 Vbias.n2472 115.576
R8499 Vbias.n2539 Vbias.n2536 115.576
R8500 Vbias.n2541 Vbias.n2539 115.576
R8501 Vbias.n2561 Vbias.n2560 115.576
R8502 Vbias.n2560 Vbias.n2458 115.576
R8503 Vbias.n2448 Vbias.n2443 115.576
R8504 Vbias.n2567 Vbias.n2443 115.576
R8505 Vbias.n2570 Vbias.n2567 115.576
R8506 Vbias.n2572 Vbias.n2570 115.576
R8507 Vbias.n5043 Vbias.n5042 115.576
R8508 Vbias.n5047 Vbias.n5043 115.576
R8509 Vbias.n5047 Vbias.n5046 115.576
R8510 Vbias.n5046 Vbias.n2419 115.576
R8511 Vbias.n4547 Vbias.n4546 115.576
R8512 Vbias.n4546 Vbias.n4545 115.576
R8513 Vbias.n4545 Vbias.n4411 115.576
R8514 Vbias.n4536 Vbias.n4411 115.576
R8515 Vbias.n3828 Vbias.n3827 115.576
R8516 Vbias.n3829 Vbias.n3828 115.576
R8517 Vbias.n3835 Vbias.n3829 115.576
R8518 Vbias.n3836 Vbias.n3835 115.576
R8519 Vbias.n3812 Vbias.n3793 115.576
R8520 Vbias.n3845 Vbias.n3812 115.576
R8521 Vbias.n3845 Vbias.n3844 115.576
R8522 Vbias.n3844 Vbias.n3843 115.576
R8523 Vbias.n3872 Vbias.n3871 115.576
R8524 Vbias.n3873 Vbias.n3872 115.576
R8525 Vbias.n3864 Vbias.n3783 115.576
R8526 Vbias.n3879 Vbias.n3783 115.576
R8527 Vbias.n3904 Vbias.n3903 115.576
R8528 Vbias.n3905 Vbias.n3904 115.576
R8529 Vbias.n3911 Vbias.n3905 115.576
R8530 Vbias.n3912 Vbias.n3911 115.576
R8531 Vbias.n3765 Vbias.n3746 115.576
R8532 Vbias.n3921 Vbias.n3765 115.576
R8533 Vbias.n3921 Vbias.n3920 115.576
R8534 Vbias.n3920 Vbias.n3919 115.576
R8535 Vbias.n3942 Vbias.n3941 115.576
R8536 Vbias.n3943 Vbias.n3942 115.576
R8537 Vbias.n3949 Vbias.n3943 115.576
R8538 Vbias.n3950 Vbias.n3949 115.576
R8539 Vbias.n3736 Vbias.n3717 115.576
R8540 Vbias.n3959 Vbias.n3736 115.576
R8541 Vbias.n3959 Vbias.n3958 115.576
R8542 Vbias.n3958 Vbias.n3957 115.576
R8543 Vbias.n3290 Vbias.n3289 115.576
R8544 Vbias.n3291 Vbias.n3290 115.576
R8545 Vbias.n3297 Vbias.n3291 115.576
R8546 Vbias.n3298 Vbias.n3297 115.576
R8547 Vbias.n3274 Vbias.n3255 115.576
R8548 Vbias.n3307 Vbias.n3274 115.576
R8549 Vbias.n3307 Vbias.n3306 115.576
R8550 Vbias.n3306 Vbias.n3305 115.576
R8551 Vbias.n3334 Vbias.n3333 115.576
R8552 Vbias.n3335 Vbias.n3334 115.576
R8553 Vbias.n3326 Vbias.n3245 115.576
R8554 Vbias.n3341 Vbias.n3245 115.576
R8555 Vbias.n3366 Vbias.n3365 115.576
R8556 Vbias.n3367 Vbias.n3366 115.576
R8557 Vbias.n3373 Vbias.n3367 115.576
R8558 Vbias.n3374 Vbias.n3373 115.576
R8559 Vbias.n3227 Vbias.n3208 115.576
R8560 Vbias.n3383 Vbias.n3227 115.576
R8561 Vbias.n3383 Vbias.n3382 115.576
R8562 Vbias.n3382 Vbias.n3381 115.576
R8563 Vbias.n3404 Vbias.n3403 115.576
R8564 Vbias.n3405 Vbias.n3404 115.576
R8565 Vbias.n3411 Vbias.n3405 115.576
R8566 Vbias.n3412 Vbias.n3411 115.576
R8567 Vbias.n3198 Vbias.n3179 115.576
R8568 Vbias.n3421 Vbias.n3198 115.576
R8569 Vbias.n3421 Vbias.n3420 115.576
R8570 Vbias.n3420 Vbias.n3419 115.576
R8571 Vbias.n3559 Vbias.n3558 115.576
R8572 Vbias.n3560 Vbias.n3559 115.576
R8573 Vbias.n3566 Vbias.n3560 115.576
R8574 Vbias.n3567 Vbias.n3566 115.576
R8575 Vbias.n3543 Vbias.n3524 115.576
R8576 Vbias.n3576 Vbias.n3543 115.576
R8577 Vbias.n3576 Vbias.n3575 115.576
R8578 Vbias.n3575 Vbias.n3574 115.576
R8579 Vbias.n3603 Vbias.n3602 115.576
R8580 Vbias.n3604 Vbias.n3603 115.576
R8581 Vbias.n3595 Vbias.n3514 115.576
R8582 Vbias.n3610 Vbias.n3514 115.576
R8583 Vbias.n3635 Vbias.n3634 115.576
R8584 Vbias.n3636 Vbias.n3635 115.576
R8585 Vbias.n3642 Vbias.n3636 115.576
R8586 Vbias.n3643 Vbias.n3642 115.576
R8587 Vbias.n3496 Vbias.n3477 115.576
R8588 Vbias.n3652 Vbias.n3496 115.576
R8589 Vbias.n3652 Vbias.n3651 115.576
R8590 Vbias.n3651 Vbias.n3650 115.576
R8591 Vbias.n3673 Vbias.n3672 115.576
R8592 Vbias.n3674 Vbias.n3673 115.576
R8593 Vbias.n3680 Vbias.n3674 115.576
R8594 Vbias.n3681 Vbias.n3680 115.576
R8595 Vbias.n3467 Vbias.n3448 115.576
R8596 Vbias.n3690 Vbias.n3467 115.576
R8597 Vbias.n3690 Vbias.n3689 115.576
R8598 Vbias.n3689 Vbias.n3688 115.576
R8599 Vbias.n4066 Vbias.n4051 115.576
R8600 Vbias.n4191 Vbias.n4066 115.576
R8601 Vbias.n4191 Vbias.n4190 115.576
R8602 Vbias.n4190 Vbias.n4189 115.576
R8603 Vbias.n4152 Vbias.n4041 115.576
R8604 Vbias.n4205 Vbias.n4041 115.576
R8605 Vbias.n4024 Vbias.n4009 115.576
R8606 Vbias.n4225 Vbias.n4024 115.576
R8607 Vbias.n4225 Vbias.n4224 115.576
R8608 Vbias.n4224 Vbias.n4223 115.576
R8609 Vbias.n4246 Vbias.n4245 115.576
R8610 Vbias.n4245 Vbias.n4244 115.576
R8611 Vbias.n4244 Vbias.n3992 115.576
R8612 Vbias.n4236 Vbias.n3992 115.576
R8613 Vbias.n4171 Vbias.n4170 115.576
R8614 Vbias.n4170 Vbias.n4169 115.576
R8615 Vbias.n4169 Vbias.n4074 115.576
R8616 Vbias.n4184 Vbias.n4074 115.576
R8617 Vbias.n4160 Vbias.n4159 115.576
R8618 Vbias.n4161 Vbias.n4160 115.576
R8619 Vbias.n4135 Vbias.n4134 115.576
R8620 Vbias.n4136 Vbias.n4135 115.576
R8621 Vbias.n4137 Vbias.n4136 115.576
R8622 Vbias.n4138 Vbias.n4137 115.576
R8623 Vbias.n4119 Vbias.n4118 115.576
R8624 Vbias.n4120 Vbias.n4119 115.576
R8625 Vbias.n4121 Vbias.n4120 115.576
R8626 Vbias.n4122 Vbias.n4121 115.576
R8627 Vbias.n2624 Vbias.n2612 115.576
R8628 Vbias.n4978 Vbias.n2612 115.576
R8629 Vbias.n4981 Vbias.n4978 115.576
R8630 Vbias.n4982 Vbias.n4981 115.576
R8631 Vbias.n4963 Vbias.n4960 115.576
R8632 Vbias.n4964 Vbias.n4963 115.576
R8633 Vbias.n4938 Vbias.n4937 115.576
R8634 Vbias.n4937 Vbias.n2635 115.576
R8635 Vbias.n4951 Vbias.n2635 115.576
R8636 Vbias.n4952 Vbias.n4951 115.576
R8637 Vbias.n4916 Vbias.n4915 115.576
R8638 Vbias.n4915 Vbias.n2649 115.576
R8639 Vbias.n4928 Vbias.n2649 115.576
R8640 Vbias.n4929 Vbias.n4928 115.576
R8641 Vbias.n3020 Vbias.n3019 115.576
R8642 Vbias.n3021 Vbias.n3020 115.576
R8643 Vbias.n3027 Vbias.n3021 115.576
R8644 Vbias.n3028 Vbias.n3027 115.576
R8645 Vbias.n3004 Vbias.n2985 115.576
R8646 Vbias.n3037 Vbias.n3004 115.576
R8647 Vbias.n3037 Vbias.n3036 115.576
R8648 Vbias.n3036 Vbias.n3035 115.576
R8649 Vbias.n3064 Vbias.n3063 115.576
R8650 Vbias.n3065 Vbias.n3064 115.576
R8651 Vbias.n3056 Vbias.n2975 115.576
R8652 Vbias.n3071 Vbias.n2975 115.576
R8653 Vbias.n3096 Vbias.n3095 115.576
R8654 Vbias.n3097 Vbias.n3096 115.576
R8655 Vbias.n3103 Vbias.n3097 115.576
R8656 Vbias.n3104 Vbias.n3103 115.576
R8657 Vbias.n2957 Vbias.n2938 115.576
R8658 Vbias.n3113 Vbias.n2957 115.576
R8659 Vbias.n3113 Vbias.n3112 115.576
R8660 Vbias.n3112 Vbias.n3111 115.576
R8661 Vbias.n3134 Vbias.n3133 115.576
R8662 Vbias.n3135 Vbias.n3134 115.576
R8663 Vbias.n3141 Vbias.n3135 115.576
R8664 Vbias.n3142 Vbias.n3141 115.576
R8665 Vbias.n2928 Vbias.n2909 115.576
R8666 Vbias.n3151 Vbias.n2928 115.576
R8667 Vbias.n3151 Vbias.n3150 115.576
R8668 Vbias.n3150 Vbias.n3149 115.576
R8669 Vbias.n4696 Vbias.n4695 115.576
R8670 Vbias.n4697 Vbias.n4696 115.576
R8671 Vbias.n4703 Vbias.n4697 115.576
R8672 Vbias.n4704 Vbias.n4703 115.576
R8673 Vbias.n2765 Vbias.n2746 115.576
R8674 Vbias.n4713 Vbias.n2765 115.576
R8675 Vbias.n4713 Vbias.n4712 115.576
R8676 Vbias.n4712 Vbias.n4711 115.576
R8677 Vbias.n4740 Vbias.n4739 115.576
R8678 Vbias.n4741 Vbias.n4740 115.576
R8679 Vbias.n4732 Vbias.n2736 115.576
R8680 Vbias.n4747 Vbias.n2736 115.576
R8681 Vbias.n4772 Vbias.n4771 115.576
R8682 Vbias.n4773 Vbias.n4772 115.576
R8683 Vbias.n4779 Vbias.n4773 115.576
R8684 Vbias.n4780 Vbias.n4779 115.576
R8685 Vbias.n2718 Vbias.n2699 115.576
R8686 Vbias.n4789 Vbias.n2718 115.576
R8687 Vbias.n4789 Vbias.n4788 115.576
R8688 Vbias.n4788 Vbias.n4787 115.576
R8689 Vbias.n4810 Vbias.n4809 115.576
R8690 Vbias.n4811 Vbias.n4810 115.576
R8691 Vbias.n4817 Vbias.n4811 115.576
R8692 Vbias.n4818 Vbias.n4817 115.576
R8693 Vbias.n2689 Vbias.n2670 115.576
R8694 Vbias.n4827 Vbias.n2689 115.576
R8695 Vbias.n4827 Vbias.n4826 115.576
R8696 Vbias.n4826 Vbias.n4825 115.576
R8697 Vbias.n4566 Vbias.n4553 115.576
R8698 Vbias.n4568 Vbias.n4566 115.576
R8699 Vbias.n4568 Vbias.n4567 115.576
R8700 Vbias.n4567 Vbias.n4559 115.576
R8701 Vbias.n2218 Vbias.n2204 115.576
R8702 Vbias.n5657 Vbias.n2204 115.576
R8703 Vbias.n5658 Vbias.n5657 115.576
R8704 Vbias.n5659 Vbias.n5658 115.576
R8705 Vbias.n5644 Vbias.n5643 115.576
R8706 Vbias.n5645 Vbias.n5644 115.576
R8707 Vbias.n5621 Vbias.n5558 115.576
R8708 Vbias.n5633 Vbias.n5558 115.576
R8709 Vbias.n5634 Vbias.n5633 115.576
R8710 Vbias.n5635 Vbias.n5634 115.576
R8711 Vbias.n5603 Vbias.n5576 115.576
R8712 Vbias.n5614 Vbias.n5576 115.576
R8713 Vbias.n5615 Vbias.n5614 115.576
R8714 Vbias.n5616 Vbias.n5615 115.576
R8715 Vbias.n2147 Vbias.n2133 115.576
R8716 Vbias.n5731 Vbias.n2133 115.576
R8717 Vbias.n5732 Vbias.n5731 115.576
R8718 Vbias.n5733 Vbias.n5732 115.576
R8719 Vbias.n5718 Vbias.n5717 115.576
R8720 Vbias.n5719 Vbias.n5718 115.576
R8721 Vbias.n5695 Vbias.n2161 115.576
R8722 Vbias.n5707 Vbias.n2161 115.576
R8723 Vbias.n5708 Vbias.n5707 115.576
R8724 Vbias.n5709 Vbias.n5708 115.576
R8725 Vbias.n5677 Vbias.n2179 115.576
R8726 Vbias.n5688 Vbias.n2179 115.576
R8727 Vbias.n5689 Vbias.n5688 115.576
R8728 Vbias.n5690 Vbias.n5689 115.576
R8729 Vbias.n5792 Vbias.n2078 115.576
R8730 Vbias.n5820 Vbias.n2078 115.576
R8731 Vbias.n5821 Vbias.n5820 115.576
R8732 Vbias.n5822 Vbias.n5821 115.576
R8733 Vbias.n5807 Vbias.n5806 115.576
R8734 Vbias.n5808 Vbias.n5807 115.576
R8735 Vbias.n2108 Vbias.n2092 115.576
R8736 Vbias.n5777 Vbias.n2092 115.576
R8737 Vbias.n5778 Vbias.n5777 115.576
R8738 Vbias.n5779 Vbias.n5778 115.576
R8739 Vbias.n5747 Vbias.n2116 115.576
R8740 Vbias.n5763 Vbias.n2116 115.576
R8741 Vbias.n5764 Vbias.n5763 115.576
R8742 Vbias.n5765 Vbias.n5764 115.576
R8743 Vbias.n1496 Vbias.n1495 115.576
R8744 Vbias.n6658 Vbias.n1496 115.576
R8745 Vbias.n6658 Vbias.n6657 115.576
R8746 Vbias.n6657 Vbias.n6656 115.576
R8747 Vbias.n6672 Vbias.n6671 115.576
R8748 Vbias.n6671 Vbias.n6670 115.576
R8749 Vbias.n5848 Vbias.n5847 115.576
R8750 Vbias.n5849 Vbias.n5848 115.576
R8751 Vbias.n5850 Vbias.n5849 115.576
R8752 Vbias.n5851 Vbias.n5850 115.576
R8753 Vbias.n6354 Vbias.n6231 115.576
R8754 Vbias.n6584 Vbias.n6231 115.576
R8755 Vbias.n6585 Vbias.n6584 115.576
R8756 Vbias.n6586 Vbias.n6585 115.576
R8757 Vbias.n6348 Vbias.n6347 115.576
R8758 Vbias.n6349 Vbias.n6348 115.576
R8759 Vbias.n6281 Vbias.n6267 115.576
R8760 Vbias.n6334 Vbias.n6267 115.576
R8761 Vbias.n6335 Vbias.n6334 115.576
R8762 Vbias.n6336 Vbias.n6335 115.576
R8763 Vbias.n6304 Vbias.n6289 115.576
R8764 Vbias.n6320 Vbias.n6289 115.576
R8765 Vbias.n6321 Vbias.n6320 115.576
R8766 Vbias.n6322 Vbias.n6321 115.576
R8767 Vbias.n852 Vbias.n851 115.576
R8768 Vbias.n7597 Vbias.n852 115.576
R8769 Vbias.n7597 Vbias.n7596 115.576
R8770 Vbias.n7596 Vbias.n7595 115.576
R8771 Vbias.n7611 Vbias.n7610 115.576
R8772 Vbias.n7610 Vbias.n7609 115.576
R8773 Vbias.n7626 Vbias.n7625 115.576
R8774 Vbias.n7625 Vbias.n7624 115.576
R8775 Vbias.n7624 Vbias.n804 115.576
R8776 Vbias.n7616 Vbias.n804 115.576
R8777 Vbias.n7641 Vbias.n7640 115.576
R8778 Vbias.n7640 Vbias.n7639 115.576
R8779 Vbias.n7639 Vbias.n785 115.576
R8780 Vbias.n7631 Vbias.n785 115.576
R8781 Vbias.n1007 Vbias.n1006 115.576
R8782 Vbias.n7475 Vbias.n1007 115.576
R8783 Vbias.n7475 Vbias.n7474 115.576
R8784 Vbias.n7474 Vbias.n7473 115.576
R8785 Vbias.n7489 Vbias.n7488 115.576
R8786 Vbias.n7488 Vbias.n7487 115.576
R8787 Vbias.n7505 Vbias.n7504 115.576
R8788 Vbias.n7504 Vbias.n7503 115.576
R8789 Vbias.n7503 Vbias.n959 115.576
R8790 Vbias.n7495 Vbias.n959 115.576
R8791 Vbias.n7520 Vbias.n7519 115.576
R8792 Vbias.n7519 Vbias.n7518 115.576
R8793 Vbias.n7518 Vbias.n936 115.576
R8794 Vbias.n7510 Vbias.n936 115.576
R8795 Vbias.n6218 Vbias.n6204 115.576
R8796 Vbias.n6220 Vbias.n6218 115.576
R8797 Vbias.n6220 Vbias.n6219 115.576
R8798 Vbias.n6219 Vbias.n6211 115.576
R8799 Vbias.n6198 Vbias.n6190 115.576
R8800 Vbias.n6198 Vbias.n6194 115.576
R8801 Vbias.n6171 Vbias.n6167 115.576
R8802 Vbias.n6180 Vbias.n6167 115.576
R8803 Vbias.n6181 Vbias.n6180 115.576
R8804 Vbias.n6182 Vbias.n6181 115.576
R8805 Vbias.n6455 Vbias.n6441 115.576
R8806 Vbias.n6457 Vbias.n6455 115.576
R8807 Vbias.n6457 Vbias.n6456 115.576
R8808 Vbias.n6456 Vbias.n6448 115.576
R8809 Vbias.n6435 Vbias.n6427 115.576
R8810 Vbias.n6435 Vbias.n6431 115.576
R8811 Vbias.n6408 Vbias.n6385 115.576
R8812 Vbias.n6417 Vbias.n6385 115.576
R8813 Vbias.n6418 Vbias.n6417 115.576
R8814 Vbias.n6419 Vbias.n6418 115.576
R8815 Vbias.n6391 Vbias.n6388 115.576
R8816 Vbias.n6400 Vbias.n6388 115.576
R8817 Vbias.n6401 Vbias.n6400 115.576
R8818 Vbias.n6402 Vbias.n6401 115.576
R8819 Vbias.n909 Vbias.n895 115.576
R8820 Vbias.n911 Vbias.n909 115.576
R8821 Vbias.n911 Vbias.n910 115.576
R8822 Vbias.n910 Vbias.n902 115.576
R8823 Vbias.n889 Vbias.n881 115.576
R8824 Vbias.n889 Vbias.n885 115.576
R8825 Vbias.n6487 Vbias.n6486 115.576
R8826 Vbias.n6486 Vbias.n6485 115.576
R8827 Vbias.n6485 Vbias.n6470 115.576
R8828 Vbias.n6479 Vbias.n6470 115.576
R8829 Vbias.n6501 Vbias.n6500 115.576
R8830 Vbias.n6500 Vbias.n6499 115.576
R8831 Vbias.n6499 Vbias.n6464 115.576
R8832 Vbias.n6493 Vbias.n6464 115.576
R8833 Vbias.n7395 Vbias.n7382 115.576
R8834 Vbias.n7406 Vbias.n7395 115.576
R8835 Vbias.n7406 Vbias.n7405 115.576
R8836 Vbias.n7405 Vbias.n7404 115.576
R8837 Vbias.n7378 Vbias.n7371 115.576
R8838 Vbias.n7420 Vbias.n7371 115.576
R8839 Vbias.n7357 Vbias.n7344 115.576
R8840 Vbias.n7440 Vbias.n7357 115.576
R8841 Vbias.n7440 Vbias.n7439 115.576
R8842 Vbias.n7439 Vbias.n7438 115.576
R8843 Vbias.n7461 Vbias.n7460 115.576
R8844 Vbias.n7460 Vbias.n7459 115.576
R8845 Vbias.n7459 Vbias.n7333 115.576
R8846 Vbias.n7451 Vbias.n7333 115.576
R8847 Vbias.n6142 Vbias.n6138 115.576
R8848 Vbias.n6641 Vbias.n6138 115.576
R8849 Vbias.n6641 Vbias.n6640 115.576
R8850 Vbias.n6640 Vbias.n6639 115.576
R8851 Vbias.n7257 Vbias.n7256 115.576
R8852 Vbias.n7269 Vbias.n7257 115.576
R8853 Vbias.n7269 Vbias.n7268 115.576
R8854 Vbias.n7268 Vbias.n7267 115.576
R8855 Vbias.n7283 Vbias.n7282 115.576
R8856 Vbias.n7282 Vbias.n7281 115.576
R8857 Vbias.n7298 Vbias.n7297 115.576
R8858 Vbias.n7297 Vbias.n7296 115.576
R8859 Vbias.n7296 Vbias.n1054 115.576
R8860 Vbias.n7288 Vbias.n1054 115.576
R8861 Vbias.n7313 Vbias.n7312 115.576
R8862 Vbias.n7312 Vbias.n7311 115.576
R8863 Vbias.n7311 Vbias.n1033 115.576
R8864 Vbias.n7303 Vbias.n1033 115.576
R8865 Vbias.n693 Vbias.n681 115.576
R8866 Vbias.n7727 Vbias.n693 115.576
R8867 Vbias.n7727 Vbias.n7726 115.576
R8868 Vbias.n7726 Vbias.n7725 115.576
R8869 Vbias.n2056 Vbias.n2055 115.576
R8870 Vbias.n2055 Vbias.n2054 115.576
R8871 Vbias.n2054 Vbias.n1708 115.576
R8872 Vbias.n2045 Vbias.n1708 115.576
R8873 Vbias.n6683 Vbias.n6682 115.576
R8874 Vbias.n6683 Vbias.n1452 115.576
R8875 Vbias.n1691 Vbias.n1684 115.576
R8876 Vbias.n5863 Vbias.n1684 115.576
R8877 Vbias.n5522 Vbias.n5511 115.576
R8878 Vbias.n5523 Vbias.n5522 115.576
R8879 Vbias.n2244 Vbias.n2237 115.576
R8880 Vbias.n5539 Vbias.n2237 115.576
R8881 Vbias.n5014 Vbias.n2589 115.576
R8882 Vbias.n5020 Vbias.n2589 115.576
R8883 Vbias.n24 Vbias.n12 115.576
R8884 Vbias.n8067 Vbias.n24 115.576
R8885 Vbias.n8067 Vbias.n8066 115.576
R8886 Vbias.n8066 Vbias.n8065 115.576
R8887 Vbias.n6754 Vbias.n6751 112.255
R8888 Vbias.n5878 Vbias.n1672 112.255
R8889 Vbias.n5080 Vbias.n2228 112.255
R8890 Vbias.n6101 Vbias.n1523 106.32
R8891 Vbias.n6676 Vbias.n1460 106.32
R8892 Vbias.n6101 Vbias.n1525 106.32
R8893 Vbias.n6676 Vbias.n1463 106.32
R8894 Vbias.n6101 Vbias.n1526 106.32
R8895 Vbias.n6676 Vbias.n1464 106.32
R8896 Vbias.n6102 Vbias.n6101 106.162
R8897 Vbias.n6676 Vbias.n1462 106.162
R8898 Vbias.t793 Vbias.t815 104.74
R8899 Vbias.n1806 Vbias.n1804 104.74
R8900 Vbias.n5858 Vbias.n1693 99.4607
R8901 Vbias.n4865 Vbias.n4864 99.0123
R8902 Vbias.n4866 Vbias.n4865 99.0123
R8903 Vbias.n4876 Vbias.n4875 99.0123
R8904 Vbias.n4875 Vbias.n4874 99.0123
R8905 Vbias.n4881 Vbias.n4850 99.0123
R8906 Vbias.n4882 Vbias.n4881 99.0123
R8907 Vbias.n6101 Vbias.n6100 88.201
R8908 Vbias.n4911 Vbias.n4910 86.184
R8909 Vbias.n4933 Vbias.n4932 86.184
R8910 Vbias.n2628 Vbias.n2627 86.184
R8911 Vbias.n606 Vbias.n605 83.5719
R8912 Vbias.t681 Vbias.n606 83.5719
R8913 Vbias.n615 Vbias.n614 83.5719
R8914 Vbias.n615 Vbias.t614 83.5719
R8915 Vbias.n598 Vbias.n596 83.5719
R8916 Vbias.n596 Vbias.t275 83.5719
R8917 Vbias.n7781 Vbias.n604 83.5719
R8918 Vbias.t681 Vbias.n604 83.5719
R8919 Vbias.n7783 Vbias.n602 83.5719
R8920 Vbias.t614 Vbias.n602 83.5719
R8921 Vbias.n7786 Vbias.n597 83.5719
R8922 Vbias.n597 Vbias.t275 83.5719
R8923 Vbias.n622 Vbias.n620 83.5719
R8924 Vbias.n620 Vbias.t817 83.5719
R8925 Vbias.n7774 Vbias.n621 83.5719
R8926 Vbias.n621 Vbias.t817 83.5719
R8927 Vbias.n631 Vbias.n630 83.5719
R8928 Vbias.t848 Vbias.n631 83.5719
R8929 Vbias.n638 Vbias.n637 83.5719
R8930 Vbias.n638 Vbias.t855 83.5719
R8931 Vbias.n7768 Vbias.n629 83.5719
R8932 Vbias.t848 Vbias.n629 83.5719
R8933 Vbias.n7770 Vbias.n627 83.5719
R8934 Vbias.t855 Vbias.n627 83.5719
R8935 Vbias.n653 Vbias.n652 83.5719
R8936 Vbias.t786 Vbias.n653 83.5719
R8937 Vbias.n662 Vbias.n661 83.5719
R8938 Vbias.n662 Vbias.t721 83.5719
R8939 Vbias.n645 Vbias.n643 83.5719
R8940 Vbias.n643 Vbias.t273 83.5719
R8941 Vbias.n7756 Vbias.n651 83.5719
R8942 Vbias.t786 Vbias.n651 83.5719
R8943 Vbias.n7758 Vbias.n649 83.5719
R8944 Vbias.t721 Vbias.n649 83.5719
R8945 Vbias.n7761 Vbias.n644 83.5719
R8946 Vbias.n644 Vbias.t273 83.5719
R8947 Vbias.n7793 Vbias.n580 83.5719
R8948 Vbias.t441 Vbias.n580 83.5719
R8949 Vbias.n7795 Vbias.n578 83.5719
R8950 Vbias.t600 Vbias.n578 83.5719
R8951 Vbias.n582 Vbias.n581 83.5719
R8952 Vbias.t441 Vbias.n582 83.5719
R8953 Vbias.n591 Vbias.n590 83.5719
R8954 Vbias.n591 Vbias.t600 83.5719
R8955 Vbias.n574 Vbias.n572 83.5719
R8956 Vbias.n572 Vbias.t50 83.5719
R8957 Vbias.n7798 Vbias.n573 83.5719
R8958 Vbias.n573 Vbias.t50 83.5719
R8959 Vbias.n492 Vbias.n491 83.5719
R8960 Vbias.t153 Vbias.n492 83.5719
R8961 Vbias.n501 Vbias.n500 83.5719
R8962 Vbias.n501 Vbias.t547 83.5719
R8963 Vbias.n484 Vbias.n482 83.5719
R8964 Vbias.n482 Vbias.t218 83.5719
R8965 Vbias.n7850 Vbias.n490 83.5719
R8966 Vbias.t153 Vbias.n490 83.5719
R8967 Vbias.n7852 Vbias.n488 83.5719
R8968 Vbias.t547 Vbias.n488 83.5719
R8969 Vbias.n7855 Vbias.n483 83.5719
R8970 Vbias.n483 Vbias.t218 83.5719
R8971 Vbias.n508 Vbias.n506 83.5719
R8972 Vbias.n506 Vbias.t397 83.5719
R8973 Vbias.n7843 Vbias.n507 83.5719
R8974 Vbias.n507 Vbias.t397 83.5719
R8975 Vbias.n517 Vbias.n516 83.5719
R8976 Vbias.t741 Vbias.n517 83.5719
R8977 Vbias.n524 Vbias.n523 83.5719
R8978 Vbias.n524 Vbias.t889 83.5719
R8979 Vbias.n7837 Vbias.n515 83.5719
R8980 Vbias.t741 Vbias.n515 83.5719
R8981 Vbias.n7839 Vbias.n513 83.5719
R8982 Vbias.t889 Vbias.n513 83.5719
R8983 Vbias.n539 Vbias.n538 83.5719
R8984 Vbias.t823 Vbias.n539 83.5719
R8985 Vbias.n548 Vbias.n547 83.5719
R8986 Vbias.n548 Vbias.t505 83.5719
R8987 Vbias.n531 Vbias.n529 83.5719
R8988 Vbias.n529 Vbias.t184 83.5719
R8989 Vbias.n7825 Vbias.n537 83.5719
R8990 Vbias.t823 Vbias.n537 83.5719
R8991 Vbias.n7827 Vbias.n535 83.5719
R8992 Vbias.t505 Vbias.n535 83.5719
R8993 Vbias.n7830 Vbias.n530 83.5719
R8994 Vbias.n530 Vbias.t184 83.5719
R8995 Vbias.n7862 Vbias.n466 83.5719
R8996 Vbias.t327 Vbias.n466 83.5719
R8997 Vbias.n7864 Vbias.n464 83.5719
R8998 Vbias.t161 Vbias.n464 83.5719
R8999 Vbias.n468 Vbias.n467 83.5719
R9000 Vbias.t327 Vbias.n468 83.5719
R9001 Vbias.n477 Vbias.n476 83.5719
R9002 Vbias.n477 Vbias.t161 83.5719
R9003 Vbias.n460 Vbias.n458 83.5719
R9004 Vbias.n458 Vbias.t112 83.5719
R9005 Vbias.n7867 Vbias.n459 83.5719
R9006 Vbias.n459 Vbias.t112 83.5719
R9007 Vbias.n386 Vbias.n385 83.5719
R9008 Vbias.t430 Vbias.n386 83.5719
R9009 Vbias.n395 Vbias.n394 83.5719
R9010 Vbias.n395 Vbias.t797 83.5719
R9011 Vbias.n378 Vbias.n376 83.5719
R9012 Vbias.n376 Vbias.t172 83.5719
R9013 Vbias.n7916 Vbias.n384 83.5719
R9014 Vbias.t430 Vbias.n384 83.5719
R9015 Vbias.n7918 Vbias.n382 83.5719
R9016 Vbias.t797 Vbias.n382 83.5719
R9017 Vbias.n7921 Vbias.n377 83.5719
R9018 Vbias.n377 Vbias.t172 83.5719
R9019 Vbias.n402 Vbias.n400 83.5719
R9020 Vbias.n400 Vbias.t590 83.5719
R9021 Vbias.n7909 Vbias.n401 83.5719
R9022 Vbias.n401 Vbias.t590 83.5719
R9023 Vbias.n411 Vbias.n410 83.5719
R9024 Vbias.t633 Vbias.n411 83.5719
R9025 Vbias.n418 Vbias.n417 83.5719
R9026 Vbias.n418 Vbias.t320 83.5719
R9027 Vbias.n7903 Vbias.n409 83.5719
R9028 Vbias.t633 Vbias.n409 83.5719
R9029 Vbias.n7905 Vbias.n407 83.5719
R9030 Vbias.t320 Vbias.n407 83.5719
R9031 Vbias.n433 Vbias.n432 83.5719
R9032 Vbias.t774 Vbias.n433 83.5719
R9033 Vbias.n442 Vbias.n441 83.5719
R9034 Vbias.n442 Vbias.t886 83.5719
R9035 Vbias.n425 Vbias.n423 83.5719
R9036 Vbias.n423 Vbias.t190 83.5719
R9037 Vbias.n7891 Vbias.n431 83.5719
R9038 Vbias.t774 Vbias.n431 83.5719
R9039 Vbias.n7893 Vbias.n429 83.5719
R9040 Vbias.t886 Vbias.n429 83.5719
R9041 Vbias.n7896 Vbias.n424 83.5719
R9042 Vbias.n424 Vbias.t190 83.5719
R9043 Vbias.n7928 Vbias.n360 83.5719
R9044 Vbias.t443 Vbias.n360 83.5719
R9045 Vbias.n7930 Vbias.n358 83.5719
R9046 Vbias.t673 Vbias.n358 83.5719
R9047 Vbias.n362 Vbias.n361 83.5719
R9048 Vbias.t443 Vbias.n362 83.5719
R9049 Vbias.n371 Vbias.n370 83.5719
R9050 Vbias.n371 Vbias.t673 83.5719
R9051 Vbias.n177 Vbias.n175 83.5719
R9052 Vbias.n175 Vbias.t86 83.5719
R9053 Vbias.n7933 Vbias.n176 83.5719
R9054 Vbias.n176 Vbias.t86 83.5719
R9055 Vbias.n216 Vbias.n215 83.5719
R9056 Vbias.t455 Vbias.n216 83.5719
R9057 Vbias.n280 Vbias.n279 83.5719
R9058 Vbias.n279 Vbias.t309 83.5719
R9059 Vbias.n277 Vbias.n222 83.5719
R9060 Vbias.n277 Vbias.t206 83.5719
R9061 Vbias.n290 Vbias.n214 83.5719
R9062 Vbias.t455 Vbias.n214 83.5719
R9063 Vbias.n229 Vbias.n228 83.5719
R9064 Vbias.n228 Vbias.t309 83.5719
R9065 Vbias.n276 Vbias.n275 83.5719
R9066 Vbias.t206 Vbias.n276 83.5719
R9067 Vbias.n210 Vbias.n208 83.5719
R9068 Vbias.n208 Vbias.t863 83.5719
R9069 Vbias.n295 Vbias.n209 83.5719
R9070 Vbias.n209 Vbias.t863 83.5719
R9071 Vbias.n202 Vbias.n201 83.5719
R9072 Vbias.t859 Vbias.n202 83.5719
R9073 Vbias.n302 Vbias.n301 83.5719
R9074 Vbias.n301 Vbias.t802 83.5719
R9075 Vbias.n310 Vbias.n200 83.5719
R9076 Vbias.t859 Vbias.n200 83.5719
R9077 Vbias.n207 Vbias.n206 83.5719
R9078 Vbias.n207 Vbias.t802 83.5719
R9079 Vbias.n183 Vbias.n182 83.5719
R9080 Vbias.t4 Vbias.n183 83.5719
R9081 Vbias.n319 Vbias.n318 83.5719
R9082 Vbias.n318 Vbias.t780 83.5719
R9083 Vbias.n316 Vbias.n189 83.5719
R9084 Vbias.n316 Vbias.t247 83.5719
R9085 Vbias.n353 Vbias.n181 83.5719
R9086 Vbias.t4 Vbias.n181 83.5719
R9087 Vbias.n196 Vbias.n195 83.5719
R9088 Vbias.n195 Vbias.t780 83.5719
R9089 Vbias.n315 Vbias.n314 83.5719
R9090 Vbias.t247 Vbias.n315 83.5719
R9091 Vbias.n271 Vbias.n233 83.5719
R9092 Vbias.t866 Vbias.n233 83.5719
R9093 Vbias.n246 Vbias.n245 83.5719
R9094 Vbias.n245 Vbias.t495 83.5719
R9095 Vbias.n235 Vbias.n234 83.5719
R9096 Vbias.t866 Vbias.n235 83.5719
R9097 Vbias.n263 Vbias.n262 83.5719
R9098 Vbias.n262 Vbias.t495 83.5719
R9099 Vbias.n260 Vbias.n241 83.5719
R9100 Vbias.n260 Vbias.t70 83.5719
R9101 Vbias.n259 Vbias.n258 83.5719
R9102 Vbias.t70 Vbias.n259 83.5719
R9103 Vbias.n1265 Vbias.n1182 83.5719
R9104 Vbias.n1265 Vbias.t188 83.5719
R9105 Vbias.n1267 Vbias.n1171 83.5719
R9106 Vbias.t704 Vbias.n1267 83.5719
R9107 Vbias.n1272 Vbias.n1170 83.5719
R9108 Vbias.t796 Vbias.n1170 83.5719
R9109 Vbias.n1264 Vbias.n1263 83.5719
R9110 Vbias.t188 Vbias.n1264 83.5719
R9111 Vbias.n1258 Vbias.n1179 83.5719
R9112 Vbias.t704 Vbias.n1179 83.5719
R9113 Vbias.n1177 Vbias.n1176 83.5719
R9114 Vbias.t796 Vbias.n1177 83.5719
R9115 Vbias.n1247 Vbias.n1246 83.5719
R9116 Vbias.t315 Vbias.n1247 83.5719
R9117 Vbias.n1185 Vbias.n1183 83.5719
R9118 Vbias.n1183 Vbias.t429 83.5719
R9119 Vbias.n1191 Vbias.n1186 83.5719
R9120 Vbias.t315 Vbias.n1191 83.5719
R9121 Vbias.n1252 Vbias.n1184 83.5719
R9122 Vbias.n1184 Vbias.t429 83.5719
R9123 Vbias.n1234 Vbias.n1213 83.5719
R9124 Vbias.n1234 Vbias.t255 83.5719
R9125 Vbias.n1236 Vbias.n1199 83.5719
R9126 Vbias.t874 Vbias.n1236 83.5719
R9127 Vbias.n1241 Vbias.n1198 83.5719
R9128 Vbias.t126 Vbias.n1198 83.5719
R9129 Vbias.n1233 Vbias.n1232 83.5719
R9130 Vbias.t255 Vbias.n1233 83.5719
R9131 Vbias.n1227 Vbias.n1208 83.5719
R9132 Vbias.t874 Vbias.n1208 83.5719
R9133 Vbias.n1206 Vbias.n1205 83.5719
R9134 Vbias.t126 Vbias.n1206 83.5719
R9135 Vbias.n1077 Vbias.n1075 83.5719
R9136 Vbias.n1075 Vbias.t104 83.5719
R9137 Vbias.n7209 Vbias.n7208 83.5719
R9138 Vbias.t298 Vbias.n7209 83.5719
R9139 Vbias.n1216 Vbias.n1214 83.5719
R9140 Vbias.n1214 Vbias.t336 83.5719
R9141 Vbias.n7214 Vbias.n1076 83.5719
R9142 Vbias.n1076 Vbias.t104 83.5719
R9143 Vbias.n1083 Vbias.n1078 83.5719
R9144 Vbias.t298 Vbias.n1083 83.5719
R9145 Vbias.n1221 Vbias.n1215 83.5719
R9146 Vbias.n1215 Vbias.t336 83.5719
R9147 Vbias.n7221 Vbias.n1073 83.5719
R9148 Vbias.n1073 Vbias.t688 83.5719
R9149 Vbias.n1074 Vbias.n1072 83.5719
R9150 Vbias.n1072 Vbias.t688 83.5719
R9151 Vbias.n1137 Vbias.n1135 83.5719
R9152 Vbias.n1135 Vbias.t32 83.5719
R9153 Vbias.n7133 Vbias.n7132 83.5719
R9154 Vbias.t776 Vbias.n7133 83.5719
R9155 Vbias.n7127 Vbias.n7126 83.5719
R9156 Vbias.n7126 Vbias.t511 83.5719
R9157 Vbias.n7139 Vbias.n1136 83.5719
R9158 Vbias.n1136 Vbias.t32 83.5719
R9159 Vbias.n7135 Vbias.n7134 83.5719
R9160 Vbias.n7134 Vbias.t776 83.5719
R9161 Vbias.n7125 Vbias.n7124 83.5719
R9162 Vbias.t511 Vbias.n7125 83.5719
R9163 Vbias.n1130 Vbias.n1128 83.5719
R9164 Vbias.n1128 Vbias.t845 83.5719
R9165 Vbias.n7150 Vbias.n7149 83.5719
R9166 Vbias.t354 Vbias.n7150 83.5719
R9167 Vbias.n7156 Vbias.n1129 83.5719
R9168 Vbias.n1129 Vbias.t845 83.5719
R9169 Vbias.n7152 Vbias.n7151 83.5719
R9170 Vbias.n7151 Vbias.t354 83.5719
R9171 Vbias.n1127 Vbias.n1126 83.5719
R9172 Vbias.t498 Vbias.n1127 83.5719
R9173 Vbias.n7165 Vbias.n1125 83.5719
R9174 Vbias.t498 Vbias.n1125 83.5719
R9175 Vbias.n1109 Vbias.n1108 83.5719
R9176 Vbias.t62 Vbias.n1109 83.5719
R9177 Vbias.n7174 Vbias.n7173 83.5719
R9178 Vbias.n7173 Vbias.t782 83.5719
R9179 Vbias.n7171 Vbias.n1115 83.5719
R9180 Vbias.n7171 Vbias.t493 83.5719
R9181 Vbias.n7182 Vbias.n1107 83.5719
R9182 Vbias.t62 Vbias.n1107 83.5719
R9183 Vbias.n1122 Vbias.n1121 83.5719
R9184 Vbias.n1121 Vbias.t782 83.5719
R9185 Vbias.n7170 Vbias.n7169 83.5719
R9186 Vbias.t493 Vbias.n7170 83.5719
R9187 Vbias.n7196 Vbias.n1090 83.5719
R9188 Vbias.n7196 Vbias.t176 83.5719
R9189 Vbias.n7191 Vbias.n7190 83.5719
R9190 Vbias.n7190 Vbias.t599 83.5719
R9191 Vbias.n7188 Vbias.n1096 83.5719
R9192 Vbias.n7188 Vbias.t658 83.5719
R9193 Vbias.n7199 Vbias.n1089 83.5719
R9194 Vbias.t176 Vbias.n1089 83.5719
R9195 Vbias.n1103 Vbias.n1102 83.5719
R9196 Vbias.n1102 Vbias.t599 83.5719
R9197 Vbias.n7187 Vbias.n7186 83.5719
R9198 Vbias.t658 Vbias.n7187 83.5719
R9199 Vbias.n6998 Vbias.n6915 83.5719
R9200 Vbias.n6998 Vbias.t40 83.5719
R9201 Vbias.n7000 Vbias.n6904 83.5719
R9202 Vbias.t606 Vbias.n7000 83.5719
R9203 Vbias.n7005 Vbias.n6903 83.5719
R9204 Vbias.t885 Vbias.n6903 83.5719
R9205 Vbias.n6997 Vbias.n6996 83.5719
R9206 Vbias.t40 Vbias.n6997 83.5719
R9207 Vbias.n6991 Vbias.n6912 83.5719
R9208 Vbias.t606 Vbias.n6912 83.5719
R9209 Vbias.n6910 Vbias.n6909 83.5719
R9210 Vbias.t885 Vbias.n6910 83.5719
R9211 Vbias.n6980 Vbias.n6979 83.5719
R9212 Vbias.t534 Vbias.n6980 83.5719
R9213 Vbias.n6918 Vbias.n6916 83.5719
R9214 Vbias.n6916 Vbias.t145 83.5719
R9215 Vbias.n6924 Vbias.n6919 83.5719
R9216 Vbias.t534 Vbias.n6924 83.5719
R9217 Vbias.n6985 Vbias.n6917 83.5719
R9218 Vbias.n6917 Vbias.t145 83.5719
R9219 Vbias.n6967 Vbias.n6946 83.5719
R9220 Vbias.n6967 Vbias.t66 83.5719
R9221 Vbias.n6969 Vbias.n6932 83.5719
R9222 Vbias.t378 Vbias.n6969 83.5719
R9223 Vbias.n6974 Vbias.n6931 83.5719
R9224 Vbias.t544 Vbias.n6931 83.5719
R9225 Vbias.n6966 Vbias.n6965 83.5719
R9226 Vbias.t66 Vbias.n6966 83.5719
R9227 Vbias.n6960 Vbias.n6941 83.5719
R9228 Vbias.t378 Vbias.n6941 83.5719
R9229 Vbias.n6939 Vbias.n6938 83.5719
R9230 Vbias.t544 Vbias.n6939 83.5719
R9231 Vbias.n1158 Vbias.n1156 83.5719
R9232 Vbias.n1156 Vbias.t196 83.5719
R9233 Vbias.n7105 Vbias.n7104 83.5719
R9234 Vbias.t842 Vbias.n7105 83.5719
R9235 Vbias.n6949 Vbias.n6947 83.5719
R9236 Vbias.n6947 Vbias.t497 83.5719
R9237 Vbias.n7110 Vbias.n1157 83.5719
R9238 Vbias.n1157 Vbias.t196 83.5719
R9239 Vbias.n1164 Vbias.n1159 83.5719
R9240 Vbias.t842 Vbias.n1164 83.5719
R9241 Vbias.n6954 Vbias.n6948 83.5719
R9242 Vbias.n6948 Vbias.t497 83.5719
R9243 Vbias.n1155 Vbias.n1153 83.5719
R9244 Vbias.n1153 Vbias.t509 83.5719
R9245 Vbias.n7117 Vbias.n1154 83.5719
R9246 Vbias.n1154 Vbias.t509 83.5719
R9247 Vbias.n1325 Vbias.n1323 83.5719
R9248 Vbias.n1323 Vbias.t239 83.5719
R9249 Vbias.n7027 Vbias.n7026 83.5719
R9250 Vbias.t496 Vbias.n7027 83.5719
R9251 Vbias.n7021 Vbias.n7020 83.5719
R9252 Vbias.n7020 Vbias.t230 83.5719
R9253 Vbias.n7033 Vbias.n1324 83.5719
R9254 Vbias.n1324 Vbias.t239 83.5719
R9255 Vbias.n7029 Vbias.n7028 83.5719
R9256 Vbias.n7028 Vbias.t496 83.5719
R9257 Vbias.n7019 Vbias.n7018 83.5719
R9258 Vbias.t230 Vbias.n7019 83.5719
R9259 Vbias.n1318 Vbias.n1316 83.5719
R9260 Vbias.n1316 Vbias.t542 83.5719
R9261 Vbias.n7044 Vbias.n7043 83.5719
R9262 Vbias.t556 Vbias.n7044 83.5719
R9263 Vbias.n7050 Vbias.n1317 83.5719
R9264 Vbias.n1317 Vbias.t542 83.5719
R9265 Vbias.n7046 Vbias.n7045 83.5719
R9266 Vbias.n7045 Vbias.t556 83.5719
R9267 Vbias.n1315 Vbias.n1314 83.5719
R9268 Vbias.t381 Vbias.n1315 83.5719
R9269 Vbias.n7059 Vbias.n1313 83.5719
R9270 Vbias.t381 Vbias.n1313 83.5719
R9271 Vbias.n1296 Vbias.n1295 83.5719
R9272 Vbias.t198 Vbias.n1296 83.5719
R9273 Vbias.n7068 Vbias.n7067 83.5719
R9274 Vbias.n7067 Vbias.t355 83.5719
R9275 Vbias.n7065 Vbias.n1302 83.5719
R9276 Vbias.n7065 Vbias.t715 83.5719
R9277 Vbias.n7076 Vbias.n1294 83.5719
R9278 Vbias.t198 Vbias.n1294 83.5719
R9279 Vbias.n1310 Vbias.n1309 83.5719
R9280 Vbias.n1309 Vbias.t355 83.5719
R9281 Vbias.n7064 Vbias.n7063 83.5719
R9282 Vbias.t715 Vbias.n7064 83.5719
R9283 Vbias.n7090 Vbias.n1277 83.5719
R9284 Vbias.n7090 Vbias.t114 83.5719
R9285 Vbias.n7085 Vbias.n7084 83.5719
R9286 Vbias.n7084 Vbias.t636 83.5719
R9287 Vbias.n7082 Vbias.n1283 83.5719
R9288 Vbias.n7082 Vbias.t593 83.5719
R9289 Vbias.n7093 Vbias.n1276 83.5719
R9290 Vbias.t114 Vbias.n1276 83.5719
R9291 Vbias.n1290 Vbias.n1289 83.5719
R9292 Vbias.n1289 Vbias.t636 83.5719
R9293 Vbias.n7081 Vbias.n7080 83.5719
R9294 Vbias.t593 Vbias.n7081 83.5719
R9295 Vbias.n6831 Vbias.n6830 83.5719
R9296 Vbias.n6830 Vbias.t118 83.5719
R9297 Vbias.n6822 Vbias.n6821 83.5719
R9298 Vbias.t160 Vbias.n6822 83.5719
R9299 Vbias.n6817 Vbias.n1400 83.5719
R9300 Vbias.t361 Vbias.n1400 83.5719
R9301 Vbias.n6829 Vbias.n6828 83.5719
R9302 Vbias.t118 Vbias.n6829 83.5719
R9303 Vbias.n6824 Vbias.n6823 83.5719
R9304 Vbias.n6823 Vbias.t160 83.5719
R9305 Vbias.n1555 Vbias.n1554 83.5719
R9306 Vbias.n1555 Vbias.t361 83.5719
R9307 Vbias.n1378 Vbias.n1376 83.5719
R9308 Vbias.n1376 Vbias.t488 83.5719
R9309 Vbias.n6838 Vbias.n6837 83.5719
R9310 Vbias.t754 Vbias.n6838 83.5719
R9311 Vbias.n6843 Vbias.n1377 83.5719
R9312 Vbias.n1377 Vbias.t488 83.5719
R9313 Vbias.n1384 Vbias.n1379 83.5719
R9314 Vbias.t754 Vbias.n1384 83.5719
R9315 Vbias.n1365 Vbias.n1363 83.5719
R9316 Vbias.n1363 Vbias.t122 83.5719
R9317 Vbias.n6861 Vbias.n6860 83.5719
R9318 Vbias.t579 Vbias.n6861 83.5719
R9319 Vbias.n6855 Vbias.n6854 83.5719
R9320 Vbias.n6854 Vbias.t492 83.5719
R9321 Vbias.n6866 Vbias.n1364 83.5719
R9322 Vbias.n1364 Vbias.t122 83.5719
R9323 Vbias.n1371 Vbias.n1366 83.5719
R9324 Vbias.t579 Vbias.n1371 83.5719
R9325 Vbias.n6853 Vbias.n6852 83.5719
R9326 Vbias.t492 Vbias.n6853 83.5719
R9327 Vbias.n1352 Vbias.n1350 83.5719
R9328 Vbias.n1350 Vbias.t222 83.5719
R9329 Vbias.n6884 Vbias.n6883 83.5719
R9330 Vbias.t1 Vbias.n6884 83.5719
R9331 Vbias.n6878 Vbias.n6877 83.5719
R9332 Vbias.n6877 Vbias.t380 83.5719
R9333 Vbias.n6889 Vbias.n1351 83.5719
R9334 Vbias.n1351 Vbias.t222 83.5719
R9335 Vbias.n1358 Vbias.n1353 83.5719
R9336 Vbias.t1 Vbias.n1358 83.5719
R9337 Vbias.n6876 Vbias.n6875 83.5719
R9338 Vbias.t380 Vbias.n6876 83.5719
R9339 Vbias.n6897 Vbias.n6896 83.5719
R9340 Vbias.n6896 Vbias.t420 83.5719
R9341 Vbias.n6895 Vbias.n6894 83.5719
R9342 Vbias.t420 Vbias.n6895 83.5719
R9343 Vbias.n6064 Vbias.n6063 83.5719
R9344 Vbias.t267 Vbias.n6064 83.5719
R9345 Vbias.n6069 Vbias.n6068 83.5719
R9346 Vbias.n6068 Vbias.t541 83.5719
R9347 Vbias.n6072 Vbias.n6071 83.5719
R9348 Vbias.n6072 Vbias.t731 83.5719
R9349 Vbias.n6808 Vbias.n1407 83.5719
R9350 Vbias.t267 Vbias.n1407 83.5719
R9351 Vbias.n6810 Vbias.n1405 83.5719
R9352 Vbias.t541 Vbias.n1405 83.5719
R9353 Vbias.n6812 Vbias.n1403 83.5719
R9354 Vbias.t731 Vbias.n1403 83.5719
R9355 Vbias.n1415 Vbias.n1414 83.5719
R9356 Vbias.t490 Vbias.n1415 83.5719
R9357 Vbias.n6058 Vbias.n6057 83.5719
R9358 Vbias.n6058 Vbias.t756 83.5719
R9359 Vbias.n6802 Vbias.n1413 83.5719
R9360 Vbias.t490 Vbias.n1413 83.5719
R9361 Vbias.n6804 Vbias.n1411 83.5719
R9362 Vbias.t756 Vbias.n1411 83.5719
R9363 Vbias.n1418 Vbias.n1416 83.5719
R9364 Vbias.n1416 Vbias.t330 83.5719
R9365 Vbias.n6795 Vbias.n1417 83.5719
R9366 Vbias.n1417 Vbias.t330 83.5719
R9367 Vbias.n6768 Vbias.n6767 83.5719
R9368 Vbias.n6768 Vbias.t265 83.5719
R9369 Vbias.n6765 Vbias.n6764 83.5719
R9370 Vbias.n6764 Vbias.t799 83.5719
R9371 Vbias.n6757 Vbias.n6756 83.5719
R9372 Vbias.t781 Vbias.n6757 83.5719
R9373 Vbias.n6787 Vbias.n1427 83.5719
R9374 Vbias.t265 Vbias.n1427 83.5719
R9375 Vbias.n6789 Vbias.n1425 83.5719
R9376 Vbias.t799 Vbias.n1425 83.5719
R9377 Vbias.n6791 Vbias.n1423 83.5719
R9378 Vbias.t781 Vbias.n1423 83.5719
R9379 Vbias.n1343 Vbias.n1341 83.5719
R9380 Vbias.n1341 Vbias.t92 83.5719
R9381 Vbias.n6779 Vbias.n6778 83.5719
R9382 Vbias.t647 Vbias.n6779 83.5719
R9383 Vbias.n6773 Vbias.n6772 83.5719
R9384 Vbias.n6772 Vbias.t340 83.5719
R9385 Vbias.n7011 Vbias.n1342 83.5719
R9386 Vbias.n1342 Vbias.t92 83.5719
R9387 Vbias.n6781 Vbias.n6780 83.5719
R9388 Vbias.n6780 Vbias.t647 83.5719
R9389 Vbias.n6783 Vbias.n1430 83.5719
R9390 Vbias.t340 Vbias.n1430 83.5719
R9391 Vbias.n5973 Vbias.n5972 83.5719
R9392 Vbias.n5972 Vbias.t60 83.5719
R9393 Vbias.n5964 Vbias.n5963 83.5719
R9394 Vbias.t569 Vbias.n5964 83.5719
R9395 Vbias.n5959 Vbias.n1611 83.5719
R9396 Vbias.t680 Vbias.n1611 83.5719
R9397 Vbias.n5971 Vbias.n5970 83.5719
R9398 Vbias.t60 Vbias.n5971 83.5719
R9399 Vbias.n5966 Vbias.n5965 83.5719
R9400 Vbias.n5965 Vbias.t569 83.5719
R9401 Vbias.n1636 Vbias.n1635 83.5719
R9402 Vbias.n1636 Vbias.t680 83.5719
R9403 Vbias.n1589 Vbias.n1587 83.5719
R9404 Vbias.n1587 Vbias.t318 83.5719
R9405 Vbias.n5980 Vbias.n5979 83.5719
R9406 Vbias.t456 Vbias.n5980 83.5719
R9407 Vbias.n5985 Vbias.n1588 83.5719
R9408 Vbias.n1588 Vbias.t318 83.5719
R9409 Vbias.n1595 Vbias.n1590 83.5719
R9410 Vbias.t456 Vbias.n1595 83.5719
R9411 Vbias.n1576 Vbias.n1574 83.5719
R9412 Vbias.n1574 Vbias.t94 83.5719
R9413 Vbias.n6003 Vbias.n6002 83.5719
R9414 Vbias.t852 Vbias.n6003 83.5719
R9415 Vbias.n5997 Vbias.n5996 83.5719
R9416 Vbias.n5996 Vbias.t752 83.5719
R9417 Vbias.n6008 Vbias.n1575 83.5719
R9418 Vbias.n1575 Vbias.t94 83.5719
R9419 Vbias.n1582 Vbias.n1577 83.5719
R9420 Vbias.t852 Vbias.n1582 83.5719
R9421 Vbias.n5995 Vbias.n5994 83.5719
R9422 Vbias.t752 Vbias.n5995 83.5719
R9423 Vbias.n1563 Vbias.n1561 83.5719
R9424 Vbias.n1561 Vbias.t243 83.5719
R9425 Vbias.n6029 Vbias.n6028 83.5719
R9426 Vbias.t732 Vbias.n6029 83.5719
R9427 Vbias.n6020 Vbias.n6019 83.5719
R9428 Vbias.n6019 Vbias.t660 83.5719
R9429 Vbias.n6034 Vbias.n1562 83.5719
R9430 Vbias.n1562 Vbias.t243 83.5719
R9431 Vbias.n1569 Vbias.n1564 83.5719
R9432 Vbias.t732 Vbias.n1569 83.5719
R9433 Vbias.n6018 Vbias.n6017 83.5719
R9434 Vbias.t660 Vbias.n6018 83.5719
R9435 Vbias.n1560 Vbias.n1558 83.5719
R9436 Vbias.n1558 Vbias.t728 83.5719
R9437 Vbias.n6041 Vbias.n1559 83.5719
R9438 Vbias.n1559 Vbias.t728 83.5719
R9439 Vbias.n1793 Vbias.n1792 83.5719
R9440 Vbias.n1793 Vbias.t182 83.5719
R9441 Vbias.n6089 Vbias.n1543 83.5719
R9442 Vbias.n1543 Vbias.t182 83.5719
R9443 Vbias.n1553 Vbias.n1552 83.5719
R9444 Vbias.t76 Vbias.n1553 83.5719
R9445 Vbias.n1784 Vbias.n1783 83.5719
R9446 Vbias.n1783 Vbias.t305 83.5719
R9447 Vbias.n1787 Vbias.n1786 83.5719
R9448 Vbias.n1787 Vbias.t500 83.5719
R9449 Vbias.n6081 Vbias.n1551 83.5719
R9450 Vbias.t76 Vbias.n1551 83.5719
R9451 Vbias.n6083 Vbias.n1549 83.5719
R9452 Vbias.n1549 Vbias.t305 83.5719
R9453 Vbias.n6085 Vbias.n1547 83.5719
R9454 Vbias.t500 Vbias.n1547 83.5719
R9455 Vbias.n1904 Vbias.n1900 83.5719
R9456 Vbias.n1904 Vbias.t644 83.5719
R9457 Vbias.n1906 Vbias.n1882 83.5719
R9458 Vbias.t883 Vbias.n1906 83.5719
R9459 Vbias.n1913 Vbias.n1912 83.5719
R9460 Vbias.n1912 Vbias.t758 83.5719
R9461 Vbias.n1903 Vbias.n1902 83.5719
R9462 Vbias.t644 Vbias.n1903 83.5719
R9463 Vbias.n1908 Vbias.n1907 83.5719
R9464 Vbias.n1907 Vbias.t883 83.5719
R9465 Vbias.n1911 Vbias.n1910 83.5719
R9466 Vbias.t758 Vbias.n1911 83.5719
R9467 Vbias.n1972 Vbias.n1971 83.5719
R9468 Vbias.t763 Vbias.n1972 83.5719
R9469 Vbias.n1981 Vbias.n1980 83.5719
R9470 Vbias.n1980 Vbias.t436 83.5719
R9471 Vbias.n1963 Vbias.n1950 83.5719
R9472 Vbias.t746 Vbias.n1963 83.5719
R9473 Vbias.n1974 Vbias.n1973 83.5719
R9474 Vbias.n1973 Vbias.t763 83.5719
R9475 Vbias.n1979 Vbias.n1978 83.5719
R9476 Vbias.t436 Vbias.n1979 83.5719
R9477 Vbias.n1965 Vbias.n1964 83.5719
R9478 Vbias.n1964 Vbias.t746 83.5719
R9479 Vbias.n6112 Vbias.n6111 83.5719
R9480 Vbias.t594 Vbias.n6112 83.5719
R9481 Vbias.n6121 Vbias.n6120 83.5719
R9482 Vbias.n6120 Vbias.t142 83.5719
R9483 Vbias.n6103 Vbias.n1510 83.5719
R9484 Vbias.t140 Vbias.n6103 83.5719
R9485 Vbias.n6114 Vbias.n6113 83.5719
R9486 Vbias.n6113 Vbias.t594 83.5719
R9487 Vbias.n6119 Vbias.n6118 83.5719
R9488 Vbias.t142 Vbias.n6119 83.5719
R9489 Vbias.n6105 Vbias.n6104 83.5719
R9490 Vbias.n6104 Vbias.t140 83.5719
R9491 Vbias.n2014 Vbias.n1986 83.5719
R9492 Vbias.t853 Vbias.n1986 83.5719
R9493 Vbias.n1998 Vbias.n1997 83.5719
R9494 Vbias.n1997 Vbias.t5 83.5719
R9495 Vbias.n2002 Vbias.n2001 83.5719
R9496 Vbias.t662 Vbias.n2002 83.5719
R9497 Vbias.n2011 Vbias.n1987 83.5719
R9498 Vbias.n2011 Vbias.t853 83.5719
R9499 Vbias.n2006 Vbias.n2005 83.5719
R9500 Vbias.n2005 Vbias.t5 83.5719
R9501 Vbias.n2003 Vbias.n1993 83.5719
R9502 Vbias.n2003 Vbias.t662 83.5719
R9503 Vbias.n1938 Vbias.n1937 83.5719
R9504 Vbias.t422 Vbias.n1938 83.5719
R9505 Vbias.n1947 Vbias.n1946 83.5719
R9506 Vbias.n1946 Vbias.t870 83.5719
R9507 Vbias.n1929 Vbias.n1916 83.5719
R9508 Vbias.t868 Vbias.n1929 83.5719
R9509 Vbias.n1940 Vbias.n1939 83.5719
R9510 Vbias.n1939 Vbias.t422 83.5719
R9511 Vbias.n1945 Vbias.n1944 83.5719
R9512 Vbias.t870 Vbias.n1945 83.5719
R9513 Vbias.n1931 Vbias.n1930 83.5719
R9514 Vbias.n1930 Vbias.t868 83.5719
R9515 Vbias.n1872 Vbias.n1871 83.5719
R9516 Vbias.t358 Vbias.n1872 83.5719
R9517 Vbias.n1879 Vbias.n1878 83.5719
R9518 Vbias.n1878 Vbias.t779 83.5719
R9519 Vbias.n1861 Vbias.n1848 83.5719
R9520 Vbias.t427 Vbias.n1861 83.5719
R9521 Vbias.n1874 Vbias.n1873 83.5719
R9522 Vbias.n1873 Vbias.t358 83.5719
R9523 Vbias.n1877 Vbias.n1876 83.5719
R9524 Vbias.t779 Vbias.n1877 83.5719
R9525 Vbias.n1863 Vbias.n1862 83.5719
R9526 Vbias.n1862 Vbias.t427 83.5719
R9527 Vbias.n1819 Vbias.n1818 83.5719
R9528 Vbias.n1818 Vbias.t560 83.5719
R9529 Vbias.n1812 Vbias.n1753 83.5719
R9530 Vbias.t795 Vbias.n1812 83.5719
R9531 Vbias.n1810 Vbias.n1754 83.5719
R9532 Vbias.n1810 Vbias.t793 83.5719
R9533 Vbias.n1817 Vbias.n1816 83.5719
R9534 Vbias.t560 Vbias.n1817 83.5719
R9535 Vbias.n1814 Vbias.n1813 83.5719
R9536 Vbias.n1813 Vbias.t795 83.5719
R9537 Vbias.n1809 Vbias.n1808 83.5719
R9538 Vbias.t793 Vbias.n1809 83.5719
R9539 Vbias.n1535 Vbias.n1533 83.5719
R9540 Vbias.t815 Vbias.n1533 83.5719
R9541 Vbias.n6097 Vbias.n1534 83.5719
R9542 Vbias.t815 Vbias.n1534 83.5719
R9543 Vbias.n1796 Vbias.n1795 83.5719
R9544 Vbias.n1795 Vbias.t414 83.5719
R9545 Vbias.n1799 Vbias.n1798 83.5719
R9546 Vbias.t317 Vbias.n1799 83.5719
R9547 Vbias.n6091 Vbias.n1541 83.5719
R9548 Vbias.t414 Vbias.n1541 83.5719
R9549 Vbias.n6093 Vbias.n1539 83.5719
R9550 Vbias.t317 Vbias.n1539 83.5719
R9551 Vbias.n5930 Vbias.n1629 83.5719
R9552 Vbias.n5930 Vbias.t212 83.5719
R9553 Vbias.n5926 Vbias.n5925 83.5719
R9554 Vbias.t730 Vbias.n5926 83.5719
R9555 Vbias.n5922 Vbias.n5921 83.5719
R9556 Vbias.n5921 Vbias.t155 83.5719
R9557 Vbias.n5950 Vbias.n1618 83.5719
R9558 Vbias.t212 Vbias.n1618 83.5719
R9559 Vbias.n5952 Vbias.n1616 83.5719
R9560 Vbias.t730 Vbias.n1616 83.5719
R9561 Vbias.n5954 Vbias.n1614 83.5719
R9562 Vbias.t155 Vbias.n1614 83.5719
R9563 Vbias.n5941 Vbias.n1626 83.5719
R9564 Vbias.n5941 Vbias.t750 83.5719
R9565 Vbias.n5937 Vbias.n5936 83.5719
R9566 Vbias.t867 Vbias.n5937 83.5719
R9567 Vbias.n5944 Vbias.n1625 83.5719
R9568 Vbias.t750 Vbias.n1625 83.5719
R9569 Vbias.n5946 Vbias.n1623 83.5719
R9570 Vbias.t867 Vbias.n1623 83.5719
R9571 Vbias.n5406 Vbias.n5286 83.5719
R9572 Vbias.n5406 Vbias.t98 83.5719
R9573 Vbias.n5408 Vbias.n5274 83.5719
R9574 Vbias.t635 Vbias.n5408 83.5719
R9575 Vbias.n5413 Vbias.n5273 83.5719
R9576 Vbias.t532 Vbias.n5273 83.5719
R9577 Vbias.n5405 Vbias.n5404 83.5719
R9578 Vbias.t98 Vbias.n5405 83.5719
R9579 Vbias.n5399 Vbias.n5283 83.5719
R9580 Vbias.t635 Vbias.n5283 83.5719
R9581 Vbias.n5281 Vbias.n5280 83.5719
R9582 Vbias.t532 Vbias.n5281 83.5719
R9583 Vbias.n5388 Vbias.n5387 83.5719
R9584 Vbias.t404 Vbias.n5388 83.5719
R9585 Vbias.n5289 Vbias.n5287 83.5719
R9586 Vbias.n5287 Vbias.t413 83.5719
R9587 Vbias.n5295 Vbias.n5290 83.5719
R9588 Vbias.t404 Vbias.n5295 83.5719
R9589 Vbias.n5393 Vbias.n5288 83.5719
R9590 Vbias.n5288 Vbias.t413 83.5719
R9591 Vbias.n5375 Vbias.n5315 83.5719
R9592 Vbias.n5375 Vbias.t22 83.5719
R9593 Vbias.n5377 Vbias.n5303 83.5719
R9594 Vbias.t642 Vbias.n5377 83.5719
R9595 Vbias.n5382 Vbias.n5302 83.5719
R9596 Vbias.t13 Vbias.n5302 83.5719
R9597 Vbias.n5374 Vbias.n5373 83.5719
R9598 Vbias.t22 Vbias.n5374 83.5719
R9599 Vbias.n5368 Vbias.n5312 83.5719
R9600 Vbias.t642 Vbias.n5312 83.5719
R9601 Vbias.n5310 Vbias.n5309 83.5719
R9602 Vbias.t13 Vbias.n5310 83.5719
R9603 Vbias.n5354 Vbias.n5353 83.5719
R9604 Vbias.n5353 Vbias.t194 83.5719
R9605 Vbias.n5358 Vbias.n5357 83.5719
R9606 Vbias.t154 Vbias.n5358 83.5719
R9607 Vbias.n5318 Vbias.n5316 83.5719
R9608 Vbias.n5316 Vbias.t814 83.5719
R9609 Vbias.n5352 Vbias.n5351 83.5719
R9610 Vbias.t194 Vbias.n5352 83.5719
R9611 Vbias.n5360 Vbias.n5359 83.5719
R9612 Vbias.n5359 Vbias.t154 83.5719
R9613 Vbias.n5362 Vbias.n5317 83.5719
R9614 Vbias.n5317 Vbias.t814 83.5719
R9615 Vbias.n5343 Vbias.n5338 83.5719
R9616 Vbias.n5338 Vbias.t742 83.5719
R9617 Vbias.n5346 Vbias.n5339 83.5719
R9618 Vbias.n5339 Vbias.t742 83.5719
R9619 Vbias.n5422 Vbias.n5421 83.5719
R9620 Vbias.t178 Vbias.n5422 83.5719
R9621 Vbias.n5431 Vbias.n5430 83.5719
R9622 Vbias.n5431 Vbias.t479 83.5719
R9623 Vbias.n2291 Vbias.n2289 83.5719
R9624 Vbias.n2289 Vbias.t710 83.5719
R9625 Vbias.n5476 Vbias.n5420 83.5719
R9626 Vbias.t178 Vbias.n5420 83.5719
R9627 Vbias.n5478 Vbias.n5418 83.5719
R9628 Vbias.t479 Vbias.n5418 83.5719
R9629 Vbias.n5481 Vbias.n2290 83.5719
R9630 Vbias.n2290 Vbias.t710 83.5719
R9631 Vbias.n5444 Vbias.n5443 83.5719
R9632 Vbias.t11 Vbias.n5444 83.5719
R9633 Vbias.n5438 Vbias.n5436 83.5719
R9634 Vbias.n5436 Vbias.t736 83.5719
R9635 Vbias.n5466 Vbias.n5442 83.5719
R9636 Vbias.t11 Vbias.n5442 83.5719
R9637 Vbias.n5469 Vbias.n5437 83.5719
R9638 Vbias.n5437 Vbias.t736 83.5719
R9639 Vbias.n5453 Vbias.n5451 83.5719
R9640 Vbias.n5451 Vbias.t395 83.5719
R9641 Vbias.n5459 Vbias.n5452 83.5719
R9642 Vbias.n5452 Vbias.t395 83.5719
R9643 Vbias.n1658 Vbias.n1656 83.5719
R9644 Vbias.n1656 Vbias.t237 83.5719
R9645 Vbias.n5888 Vbias.n5887 83.5719
R9646 Vbias.t449 Vbias.n5888 83.5719
R9647 Vbias.n5882 Vbias.n5881 83.5719
R9648 Vbias.n5881 Vbias.t403 83.5719
R9649 Vbias.n5894 Vbias.n1657 83.5719
R9650 Vbias.n1657 Vbias.t237 83.5719
R9651 Vbias.n5890 Vbias.n5889 83.5719
R9652 Vbias.n5889 Vbias.t449 83.5719
R9653 Vbias.n5880 Vbias.n5879 83.5719
R9654 Vbias.t403 Vbias.n5880 83.5719
R9655 Vbias.n1642 Vbias.n1640 83.5719
R9656 Vbias.n1640 Vbias.t26 83.5719
R9657 Vbias.n5908 Vbias.n5907 83.5719
R9658 Vbias.t757 Vbias.n5908 83.5719
R9659 Vbias.n5902 Vbias.n5901 83.5719
R9660 Vbias.n5901 Vbias.t592 83.5719
R9661 Vbias.n5914 Vbias.n1641 83.5719
R9662 Vbias.n1641 Vbias.t26 83.5719
R9663 Vbias.n5910 Vbias.n5909 83.5719
R9664 Vbias.n5909 Vbias.t757 83.5719
R9665 Vbias.n5900 Vbias.n5899 83.5719
R9666 Vbias.t592 Vbias.n5900 83.5719
R9667 Vbias.n5200 Vbias.n5199 83.5719
R9668 Vbias.n5199 Vbias.t54 83.5719
R9669 Vbias.n5191 Vbias.n5190 83.5719
R9670 Vbias.t347 Vbias.n5191 83.5719
R9671 Vbias.n5186 Vbias.n2348 83.5719
R9672 Vbias.t765 Vbias.n2348 83.5719
R9673 Vbias.n5198 Vbias.n5197 83.5719
R9674 Vbias.t54 Vbias.n5198 83.5719
R9675 Vbias.n5193 Vbias.n5192 83.5719
R9676 Vbias.n5192 Vbias.t347 83.5719
R9677 Vbias.n2368 Vbias.n2367 83.5719
R9678 Vbias.n2368 Vbias.t765 83.5719
R9679 Vbias.n2326 Vbias.n2324 83.5719
R9680 Vbias.n2324 Vbias.t664 83.5719
R9681 Vbias.n5207 Vbias.n5206 83.5719
R9682 Vbias.t711 Vbias.n5207 83.5719
R9683 Vbias.n5212 Vbias.n2325 83.5719
R9684 Vbias.n2325 Vbias.t664 83.5719
R9685 Vbias.n2332 Vbias.n2327 83.5719
R9686 Vbias.t711 Vbias.n2332 83.5719
R9687 Vbias.n2313 Vbias.n2311 83.5719
R9688 Vbias.n2311 Vbias.t28 83.5719
R9689 Vbias.n5230 Vbias.n5229 83.5719
R9690 Vbias.t531 Vbias.n5230 83.5719
R9691 Vbias.n5224 Vbias.n5223 83.5719
R9692 Vbias.n5223 Vbias.t685 83.5719
R9693 Vbias.n5235 Vbias.n2312 83.5719
R9694 Vbias.n2312 Vbias.t28 83.5719
R9695 Vbias.n2319 Vbias.n2314 83.5719
R9696 Vbias.t531 Vbias.n2319 83.5719
R9697 Vbias.n5222 Vbias.n5221 83.5719
R9698 Vbias.t685 Vbias.n5222 83.5719
R9699 Vbias.n2300 Vbias.n2298 83.5719
R9700 Vbias.n2298 Vbias.t216 83.5719
R9701 Vbias.n5253 Vbias.n5252 83.5719
R9702 Vbias.t139 Vbias.n5253 83.5719
R9703 Vbias.n5247 Vbias.n5246 83.5719
R9704 Vbias.n5246 Vbias.t394 83.5719
R9705 Vbias.n5258 Vbias.n2299 83.5719
R9706 Vbias.n2299 Vbias.t216 83.5719
R9707 Vbias.n2306 Vbias.n2301 83.5719
R9708 Vbias.t139 Vbias.n2306 83.5719
R9709 Vbias.n5245 Vbias.n5244 83.5719
R9710 Vbias.t394 Vbias.n5245 83.5719
R9711 Vbias.n5267 Vbias.n5266 83.5719
R9712 Vbias.n5266 Vbias.t707 83.5719
R9713 Vbias.n5265 Vbias.n5264 83.5719
R9714 Vbias.t707 Vbias.n5265 83.5719
R9715 Vbias.n5137 Vbias.n5136 83.5719
R9716 Vbias.n5137 Vbias.t220 83.5719
R9717 Vbias.n5134 Vbias.n5133 83.5719
R9718 Vbias.n5133 Vbias.t520 83.5719
R9719 Vbias.n5126 Vbias.n5125 83.5719
R9720 Vbias.t605 Vbias.n5126 83.5719
R9721 Vbias.n5177 Vbias.n2355 83.5719
R9722 Vbias.t220 Vbias.n2355 83.5719
R9723 Vbias.n5179 Vbias.n2353 83.5719
R9724 Vbias.t520 Vbias.n2353 83.5719
R9725 Vbias.n5181 Vbias.n2351 83.5719
R9726 Vbias.t605 Vbias.n2351 83.5719
R9727 Vbias.n2363 Vbias.n2362 83.5719
R9728 Vbias.t686 Vbias.n2363 83.5719
R9729 Vbias.n5144 Vbias.n5143 83.5719
R9730 Vbias.n5144 Vbias.t406 83.5719
R9731 Vbias.n5171 Vbias.n2361 83.5719
R9732 Vbias.t686 Vbias.n2361 83.5719
R9733 Vbias.n5173 Vbias.n2359 83.5719
R9734 Vbias.t406 Vbias.n2359 83.5719
R9735 Vbias.n5151 Vbias.n5149 83.5719
R9736 Vbias.n5149 Vbias.t586 83.5719
R9737 Vbias.n5164 Vbias.n5150 83.5719
R9738 Vbias.n5150 Vbias.t586 83.5719
R9739 Vbias.n2256 Vbias.n2255 83.5719
R9740 Vbias.t259 Vbias.n2256 83.5719
R9741 Vbias.n2260 Vbias.n2259 83.5719
R9742 Vbias.n2259 Vbias.t554 83.5719
R9743 Vbias.n5154 Vbias.n5152 83.5719
R9744 Vbias.n5152 Vbias.t666 83.5719
R9745 Vbias.n5501 Vbias.n2254 83.5719
R9746 Vbias.t259 Vbias.n2254 83.5719
R9747 Vbias.n5504 Vbias.n2250 83.5719
R9748 Vbias.n2250 Vbias.t554 83.5719
R9749 Vbias.n5153 Vbias.n2249 83.5719
R9750 Vbias.n5153 Vbias.t666 83.5719
R9751 Vbias.n2274 Vbias.n2273 83.5719
R9752 Vbias.t100 Vbias.n2274 83.5719
R9753 Vbias.n2283 Vbias.n2282 83.5719
R9754 Vbias.n2283 Vbias.t894 83.5719
R9755 Vbias.n2267 Vbias.n2265 83.5719
R9756 Vbias.n2265 Vbias.t339 83.5719
R9757 Vbias.n5489 Vbias.n2272 83.5719
R9758 Vbias.t100 Vbias.n2272 83.5719
R9759 Vbias.n5491 Vbias.n2270 83.5719
R9760 Vbias.t894 Vbias.n2270 83.5719
R9761 Vbias.n5494 Vbias.n2266 83.5719
R9762 Vbias.n2266 Vbias.t339 83.5719
R9763 Vbias.n2574 Vbias.n2454 83.5719
R9764 Vbias.n2574 Vbias.t38 83.5719
R9765 Vbias.n2576 Vbias.n2442 83.5719
R9766 Vbias.t762 Vbias.n2576 83.5719
R9767 Vbias.n2581 Vbias.n2441 83.5719
R9768 Vbias.t851 Vbias.n2441 83.5719
R9769 Vbias.n2573 Vbias.n2572 83.5719
R9770 Vbias.t38 Vbias.n2573 83.5719
R9771 Vbias.n2567 Vbias.n2451 83.5719
R9772 Vbias.t762 Vbias.n2451 83.5719
R9773 Vbias.n2449 Vbias.n2448 83.5719
R9774 Vbias.t851 Vbias.n2449 83.5719
R9775 Vbias.n2556 Vbias.n2555 83.5719
R9776 Vbias.t690 Vbias.n2556 83.5719
R9777 Vbias.n2457 Vbias.n2455 83.5719
R9778 Vbias.n2455 Vbias.t546 83.5719
R9779 Vbias.n2463 Vbias.n2458 83.5719
R9780 Vbias.t690 Vbias.n2463 83.5719
R9781 Vbias.n2561 Vbias.n2456 83.5719
R9782 Vbias.n2456 Vbias.t546 83.5719
R9783 Vbias.n2543 Vbias.n2483 83.5719
R9784 Vbias.n2543 Vbias.t108 83.5719
R9785 Vbias.n2545 Vbias.n2471 83.5719
R9786 Vbias.t598 Vbias.n2545 83.5719
R9787 Vbias.n2550 Vbias.n2470 83.5719
R9788 Vbias.t9 Vbias.n2470 83.5719
R9789 Vbias.n2542 Vbias.n2541 83.5719
R9790 Vbias.t108 Vbias.n2542 83.5719
R9791 Vbias.n2536 Vbias.n2480 83.5719
R9792 Vbias.t598 Vbias.n2480 83.5719
R9793 Vbias.n2478 Vbias.n2477 83.5719
R9794 Vbias.t9 Vbias.n2478 83.5719
R9795 Vbias.n2522 Vbias.n2521 83.5719
R9796 Vbias.n2521 Vbias.t263 83.5719
R9797 Vbias.n2526 Vbias.n2525 83.5719
R9798 Vbias.t603 Vbias.n2526 83.5719
R9799 Vbias.n2486 Vbias.n2484 83.5719
R9800 Vbias.n2484 Vbias.t480 83.5719
R9801 Vbias.n2520 Vbias.n2519 83.5719
R9802 Vbias.t263 Vbias.n2520 83.5719
R9803 Vbias.n2528 Vbias.n2527 83.5719
R9804 Vbias.n2527 Vbias.t603 83.5719
R9805 Vbias.n2530 Vbias.n2485 83.5719
R9806 Vbias.n2485 Vbias.t480 83.5719
R9807 Vbias.n2511 Vbias.n2506 83.5719
R9808 Vbias.n2506 Vbias.t601 83.5719
R9809 Vbias.n2514 Vbias.n2507 83.5719
R9810 Vbias.n2507 Vbias.t601 83.5719
R9811 Vbias.n2411 Vbias.n2410 83.5719
R9812 Vbias.t640 Vbias.n2411 83.5719
R9813 Vbias.n5061 Vbias.n5060 83.5719
R9814 Vbias.n5060 Vbias.t892 83.5719
R9815 Vbias.n5071 Vbias.n2409 83.5719
R9816 Vbias.t640 Vbias.n2409 83.5719
R9817 Vbias.n2416 Vbias.n2415 83.5719
R9818 Vbias.n2416 Vbias.t892 83.5719
R9819 Vbias.n2405 Vbias.n2403 83.5719
R9820 Vbias.n2403 Vbias.t385 83.5719
R9821 Vbias.n5076 Vbias.n2404 83.5719
R9822 Vbias.n2404 Vbias.t385 83.5719
R9823 Vbias.n2390 Vbias.n2388 83.5719
R9824 Vbias.n2388 Vbias.t271 83.5719
R9825 Vbias.n5091 Vbias.n5090 83.5719
R9826 Vbias.t722 Vbias.n5091 83.5719
R9827 Vbias.n5085 Vbias.n5084 83.5719
R9828 Vbias.n5084 Vbias.t287 83.5719
R9829 Vbias.n5097 Vbias.n2389 83.5719
R9830 Vbias.n2389 Vbias.t271 83.5719
R9831 Vbias.n5093 Vbias.n5092 83.5719
R9832 Vbias.n5092 Vbias.t722 83.5719
R9833 Vbias.n5083 Vbias.n5082 83.5719
R9834 Vbias.t287 Vbias.n5083 83.5719
R9835 Vbias.n2374 Vbias.n2372 83.5719
R9836 Vbias.n2372 Vbias.t56 83.5719
R9837 Vbias.n5111 Vbias.n5110 83.5719
R9838 Vbias.t627 Vbias.n5111 83.5719
R9839 Vbias.n5105 Vbias.n5104 83.5719
R9840 Vbias.n5104 Vbias.t411 83.5719
R9841 Vbias.n5117 Vbias.n2373 83.5719
R9842 Vbias.n2373 Vbias.t56 83.5719
R9843 Vbias.n5113 Vbias.n5112 83.5719
R9844 Vbias.n5112 Vbias.t627 83.5719
R9845 Vbias.n5103 Vbias.n5102 83.5719
R9846 Vbias.t411 Vbias.n5103 83.5719
R9847 Vbias.n5054 Vbias.n2418 83.5719
R9848 Vbias.n2418 Vbias.t241 83.5719
R9849 Vbias.n5050 Vbias.n5049 83.5719
R9850 Vbias.n5049 Vbias.t325 83.5719
R9851 Vbias.n2419 Vbias.n2417 83.5719
R9852 Vbias.n2417 Vbias.t241 83.5719
R9853 Vbias.n5048 Vbias.n5047 83.5719
R9854 Vbias.t325 Vbias.n5048 83.5719
R9855 Vbias.n5042 Vbias.n5041 83.5719
R9856 Vbias.n5041 Vbias.t828 83.5719
R9857 Vbias.n5040 Vbias.n5039 83.5719
R9858 Vbias.t828 Vbias.n5040 83.5719
R9859 Vbias.n4111 Vbias.n4110 83.5719
R9860 Vbias.n4110 Vbias.t573 83.5719
R9861 Vbias.n4109 Vbias.n4108 83.5719
R9862 Vbias.t573 Vbias.n4109 83.5719
R9863 Vbias.n4124 Vbias.n4003 83.5719
R9864 Vbias.t131 Vbias.n4003 83.5719
R9865 Vbias.n4099 Vbias.n3994 83.5719
R9866 Vbias.t286 Vbias.n3994 83.5719
R9867 Vbias.n4115 Vbias.n3986 83.5719
R9868 Vbias.t528 Vbias.n3986 83.5719
R9869 Vbias.n4122 Vbias.n4004 83.5719
R9870 Vbias.t131 Vbias.n4004 83.5719
R9871 Vbias.n4120 Vbias.n3995 83.5719
R9872 Vbias.t286 Vbias.n3995 83.5719
R9873 Vbias.n4118 Vbias.n3987 83.5719
R9874 Vbias.t528 Vbias.n3987 83.5719
R9875 Vbias.n4140 Vbias.n4029 83.5719
R9876 Vbias.t296 Vbias.n4029 83.5719
R9877 Vbias.n4087 Vbias.n4017 83.5719
R9878 Vbias.t163 Vbias.n4017 83.5719
R9879 Vbias.n4129 Vbias.n4128 83.5719
R9880 Vbias.n4129 Vbias.t82 83.5719
R9881 Vbias.n4138 Vbias.n4030 83.5719
R9882 Vbias.t296 Vbias.n4030 83.5719
R9883 Vbias.n4136 Vbias.n4018 83.5719
R9884 Vbias.t163 Vbias.n4018 83.5719
R9885 Vbias.n4134 Vbias.n4133 83.5719
R9886 Vbias.n4133 Vbias.t82 83.5719
R9887 Vbias.n4163 Vbias.n4045 83.5719
R9888 Vbias.t467 Vbias.n4045 83.5719
R9889 Vbias.n4149 Vbias.n4148 83.5719
R9890 Vbias.n4149 Vbias.t289 83.5719
R9891 Vbias.n4161 Vbias.n4046 83.5719
R9892 Vbias.t467 Vbias.n4046 83.5719
R9893 Vbias.n4159 Vbias.n4158 83.5719
R9894 Vbias.n4158 Vbias.t289 83.5719
R9895 Vbias.n4182 Vbias.n4071 83.5719
R9896 Vbias.t783 Vbias.n4071 83.5719
R9897 Vbias.n4179 Vbias.n4059 83.5719
R9898 Vbias.t10 Vbias.n4059 83.5719
R9899 Vbias.n4177 Vbias.n4176 83.5719
R9900 Vbias.n4176 Vbias.t36 83.5719
R9901 Vbias.n4185 Vbias.n4184 83.5719
R9902 Vbias.t783 Vbias.n4185 83.5719
R9903 Vbias.n4169 Vbias.n4060 83.5719
R9904 Vbias.t10 Vbias.n4060 83.5719
R9905 Vbias.n4172 Vbias.n4171 83.5719
R9906 Vbias.n4172 Vbias.t36 83.5719
R9907 Vbias.n4237 Vbias.n4236 83.5719
R9908 Vbias.t131 Vbias.n4237 83.5719
R9909 Vbias.n4244 Vbias.n4243 83.5719
R9910 Vbias.n4243 Vbias.t286 83.5719
R9911 Vbias.n4247 Vbias.n4246 83.5719
R9912 Vbias.t528 Vbias.n4247 83.5719
R9913 Vbias.n4239 Vbias.n4238 83.5719
R9914 Vbias.n4238 Vbias.t131 83.5719
R9915 Vbias.n4242 Vbias.n4241 83.5719
R9916 Vbias.t286 Vbias.n4242 83.5719
R9917 Vbias.n4249 Vbias.n4248 83.5719
R9918 Vbias.n4248 Vbias.t528 83.5719
R9919 Vbias.n4223 Vbias.n4222 83.5719
R9920 Vbias.n4222 Vbias.t296 83.5719
R9921 Vbias.n4226 Vbias.n4225 83.5719
R9922 Vbias.t163 Vbias.n4226 83.5719
R9923 Vbias.n4009 Vbias.n4007 83.5719
R9924 Vbias.n4007 Vbias.t82 83.5719
R9925 Vbias.n4221 Vbias.n4220 83.5719
R9926 Vbias.t296 Vbias.n4221 83.5719
R9927 Vbias.n4228 Vbias.n4227 83.5719
R9928 Vbias.n4227 Vbias.t163 83.5719
R9929 Vbias.n4231 Vbias.n4008 83.5719
R9930 Vbias.n4008 Vbias.t82 83.5719
R9931 Vbias.n4034 Vbias.n4032 83.5719
R9932 Vbias.n4032 Vbias.t503 83.5719
R9933 Vbias.n4215 Vbias.n4033 83.5719
R9934 Vbias.n4033 Vbias.t503 83.5719
R9935 Vbias.n4206 Vbias.n4205 83.5719
R9936 Vbias.t467 Vbias.n4206 83.5719
R9937 Vbias.n4153 Vbias.n4152 83.5719
R9938 Vbias.n4153 Vbias.t289 83.5719
R9939 Vbias.n4202 Vbias.n4040 83.5719
R9940 Vbias.t467 Vbias.n4202 83.5719
R9941 Vbias.n4211 Vbias.n4039 83.5719
R9942 Vbias.t289 Vbias.n4039 83.5719
R9943 Vbias.n4189 Vbias.n4188 83.5719
R9944 Vbias.n4188 Vbias.t783 83.5719
R9945 Vbias.n4192 Vbias.n4191 83.5719
R9946 Vbias.t10 Vbias.n4192 83.5719
R9947 Vbias.n4051 Vbias.n4049 83.5719
R9948 Vbias.n4049 Vbias.t36 83.5719
R9949 Vbias.n4187 Vbias.n4186 83.5719
R9950 Vbias.t783 Vbias.n4187 83.5719
R9951 Vbias.n4194 Vbias.n4193 83.5719
R9952 Vbias.n4193 Vbias.t10 83.5719
R9953 Vbias.n4197 Vbias.n4050 83.5719
R9954 Vbias.n4050 Vbias.t36 83.5719
R9955 Vbias.n3705 Vbias.n3704 83.5719
R9956 Vbias.n3704 Vbias.t835 83.5719
R9957 Vbias.n3703 Vbias.n3702 83.5719
R9958 Vbias.t835 Vbias.n3703 83.5719
R9959 Vbias.n3685 Vbias.n3472 83.5719
R9960 Vbias.t389 Vbias.n3472 83.5719
R9961 Vbias.n3693 Vbias.n3455 83.5719
R9962 Vbias.t575 Vbias.n3455 83.5719
R9963 Vbias.n3696 Vbias.n3450 83.5719
R9964 Vbias.n3450 Vbias.t170 83.5719
R9965 Vbias.n3681 Vbias.n3473 83.5719
R9966 Vbias.t389 Vbias.n3473 83.5719
R9967 Vbias.n3674 Vbias.n3460 83.5719
R9968 Vbias.t575 Vbias.n3460 83.5719
R9969 Vbias.n3672 Vbias.n3671 83.5719
R9970 Vbias.n3671 Vbias.t170 83.5719
R9971 Vbias.n3647 Vbias.n3501 83.5719
R9972 Vbias.t417 Vbias.n3501 83.5719
R9973 Vbias.n3655 Vbias.n3484 83.5719
R9974 Vbias.t624 Vbias.n3484 83.5719
R9975 Vbias.n3658 Vbias.n3479 83.5719
R9976 Vbias.n3479 Vbias.t462 83.5719
R9977 Vbias.n3643 Vbias.n3502 83.5719
R9978 Vbias.t417 Vbias.n3502 83.5719
R9979 Vbias.n3636 Vbias.n3489 83.5719
R9980 Vbias.t624 Vbias.n3489 83.5719
R9981 Vbias.n3634 Vbias.n3633 83.5719
R9982 Vbias.n3633 Vbias.t462 83.5719
R9983 Vbias.n3607 Vbias.n3519 83.5719
R9984 Vbias.t693 Vbias.n3519 83.5719
R9985 Vbias.n3617 Vbias.n3511 83.5719
R9986 Vbias.t148 Vbias.n3511 83.5719
R9987 Vbias.n3604 Vbias.n3520 83.5719
R9988 Vbias.t693 Vbias.n3520 83.5719
R9989 Vbias.n3602 Vbias.n3601 83.5719
R9990 Vbias.n3601 Vbias.t148 83.5719
R9991 Vbias.n3571 Vbias.n3548 83.5719
R9992 Vbias.t6 Vbias.n3548 83.5719
R9993 Vbias.n3579 Vbias.n3531 83.5719
R9994 Vbias.t684 Vbias.n3531 83.5719
R9995 Vbias.n3582 Vbias.n3526 83.5719
R9996 Vbias.n3526 Vbias.t609 83.5719
R9997 Vbias.n3567 Vbias.n3549 83.5719
R9998 Vbias.t6 Vbias.n3549 83.5719
R9999 Vbias.n3560 Vbias.n3536 83.5719
R10000 Vbias.t684 Vbias.n3536 83.5719
R10001 Vbias.n3558 Vbias.n3557 83.5719
R10002 Vbias.n3557 Vbias.t609 83.5719
R10003 Vbias.n3688 Vbias.n3687 83.5719
R10004 Vbias.n3687 Vbias.t389 83.5719
R10005 Vbias.n3691 Vbias.n3690 83.5719
R10006 Vbias.t575 Vbias.n3691 83.5719
R10007 Vbias.n3448 Vbias.n3446 83.5719
R10008 Vbias.n3446 Vbias.t170 83.5719
R10009 Vbias.n3686 Vbias.n3685 83.5719
R10010 Vbias.t389 Vbias.n3686 83.5719
R10011 Vbias.n3693 Vbias.n3692 83.5719
R10012 Vbias.n3692 Vbias.t575 83.5719
R10013 Vbias.n3696 Vbias.n3447 83.5719
R10014 Vbias.n3447 Vbias.t170 83.5719
R10015 Vbias.n3650 Vbias.n3649 83.5719
R10016 Vbias.n3649 Vbias.t417 83.5719
R10017 Vbias.n3653 Vbias.n3652 83.5719
R10018 Vbias.t624 Vbias.n3653 83.5719
R10019 Vbias.n3477 Vbias.n3475 83.5719
R10020 Vbias.n3475 Vbias.t462 83.5719
R10021 Vbias.n3648 Vbias.n3647 83.5719
R10022 Vbias.t417 Vbias.n3648 83.5719
R10023 Vbias.n3655 Vbias.n3654 83.5719
R10024 Vbias.n3654 Vbias.t624 83.5719
R10025 Vbias.n3658 Vbias.n3476 83.5719
R10026 Vbias.n3476 Vbias.t462 83.5719
R10027 Vbias.n3505 Vbias.n3503 83.5719
R10028 Vbias.n3503 Vbias.t809 83.5719
R10029 Vbias.n3621 Vbias.n3504 83.5719
R10030 Vbias.n3504 Vbias.t809 83.5719
R10031 Vbias.n3611 Vbias.n3610 83.5719
R10032 Vbias.t693 Vbias.n3611 83.5719
R10033 Vbias.n3595 Vbias.n3594 83.5719
R10034 Vbias.n3594 Vbias.t148 83.5719
R10035 Vbias.n3607 Vbias.n3588 83.5719
R10036 Vbias.t693 Vbias.n3588 83.5719
R10037 Vbias.n3617 Vbias.n3510 83.5719
R10038 Vbias.t148 Vbias.n3510 83.5719
R10039 Vbias.n3574 Vbias.n3573 83.5719
R10040 Vbias.n3573 Vbias.t6 83.5719
R10041 Vbias.n3577 Vbias.n3576 83.5719
R10042 Vbias.t684 Vbias.n3577 83.5719
R10043 Vbias.n3524 Vbias.n3522 83.5719
R10044 Vbias.n3522 Vbias.t609 83.5719
R10045 Vbias.n3572 Vbias.n3571 83.5719
R10046 Vbias.t6 Vbias.n3572 83.5719
R10047 Vbias.n3579 Vbias.n3578 83.5719
R10048 Vbias.n3578 Vbias.t684 83.5719
R10049 Vbias.n3582 Vbias.n3523 83.5719
R10050 Vbias.n3523 Vbias.t609 83.5719
R10051 Vbias.n3436 Vbias.n3435 83.5719
R10052 Vbias.n3435 Vbias.t877 83.5719
R10053 Vbias.n3434 Vbias.n3433 83.5719
R10054 Vbias.t877 Vbias.n3434 83.5719
R10055 Vbias.n3416 Vbias.n3203 83.5719
R10056 Vbias.t314 Vbias.n3203 83.5719
R10057 Vbias.n3424 Vbias.n3186 83.5719
R10058 Vbias.t653 Vbias.n3186 83.5719
R10059 Vbias.n3427 Vbias.n3181 83.5719
R10060 Vbias.n3181 Vbias.t550 83.5719
R10061 Vbias.n3412 Vbias.n3204 83.5719
R10062 Vbias.t314 Vbias.n3204 83.5719
R10063 Vbias.n3405 Vbias.n3191 83.5719
R10064 Vbias.t653 Vbias.n3191 83.5719
R10065 Vbias.n3403 Vbias.n3402 83.5719
R10066 Vbias.n3402 Vbias.t550 83.5719
R10067 Vbias.n3378 Vbias.n3232 83.5719
R10068 Vbias.t150 Vbias.n3232 83.5719
R10069 Vbias.n3386 Vbias.n3215 83.5719
R10070 Vbias.t692 Vbias.n3215 83.5719
R10071 Vbias.n3389 Vbias.n3210 83.5719
R10072 Vbias.n3210 Vbias.t374 83.5719
R10073 Vbias.n3374 Vbias.n3233 83.5719
R10074 Vbias.t150 Vbias.n3233 83.5719
R10075 Vbias.n3367 Vbias.n3220 83.5719
R10076 Vbias.t692 Vbias.n3220 83.5719
R10077 Vbias.n3365 Vbias.n3364 83.5719
R10078 Vbias.n3364 Vbias.t374 83.5719
R10079 Vbias.n3338 Vbias.n3250 83.5719
R10080 Vbias.t308 Vbias.n3250 83.5719
R10081 Vbias.n3348 Vbias.n3242 83.5719
R10082 Vbias.t583 Vbias.n3242 83.5719
R10083 Vbias.n3335 Vbias.n3251 83.5719
R10084 Vbias.t308 Vbias.n3251 83.5719
R10085 Vbias.n3333 Vbias.n3332 83.5719
R10086 Vbias.n3332 Vbias.t583 83.5719
R10087 Vbias.n3302 Vbias.n3279 83.5719
R10088 Vbias.t363 Vbias.n3279 83.5719
R10089 Vbias.n3310 Vbias.n3262 83.5719
R10090 Vbias.t514 Vbias.n3262 83.5719
R10091 Vbias.n3313 Vbias.n3257 83.5719
R10092 Vbias.n3257 Vbias.t881 83.5719
R10093 Vbias.n3298 Vbias.n3280 83.5719
R10094 Vbias.t363 Vbias.n3280 83.5719
R10095 Vbias.n3291 Vbias.n3267 83.5719
R10096 Vbias.t514 Vbias.n3267 83.5719
R10097 Vbias.n3289 Vbias.n3288 83.5719
R10098 Vbias.n3288 Vbias.t881 83.5719
R10099 Vbias.n3419 Vbias.n3418 83.5719
R10100 Vbias.n3418 Vbias.t314 83.5719
R10101 Vbias.n3422 Vbias.n3421 83.5719
R10102 Vbias.t653 Vbias.n3422 83.5719
R10103 Vbias.n3179 Vbias.n3177 83.5719
R10104 Vbias.n3177 Vbias.t550 83.5719
R10105 Vbias.n3417 Vbias.n3416 83.5719
R10106 Vbias.t314 Vbias.n3417 83.5719
R10107 Vbias.n3424 Vbias.n3423 83.5719
R10108 Vbias.n3423 Vbias.t653 83.5719
R10109 Vbias.n3427 Vbias.n3178 83.5719
R10110 Vbias.n3178 Vbias.t550 83.5719
R10111 Vbias.n3381 Vbias.n3380 83.5719
R10112 Vbias.n3380 Vbias.t150 83.5719
R10113 Vbias.n3384 Vbias.n3383 83.5719
R10114 Vbias.t692 Vbias.n3384 83.5719
R10115 Vbias.n3208 Vbias.n3206 83.5719
R10116 Vbias.n3206 Vbias.t374 83.5719
R10117 Vbias.n3379 Vbias.n3378 83.5719
R10118 Vbias.t150 Vbias.n3379 83.5719
R10119 Vbias.n3386 Vbias.n3385 83.5719
R10120 Vbias.n3385 Vbias.t692 83.5719
R10121 Vbias.n3389 Vbias.n3207 83.5719
R10122 Vbias.n3207 Vbias.t374 83.5719
R10123 Vbias.n3236 Vbias.n3234 83.5719
R10124 Vbias.n3234 Vbias.t387 83.5719
R10125 Vbias.n3352 Vbias.n3235 83.5719
R10126 Vbias.n3235 Vbias.t387 83.5719
R10127 Vbias.n3342 Vbias.n3341 83.5719
R10128 Vbias.t308 Vbias.n3342 83.5719
R10129 Vbias.n3326 Vbias.n3325 83.5719
R10130 Vbias.n3325 Vbias.t583 83.5719
R10131 Vbias.n3338 Vbias.n3319 83.5719
R10132 Vbias.t308 Vbias.n3319 83.5719
R10133 Vbias.n3348 Vbias.n3241 83.5719
R10134 Vbias.t583 Vbias.n3241 83.5719
R10135 Vbias.n3305 Vbias.n3304 83.5719
R10136 Vbias.n3304 Vbias.t363 83.5719
R10137 Vbias.n3308 Vbias.n3307 83.5719
R10138 Vbias.t514 Vbias.n3308 83.5719
R10139 Vbias.n3255 Vbias.n3253 83.5719
R10140 Vbias.n3253 Vbias.t881 83.5719
R10141 Vbias.n3303 Vbias.n3302 83.5719
R10142 Vbias.t363 Vbias.n3303 83.5719
R10143 Vbias.n3310 Vbias.n3309 83.5719
R10144 Vbias.n3309 Vbias.t514 83.5719
R10145 Vbias.n3313 Vbias.n3254 83.5719
R10146 Vbias.n3254 Vbias.t881 83.5719
R10147 Vbias.n3974 Vbias.n3973 83.5719
R10148 Vbias.n3973 Vbias.t651 83.5719
R10149 Vbias.n3972 Vbias.n3971 83.5719
R10150 Vbias.t651 Vbias.n3972 83.5719
R10151 Vbias.n3954 Vbias.n3741 83.5719
R10152 Vbias.t127 Vbias.n3741 83.5719
R10153 Vbias.n3962 Vbias.n3724 83.5719
R10154 Vbias.t310 Vbias.n3724 83.5719
R10155 Vbias.n3965 Vbias.n3719 83.5719
R10156 Vbias.n3719 Vbias.t458 83.5719
R10157 Vbias.n3950 Vbias.n3742 83.5719
R10158 Vbias.t127 Vbias.n3742 83.5719
R10159 Vbias.n3943 Vbias.n3729 83.5719
R10160 Vbias.t310 Vbias.n3729 83.5719
R10161 Vbias.n3941 Vbias.n3940 83.5719
R10162 Vbias.n3940 Vbias.t458 83.5719
R10163 Vbias.n3916 Vbias.n3770 83.5719
R10164 Vbias.t435 Vbias.n3770 83.5719
R10165 Vbias.n3924 Vbias.n3753 83.5719
R10166 Vbias.t696 Vbias.n3753 83.5719
R10167 Vbias.n3927 Vbias.n3748 83.5719
R10168 Vbias.n3748 Vbias.t351 83.5719
R10169 Vbias.n3912 Vbias.n3771 83.5719
R10170 Vbias.t435 Vbias.n3771 83.5719
R10171 Vbias.n3905 Vbias.n3758 83.5719
R10172 Vbias.t696 Vbias.n3758 83.5719
R10173 Vbias.n3903 Vbias.n3902 83.5719
R10174 Vbias.n3902 Vbias.t351 83.5719
R10175 Vbias.n3876 Vbias.n3788 83.5719
R10176 Vbias.t545 Vbias.n3788 83.5719
R10177 Vbias.n3886 Vbias.n3780 83.5719
R10178 Vbias.t124 Vbias.n3780 83.5719
R10179 Vbias.n3873 Vbias.n3789 83.5719
R10180 Vbias.t545 Vbias.n3789 83.5719
R10181 Vbias.n3871 Vbias.n3870 83.5719
R10182 Vbias.n3870 Vbias.t124 83.5719
R10183 Vbias.n3840 Vbias.n3817 83.5719
R10184 Vbias.t438 Vbias.n3817 83.5719
R10185 Vbias.n3848 Vbias.n3800 83.5719
R10186 Vbias.t620 Vbias.n3800 83.5719
R10187 Vbias.n3851 Vbias.n3795 83.5719
R10188 Vbias.n3795 Vbias.t524 83.5719
R10189 Vbias.n3836 Vbias.n3818 83.5719
R10190 Vbias.t438 Vbias.n3818 83.5719
R10191 Vbias.n3829 Vbias.n3805 83.5719
R10192 Vbias.t620 Vbias.n3805 83.5719
R10193 Vbias.n3827 Vbias.n3826 83.5719
R10194 Vbias.n3826 Vbias.t524 83.5719
R10195 Vbias.n3957 Vbias.n3956 83.5719
R10196 Vbias.n3956 Vbias.t127 83.5719
R10197 Vbias.n3960 Vbias.n3959 83.5719
R10198 Vbias.t310 Vbias.n3960 83.5719
R10199 Vbias.n3717 Vbias.n3715 83.5719
R10200 Vbias.n3715 Vbias.t458 83.5719
R10201 Vbias.n3955 Vbias.n3954 83.5719
R10202 Vbias.t127 Vbias.n3955 83.5719
R10203 Vbias.n3962 Vbias.n3961 83.5719
R10204 Vbias.n3961 Vbias.t310 83.5719
R10205 Vbias.n3965 Vbias.n3716 83.5719
R10206 Vbias.n3716 Vbias.t458 83.5719
R10207 Vbias.n3919 Vbias.n3918 83.5719
R10208 Vbias.n3918 Vbias.t435 83.5719
R10209 Vbias.n3922 Vbias.n3921 83.5719
R10210 Vbias.t696 Vbias.n3922 83.5719
R10211 Vbias.n3746 Vbias.n3744 83.5719
R10212 Vbias.n3744 Vbias.t351 83.5719
R10213 Vbias.n3917 Vbias.n3916 83.5719
R10214 Vbias.t435 Vbias.n3917 83.5719
R10215 Vbias.n3924 Vbias.n3923 83.5719
R10216 Vbias.n3923 Vbias.t696 83.5719
R10217 Vbias.n3927 Vbias.n3745 83.5719
R10218 Vbias.n3745 Vbias.t351 83.5719
R10219 Vbias.n3774 Vbias.n3772 83.5719
R10220 Vbias.n3772 Vbias.t450 83.5719
R10221 Vbias.n3890 Vbias.n3773 83.5719
R10222 Vbias.n3773 Vbias.t450 83.5719
R10223 Vbias.n3880 Vbias.n3879 83.5719
R10224 Vbias.t545 Vbias.n3880 83.5719
R10225 Vbias.n3864 Vbias.n3863 83.5719
R10226 Vbias.n3863 Vbias.t124 83.5719
R10227 Vbias.n3876 Vbias.n3857 83.5719
R10228 Vbias.t545 Vbias.n3857 83.5719
R10229 Vbias.n3886 Vbias.n3779 83.5719
R10230 Vbias.t124 Vbias.n3779 83.5719
R10231 Vbias.n3843 Vbias.n3842 83.5719
R10232 Vbias.n3842 Vbias.t438 83.5719
R10233 Vbias.n3846 Vbias.n3845 83.5719
R10234 Vbias.t620 Vbias.n3846 83.5719
R10235 Vbias.n3793 Vbias.n3791 83.5719
R10236 Vbias.n3791 Vbias.t524 83.5719
R10237 Vbias.n3841 Vbias.n3840 83.5719
R10238 Vbias.t438 Vbias.n3841 83.5719
R10239 Vbias.n3848 Vbias.n3847 83.5719
R10240 Vbias.n3847 Vbias.t620 83.5719
R10241 Vbias.n3851 Vbias.n3792 83.5719
R10242 Vbias.n3792 Vbias.t524 83.5719
R10243 Vbias.n3166 Vbias.n3165 83.5719
R10244 Vbias.n3165 Vbias.t833 83.5719
R10245 Vbias.n3164 Vbias.n3163 83.5719
R10246 Vbias.t833 Vbias.n3164 83.5719
R10247 Vbias.n3146 Vbias.n2933 83.5719
R10248 Vbias.t639 Vbias.n2933 83.5719
R10249 Vbias.n3154 Vbias.n2916 83.5719
R10250 Vbias.t365 Vbias.n2916 83.5719
R10251 Vbias.n3157 Vbias.n2911 83.5719
R10252 Vbias.n2911 Vbias.t137 83.5719
R10253 Vbias.n3142 Vbias.n2934 83.5719
R10254 Vbias.t639 Vbias.n2934 83.5719
R10255 Vbias.n3135 Vbias.n2921 83.5719
R10256 Vbias.t365 Vbias.n2921 83.5719
R10257 Vbias.n3133 Vbias.n3132 83.5719
R10258 Vbias.n3132 Vbias.t137 83.5719
R10259 Vbias.n3108 Vbias.n2962 83.5719
R10260 Vbias.t130 Vbias.n2962 83.5719
R10261 Vbias.n3116 Vbias.n2945 83.5719
R10262 Vbias.t147 Vbias.n2945 83.5719
R10263 Vbias.n3119 Vbias.n2940 83.5719
R10264 Vbias.n2940 Vbias.t726 83.5719
R10265 Vbias.n3104 Vbias.n2963 83.5719
R10266 Vbias.t130 Vbias.n2963 83.5719
R10267 Vbias.n3097 Vbias.n2950 83.5719
R10268 Vbias.t147 Vbias.n2950 83.5719
R10269 Vbias.n3095 Vbias.n3094 83.5719
R10270 Vbias.n3094 Vbias.t726 83.5719
R10271 Vbias.n3068 Vbias.n2980 83.5719
R10272 Vbias.t311 Vbias.n2980 83.5719
R10273 Vbias.n3078 Vbias.n2972 83.5719
R10274 Vbias.t280 Vbias.n2972 83.5719
R10275 Vbias.n3065 Vbias.n2981 83.5719
R10276 Vbias.t311 Vbias.n2981 83.5719
R10277 Vbias.n3063 Vbias.n3062 83.5719
R10278 Vbias.n3062 Vbias.t280 83.5719
R10279 Vbias.n3032 Vbias.n3009 83.5719
R10280 Vbias.t775 Vbias.n3009 83.5719
R10281 Vbias.n3040 Vbias.n2992 83.5719
R10282 Vbias.t362 Vbias.n2992 83.5719
R10283 Vbias.n3043 Vbias.n2987 83.5719
R10284 Vbias.n2987 Vbias.t165 83.5719
R10285 Vbias.n3028 Vbias.n3010 83.5719
R10286 Vbias.t775 Vbias.n3010 83.5719
R10287 Vbias.n3021 Vbias.n2997 83.5719
R10288 Vbias.t362 Vbias.n2997 83.5719
R10289 Vbias.n3019 Vbias.n3018 83.5719
R10290 Vbias.n3018 Vbias.t165 83.5719
R10291 Vbias.n3149 Vbias.n3148 83.5719
R10292 Vbias.n3148 Vbias.t639 83.5719
R10293 Vbias.n3152 Vbias.n3151 83.5719
R10294 Vbias.t365 Vbias.n3152 83.5719
R10295 Vbias.n2909 Vbias.n2907 83.5719
R10296 Vbias.n2907 Vbias.t137 83.5719
R10297 Vbias.n3147 Vbias.n3146 83.5719
R10298 Vbias.t639 Vbias.n3147 83.5719
R10299 Vbias.n3154 Vbias.n3153 83.5719
R10300 Vbias.n3153 Vbias.t365 83.5719
R10301 Vbias.n3157 Vbias.n2908 83.5719
R10302 Vbias.n2908 Vbias.t137 83.5719
R10303 Vbias.n3111 Vbias.n3110 83.5719
R10304 Vbias.n3110 Vbias.t130 83.5719
R10305 Vbias.n3114 Vbias.n3113 83.5719
R10306 Vbias.t147 Vbias.n3114 83.5719
R10307 Vbias.n2938 Vbias.n2936 83.5719
R10308 Vbias.n2936 Vbias.t726 83.5719
R10309 Vbias.n3109 Vbias.n3108 83.5719
R10310 Vbias.t130 Vbias.n3109 83.5719
R10311 Vbias.n3116 Vbias.n3115 83.5719
R10312 Vbias.n3115 Vbias.t147 83.5719
R10313 Vbias.n3119 Vbias.n2937 83.5719
R10314 Vbias.n2937 Vbias.t726 83.5719
R10315 Vbias.n2966 Vbias.n2964 83.5719
R10316 Vbias.n2964 Vbias.t871 83.5719
R10317 Vbias.n3082 Vbias.n2965 83.5719
R10318 Vbias.n2965 Vbias.t871 83.5719
R10319 Vbias.n3072 Vbias.n3071 83.5719
R10320 Vbias.t311 Vbias.n3072 83.5719
R10321 Vbias.n3056 Vbias.n3055 83.5719
R10322 Vbias.n3055 Vbias.t280 83.5719
R10323 Vbias.n3068 Vbias.n3049 83.5719
R10324 Vbias.t311 Vbias.n3049 83.5719
R10325 Vbias.n3078 Vbias.n2971 83.5719
R10326 Vbias.t280 Vbias.n2971 83.5719
R10327 Vbias.n3035 Vbias.n3034 83.5719
R10328 Vbias.n3034 Vbias.t775 83.5719
R10329 Vbias.n3038 Vbias.n3037 83.5719
R10330 Vbias.t362 Vbias.n3038 83.5719
R10331 Vbias.n2985 Vbias.n2983 83.5719
R10332 Vbias.n2983 Vbias.t165 83.5719
R10333 Vbias.n3033 Vbias.n3032 83.5719
R10334 Vbias.t775 Vbias.n3033 83.5719
R10335 Vbias.n3040 Vbias.n3039 83.5719
R10336 Vbias.n3039 Vbias.t362 83.5719
R10337 Vbias.n3043 Vbias.n2984 83.5719
R10338 Vbias.n2984 Vbias.t165 83.5719
R10339 Vbias.n2666 Vbias.n2664 83.5719
R10340 Vbias.n2664 Vbias.t875 83.5719
R10341 Vbias.n4841 Vbias.n2665 83.5719
R10342 Vbias.n2665 Vbias.t875 83.5719
R10343 Vbias.n4822 Vbias.n2694 83.5719
R10344 Vbias.t448 Vbias.n2694 83.5719
R10345 Vbias.n4830 Vbias.n2677 83.5719
R10346 Vbias.t400 Vbias.n2677 83.5719
R10347 Vbias.n4833 Vbias.n2672 83.5719
R10348 Vbias.n2672 Vbias.t227 83.5719
R10349 Vbias.n4818 Vbias.n2695 83.5719
R10350 Vbias.t448 Vbias.n2695 83.5719
R10351 Vbias.n4811 Vbias.n2682 83.5719
R10352 Vbias.t400 Vbias.n2682 83.5719
R10353 Vbias.n4809 Vbias.n4808 83.5719
R10354 Vbias.n4808 Vbias.t227 83.5719
R10355 Vbias.n4784 Vbias.n2723 83.5719
R10356 Vbias.t282 Vbias.n2723 83.5719
R10357 Vbias.n4792 Vbias.n2706 83.5719
R10358 Vbias.t626 Vbias.n2706 83.5719
R10359 Vbias.n4795 Vbias.n2701 83.5719
R10360 Vbias.n2701 Vbias.t133 83.5719
R10361 Vbias.n4780 Vbias.n2724 83.5719
R10362 Vbias.t282 Vbias.n2724 83.5719
R10363 Vbias.n4773 Vbias.n2711 83.5719
R10364 Vbias.t626 Vbias.n2711 83.5719
R10365 Vbias.n4771 Vbias.n4770 83.5719
R10366 Vbias.n4770 Vbias.t133 83.5719
R10367 Vbias.n4744 Vbias.n2741 83.5719
R10368 Vbias.t312 Vbias.n2741 83.5719
R10369 Vbias.n4754 Vbias.n2733 83.5719
R10370 Vbias.t348 Vbias.n2733 83.5719
R10371 Vbias.n4741 Vbias.n2742 83.5719
R10372 Vbias.t312 Vbias.n2742 83.5719
R10373 Vbias.n4739 Vbias.n4738 83.5719
R10374 Vbias.n4738 Vbias.t348 83.5719
R10375 Vbias.n4708 Vbias.n2770 83.5719
R10376 Vbias.t297 Vbias.n2770 83.5719
R10377 Vbias.n4716 Vbias.n2753 83.5719
R10378 Vbias.t304 Vbias.n2753 83.5719
R10379 Vbias.n4719 Vbias.n2748 83.5719
R10380 Vbias.n2748 Vbias.t460 83.5719
R10381 Vbias.n4704 Vbias.n2771 83.5719
R10382 Vbias.t297 Vbias.n2771 83.5719
R10383 Vbias.n4697 Vbias.n2758 83.5719
R10384 Vbias.t304 Vbias.n2758 83.5719
R10385 Vbias.n4695 Vbias.n4694 83.5719
R10386 Vbias.n4694 Vbias.t460 83.5719
R10387 Vbias.n4825 Vbias.n4824 83.5719
R10388 Vbias.n4824 Vbias.t448 83.5719
R10389 Vbias.n4828 Vbias.n4827 83.5719
R10390 Vbias.t400 Vbias.n4828 83.5719
R10391 Vbias.n2670 Vbias.n2668 83.5719
R10392 Vbias.n2668 Vbias.t227 83.5719
R10393 Vbias.n4823 Vbias.n4822 83.5719
R10394 Vbias.t448 Vbias.n4823 83.5719
R10395 Vbias.n4830 Vbias.n4829 83.5719
R10396 Vbias.n4829 Vbias.t400 83.5719
R10397 Vbias.n4833 Vbias.n2669 83.5719
R10398 Vbias.n2669 Vbias.t227 83.5719
R10399 Vbias.n4787 Vbias.n4786 83.5719
R10400 Vbias.n4786 Vbias.t282 83.5719
R10401 Vbias.n4790 Vbias.n4789 83.5719
R10402 Vbias.t626 Vbias.n4790 83.5719
R10403 Vbias.n2699 Vbias.n2697 83.5719
R10404 Vbias.n2697 Vbias.t133 83.5719
R10405 Vbias.n4785 Vbias.n4784 83.5719
R10406 Vbias.t282 Vbias.n4785 83.5719
R10407 Vbias.n4792 Vbias.n4791 83.5719
R10408 Vbias.n4791 Vbias.t626 83.5719
R10409 Vbias.n4795 Vbias.n2698 83.5719
R10410 Vbias.n2698 Vbias.t133 83.5719
R10411 Vbias.n2727 Vbias.n2725 83.5719
R10412 Vbias.n2725 Vbias.t446 83.5719
R10413 Vbias.n4758 Vbias.n2726 83.5719
R10414 Vbias.n2726 Vbias.t446 83.5719
R10415 Vbias.n4748 Vbias.n4747 83.5719
R10416 Vbias.t312 Vbias.n4748 83.5719
R10417 Vbias.n4732 Vbias.n4731 83.5719
R10418 Vbias.n4731 Vbias.t348 83.5719
R10419 Vbias.n4744 Vbias.n4725 83.5719
R10420 Vbias.t312 Vbias.n4725 83.5719
R10421 Vbias.n4754 Vbias.n2732 83.5719
R10422 Vbias.t348 Vbias.n2732 83.5719
R10423 Vbias.n4711 Vbias.n4710 83.5719
R10424 Vbias.n4710 Vbias.t297 83.5719
R10425 Vbias.n4714 Vbias.n4713 83.5719
R10426 Vbias.t304 Vbias.n4714 83.5719
R10427 Vbias.n2746 Vbias.n2744 83.5719
R10428 Vbias.n2744 Vbias.t460 83.5719
R10429 Vbias.n4709 Vbias.n4708 83.5719
R10430 Vbias.t297 Vbias.n4709 83.5719
R10431 Vbias.n4716 Vbias.n4715 83.5719
R10432 Vbias.n4715 Vbias.t304 83.5719
R10433 Vbias.n4719 Vbias.n2745 83.5719
R10434 Vbias.n2745 Vbias.t460 83.5719
R10435 Vbias.n2662 Vbias.n2660 83.5719
R10436 Vbias.n2660 Vbias.t839 83.5719
R10437 Vbias.n4907 Vbias.n2661 83.5719
R10438 Vbias.n2661 Vbias.t839 83.5719
R10439 Vbias.n2648 Vbias.n2646 83.5719
R10440 Vbias.n2646 Vbias.t445 83.5719
R10441 Vbias.n4924 Vbias.n4923 83.5719
R10442 Vbias.t577 Vbias.n4924 83.5719
R10443 Vbias.n4919 Vbias.n4918 83.5719
R10444 Vbias.n4918 Vbias.t526 83.5719
R10445 Vbias.n4929 Vbias.n2647 83.5719
R10446 Vbias.n2647 Vbias.t445 83.5719
R10447 Vbias.n2654 Vbias.n2649 83.5719
R10448 Vbias.t577 Vbias.n2654 83.5719
R10449 Vbias.n4917 Vbias.n4916 83.5719
R10450 Vbias.t526 Vbias.n4917 83.5719
R10451 Vbias.n2634 Vbias.n2632 83.5719
R10452 Vbias.n2632 Vbias.t517 83.5719
R10453 Vbias.n4947 Vbias.n4946 83.5719
R10454 Vbias.t632 Vbias.n4947 83.5719
R10455 Vbias.n4941 Vbias.n4940 83.5719
R10456 Vbias.n4940 Vbias.t831 83.5719
R10457 Vbias.n4952 Vbias.n2633 83.5719
R10458 Vbias.n2633 Vbias.t517 83.5719
R10459 Vbias.n2640 Vbias.n2635 83.5719
R10460 Vbias.t632 Vbias.n2640 83.5719
R10461 Vbias.n4939 Vbias.n4938 83.5719
R10462 Vbias.t831 Vbias.n4939 83.5719
R10463 Vbias.n4967 Vbias.n4966 83.5719
R10464 Vbias.n4966 Vbias.t650 83.5719
R10465 Vbias.n4958 Vbias.n4957 83.5719
R10466 Vbias.t424 Vbias.n4958 83.5719
R10467 Vbias.n4965 Vbias.n4964 83.5719
R10468 Vbias.t650 Vbias.n4965 83.5719
R10469 Vbias.n4960 Vbias.n4959 83.5719
R10470 Vbias.n4959 Vbias.t424 83.5719
R10471 Vbias.n4985 Vbias.n4984 83.5719
R10472 Vbias.n4984 Vbias.t283 83.5719
R10473 Vbias.n4976 Vbias.n4975 83.5719
R10474 Vbias.t164 Vbias.n4976 83.5719
R10475 Vbias.n4971 Vbias.n2617 83.5719
R10476 Vbias.t826 Vbias.n2617 83.5719
R10477 Vbias.n4983 Vbias.n4982 83.5719
R10478 Vbias.t283 Vbias.n4983 83.5719
R10479 Vbias.n4978 Vbias.n4977 83.5719
R10480 Vbias.n4977 Vbias.t164 83.5719
R10481 Vbias.n2625 Vbias.n2624 83.5719
R10482 Vbias.n2625 Vbias.t826 83.5719
R10483 Vbias.n4539 Vbias.n4538 83.5719
R10484 Vbias.n4538 Vbias.t110 83.5719
R10485 Vbias.n4543 Vbias.n4542 83.5719
R10486 Vbias.t303 Vbias.n4543 83.5719
R10487 Vbias.n4409 Vbias.n4407 83.5719
R10488 Vbias.n4407 Vbias.t536 83.5719
R10489 Vbias.n4537 Vbias.n4536 83.5719
R10490 Vbias.t110 Vbias.n4537 83.5719
R10491 Vbias.n4545 Vbias.n4544 83.5719
R10492 Vbias.n4544 Vbias.t303 83.5719
R10493 Vbias.n4547 Vbias.n4408 83.5719
R10494 Vbias.n4408 Vbias.t536 83.5719
R10495 Vbias.n4527 Vbias.n4526 83.5719
R10496 Vbias.t300 Vbias.n4527 83.5719
R10497 Vbias.n4428 Vbias.n4426 83.5719
R10498 Vbias.n4426 Vbias.t804 83.5719
R10499 Vbias.n4529 Vbias.n4528 83.5719
R10500 Vbias.n4528 Vbias.t300 83.5719
R10501 Vbias.n4531 Vbias.n4427 83.5719
R10502 Vbias.n4427 Vbias.t804 83.5719
R10503 Vbias.n4513 Vbias.n4512 83.5719
R10504 Vbias.t58 Vbias.n4513 83.5719
R10505 Vbias.n4520 Vbias.n4519 83.5719
R10506 Vbias.n4519 Vbias.t474 83.5719
R10507 Vbias.n4522 Vbias.n4441 83.5719
R10508 Vbias.t454 Vbias.n4441 83.5719
R10509 Vbias.n4515 Vbias.n4514 83.5719
R10510 Vbias.n4514 Vbias.t58 83.5719
R10511 Vbias.n4518 Vbias.n4517 83.5719
R10512 Vbias.t474 Vbias.n4518 83.5719
R10513 Vbias.n4454 Vbias.n4453 83.5719
R10514 Vbias.n4453 Vbias.t454 83.5719
R10515 Vbias.n4499 Vbias.n4498 83.5719
R10516 Vbias.t180 Vbias.n4499 83.5719
R10517 Vbias.n4506 Vbias.n4505 83.5719
R10518 Vbias.n4505 Vbias.t226 83.5719
R10519 Vbias.n4508 Vbias.n4463 83.5719
R10520 Vbias.t408 Vbias.n4463 83.5719
R10521 Vbias.n4501 Vbias.n4500 83.5719
R10522 Vbias.n4500 Vbias.t180 83.5719
R10523 Vbias.n4504 Vbias.n4503 83.5719
R10524 Vbias.t226 Vbias.n4504 83.5719
R10525 Vbias.n4476 Vbias.n4475 83.5719
R10526 Vbias.n4475 Vbias.t408 83.5719
R10527 Vbias.n4494 Vbias.n4486 83.5719
R10528 Vbias.t824 Vbias.n4486 83.5719
R10529 Vbias.n4488 Vbias.n4487 83.5719
R10530 Vbias.t824 Vbias.n4488 83.5719
R10531 Vbias.n4582 Vbias.n4581 83.5719
R10532 Vbias.t452 Vbias.n4582 83.5719
R10533 Vbias.n4576 Vbias.n4574 83.5719
R10534 Vbias.n4574 Vbias.t679 83.5719
R10535 Vbias.n4664 Vbias.n4580 83.5719
R10536 Vbias.t452 Vbias.n4580 83.5719
R10537 Vbias.n4667 Vbias.n4575 83.5719
R10538 Vbias.n4575 Vbias.t679 83.5719
R10539 Vbias.n4591 Vbias.n4589 83.5719
R10540 Vbias.n4589 Vbias.t334 83.5719
R10541 Vbias.n4657 Vbias.n4590 83.5719
R10542 Vbias.n4590 Vbias.t334 83.5719
R10543 Vbias.n4630 Vbias.n4629 83.5719
R10544 Vbias.n4630 Vbias.t214 83.5719
R10545 Vbias.n4627 Vbias.n4626 83.5719
R10546 Vbias.n4626 Vbias.t716 83.5719
R10547 Vbias.n4621 Vbias.n4620 83.5719
R10548 Vbias.n4621 Vbias.t285 83.5719
R10549 Vbias.n4649 Vbias.n4599 83.5719
R10550 Vbias.t214 Vbias.n4599 83.5719
R10551 Vbias.n4651 Vbias.n4597 83.5719
R10552 Vbias.t716 Vbias.n4597 83.5719
R10553 Vbias.n4653 Vbias.n4595 83.5719
R10554 Vbias.n4595 Vbias.t285 83.5719
R10555 Vbias.n2436 Vbias.n2434 83.5719
R10556 Vbias.n2434 Vbias.t42 83.5719
R10557 Vbias.n4641 Vbias.n4640 83.5719
R10558 Vbias.t439 Vbias.n4641 83.5719
R10559 Vbias.n4635 Vbias.n4634 83.5719
R10560 Vbias.n4634 Vbias.t861 83.5719
R10561 Vbias.n5033 Vbias.n2435 83.5719
R10562 Vbias.n2435 Vbias.t42 83.5719
R10563 Vbias.n4643 Vbias.n4642 83.5719
R10564 Vbias.n4642 Vbias.t439 83.5719
R10565 Vbias.n4645 Vbias.n4602 83.5719
R10566 Vbias.t861 Vbias.n4602 83.5719
R10567 Vbias.n4674 Vbias.n4558 83.5719
R10568 Vbias.t269 Vbias.n4558 83.5719
R10569 Vbias.n4676 Vbias.n4556 83.5719
R10570 Vbias.t513 Vbias.n4556 83.5719
R10571 Vbias.n4560 Vbias.n4559 83.5719
R10572 Vbias.t269 Vbias.n4560 83.5719
R10573 Vbias.n4569 Vbias.n4568 83.5719
R10574 Vbias.n4569 Vbias.t513 83.5719
R10575 Vbias.n4553 Vbias.n4551 83.5719
R10576 Vbias.n4551 Vbias.t789 83.5719
R10577 Vbias.n4678 Vbias.n4552 83.5719
R10578 Vbias.n4552 Vbias.t789 83.5719
R10579 Vbias.n7452 Vbias.n7451 83.5719
R10580 Vbias.t393 Vbias.n7452 83.5719
R10581 Vbias.n7459 Vbias.n7458 83.5719
R10582 Vbias.n7458 Vbias.t873 83.5719
R10583 Vbias.n7462 Vbias.n7461 83.5719
R10584 Vbias.t64 Vbias.n7462 83.5719
R10585 Vbias.n7454 Vbias.n7453 83.5719
R10586 Vbias.n7453 Vbias.t393 83.5719
R10587 Vbias.n7457 Vbias.n7456 83.5719
R10588 Vbias.t873 Vbias.n7457 83.5719
R10589 Vbias.n7464 Vbias.n7463 83.5719
R10590 Vbias.n7463 Vbias.t64 83.5719
R10591 Vbias.n7438 Vbias.n7437 83.5719
R10592 Vbias.n7437 Vbias.t302 83.5719
R10593 Vbias.n7441 Vbias.n7440 83.5719
R10594 Vbias.t146 Vbias.n7441 83.5719
R10595 Vbias.n7344 Vbias.n7342 83.5719
R10596 Vbias.n7342 Vbias.t192 83.5719
R10597 Vbias.n7436 Vbias.n7435 83.5719
R10598 Vbias.t302 Vbias.n7436 83.5719
R10599 Vbias.n7443 Vbias.n7442 83.5719
R10600 Vbias.n7442 Vbias.t146 83.5719
R10601 Vbias.n7446 Vbias.n7343 83.5719
R10602 Vbias.n7343 Vbias.t192 83.5719
R10603 Vbias.n7364 Vbias.n7362 83.5719
R10604 Vbias.n7362 Vbias.t588 83.5719
R10605 Vbias.n7430 Vbias.n7363 83.5719
R10606 Vbias.n7363 Vbias.t588 83.5719
R10607 Vbias.n7421 Vbias.n7420 83.5719
R10608 Vbias.t581 Vbias.n7421 83.5719
R10609 Vbias.n7379 Vbias.n7378 83.5719
R10610 Vbias.t667 Vbias.n7379 83.5719
R10611 Vbias.n7417 Vbias.n7370 83.5719
R10612 Vbias.t581 Vbias.n7417 83.5719
R10613 Vbias.n7426 Vbias.n7369 83.5719
R10614 Vbias.t667 Vbias.n7369 83.5719
R10615 Vbias.n7404 Vbias.n7403 83.5719
R10616 Vbias.n7403 Vbias.t299 83.5719
R10617 Vbias.n7407 Vbias.n7406 83.5719
R10618 Vbias.t705 Vbias.n7407 83.5719
R10619 Vbias.n7382 Vbias.n7380 83.5719
R10620 Vbias.n7380 Vbias.t251 83.5719
R10621 Vbias.n7401 Vbias.n7400 83.5719
R10622 Vbias.n7409 Vbias.n7408 83.5719
R10623 Vbias.n7408 Vbias.t705 83.5719
R10624 Vbias.n7412 Vbias.n7381 83.5719
R10625 Vbias.n7381 Vbias.t251 83.5719
R10626 Vbias.n6494 Vbias.n6493 83.5719
R10627 Vbias.t326 Vbias.n6494 83.5719
R10628 Vbias.n6499 Vbias.n6498 83.5719
R10629 Vbias.n6498 Vbias.t578 83.5719
R10630 Vbias.n6502 Vbias.n6501 83.5719
R10631 Vbias.n6502 Vbias.t120 83.5719
R10632 Vbias.n7582 Vbias.n865 83.5719
R10633 Vbias.t326 Vbias.n865 83.5719
R10634 Vbias.n7584 Vbias.n863 83.5719
R10635 Vbias.t578 Vbias.n863 83.5719
R10636 Vbias.n7586 Vbias.n861 83.5719
R10637 Vbias.t120 Vbias.n861 83.5719
R10638 Vbias.n6480 Vbias.n6479 83.5719
R10639 Vbias.t570 Vbias.n6480 83.5719
R10640 Vbias.n6485 Vbias.n6484 83.5719
R10641 Vbias.n6484 Vbias.t476 83.5719
R10642 Vbias.n6488 Vbias.n6487 83.5719
R10643 Vbias.n6488 Vbias.t249 83.5719
R10644 Vbias.n7574 Vbias.n873 83.5719
R10645 Vbias.t570 Vbias.n873 83.5719
R10646 Vbias.n7576 Vbias.n871 83.5719
R10647 Vbias.t476 Vbias.n871 83.5719
R10648 Vbias.n7578 Vbias.n869 83.5719
R10649 Vbias.t249 Vbias.n869 83.5719
R10650 Vbias.n878 Vbias.n877 83.5719
R10651 Vbias.t337 Vbias.n878 83.5719
R10652 Vbias.n7570 Vbias.n876 83.5719
R10653 Vbias.t337 Vbias.n876 83.5719
R10654 Vbias.n886 Vbias.n885 83.5719
R10655 Vbias.t391 Vbias.n886 83.5719
R10656 Vbias.n881 Vbias.n879 83.5719
R10657 Vbias.n879 Vbias.t807 83.5719
R10658 Vbias.n7560 Vbias.n884 83.5719
R10659 Vbias.t391 Vbias.n884 83.5719
R10660 Vbias.n7563 Vbias.n880 83.5719
R10661 Vbias.n880 Vbias.t807 83.5719
R10662 Vbias.n903 Vbias.n902 83.5719
R10663 Vbias.t582 Vbias.n903 83.5719
R10664 Vbias.n912 Vbias.n911 83.5719
R10665 Vbias.n912 Vbias.t506 83.5719
R10666 Vbias.n895 Vbias.n893 83.5719
R10667 Vbias.n893 Vbias.t204 83.5719
R10668 Vbias.n7548 Vbias.n901 83.5719
R10669 Vbias.t582 Vbias.n901 83.5719
R10670 Vbias.n7550 Vbias.n899 83.5719
R10671 Vbias.t506 Vbias.n899 83.5719
R10672 Vbias.n7553 Vbias.n894 83.5719
R10673 Vbias.n894 Vbias.t204 83.5719
R10674 Vbias.n6403 Vbias.n6402 83.5719
R10675 Vbias.n6403 Vbias.t442 83.5719
R10676 Vbias.n6400 Vbias.n6399 83.5719
R10677 Vbias.n6399 Vbias.t654 83.5719
R10678 Vbias.n6392 Vbias.n6391 83.5719
R10679 Vbias.t88 Vbias.n6392 83.5719
R10680 Vbias.n6569 Vbias.n6370 83.5719
R10681 Vbias.t442 Vbias.n6370 83.5719
R10682 Vbias.n6571 Vbias.n6368 83.5719
R10683 Vbias.t654 Vbias.n6368 83.5719
R10684 Vbias.n6573 Vbias.n6366 83.5719
R10685 Vbias.t88 Vbias.n6366 83.5719
R10686 Vbias.n6420 Vbias.n6419 83.5719
R10687 Vbias.n6420 Vbias.t555 83.5719
R10688 Vbias.n6417 Vbias.n6416 83.5719
R10689 Vbias.n6416 Vbias.t800 83.5719
R10690 Vbias.n6409 Vbias.n6408 83.5719
R10691 Vbias.t277 Vbias.n6409 83.5719
R10692 Vbias.n6561 Vbias.n6378 83.5719
R10693 Vbias.t555 Vbias.n6378 83.5719
R10694 Vbias.n6563 Vbias.n6376 83.5719
R10695 Vbias.t800 Vbias.n6376 83.5719
R10696 Vbias.n6565 Vbias.n6374 83.5719
R10697 Vbias.t277 Vbias.n6374 83.5719
R10698 Vbias.n6383 Vbias.n6382 83.5719
R10699 Vbias.t483 Vbias.n6383 83.5719
R10700 Vbias.n6557 Vbias.n6381 83.5719
R10701 Vbias.t483 Vbias.n6381 83.5719
R10702 Vbias.n6432 Vbias.n6431 83.5719
R10703 Vbias.t745 Vbias.n6432 83.5719
R10704 Vbias.n6427 Vbias.n6425 83.5719
R10705 Vbias.n6425 Vbias.t344 83.5719
R10706 Vbias.n6547 Vbias.n6430 83.5719
R10707 Vbias.t745 Vbias.n6430 83.5719
R10708 Vbias.n6550 Vbias.n6426 83.5719
R10709 Vbias.n6426 Vbias.t344 83.5719
R10710 Vbias.n6449 Vbias.n6448 83.5719
R10711 Vbias.t373 Vbias.n6449 83.5719
R10712 Vbias.n6458 Vbias.n6457 83.5719
R10713 Vbias.n6458 Vbias.t753 83.5719
R10714 Vbias.n6441 Vbias.n6439 83.5719
R10715 Vbias.n6439 Vbias.t231 83.5719
R10716 Vbias.n6535 Vbias.n6447 83.5719
R10717 Vbias.t373 Vbias.n6447 83.5719
R10718 Vbias.n6537 Vbias.n6445 83.5719
R10719 Vbias.t753 Vbias.n6445 83.5719
R10720 Vbias.n6540 Vbias.n6440 83.5719
R10721 Vbias.n6440 Vbias.t231 83.5719
R10722 Vbias.n6183 Vbias.n6182 83.5719
R10723 Vbias.n6183 Vbias.t132 83.5719
R10724 Vbias.n6180 Vbias.n6179 83.5719
R10725 Vbias.n6179 Vbias.t860 83.5719
R10726 Vbias.n6172 Vbias.n6171 83.5719
R10727 Vbias.t224 Vbias.n6172 83.5719
R10728 Vbias.n6628 Vbias.n6160 83.5719
R10729 Vbias.t132 Vbias.n6160 83.5719
R10730 Vbias.n6630 Vbias.n6158 83.5719
R10731 Vbias.t860 Vbias.n6158 83.5719
R10732 Vbias.n6632 Vbias.n6156 83.5719
R10733 Vbias.t224 Vbias.n6156 83.5719
R10734 Vbias.n6165 Vbias.n6164 83.5719
R10735 Vbias.t383 Vbias.n6165 83.5719
R10736 Vbias.n6624 Vbias.n6163 83.5719
R10737 Vbias.t383 Vbias.n6163 83.5719
R10738 Vbias.n6195 Vbias.n6194 83.5719
R10739 Vbias.t749 Vbias.n6195 83.5719
R10740 Vbias.n6190 Vbias.n6188 83.5719
R10741 Vbias.n6188 Vbias.t733 83.5719
R10742 Vbias.n6614 Vbias.n6193 83.5719
R10743 Vbias.t749 Vbias.n6193 83.5719
R10744 Vbias.n6617 Vbias.n6189 83.5719
R10745 Vbias.n6189 Vbias.t733 83.5719
R10746 Vbias.n6212 Vbias.n6211 83.5719
R10747 Vbias.t770 Vbias.n6212 83.5719
R10748 Vbias.n6221 Vbias.n6220 83.5719
R10749 Vbias.n6221 Vbias.t515 83.5719
R10750 Vbias.n6204 Vbias.n6202 83.5719
R10751 Vbias.n6202 Vbias.t186 83.5719
R10752 Vbias.n6602 Vbias.n6210 83.5719
R10753 Vbias.t770 Vbias.n6210 83.5719
R10754 Vbias.n6604 Vbias.n6208 83.5719
R10755 Vbias.t515 Vbias.n6208 83.5719
R10756 Vbias.n6607 Vbias.n6203 83.5719
R10757 Vbias.n6203 Vbias.t186 83.5719
R10758 Vbias.n6637 Vbias.n6636 83.5719
R10759 Vbias.t865 Vbias.n6637 83.5719
R10760 Vbias.n6145 Vbias.n6137 83.5719
R10761 Vbias.t625 Vbias.n6145 83.5719
R10762 Vbias.n6639 Vbias.n6638 83.5719
R10763 Vbias.n6638 Vbias.t865 83.5719
R10764 Vbias.n6642 Vbias.n6641 83.5719
R10765 Vbias.t625 Vbias.n6642 83.5719
R10766 Vbias.n6143 Vbias.n6142 83.5719
R10767 Vbias.t74 Vbias.n6143 83.5719
R10768 Vbias.n6647 Vbias.n6136 83.5719
R10769 Vbias.t74 Vbias.n6136 83.5719
R10770 Vbias.n7725 Vbias.n7724 83.5719
R10771 Vbias.n7724 Vbias.t487 83.5719
R10772 Vbias.n7728 Vbias.n7727 83.5719
R10773 Vbias.t623 Vbias.n7728 83.5719
R10774 Vbias.n681 Vbias.n679 83.5719
R10775 Vbias.n679 Vbias.t24 83.5719
R10776 Vbias.n7723 Vbias.n7722 83.5719
R10777 Vbias.t487 Vbias.n7723 83.5719
R10778 Vbias.n7730 Vbias.n7729 83.5719
R10779 Vbias.n7729 Vbias.t623 83.5719
R10780 Vbias.n7732 Vbias.n680 83.5719
R10781 Vbias.n680 Vbias.t24 83.5719
R10782 Vbias.n7710 Vbias.n7709 83.5719
R10783 Vbias.n7709 Vbias.t292 83.5719
R10784 Vbias.n7713 Vbias.n7712 83.5719
R10785 Vbias.t778 Vbias.n7713 83.5719
R10786 Vbias.n709 Vbias.n708 83.5719
R10787 Vbias.t245 Vbias.n709 83.5719
R10788 Vbias.n7708 Vbias.n7707 83.5719
R10789 Vbias.t292 Vbias.n7708 83.5719
R10790 Vbias.n711 Vbias.n702 83.5719
R10791 Vbias.t778 Vbias.n711 83.5719
R10792 Vbias.n7718 Vbias.n701 83.5719
R10793 Vbias.t245 Vbias.n701 83.5719
R10794 Vbias.n723 Vbias.n722 83.5719
R10795 Vbias.t332 Vbias.n723 83.5719
R10796 Vbias.n7703 Vbias.n721 83.5719
R10797 Vbias.t332 Vbias.n721 83.5719
R10798 Vbias.n7691 Vbias.n7690 83.5719
R10799 Vbias.t540 Vbias.n7691 83.5719
R10800 Vbias.n728 Vbias.n726 83.5719
R10801 Vbias.n726 Vbias.t671 83.5719
R10802 Vbias.n7693 Vbias.n7692 83.5719
R10803 Vbias.n7692 Vbias.t540 83.5719
R10804 Vbias.n7696 Vbias.n727 83.5719
R10805 Vbias.n727 Vbias.t671 83.5719
R10806 Vbias.n7673 Vbias.n7672 83.5719
R10807 Vbias.n7672 Vbias.t552 83.5719
R10808 Vbias.n7676 Vbias.n7675 83.5719
R10809 Vbias.t706 Vbias.n7676 83.5719
R10810 Vbias.n737 Vbias.n735 83.5719
R10811 Vbias.n735 Vbias.t200 83.5719
R10812 Vbias.n7671 Vbias.n7670 83.5719
R10813 Vbias.t552 Vbias.n7671 83.5719
R10814 Vbias.n7678 Vbias.n7677 83.5719
R10815 Vbias.n7677 Vbias.t706 83.5719
R10816 Vbias.n7681 Vbias.n736 83.5719
R10817 Vbias.n736 Vbias.t200 83.5719
R10818 Vbias.n6668 Vbias.n6667 83.5719
R10819 Vbias.t539 Vbias.n6668 83.5719
R10820 Vbias.n1470 Vbias.n1468 83.5719
R10821 Vbias.n1468 Vbias.t293 83.5719
R10822 Vbias.n6670 Vbias.n6669 83.5719
R10823 Vbias.n6669 Vbias.t539 83.5719
R10824 Vbias.n6672 Vbias.n1469 83.5719
R10825 Vbias.n1469 Vbias.t293 83.5719
R10826 Vbias.n6654 Vbias.n6653 83.5719
R10827 Vbias.t549 Vbias.n6654 83.5719
R10828 Vbias.n6661 Vbias.n6660 83.5719
R10829 Vbias.n6660 Vbias.t537 83.5719
R10830 Vbias.n6663 Vbias.n1483 83.5719
R10831 Vbias.n1483 Vbias.t52 83.5719
R10832 Vbias.n6656 Vbias.n6655 83.5719
R10833 Vbias.n6655 Vbias.t549 83.5719
R10834 Vbias.n6659 Vbias.n6658 83.5719
R10835 Vbias.t537 Vbias.n6659 83.5719
R10836 Vbias.n1495 Vbias.n1494 83.5719
R10837 Vbias.n1494 Vbias.t52 83.5719
R10838 Vbias.n6311 Vbias.n6299 83.5719
R10839 Vbias.t611 Vbias.n6299 83.5719
R10840 Vbias.n6301 Vbias.n6300 83.5719
R10841 Vbias.t611 Vbias.n6301 83.5719
R10842 Vbias.n6325 Vbias.n6324 83.5719
R10843 Vbias.n6324 Vbias.t444 83.5719
R10844 Vbias.n6318 Vbias.n6317 83.5719
R10845 Vbias.t608 Vbias.n6318 83.5719
R10846 Vbias.n6315 Vbias.n6296 83.5719
R10847 Vbias.t253 Vbias.n6296 83.5719
R10848 Vbias.n6323 Vbias.n6322 83.5719
R10849 Vbias.t444 Vbias.n6323 83.5719
R10850 Vbias.n6320 Vbias.n6319 83.5719
R10851 Vbias.n6319 Vbias.t608 83.5719
R10852 Vbias.n6305 Vbias.n6304 83.5719
R10853 Vbias.n6305 Vbias.t253 83.5719
R10854 Vbias.n6339 Vbias.n6338 83.5719
R10855 Vbias.n6338 Vbias.t735 83.5719
R10856 Vbias.n6332 Vbias.n6331 83.5719
R10857 Vbias.t755 Vbias.n6332 83.5719
R10858 Vbias.n6329 Vbias.n6274 83.5719
R10859 Vbias.t18 Vbias.n6274 83.5719
R10860 Vbias.n6337 Vbias.n6336 83.5719
R10861 Vbias.t735 Vbias.n6337 83.5719
R10862 Vbias.n6334 Vbias.n6333 83.5719
R10863 Vbias.n6333 Vbias.t755 83.5719
R10864 Vbias.n6282 Vbias.n6281 83.5719
R10865 Vbias.n6282 Vbias.t18 83.5719
R10866 Vbias.n6247 Vbias.n6245 83.5719
R10867 Vbias.n6245 Vbias.t748 83.5719
R10868 Vbias.n6345 Vbias.n6344 83.5719
R10869 Vbias.t464 Vbias.n6345 83.5719
R10870 Vbias.n6349 Vbias.n6246 83.5719
R10871 Vbias.n6246 Vbias.t748 83.5719
R10872 Vbias.n6347 Vbias.n6346 83.5719
R10873 Vbias.n6346 Vbias.t464 83.5719
R10874 Vbias.n6229 Vbias.n6227 83.5719
R10875 Vbias.n6227 Vbias.t501 83.5719
R10876 Vbias.n6582 Vbias.n6581 83.5719
R10877 Vbias.t521 Vbias.n6582 83.5719
R10878 Vbias.n6357 Vbias.n6356 83.5719
R10879 Vbias.n6356 Vbias.t78 83.5719
R10880 Vbias.n6586 Vbias.n6228 83.5719
R10881 Vbias.n6228 Vbias.t501 83.5719
R10882 Vbias.n6584 Vbias.n6583 83.5719
R10883 Vbias.n6583 Vbias.t521 83.5719
R10884 Vbias.n6355 Vbias.n6354 83.5719
R10885 Vbias.t78 Vbias.n6355 83.5719
R10886 Vbias.n780 Vbias.n778 83.5719
R10887 Vbias.n778 Vbias.t366 83.5719
R10888 Vbias.n7648 Vbias.n779 83.5719
R10889 Vbias.n779 Vbias.t366 83.5719
R10890 Vbias.n7634 Vbias.n7633 83.5719
R10891 Vbias.n7633 Vbias.t657 83.5719
R10892 Vbias.n7637 Vbias.n7636 83.5719
R10893 Vbias.t769 Vbias.n7637 83.5719
R10894 Vbias.n783 Vbias.n781 83.5719
R10895 Vbias.n781 Vbias.t233 83.5719
R10896 Vbias.n7632 Vbias.n7631 83.5719
R10897 Vbias.t657 Vbias.n7632 83.5719
R10898 Vbias.n7639 Vbias.n7638 83.5719
R10899 Vbias.n7638 Vbias.t769 83.5719
R10900 Vbias.n7641 Vbias.n782 83.5719
R10901 Vbias.n782 Vbias.t233 83.5719
R10902 Vbias.n7619 Vbias.n7618 83.5719
R10903 Vbias.n7618 Vbias.t346 83.5719
R10904 Vbias.n7622 Vbias.n7621 83.5719
R10905 Vbias.t847 Vbias.n7622 83.5719
R10906 Vbias.n802 Vbias.n800 83.5719
R10907 Vbias.n800 Vbias.t96 83.5719
R10908 Vbias.n7617 Vbias.n7616 83.5719
R10909 Vbias.t346 Vbias.n7617 83.5719
R10910 Vbias.n7624 Vbias.n7623 83.5719
R10911 Vbias.n7623 Vbias.t847 83.5719
R10912 Vbias.n7626 Vbias.n801 83.5719
R10913 Vbias.n801 Vbias.t96 83.5719
R10914 Vbias.n7607 Vbias.n7606 83.5719
R10915 Vbias.t353 Vbias.n7607 83.5719
R10916 Vbias.n824 Vbias.n822 83.5719
R10917 Vbias.n822 Vbias.t564 83.5719
R10918 Vbias.n7609 Vbias.n7608 83.5719
R10919 Vbias.n7608 Vbias.t353 83.5719
R10920 Vbias.n7611 Vbias.n823 83.5719
R10921 Vbias.n823 Vbias.t564 83.5719
R10922 Vbias.n7593 Vbias.n7592 83.5719
R10923 Vbias.t649 Vbias.n7593 83.5719
R10924 Vbias.n7600 Vbias.n7599 83.5719
R10925 Vbias.n7599 Vbias.t0 83.5719
R10926 Vbias.n7602 Vbias.n838 83.5719
R10927 Vbias.t34 Vbias.n838 83.5719
R10928 Vbias.n7595 Vbias.n7594 83.5719
R10929 Vbias.n7594 Vbias.t649 83.5719
R10930 Vbias.n7598 Vbias.n7597 83.5719
R10931 Vbias.t0 Vbias.n7598 83.5719
R10932 Vbias.n851 Vbias.n850 83.5719
R10933 Vbias.n850 Vbias.t34 83.5719
R10934 Vbias.n931 Vbias.n929 83.5719
R10935 Vbias.n929 Vbias.t156 83.5719
R10936 Vbias.n7527 Vbias.n930 83.5719
R10937 Vbias.n930 Vbias.t156 83.5719
R10938 Vbias.n7513 Vbias.n7512 83.5719
R10939 Vbias.n7512 Vbias.t399 83.5719
R10940 Vbias.n7516 Vbias.n7515 83.5719
R10941 Vbias.t376 Vbias.n7516 83.5719
R10942 Vbias.n934 Vbias.n932 83.5719
R10943 Vbias.n932 Vbias.t208 83.5719
R10944 Vbias.n7511 Vbias.n7510 83.5719
R10945 Vbias.t399 Vbias.n7511 83.5719
R10946 Vbias.n7518 Vbias.n7517 83.5719
R10947 Vbias.n7517 Vbias.t376 83.5719
R10948 Vbias.n7520 Vbias.n933 83.5719
R10949 Vbias.n933 Vbias.t208 83.5719
R10950 Vbias.n7498 Vbias.n7497 83.5719
R10951 Vbias.n7497 Vbias.t806 83.5719
R10952 Vbias.n7501 Vbias.n7500 83.5719
R10953 Vbias.t377 Vbias.n7501 83.5719
R10954 Vbias.n957 Vbias.n955 83.5719
R10955 Vbias.n955 Vbias.t16 83.5719
R10956 Vbias.n7496 Vbias.n7495 83.5719
R10957 Vbias.t806 Vbias.n7496 83.5719
R10958 Vbias.n7503 Vbias.n7502 83.5719
R10959 Vbias.n7502 Vbias.t377 83.5719
R10960 Vbias.n7505 Vbias.n956 83.5719
R10961 Vbias.n956 Vbias.t16 83.5719
R10962 Vbias.n7485 Vbias.n7484 83.5719
R10963 Vbias.t390 Vbias.n7485 83.5719
R10964 Vbias.n979 Vbias.n977 83.5719
R10965 Vbias.n977 Vbias.t571 83.5719
R10966 Vbias.n7487 Vbias.n7486 83.5719
R10967 Vbias.n7486 Vbias.t390 83.5719
R10968 Vbias.n7489 Vbias.n978 83.5719
R10969 Vbias.n978 Vbias.t571 83.5719
R10970 Vbias.n7471 Vbias.n7470 83.5719
R10971 Vbias.t699 Vbias.n7471 83.5719
R10972 Vbias.n7478 Vbias.n7477 83.5719
R10973 Vbias.n7477 Vbias.t703 83.5719
R10974 Vbias.n7480 Vbias.n993 83.5719
R10975 Vbias.t48 Vbias.n993 83.5719
R10976 Vbias.n7473 Vbias.n7472 83.5719
R10977 Vbias.n7472 Vbias.t699 83.5719
R10978 Vbias.n7476 Vbias.n7475 83.5719
R10979 Vbias.t703 Vbias.n7476 83.5719
R10980 Vbias.n1006 Vbias.n1005 83.5719
R10981 Vbias.n1005 Vbias.t48 83.5719
R10982 Vbias.n7320 Vbias.n1020 83.5719
R10983 Vbias.t477 Vbias.n1020 83.5719
R10984 Vbias.n1022 Vbias.n1021 83.5719
R10985 Vbias.t477 Vbias.n1022 83.5719
R10986 Vbias.n7306 Vbias.n7305 83.5719
R10987 Vbias.n7305 Vbias.t819 83.5719
R10988 Vbias.n7309 Vbias.n7308 83.5719
R10989 Vbias.t475 Vbias.n7309 83.5719
R10990 Vbias.n1031 Vbias.n1029 83.5719
R10991 Vbias.n1029 Vbias.t261 83.5719
R10992 Vbias.n7304 Vbias.n7303 83.5719
R10993 Vbias.t819 Vbias.n7304 83.5719
R10994 Vbias.n7311 Vbias.n7310 83.5719
R10995 Vbias.n7310 Vbias.t475 83.5719
R10996 Vbias.n7313 Vbias.n1030 83.5719
R10997 Vbias.n1030 Vbias.t261 83.5719
R10998 Vbias.n7291 Vbias.n7290 83.5719
R10999 Vbias.n7290 Vbias.t669 83.5719
R11000 Vbias.n7294 Vbias.n7293 83.5719
R11001 Vbias.t619 Vbias.n7294 83.5719
R11002 Vbias.n1052 Vbias.n1050 83.5719
R11003 Vbias.n1050 Vbias.t68 83.5719
R11004 Vbias.n7289 Vbias.n7288 83.5719
R11005 Vbias.t669 Vbias.n7289 83.5719
R11006 Vbias.n7296 Vbias.n7295 83.5719
R11007 Vbias.n7295 Vbias.t619 83.5719
R11008 Vbias.n7298 Vbias.n1051 83.5719
R11009 Vbias.n1051 Vbias.t68 83.5719
R11010 Vbias.n7279 Vbias.n7278 83.5719
R11011 Vbias.t580 Vbias.n7279 83.5719
R11012 Vbias.n7229 Vbias.n7227 83.5719
R11013 Vbias.n7227 Vbias.t143 83.5719
R11014 Vbias.n7281 Vbias.n7280 83.5719
R11015 Vbias.n7280 Vbias.t580 83.5719
R11016 Vbias.n7283 Vbias.n7228 83.5719
R11017 Vbias.n7228 Vbias.t143 83.5719
R11018 Vbias.n7264 Vbias.n7263 83.5719
R11019 Vbias.t566 Vbias.n7264 83.5719
R11020 Vbias.n7272 Vbias.n7271 83.5719
R11021 Vbias.n7271 Vbias.t788 83.5719
R11022 Vbias.n7274 Vbias.n7243 83.5719
R11023 Vbias.t116 Vbias.n7243 83.5719
R11024 Vbias.n7267 Vbias.n7266 83.5719
R11025 Vbias.n7270 Vbias.n7269 83.5719
R11026 Vbias.t788 Vbias.n7270 83.5719
R11027 Vbias.n7256 Vbias.n7255 83.5719
R11028 Vbias.n7255 Vbias.t116 83.5719
R11029 Vbias.n7664 Vbias.n7663 83.5719
R11030 Vbias.n7663 Vbias.t481 83.5719
R11031 Vbias.n7667 Vbias.n7666 83.5719
R11032 Vbias.t646 Vbias.n7667 83.5719
R11033 Vbias.n7662 Vbias.n7661 83.5719
R11034 Vbias.t481 Vbias.n7662 83.5719
R11035 Vbias.n769 Vbias.n758 83.5719
R11036 Vbias.t646 Vbias.n758 83.5719
R11037 Vbias.n777 Vbias.n776 83.5719
R11038 Vbias.t14 Vbias.n777 83.5719
R11039 Vbias.n6594 Vbias.n6593 83.5719
R11040 Vbias.n6594 Vbias.t607 83.5719
R11041 Vbias.n7655 Vbias.n775 83.5719
R11042 Vbias.t14 Vbias.n775 83.5719
R11043 Vbias.n7657 Vbias.n773 83.5719
R11044 Vbias.t607 Vbias.n773 83.5719
R11045 Vbias.n6507 Vbias.n6505 83.5719
R11046 Vbias.n6505 Vbias.t368 83.5719
R11047 Vbias.n6514 Vbias.n6506 83.5719
R11048 Vbias.n6506 Vbias.t368 83.5719
R11049 Vbias.n928 Vbias.n927 83.5719
R11050 Vbias.t328 Vbias.n928 83.5719
R11051 Vbias.n6530 Vbias.n6529 83.5719
R11052 Vbias.t402 Vbias.n6530 83.5719
R11053 Vbias.n7534 Vbias.n926 83.5719
R11054 Vbias.t328 Vbias.n926 83.5719
R11055 Vbias.n6523 Vbias.n6520 83.5719
R11056 Vbias.t402 Vbias.n6520 83.5719
R11057 Vbias.n1024 Vbias.n1023 83.5719
R11058 Vbias.n1024 Vbias.t717 83.5719
R11059 Vbias.n1014 Vbias.n1012 83.5719
R11060 Vbias.n1012 Vbias.t888 83.5719
R11061 Vbias.n7540 Vbias.n922 83.5719
R11062 Vbias.n922 Vbias.t717 83.5719
R11063 Vbias.n1013 Vbias.n921 83.5719
R11064 Vbias.n1013 Vbias.t888 83.5719
R11065 Vbias.n1503 Vbias.n1501 83.5719
R11066 Vbias.n1501 Vbias.t615 83.5719
R11067 Vbias.n6128 Vbias.n1502 83.5719
R11068 Vbias.n1502 Vbias.t615 83.5719
R11069 Vbias.n326 Vbias.n324 83.5719
R11070 Vbias.n324 Vbias.t621 83.5719
R11071 Vbias.n345 Vbias.n325 83.5719
R11072 Vbias.n325 Vbias.t621 83.5719
R11073 Vbias.n173 Vbias.n172 83.5719
R11074 Vbias.t811 Vbias.n173 83.5719
R11075 Vbias.n336 Vbias.n328 83.5719
R11076 Vbias.n328 Vbias.t440 83.5719
R11077 Vbias.n7941 Vbias.n171 83.5719
R11078 Vbias.t811 Vbias.n171 83.5719
R11079 Vbias.n338 Vbias.n329 83.5719
R11080 Vbias.n329 Vbias.t440 83.5719
R11081 Vbias.n5595 Vbias.n5590 83.5719
R11082 Vbias.n5590 Vbias.t415 83.5719
R11083 Vbias.n5598 Vbias.n5591 83.5719
R11084 Vbias.n5591 Vbias.t415 83.5719
R11085 Vbias.n5574 Vbias.n5572 83.5719
R11086 Vbias.n5572 Vbias.t659 83.5719
R11087 Vbias.n5612 Vbias.n5611 83.5719
R11088 Vbias.t2 Vbias.n5612 83.5719
R11089 Vbias.n5606 Vbias.n5605 83.5719
R11090 Vbias.n5605 Vbias.t235 83.5719
R11091 Vbias.n5616 Vbias.n5573 83.5719
R11092 Vbias.n5573 Vbias.t659 83.5719
R11093 Vbias.n5614 Vbias.n5613 83.5719
R11094 Vbias.n5613 Vbias.t2 83.5719
R11095 Vbias.n5604 Vbias.n5603 83.5719
R11096 Vbias.t235 Vbias.n5604 83.5719
R11097 Vbias.n5556 Vbias.n5554 83.5719
R11098 Vbias.t322 Vbias.n5554 83.5719
R11099 Vbias.n5631 Vbias.n5630 83.5719
R11100 Vbias.t306 Vbias.n5631 83.5719
R11101 Vbias.n5624 Vbias.n5623 83.5719
R11102 Vbias.n5623 Vbias.t90 83.5719
R11103 Vbias.n5635 Vbias.n5555 83.5719
R11104 Vbias.t322 Vbias.n5555 83.5719
R11105 Vbias.n5633 Vbias.n5632 83.5719
R11106 Vbias.n5632 Vbias.t306 83.5719
R11107 Vbias.n5622 Vbias.n5621 83.5719
R11108 Vbias.t90 Vbias.n5622 83.5719
R11109 Vbias.n5648 Vbias.n5647 83.5719
R11110 Vbias.n5647 Vbias.t634 83.5719
R11111 Vbias.n5641 Vbias.n5640 83.5719
R11112 Vbias.t431 Vbias.n5641 83.5719
R11113 Vbias.n5646 Vbias.n5645 83.5719
R11114 Vbias.t634 Vbias.n5646 83.5719
R11115 Vbias.n5643 Vbias.n5642 83.5719
R11116 Vbias.n5642 Vbias.t431 83.5719
R11117 Vbias.n5662 Vbias.n5661 83.5719
R11118 Vbias.n5661 Vbias.t630 83.5719
R11119 Vbias.n5655 Vbias.n5654 83.5719
R11120 Vbias.t291 Vbias.n5655 83.5719
R11121 Vbias.n5652 Vbias.n2211 83.5719
R11122 Vbias.t72 Vbias.n2211 83.5719
R11123 Vbias.n5660 Vbias.n5659 83.5719
R11124 Vbias.t630 Vbias.n5660 83.5719
R11125 Vbias.n5657 Vbias.n5656 83.5719
R11126 Vbias.n5656 Vbias.t291 83.5719
R11127 Vbias.n2219 Vbias.n2218 83.5719
R11128 Vbias.n2219 Vbias.t72 83.5719
R11129 Vbias.n7878 Vbias.n7877 83.5719
R11130 Vbias.t767 Vbias.n7878 83.5719
R11131 Vbias.n450 Vbias.n448 83.5719
R11132 Vbias.n448 Vbias.t3 83.5719
R11133 Vbias.n7880 Vbias.n7879 83.5719
R11134 Vbias.n7879 Vbias.t767 83.5719
R11135 Vbias.n7883 Vbias.n449 83.5719
R11136 Vbias.n449 Vbias.t3 83.5719
R11137 Vbias.n5669 Vbias.n2193 83.5719
R11138 Vbias.n2193 Vbias.t772 83.5719
R11139 Vbias.n5672 Vbias.n2194 83.5719
R11140 Vbias.n2194 Vbias.t772 83.5719
R11141 Vbias.n2177 Vbias.n2175 83.5719
R11142 Vbias.n2175 Vbias.t379 83.5719
R11143 Vbias.n5686 Vbias.n5685 83.5719
R11144 Vbias.t766 Vbias.n5686 83.5719
R11145 Vbias.n5680 Vbias.n5679 83.5719
R11146 Vbias.n5679 Vbias.t210 83.5719
R11147 Vbias.n5690 Vbias.n2176 83.5719
R11148 Vbias.n2176 Vbias.t379 83.5719
R11149 Vbias.n5688 Vbias.n5687 83.5719
R11150 Vbias.n5687 Vbias.t766 83.5719
R11151 Vbias.n5678 Vbias.n5677 83.5719
R11152 Vbias.t210 Vbias.n5678 83.5719
R11153 Vbias.n2159 Vbias.n2157 83.5719
R11154 Vbias.n2157 Vbias.t457 83.5719
R11155 Vbias.n5705 Vbias.n5704 83.5719
R11156 Vbias.t849 Vbias.n5705 83.5719
R11157 Vbias.n5698 Vbias.n5697 83.5719
R11158 Vbias.n5697 Vbias.t44 83.5719
R11159 Vbias.n5709 Vbias.n2158 83.5719
R11160 Vbias.n2158 Vbias.t457 83.5719
R11161 Vbias.n5707 Vbias.n5706 83.5719
R11162 Vbias.n5706 Vbias.t849 83.5719
R11163 Vbias.n5696 Vbias.n5695 83.5719
R11164 Vbias.t44 Vbias.n5696 83.5719
R11165 Vbias.n5722 Vbias.n5721 83.5719
R11166 Vbias.n5721 Vbias.t697 83.5719
R11167 Vbias.n5715 Vbias.n5714 83.5719
R11168 Vbias.t151 Vbias.n5715 83.5719
R11169 Vbias.n5720 Vbias.n5719 83.5719
R11170 Vbias.t697 Vbias.n5720 83.5719
R11171 Vbias.n5717 Vbias.n5716 83.5719
R11172 Vbias.n5716 Vbias.t151 83.5719
R11173 Vbias.n5736 Vbias.n5735 83.5719
R11174 Vbias.n5735 Vbias.t643 83.5719
R11175 Vbias.n5729 Vbias.n5728 83.5719
R11176 Vbias.t568 Vbias.n5729 83.5719
R11177 Vbias.n5726 Vbias.n2140 83.5719
R11178 Vbias.t80 Vbias.n2140 83.5719
R11179 Vbias.n5734 Vbias.n5733 83.5719
R11180 Vbias.t643 Vbias.n5734 83.5719
R11181 Vbias.n5731 Vbias.n5730 83.5719
R11182 Vbias.n5730 Vbias.t568 83.5719
R11183 Vbias.n2148 Vbias.n2147 83.5719
R11184 Vbias.n2148 Vbias.t80 83.5719
R11185 Vbias.n556 Vbias.n554 83.5719
R11186 Vbias.n554 Vbias.t628 83.5719
R11187 Vbias.n7817 Vbias.n555 83.5719
R11188 Vbias.n555 Vbias.t628 83.5719
R11189 Vbias.n7808 Vbias.n7807 83.5719
R11190 Vbias.t485 Vbias.n7808 83.5719
R11191 Vbias.n570 Vbias.n569 83.5719
R11192 Vbias.t850 Vbias.n570 83.5719
R11193 Vbias.n7804 Vbias.n561 83.5719
R11194 Vbias.t485 Vbias.n7804 83.5719
R11195 Vbias.n7813 Vbias.n560 83.5719
R11196 Vbias.t850 Vbias.n560 83.5719
R11197 Vbias.n5754 Vbias.n5743 83.5719
R11198 Vbias.t821 Vbias.n5743 83.5719
R11199 Vbias.n5746 Vbias.n5744 83.5719
R11200 Vbias.t821 Vbias.n5746 83.5719
R11201 Vbias.n5768 Vbias.n5767 83.5719
R11202 Vbias.n5767 Vbias.t585 83.5719
R11203 Vbias.n5761 Vbias.n5760 83.5719
R11204 Vbias.t350 Vbias.n5761 83.5719
R11205 Vbias.n5758 Vbias.n2123 83.5719
R11206 Vbias.t174 Vbias.n2123 83.5719
R11207 Vbias.n5766 Vbias.n5765 83.5719
R11208 Vbias.t585 Vbias.n5766 83.5719
R11209 Vbias.n5763 Vbias.n5762 83.5719
R11210 Vbias.n5762 Vbias.t350 83.5719
R11211 Vbias.n5748 Vbias.n5747 83.5719
R11212 Vbias.n5748 Vbias.t174 83.5719
R11213 Vbias.n5783 Vbias.n5782 83.5719
R11214 Vbias.n5782 Vbias.t857 83.5719
R11215 Vbias.n5775 Vbias.n5774 83.5719
R11216 Vbias.t805 Vbias.n5775 83.5719
R11217 Vbias.n5772 Vbias.n2101 83.5719
R11218 Vbias.t102 Vbias.n2101 83.5719
R11219 Vbias.n5780 Vbias.n5779 83.5719
R11220 Vbias.n5780 Vbias.t857 83.5719
R11221 Vbias.n5777 Vbias.n5776 83.5719
R11222 Vbias.n5776 Vbias.t805 83.5719
R11223 Vbias.n2109 Vbias.n2108 83.5719
R11224 Vbias.n2109 Vbias.t102 83.5719
R11225 Vbias.n5811 Vbias.n5810 83.5719
R11226 Vbias.n5810 Vbias.t401 83.5719
R11227 Vbias.n5804 Vbias.n5803 83.5719
R11228 Vbias.t682 Vbias.n5804 83.5719
R11229 Vbias.n5809 Vbias.n5808 83.5719
R11230 Vbias.t401 Vbias.n5809 83.5719
R11231 Vbias.n5806 Vbias.n5805 83.5719
R11232 Vbias.n5805 Vbias.t682 83.5719
R11233 Vbias.n5825 Vbias.n5824 83.5719
R11234 Vbias.n5824 Vbias.t494 83.5719
R11235 Vbias.n5818 Vbias.n5817 83.5719
R11236 Vbias.t648 Vbias.n5818 83.5719
R11237 Vbias.n5815 Vbias.n2085 83.5719
R11238 Vbias.t106 Vbias.n2085 83.5719
R11239 Vbias.n5823 Vbias.n5822 83.5719
R11240 Vbias.t494 Vbias.n5823 83.5719
R11241 Vbias.n5820 Vbias.n5819 83.5719
R11242 Vbias.n5819 Vbias.t648 83.5719
R11243 Vbias.n5793 Vbias.n5792 83.5719
R11244 Vbias.n5793 Vbias.t106 83.5719
R11245 Vbias.n7743 Vbias.n7742 83.5719
R11246 Vbias.t713 Vbias.n7743 83.5719
R11247 Vbias.n670 Vbias.n668 83.5719
R11248 Vbias.n668 Vbias.t820 83.5719
R11249 Vbias.n7745 Vbias.n7744 83.5719
R11250 Vbias.n7744 Vbias.t713 83.5719
R11251 Vbias.n7748 Vbias.n669 83.5719
R11252 Vbias.n669 Vbias.t820 83.5719
R11253 Vbias.n5840 Vbias.n5833 83.5719
R11254 Vbias.t784 Vbias.n5833 83.5719
R11255 Vbias.n5836 Vbias.n5834 83.5719
R11256 Vbias.t784 Vbias.n5836 83.5719
R11257 Vbias.n5854 Vbias.n5853 83.5719
R11258 Vbias.n5853 Vbias.t392 83.5719
R11259 Vbias.n5857 Vbias.n5856 83.5719
R11260 Vbias.t712 Vbias.n5857 83.5719
R11261 Vbias.n5845 Vbias.n5844 83.5719
R11262 Vbias.t202 Vbias.n5845 83.5719
R11263 Vbias.n5852 Vbias.n5851 83.5719
R11264 Vbias.t392 Vbias.n5852 83.5719
R11265 Vbias.n5849 Vbias.n1695 83.5719
R11266 Vbias.t712 Vbias.n1695 83.5719
R11267 Vbias.n5847 Vbias.n5846 83.5719
R11268 Vbias.n5846 Vbias.t202 83.5719
R11269 Vbias.n1706 Vbias.n1704 83.5719
R11270 Vbias.n1704 Vbias.t30 83.5719
R11271 Vbias.n2056 Vbias.n1705 83.5719
R11272 Vbias.n1705 Vbias.t30 83.5719
R11273 Vbias.n2048 Vbias.n2047 83.5719
R11274 Vbias.n2047 Vbias.t670 83.5719
R11275 Vbias.n2052 Vbias.n2051 83.5719
R11276 Vbias.t777 Vbias.n2052 83.5719
R11277 Vbias.n2046 Vbias.n2045 83.5719
R11278 Vbias.t670 Vbias.n2046 83.5719
R11279 Vbias.n2054 Vbias.n2053 83.5719
R11280 Vbias.n2053 Vbias.t777 83.5719
R11281 Vbias.n2038 Vbias.n1730 83.5719
R11282 Vbias.t341 Vbias.n2038 83.5719
R11283 Vbias.n2044 Vbias.n2043 83.5719
R11284 Vbias.t559 Vbias.n2044 83.5719
R11285 Vbias.n1738 Vbias.n1737 83.5719
R11286 Vbias.n1738 Vbias.t557 83.5719
R11287 Vbias.n2035 Vbias.n1733 83.5719
R11288 Vbias.t341 Vbias.n1733 83.5719
R11289 Vbias.n1745 Vbias.n1726 83.5719
R11290 Vbias.t559 Vbias.n1726 83.5719
R11291 Vbias.n1743 Vbias.n1742 83.5719
R11292 Vbias.n1742 Vbias.t557 83.5719
R11293 Vbias.n1447 Vbias.n1445 83.5719
R11294 Vbias.n1445 Vbias.t760 83.5719
R11295 Vbias.n6746 Vbias.n1446 83.5719
R11296 Vbias.n1446 Vbias.t760 83.5719
R11297 Vbias.n6724 Vbias.n6723 83.5719
R11298 Vbias.t737 Vbias.n6724 83.5719
R11299 Vbias.n6731 Vbias.n6730 83.5719
R11300 Vbias.n6731 Vbias.t407 83.5719
R11301 Vbias.n6740 Vbias.n6722 83.5719
R11302 Vbias.t737 Vbias.n6722 83.5719
R11303 Vbias.n6742 Vbias.n6720 83.5719
R11304 Vbias.t407 Vbias.n6720 83.5719
R11305 Vbias.n6700 Vbias.n6699 83.5719
R11306 Vbias.t677 Vbias.n6700 83.5719
R11307 Vbias.n6705 Vbias.n6704 83.5719
R11308 Vbias.n6705 Vbias.t229 83.5719
R11309 Vbias.n6713 Vbias.n6698 83.5719
R11310 Vbias.t677 Vbias.n6698 83.5719
R11311 Vbias.n6715 Vbias.n6696 83.5719
R11312 Vbias.t229 Vbias.n6696 83.5719
R11313 Vbias.n6690 Vbias.n1451 83.5719
R11314 Vbias.t723 Vbias.n1451 83.5719
R11315 Vbias.n6687 Vbias.n1452 83.5719
R11316 Vbias.n6687 Vbias.t723 83.5719
R11317 Vbias.n6682 Vbias.n6681 83.5719
R11318 Vbias.n6681 Vbias.t744 83.5719
R11319 Vbias.n1457 Vbias.n1456 83.5719
R11320 Vbias.n1457 Vbias.t744 83.5719
R11321 Vbias.n8065 Vbias.n8064 83.5719
R11322 Vbias.n8064 Vbias.t313 83.5719
R11323 Vbias.n8068 Vbias.n8067 83.5719
R11324 Vbias.t631 Vbias.n8068 83.5719
R11325 Vbias.n12 Vbias.n10 83.5719
R11326 Vbias.n10 Vbias.t158 83.5719
R11327 Vbias.n8063 Vbias.n8062 83.5719
R11328 Vbias.t313 Vbias.n8063 83.5719
R11329 Vbias.n8070 Vbias.n8069 83.5719
R11330 Vbias.n8069 Vbias.t631 83.5719
R11331 Vbias.n8072 Vbias.n11 83.5719
R11332 Vbias.n11 Vbias.t158 83.5719
R11333 Vbias.n8050 Vbias.n8049 83.5719
R11334 Vbias.n8049 Vbias.t798 83.5719
R11335 Vbias.n8053 Vbias.n8052 83.5719
R11336 Vbias.t360 Vbias.n8053 83.5719
R11337 Vbias.n40 Vbias.n39 83.5719
R11338 Vbias.t674 Vbias.n40 83.5719
R11339 Vbias.n8048 Vbias.n8047 83.5719
R11340 Vbias.t798 Vbias.n8048 83.5719
R11341 Vbias.n42 Vbias.n33 83.5719
R11342 Vbias.t360 Vbias.n42 83.5719
R11343 Vbias.n8058 Vbias.n32 83.5719
R11344 Vbias.t674 Vbias.n32 83.5719
R11345 Vbias.n54 Vbias.n53 83.5719
R11346 Vbias.t323 Vbias.n54 83.5719
R11347 Vbias.n8043 Vbias.n52 83.5719
R11348 Vbias.t323 Vbias.n52 83.5719
R11349 Vbias.n8031 Vbias.n8030 83.5719
R11350 Vbias.t307 Vbias.n8031 83.5719
R11351 Vbias.n59 Vbias.n57 83.5719
R11352 Vbias.n57 Vbias.t418 83.5719
R11353 Vbias.n8033 Vbias.n8032 83.5719
R11354 Vbias.n8032 Vbias.t307 83.5719
R11355 Vbias.n8036 Vbias.n58 83.5719
R11356 Vbias.n58 Vbias.t418 83.5719
R11357 Vbias.n8013 Vbias.n8012 83.5719
R11358 Vbias.n8012 Vbias.t694 83.5719
R11359 Vbias.n8016 Vbias.n8015 83.5719
R11360 Vbias.t533 Vbias.n8016 83.5719
R11361 Vbias.n68 Vbias.n66 83.5719
R11362 Vbias.n66 Vbias.t522 83.5719
R11363 Vbias.n8011 Vbias.n8010 83.5719
R11364 Vbias.t694 Vbias.n8011 83.5719
R11365 Vbias.n8018 Vbias.n8017 83.5719
R11366 Vbias.n8017 Vbias.t533 83.5719
R11367 Vbias.n8021 Vbias.n67 83.5719
R11368 Vbias.n67 Vbias.t522 83.5719
R11369 Vbias.n89 Vbias.n87 83.5719
R11370 Vbias.n87 Vbias.t791 83.5719
R11371 Vbias.n8004 Vbias.n88 83.5719
R11372 Vbias.n88 Vbias.t791 83.5719
R11373 Vbias.n7990 Vbias.n7989 83.5719
R11374 Vbias.n7989 Vbias.t813 83.5719
R11375 Vbias.n7993 Vbias.n7992 83.5719
R11376 Vbias.t790 Vbias.n7993 83.5719
R11377 Vbias.n92 Vbias.n90 83.5719
R11378 Vbias.n90 Vbias.t257 83.5719
R11379 Vbias.n7988 Vbias.n7987 83.5719
R11380 Vbias.t813 Vbias.n7988 83.5719
R11381 Vbias.n7995 Vbias.n7994 83.5719
R11382 Vbias.n7994 Vbias.t790 83.5719
R11383 Vbias.n7997 Vbias.n91 83.5719
R11384 Vbias.n91 Vbias.t257 83.5719
R11385 Vbias.n7975 Vbias.n7974 83.5719
R11386 Vbias.n7974 Vbias.t538 83.5719
R11387 Vbias.n7978 Vbias.n7977 83.5719
R11388 Vbias.t288 Vbias.n7978 83.5719
R11389 Vbias.n111 Vbias.n109 83.5719
R11390 Vbias.n109 Vbias.t46 83.5719
R11391 Vbias.n7973 Vbias.n7972 83.5719
R11392 Vbias.t538 Vbias.n7973 83.5719
R11393 Vbias.n7980 Vbias.n7979 83.5719
R11394 Vbias.n7979 Vbias.t288 83.5719
R11395 Vbias.n7982 Vbias.n110 83.5719
R11396 Vbias.n110 Vbias.t46 83.5719
R11397 Vbias.n7963 Vbias.n7962 83.5719
R11398 Vbias.t858 Vbias.n7963 83.5719
R11399 Vbias.n132 Vbias.n130 83.5719
R11400 Vbias.n130 Vbias.t356 83.5719
R11401 Vbias.n7965 Vbias.n7964 83.5719
R11402 Vbias.n7964 Vbias.t858 83.5719
R11403 Vbias.n7967 Vbias.n131 83.5719
R11404 Vbias.n131 Vbias.t356 83.5719
R11405 Vbias.n7949 Vbias.n7948 83.5719
R11406 Vbias.t518 Vbias.n7949 83.5719
R11407 Vbias.n7956 Vbias.n7955 83.5719
R11408 Vbias.n7955 Vbias.t801 83.5719
R11409 Vbias.n7958 Vbias.n146 83.5719
R11410 Vbias.t20 Vbias.n146 83.5719
R11411 Vbias.n7951 Vbias.n7950 83.5719
R11412 Vbias.n7950 Vbias.t518 83.5719
R11413 Vbias.n7954 Vbias.n7953 83.5719
R11414 Vbias.t801 Vbias.n7954 83.5719
R11415 Vbias.n159 Vbias.n158 83.5719
R11416 Vbias.n158 Vbias.t20 83.5719
R11417 Vbias.n2602 Vbias.n2600 83.5719
R11418 Vbias.n2600 Vbias.t739 83.5719
R11419 Vbias.n4989 Vbias.n2601 83.5719
R11420 Vbias.n2601 Vbias.t739 83.5719
R11421 Vbias.n2595 Vbias.n2593 83.5719
R11422 Vbias.n2593 Vbias.t700 83.5719
R11423 Vbias.n5000 Vbias.n4999 83.5719
R11424 Vbias.t410 Vbias.n5000 83.5719
R11425 Vbias.n5006 Vbias.n2594 83.5719
R11426 Vbias.n2594 Vbias.t700 83.5719
R11427 Vbias.n5002 Vbias.n5001 83.5719
R11428 Vbias.n5001 Vbias.t410 83.5719
R11429 Vbias.n5021 Vbias.n5020 83.5719
R11430 Vbias.t829 Vbias.n5021 83.5719
R11431 Vbias.n5015 Vbias.n5014 83.5719
R11432 Vbias.t787 Vbias.n5015 83.5719
R11433 Vbias.n5017 Vbias.n2588 83.5719
R11434 Vbias.t829 Vbias.n5017 83.5719
R11435 Vbias.n5026 Vbias.n2587 83.5719
R11436 Vbias.t787 Vbias.n2587 83.5719
R11437 Vbias.n2231 Vbias.n2229 83.5719
R11438 Vbias.n2229 Vbias.t655 83.5719
R11439 Vbias.n5549 Vbias.n2230 83.5719
R11440 Vbias.n2230 Vbias.t655 83.5719
R11441 Vbias.n5540 Vbias.n5539 83.5719
R11442 Vbias.t719 Vbias.n5540 83.5719
R11443 Vbias.n2245 Vbias.n2244 83.5719
R11444 Vbias.t862 Vbias.n2245 83.5719
R11445 Vbias.n5536 Vbias.n2236 83.5719
R11446 Vbias.t719 Vbias.n5536 83.5719
R11447 Vbias.n5545 Vbias.n2235 83.5719
R11448 Vbias.t862 Vbias.n2235 83.5719
R11449 Vbias.n5524 Vbias.n5523 83.5719
R11450 Vbias.t135 Vbias.n5524 83.5719
R11451 Vbias.n5511 Vbias.n5509 83.5719
R11452 Vbias.n5509 Vbias.t604 83.5719
R11453 Vbias.n5526 Vbias.n5525 83.5719
R11454 Vbias.n5525 Vbias.t135 83.5719
R11455 Vbias.n5529 Vbias.n5510 83.5719
R11456 Vbias.n5510 Vbias.t604 83.5719
R11457 Vbias.n1677 Vbias.n1675 83.5719
R11458 Vbias.n1675 Vbias.t370 83.5719
R11459 Vbias.n5873 Vbias.n1676 83.5719
R11460 Vbias.n1676 Vbias.t370 83.5719
R11461 Vbias.n5864 Vbias.n5863 83.5719
R11462 Vbias.t7 Vbias.n5864 83.5719
R11463 Vbias.n1692 Vbias.n1691 83.5719
R11464 Vbias.t409 Vbias.n1692 83.5719
R11465 Vbias.n5860 Vbias.n1683 83.5719
R11466 Vbias.t7 Vbias.n5860 83.5719
R11467 Vbias.n5869 Vbias.n1682 83.5719
R11468 Vbias.t409 Vbias.n1682 83.5719
R11469 Vbias.n4265 Vbias.n4257 83.5719
R11470 Vbias.t837 Vbias.n4257 83.5719
R11471 Vbias.n4259 Vbias.n4258 83.5719
R11472 Vbias.t837 Vbias.n4259 83.5719
R11473 Vbias.n4298 Vbias.n2862 83.5719
R11474 Vbias.t502 Vbias.n2862 83.5719
R11475 Vbias.n4289 Vbias.n2875 83.5719
R11476 Vbias.t576 Vbias.n2875 83.5719
R11477 Vbias.n4269 Vbias.n2886 83.5719
R11478 Vbias.t84 Vbias.n2886 83.5719
R11479 Vbias.n4280 Vbias.n2867 83.5719
R11480 Vbias.t502 Vbias.n2867 83.5719
R11481 Vbias.n4277 Vbias.n2876 83.5719
R11482 Vbias.t576 Vbias.n2876 83.5719
R11483 Vbias.n4275 Vbias.n4274 83.5719
R11484 Vbias.n4274 Vbias.t84 83.5719
R11485 Vbias.n4331 Vbias.n2826 83.5719
R11486 Vbias.t343 Vbias.n2826 83.5719
R11487 Vbias.n4322 Vbias.n2841 83.5719
R11488 Vbias.t596 Vbias.n2841 83.5719
R11489 Vbias.n4302 Vbias.n2852 83.5719
R11490 Vbias.t167 Vbias.n2852 83.5719
R11491 Vbias.n4313 Vbias.n2831 83.5719
R11492 Vbias.t343 Vbias.n2831 83.5719
R11493 Vbias.n4310 Vbias.n2842 83.5719
R11494 Vbias.t596 Vbias.n2842 83.5719
R11495 Vbias.n4308 Vbias.n4307 83.5719
R11496 Vbias.n4307 Vbias.t167 83.5719
R11497 Vbias.n4360 Vbias.n2808 83.5719
R11498 Vbias.n2808 Vbias.t466 83.5719
R11499 Vbias.n4357 Vbias.n2812 83.5719
R11500 Vbias.t128 Vbias.n2812 83.5719
R11501 Vbias.n4348 Vbias.n4347 83.5719
R11502 Vbias.n4347 Vbias.t466 83.5719
R11503 Vbias.n4346 Vbias.n4345 83.5719
R11504 Vbias.n4345 Vbias.t128 83.5719
R11505 Vbias.n2787 Vbias.n2781 83.5719
R11506 Vbias.n2787 Vbias.t162 83.5719
R11507 Vbias.n4386 Vbias.n2789 83.5719
R11508 Vbias.t372 Vbias.n2789 83.5719
R11509 Vbias.n4382 Vbias.n2799 83.5719
R11510 Vbias.t507 Vbias.n2799 83.5719
R11511 Vbias.n4401 Vbias.n4400 83.5719
R11512 Vbias.n4400 Vbias.t162 83.5719
R11513 Vbias.n4398 Vbias.n2785 83.5719
R11514 Vbias.n4398 Vbias.t372 83.5719
R11515 Vbias.n4371 Vbias.n4370 83.5719
R11516 Vbias.n4370 Vbias.t507 83.5719
R11517 Vbias.n4296 Vbias.n4295 83.5719
R11518 Vbias.t502 Vbias.n4296 83.5719
R11519 Vbias.n4292 Vbias.n4291 83.5719
R11520 Vbias.n4291 Vbias.t576 83.5719
R11521 Vbias.n4273 Vbias.n4272 83.5719
R11522 Vbias.t84 Vbias.n4273 83.5719
R11523 Vbias.n4298 Vbias.n4297 83.5719
R11524 Vbias.n4297 Vbias.t502 83.5719
R11525 Vbias.n4290 Vbias.n4289 83.5719
R11526 Vbias.t576 Vbias.n4290 83.5719
R11527 Vbias.n4269 Vbias.n2887 83.5719
R11528 Vbias.t84 Vbias.n2887 83.5719
R11529 Vbias.n4329 Vbias.n4328 83.5719
R11530 Vbias.t343 Vbias.n4329 83.5719
R11531 Vbias.n4325 Vbias.n4324 83.5719
R11532 Vbias.n4324 Vbias.t596 83.5719
R11533 Vbias.n4306 Vbias.n4305 83.5719
R11534 Vbias.t167 Vbias.n4306 83.5719
R11535 Vbias.n4331 Vbias.n4330 83.5719
R11536 Vbias.n4330 Vbias.t343 83.5719
R11537 Vbias.n4323 Vbias.n4322 83.5719
R11538 Vbias.t596 Vbias.n4323 83.5719
R11539 Vbias.n4302 Vbias.n2853 83.5719
R11540 Vbias.t167 Vbias.n2853 83.5719
R11541 Vbias.n2822 Vbias.n2820 83.5719
R11542 Vbias.n2820 Vbias.t637 83.5719
R11543 Vbias.n4335 Vbias.n2821 83.5719
R11544 Vbias.n2821 Vbias.t637 83.5719
R11545 Vbias.n2805 Vbias.n2803 83.5719
R11546 Vbias.n2803 Vbias.t466 83.5719
R11547 Vbias.n4340 Vbias.n4339 83.5719
R11548 Vbias.n4339 Vbias.t128 83.5719
R11549 Vbias.n4360 Vbias.n2804 83.5719
R11550 Vbias.n2804 Vbias.t466 83.5719
R11551 Vbias.n4357 Vbias.n2811 83.5719
R11552 Vbias.t128 Vbias.n2811 83.5719
R11553 Vbias.n2780 Vbias.n2778 83.5719
R11554 Vbias.n2778 Vbias.t162 83.5719
R11555 Vbias.n4397 Vbias.n4396 83.5719
R11556 Vbias.t372 Vbias.n4397 83.5719
R11557 Vbias.n4369 Vbias.n4368 83.5719
R11558 Vbias.t507 Vbias.n4369 83.5719
R11559 Vbias.n2781 Vbias.n2779 83.5719
R11560 Vbias.n2779 Vbias.t162 83.5719
R11561 Vbias.n4386 Vbias.n2791 83.5719
R11562 Vbias.t372 Vbias.n2791 83.5719
R11563 Vbias.n4382 Vbias.n2798 83.5719
R11564 Vbias.t507 Vbias.n2798 83.5719
R11565 Vbias.n5638 Vbias.n5553 83.1314
R11566 Vbias.n5877 Vbias.n1674 83.1314
R11567 Vbias.n8076 Vbias.n6 73.9214
R11568 Vbias.n4685 Vbias.n2772 73.9214
R11569 Vbias.n7788 Vbias.n7787 73.1255
R11570 Vbias.n7789 Vbias.n7788 73.1255
R11571 Vbias.n611 Vbias.n610 73.1255
R11572 Vbias.n610 Vbias.n609 73.1255
R11573 Vbias.n618 Vbias.n603 73.1255
R11574 Vbias.n619 Vbias.n618 73.1255
R11575 Vbias.n7780 Vbias.n7779 73.1255
R11576 Vbias.n7779 Vbias.n7778 73.1255
R11577 Vbias.n7776 Vbias.n7775 73.1255
R11578 Vbias.n7777 Vbias.n7776 73.1255
R11579 Vbias.n632 Vbias.n623 73.1255
R11580 Vbias.n633 Vbias.n632 73.1255
R11581 Vbias.n635 Vbias.n626 73.1255
R11582 Vbias.n635 Vbias.n634 73.1255
R11583 Vbias.n641 Vbias.n628 73.1255
R11584 Vbias.n642 Vbias.n641 73.1255
R11585 Vbias.n7767 Vbias.n7766 73.1255
R11586 Vbias.n7766 Vbias.n7765 73.1255
R11587 Vbias.n7763 Vbias.n7762 73.1255
R11588 Vbias.n7764 Vbias.n7763 73.1255
R11589 Vbias.n658 Vbias.n657 73.1255
R11590 Vbias.n657 Vbias.n656 73.1255
R11591 Vbias.n665 Vbias.n650 73.1255
R11592 Vbias.n666 Vbias.n665 73.1255
R11593 Vbias.n7755 Vbias.n7754 73.1255
R11594 Vbias.n7754 Vbias.n7753 73.1255
R11595 Vbias.n7792 Vbias.n7791 73.1255
R11596 Vbias.n7791 Vbias.n7790 73.1255
R11597 Vbias.n594 Vbias.n579 73.1255
R11598 Vbias.n595 Vbias.n594 73.1255
R11599 Vbias.n587 Vbias.n586 73.1255
R11600 Vbias.n586 Vbias.n585 73.1255
R11601 Vbias.n7800 Vbias.n7799 73.1255
R11602 Vbias.n7801 Vbias.n7800 73.1255
R11603 Vbias.n7857 Vbias.n7856 73.1255
R11604 Vbias.n7858 Vbias.n7857 73.1255
R11605 Vbias.n497 Vbias.n496 73.1255
R11606 Vbias.n496 Vbias.n495 73.1255
R11607 Vbias.n504 Vbias.n489 73.1255
R11608 Vbias.n505 Vbias.n504 73.1255
R11609 Vbias.n7849 Vbias.n7848 73.1255
R11610 Vbias.n7848 Vbias.n7847 73.1255
R11611 Vbias.n7845 Vbias.n7844 73.1255
R11612 Vbias.n7846 Vbias.n7845 73.1255
R11613 Vbias.n518 Vbias.n509 73.1255
R11614 Vbias.n519 Vbias.n518 73.1255
R11615 Vbias.n521 Vbias.n512 73.1255
R11616 Vbias.n521 Vbias.n520 73.1255
R11617 Vbias.n527 Vbias.n514 73.1255
R11618 Vbias.n528 Vbias.n527 73.1255
R11619 Vbias.n7836 Vbias.n7835 73.1255
R11620 Vbias.n7835 Vbias.n7834 73.1255
R11621 Vbias.n7832 Vbias.n7831 73.1255
R11622 Vbias.n7833 Vbias.n7832 73.1255
R11623 Vbias.n544 Vbias.n543 73.1255
R11624 Vbias.n543 Vbias.n542 73.1255
R11625 Vbias.n551 Vbias.n536 73.1255
R11626 Vbias.n552 Vbias.n551 73.1255
R11627 Vbias.n7824 Vbias.n7823 73.1255
R11628 Vbias.n7823 Vbias.n7822 73.1255
R11629 Vbias.n7861 Vbias.n7860 73.1255
R11630 Vbias.n7860 Vbias.n7859 73.1255
R11631 Vbias.n480 Vbias.n465 73.1255
R11632 Vbias.n481 Vbias.n480 73.1255
R11633 Vbias.n473 Vbias.n472 73.1255
R11634 Vbias.n472 Vbias.n471 73.1255
R11635 Vbias.n7869 Vbias.n7868 73.1255
R11636 Vbias.n7870 Vbias.n7869 73.1255
R11637 Vbias.n7923 Vbias.n7922 73.1255
R11638 Vbias.n7924 Vbias.n7923 73.1255
R11639 Vbias.n391 Vbias.n390 73.1255
R11640 Vbias.n390 Vbias.n389 73.1255
R11641 Vbias.n398 Vbias.n383 73.1255
R11642 Vbias.n399 Vbias.n398 73.1255
R11643 Vbias.n7915 Vbias.n7914 73.1255
R11644 Vbias.n7914 Vbias.n7913 73.1255
R11645 Vbias.n7911 Vbias.n7910 73.1255
R11646 Vbias.n7912 Vbias.n7911 73.1255
R11647 Vbias.n412 Vbias.n403 73.1255
R11648 Vbias.n413 Vbias.n412 73.1255
R11649 Vbias.n415 Vbias.n406 73.1255
R11650 Vbias.n415 Vbias.n414 73.1255
R11651 Vbias.n421 Vbias.n408 73.1255
R11652 Vbias.n422 Vbias.n421 73.1255
R11653 Vbias.n7902 Vbias.n7901 73.1255
R11654 Vbias.n7901 Vbias.n7900 73.1255
R11655 Vbias.n7898 Vbias.n7897 73.1255
R11656 Vbias.n7899 Vbias.n7898 73.1255
R11657 Vbias.n438 Vbias.n437 73.1255
R11658 Vbias.n437 Vbias.n436 73.1255
R11659 Vbias.n445 Vbias.n430 73.1255
R11660 Vbias.n446 Vbias.n445 73.1255
R11661 Vbias.n7890 Vbias.n7889 73.1255
R11662 Vbias.n7889 Vbias.n7888 73.1255
R11663 Vbias.n7927 Vbias.n7926 73.1255
R11664 Vbias.n7926 Vbias.n7925 73.1255
R11665 Vbias.n374 Vbias.n359 73.1255
R11666 Vbias.n375 Vbias.n374 73.1255
R11667 Vbias.n367 Vbias.n366 73.1255
R11668 Vbias.n366 Vbias.n365 73.1255
R11669 Vbias.n7935 Vbias.n7934 73.1255
R11670 Vbias.n7936 Vbias.n7935 73.1255
R11671 Vbias.n226 Vbias.n221 73.1255
R11672 Vbias.n223 Vbias.n221 73.1255
R11673 Vbias.n227 Vbias.n220 73.1255
R11674 Vbias.n224 Vbias.n220 73.1255
R11675 Vbias.n283 Vbias.n282 73.1255
R11676 Vbias.n284 Vbias.n283 73.1255
R11677 Vbias.n289 Vbias.n288 73.1255
R11678 Vbias.n288 Vbias.n287 73.1255
R11679 Vbias.n285 Vbias.n211 73.1255
R11680 Vbias.n286 Vbias.n285 73.1255
R11681 Vbias.n297 Vbias.n296 73.1255
R11682 Vbias.n298 Vbias.n297 73.1255
R11683 Vbias.n300 Vbias.n205 73.1255
R11684 Vbias.n300 Vbias.n299 73.1255
R11685 Vbias.n305 Vbias.n304 73.1255
R11686 Vbias.n306 Vbias.n305 73.1255
R11687 Vbias.n309 Vbias.n308 73.1255
R11688 Vbias.n308 Vbias.n307 73.1255
R11689 Vbias.n193 Vbias.n188 73.1255
R11690 Vbias.n190 Vbias.n188 73.1255
R11691 Vbias.n194 Vbias.n187 73.1255
R11692 Vbias.n191 Vbias.n187 73.1255
R11693 Vbias.n322 Vbias.n321 73.1255
R11694 Vbias.n323 Vbias.n322 73.1255
R11695 Vbias.n352 Vbias.n351 73.1255
R11696 Vbias.n351 Vbias.n350 73.1255
R11697 Vbias.n270 Vbias.n269 73.1255
R11698 Vbias.n269 Vbias.n268 73.1255
R11699 Vbias.n266 Vbias.n265 73.1255
R11700 Vbias.n267 Vbias.n266 73.1255
R11701 Vbias.n247 Vbias.n239 73.1255
R11702 Vbias.n242 Vbias.n239 73.1255
R11703 Vbias.n244 Vbias.n240 73.1255
R11704 Vbias.n240 Vbias.n86 73.1255
R11705 Vbias.n1175 Vbias.n1169 73.1255
R11706 Vbias.n1175 Vbias.n1152 73.1255
R11707 Vbias.n1270 Vbias.n1269 73.1255
R11708 Vbias.n1269 Vbias.n1268 73.1255
R11709 Vbias.n1260 Vbias.n1180 73.1255
R11710 Vbias.n1180 Vbias.n1178 73.1255
R11711 Vbias.n1262 Vbias.n1181 73.1255
R11712 Vbias.n1256 Vbias.n1181 73.1255
R11713 Vbias.n1254 Vbias.n1253 73.1255
R11714 Vbias.n1255 Vbias.n1254 73.1255
R11715 Vbias.n1250 Vbias.n1249 73.1255
R11716 Vbias.n1249 Vbias.n1248 73.1255
R11717 Vbias.n1245 Vbias.n1192 73.1255
R11718 Vbias.n1192 Vbias.n1190 73.1255
R11719 Vbias.n1204 Vbias.n1197 73.1255
R11720 Vbias.n1204 Vbias.n1203 73.1255
R11721 Vbias.n1239 Vbias.n1238 73.1255
R11722 Vbias.n1238 Vbias.n1237 73.1255
R11723 Vbias.n1229 Vbias.n1209 73.1255
R11724 Vbias.n1209 Vbias.n1207 73.1255
R11725 Vbias.n1231 Vbias.n1210 73.1255
R11726 Vbias.n1225 Vbias.n1210 73.1255
R11727 Vbias.n1223 Vbias.n1222 73.1255
R11728 Vbias.n1224 Vbias.n1223 73.1255
R11729 Vbias.n1219 Vbias.n1218 73.1255
R11730 Vbias.n1218 Vbias.n1082 73.1255
R11731 Vbias.n7212 Vbias.n7211 73.1255
R11732 Vbias.n7211 Vbias.n7210 73.1255
R11733 Vbias.n7216 Vbias.n7215 73.1255
R11734 Vbias.n7217 Vbias.n7216 73.1255
R11735 Vbias.n7220 Vbias.n7219 73.1255
R11736 Vbias.n7219 Vbias.n7218 73.1255
R11737 Vbias.n7223 Vbias.n7222 73.1255
R11738 Vbias.n7224 Vbias.n7223 73.1255
R11739 Vbias.n1150 Vbias.n1149 73.1255
R11740 Vbias.n7123 Vbias.n1150 73.1255
R11741 Vbias.n1148 Vbias.n1147 73.1255
R11742 Vbias.n1147 Vbias.n1143 73.1255
R11743 Vbias.n7130 Vbias.n7129 73.1255
R11744 Vbias.n7129 Vbias.n1144 73.1255
R11745 Vbias.n7141 Vbias.n7140 73.1255
R11746 Vbias.n7142 Vbias.n7141 73.1255
R11747 Vbias.n1133 Vbias.n1132 73.1255
R11748 Vbias.n7143 Vbias.n1133 73.1255
R11749 Vbias.n7147 Vbias.n7146 73.1255
R11750 Vbias.n7146 Vbias.n7144 73.1255
R11751 Vbias.n7158 Vbias.n7157 73.1255
R11752 Vbias.n7159 Vbias.n7158 73.1255
R11753 Vbias.n7160 Vbias.n1124 73.1255
R11754 Vbias.n7161 Vbias.n7160 73.1255
R11755 Vbias.n7164 Vbias.n7163 73.1255
R11756 Vbias.n7163 Vbias.n7162 73.1255
R11757 Vbias.n1119 Vbias.n1114 73.1255
R11758 Vbias.n1116 Vbias.n1114 73.1255
R11759 Vbias.n1120 Vbias.n1113 73.1255
R11760 Vbias.n1117 Vbias.n1113 73.1255
R11761 Vbias.n7177 Vbias.n7176 73.1255
R11762 Vbias.n7178 Vbias.n7177 73.1255
R11763 Vbias.n7181 Vbias.n7180 73.1255
R11764 Vbias.n7180 Vbias.n7179 73.1255
R11765 Vbias.n1100 Vbias.n1095 73.1255
R11766 Vbias.n1097 Vbias.n1095 73.1255
R11767 Vbias.n1101 Vbias.n1094 73.1255
R11768 Vbias.n1098 Vbias.n1094 73.1255
R11769 Vbias.n7194 Vbias.n7193 73.1255
R11770 Vbias.n7195 Vbias.n7194 73.1255
R11771 Vbias.n7198 Vbias.n7197 73.1255
R11772 Vbias.n7197 Vbias.n1071 73.1255
R11773 Vbias.n6908 Vbias.n6902 73.1255
R11774 Vbias.n6908 Vbias.n1339 73.1255
R11775 Vbias.n7003 Vbias.n7002 73.1255
R11776 Vbias.n7002 Vbias.n7001 73.1255
R11777 Vbias.n6993 Vbias.n6913 73.1255
R11778 Vbias.n6913 Vbias.n6911 73.1255
R11779 Vbias.n6995 Vbias.n6914 73.1255
R11780 Vbias.n6989 Vbias.n6914 73.1255
R11781 Vbias.n6987 Vbias.n6986 73.1255
R11782 Vbias.n6988 Vbias.n6987 73.1255
R11783 Vbias.n6983 Vbias.n6982 73.1255
R11784 Vbias.n6982 Vbias.n6981 73.1255
R11785 Vbias.n6978 Vbias.n6925 73.1255
R11786 Vbias.n6925 Vbias.n6923 73.1255
R11787 Vbias.n6937 Vbias.n6930 73.1255
R11788 Vbias.n6937 Vbias.n6936 73.1255
R11789 Vbias.n6972 Vbias.n6971 73.1255
R11790 Vbias.n6971 Vbias.n6970 73.1255
R11791 Vbias.n6962 Vbias.n6942 73.1255
R11792 Vbias.n6942 Vbias.n6940 73.1255
R11793 Vbias.n6964 Vbias.n6943 73.1255
R11794 Vbias.n6958 Vbias.n6943 73.1255
R11795 Vbias.n6956 Vbias.n6955 73.1255
R11796 Vbias.n6957 Vbias.n6956 73.1255
R11797 Vbias.n6952 Vbias.n6951 73.1255
R11798 Vbias.n6951 Vbias.n1163 73.1255
R11799 Vbias.n7108 Vbias.n7107 73.1255
R11800 Vbias.n7107 Vbias.n7106 73.1255
R11801 Vbias.n7112 Vbias.n7111 73.1255
R11802 Vbias.n7113 Vbias.n7112 73.1255
R11803 Vbias.n7116 Vbias.n7115 73.1255
R11804 Vbias.n7115 Vbias.n7114 73.1255
R11805 Vbias.n7119 Vbias.n7118 73.1255
R11806 Vbias.n7120 Vbias.n7119 73.1255
R11807 Vbias.n1338 Vbias.n1337 73.1255
R11808 Vbias.n7017 Vbias.n1338 73.1255
R11809 Vbias.n1336 Vbias.n1335 73.1255
R11810 Vbias.n1335 Vbias.n1331 73.1255
R11811 Vbias.n7024 Vbias.n7023 73.1255
R11812 Vbias.n7023 Vbias.n1332 73.1255
R11813 Vbias.n7035 Vbias.n7034 73.1255
R11814 Vbias.n7036 Vbias.n7035 73.1255
R11815 Vbias.n1321 Vbias.n1320 73.1255
R11816 Vbias.n7037 Vbias.n1321 73.1255
R11817 Vbias.n7041 Vbias.n7040 73.1255
R11818 Vbias.n7040 Vbias.n7038 73.1255
R11819 Vbias.n7052 Vbias.n7051 73.1255
R11820 Vbias.n7053 Vbias.n7052 73.1255
R11821 Vbias.n7054 Vbias.n1312 73.1255
R11822 Vbias.n7055 Vbias.n7054 73.1255
R11823 Vbias.n7058 Vbias.n7057 73.1255
R11824 Vbias.n7057 Vbias.n7056 73.1255
R11825 Vbias.n1307 Vbias.n1301 73.1255
R11826 Vbias.n1303 Vbias.n1301 73.1255
R11827 Vbias.n1308 Vbias.n1300 73.1255
R11828 Vbias.n1304 Vbias.n1300 73.1255
R11829 Vbias.n7071 Vbias.n7070 73.1255
R11830 Vbias.n7072 Vbias.n7071 73.1255
R11831 Vbias.n7075 Vbias.n7074 73.1255
R11832 Vbias.n7074 Vbias.n7073 73.1255
R11833 Vbias.n1287 Vbias.n1282 73.1255
R11834 Vbias.n1284 Vbias.n1282 73.1255
R11835 Vbias.n1288 Vbias.n1281 73.1255
R11836 Vbias.n1285 Vbias.n1281 73.1255
R11837 Vbias.n7088 Vbias.n7087 73.1255
R11838 Vbias.n7089 Vbias.n7088 73.1255
R11839 Vbias.n7092 Vbias.n7091 73.1255
R11840 Vbias.n7091 Vbias.n1151 73.1255
R11841 Vbias.n1556 Vbias.n1399 73.1255
R11842 Vbias.n1557 Vbias.n1556 73.1255
R11843 Vbias.n6819 Vbias.n6818 73.1255
R11844 Vbias.n6818 Vbias.n1397 73.1255
R11845 Vbias.n6826 Vbias.n6825 73.1255
R11846 Vbias.n6825 Vbias.n1392 73.1255
R11847 Vbias.n1391 Vbias.n1389 73.1255
R11848 Vbias.n1393 Vbias.n1391 73.1255
R11849 Vbias.n1386 Vbias.n1385 73.1255
R11850 Vbias.n1385 Vbias.n1383 73.1255
R11851 Vbias.n6841 Vbias.n6840 73.1255
R11852 Vbias.n6840 Vbias.n6839 73.1255
R11853 Vbias.n6845 Vbias.n6844 73.1255
R11854 Vbias.n6846 Vbias.n6845 73.1255
R11855 Vbias.n1375 Vbias.n1374 73.1255
R11856 Vbias.n6847 Vbias.n1375 73.1255
R11857 Vbias.n6850 Vbias.n6849 73.1255
R11858 Vbias.n6849 Vbias.n1370 73.1255
R11859 Vbias.n6864 Vbias.n6863 73.1255
R11860 Vbias.n6863 Vbias.n6862 73.1255
R11861 Vbias.n6868 Vbias.n6867 73.1255
R11862 Vbias.n6869 Vbias.n6868 73.1255
R11863 Vbias.n1362 Vbias.n1361 73.1255
R11864 Vbias.n6870 Vbias.n1362 73.1255
R11865 Vbias.n6873 Vbias.n6872 73.1255
R11866 Vbias.n6872 Vbias.n1357 73.1255
R11867 Vbias.n6887 Vbias.n6886 73.1255
R11868 Vbias.n6886 Vbias.n6885 73.1255
R11869 Vbias.n6891 Vbias.n6890 73.1255
R11870 Vbias.n6892 Vbias.n6891 73.1255
R11871 Vbias.n1348 Vbias.n1346 73.1255
R11872 Vbias.n6893 Vbias.n1348 73.1255
R11873 Vbias.n1349 Vbias.n1347 73.1255
R11874 Vbias.n1349 Vbias.n1340 73.1255
R11875 Vbias.n6073 Vbias.n1402 73.1255
R11876 Vbias.n6074 Vbias.n6073 73.1255
R11877 Vbias.n6050 Vbias.n1404 73.1255
R11878 Vbias.n6051 Vbias.n6050 73.1255
R11879 Vbias.n6066 Vbias.n1406 73.1255
R11880 Vbias.n6067 Vbias.n6066 73.1255
R11881 Vbias.n6062 Vbias.n1408 73.1255
R11882 Vbias.n6062 Vbias.n6061 73.1255
R11883 Vbias.n6059 Vbias.n1410 73.1255
R11884 Vbias.n6060 Vbias.n6059 73.1255
R11885 Vbias.n6054 Vbias.n1412 73.1255
R11886 Vbias.n6054 Vbias.n6053 73.1255
R11887 Vbias.n6801 Vbias.n6800 73.1255
R11888 Vbias.n6800 Vbias.n6799 73.1255
R11889 Vbias.n6797 Vbias.n6796 73.1255
R11890 Vbias.n6798 Vbias.n6797 73.1255
R11891 Vbias.n6752 Vbias.n1419 73.1255
R11892 Vbias.n6753 Vbias.n6752 73.1255
R11893 Vbias.n6755 Vbias.n1422 73.1255
R11894 Vbias.n6755 Vbias.n6754 73.1255
R11895 Vbias.n6759 Vbias.n1424 73.1255
R11896 Vbias.n6760 Vbias.n6759 73.1255
R11897 Vbias.n6762 Vbias.n1426 73.1255
R11898 Vbias.n6763 Vbias.n6762 73.1255
R11899 Vbias.n6769 Vbias.n1428 73.1255
R11900 Vbias.n6770 Vbias.n6769 73.1255
R11901 Vbias.n1439 Vbias.n1429 73.1255
R11902 Vbias.n6771 Vbias.n1439 73.1255
R11903 Vbias.n1436 Vbias.n1431 73.1255
R11904 Vbias.n1436 Vbias.n1434 73.1255
R11905 Vbias.n6776 Vbias.n6775 73.1255
R11906 Vbias.n6775 Vbias.n1435 73.1255
R11907 Vbias.n7013 Vbias.n7012 73.1255
R11908 Vbias.n7014 Vbias.n7013 73.1255
R11909 Vbias.n1637 Vbias.n1610 73.1255
R11910 Vbias.n1638 Vbias.n1637 73.1255
R11911 Vbias.n5961 Vbias.n5960 73.1255
R11912 Vbias.n5960 Vbias.n1608 73.1255
R11913 Vbias.n5968 Vbias.n5967 73.1255
R11914 Vbias.n5967 Vbias.n1603 73.1255
R11915 Vbias.n1602 Vbias.n1600 73.1255
R11916 Vbias.n1604 Vbias.n1602 73.1255
R11917 Vbias.n1597 Vbias.n1596 73.1255
R11918 Vbias.n1596 Vbias.n1594 73.1255
R11919 Vbias.n5983 Vbias.n5982 73.1255
R11920 Vbias.n5982 Vbias.n5981 73.1255
R11921 Vbias.n5987 Vbias.n5986 73.1255
R11922 Vbias.n5988 Vbias.n5987 73.1255
R11923 Vbias.n1586 Vbias.n1585 73.1255
R11924 Vbias.n5989 Vbias.n1586 73.1255
R11925 Vbias.n5992 Vbias.n5991 73.1255
R11926 Vbias.n5991 Vbias.n1581 73.1255
R11927 Vbias.n6006 Vbias.n6005 73.1255
R11928 Vbias.n6005 Vbias.n6004 73.1255
R11929 Vbias.n6010 Vbias.n6009 73.1255
R11930 Vbias.n6011 Vbias.n6010 73.1255
R11931 Vbias.n1573 Vbias.n1572 73.1255
R11932 Vbias.n6012 Vbias.n1573 73.1255
R11933 Vbias.n6015 Vbias.n6014 73.1255
R11934 Vbias.n6014 Vbias.n1568 73.1255
R11935 Vbias.n6032 Vbias.n6031 73.1255
R11936 Vbias.n6031 Vbias.n6030 73.1255
R11937 Vbias.n6036 Vbias.n6035 73.1255
R11938 Vbias.n6037 Vbias.n6036 73.1255
R11939 Vbias.n6040 Vbias.n6039 73.1255
R11940 Vbias.n6039 Vbias.n6038 73.1255
R11941 Vbias.n6043 Vbias.n6042 73.1255
R11942 Vbias.n6044 Vbias.n6043 73.1255
R11943 Vbias.n1791 Vbias.n1544 73.1255
R11944 Vbias.n1791 Vbias.n1790 73.1255
R11945 Vbias.n1788 Vbias.n1546 73.1255
R11946 Vbias.n1789 Vbias.n1788 73.1255
R11947 Vbias.n1777 Vbias.n1548 73.1255
R11948 Vbias.n1777 Vbias.n1776 73.1255
R11949 Vbias.n1781 Vbias.n1550 73.1255
R11950 Vbias.n1781 Vbias.n1458 73.1255
R11951 Vbias.n6078 Vbias.n6077 73.1255
R11952 Vbias.n6077 Vbias.n6076 73.1255
R11953 Vbias.n1885 Vbias.n1883 73.1255
R11954 Vbias.n1885 Vbias.n1523 73.1255
R11955 Vbias.n1890 Vbias.n1889 73.1255
R11956 Vbias.n1889 Vbias.n1887 73.1255
R11957 Vbias.n1896 Vbias.n1894 73.1255
R11958 Vbias.n1894 Vbias.n1893 73.1255
R11959 Vbias.n1901 Vbias.n1895 73.1255
R11960 Vbias.n1895 Vbias.n1460 73.1255
R11961 Vbias.n1962 Vbias.n1961 73.1255
R11962 Vbias.n1962 Vbias.n1524 73.1255
R11963 Vbias.n1960 Vbias.n1959 73.1255
R11964 Vbias.n1959 Vbias.n1955 73.1255
R11965 Vbias.n1976 Vbias.n1975 73.1255
R11966 Vbias.n1975 Vbias.n1956 73.1255
R11967 Vbias.n1968 Vbias.n1967 73.1255
R11968 Vbias.n1968 Vbias.n1461 73.1255
R11969 Vbias.n1522 Vbias.n1521 73.1255
R11970 Vbias.n6102 Vbias.n1522 73.1255
R11971 Vbias.n1520 Vbias.n1519 73.1255
R11972 Vbias.n1519 Vbias.n1515 73.1255
R11973 Vbias.n6116 Vbias.n6115 73.1255
R11974 Vbias.n6115 Vbias.n1516 73.1255
R11975 Vbias.n6108 Vbias.n6107 73.1255
R11976 Vbias.n6108 Vbias.n1462 73.1255
R11977 Vbias.n1996 Vbias.n1992 73.1255
R11978 Vbias.n1992 Vbias.n1525 73.1255
R11979 Vbias.n1999 Vbias.n1991 73.1255
R11980 Vbias.n1994 Vbias.n1991 73.1255
R11981 Vbias.n2009 Vbias.n2008 73.1255
R11982 Vbias.n2010 Vbias.n2009 73.1255
R11983 Vbias.n2013 Vbias.n2012 73.1255
R11984 Vbias.n2012 Vbias.n1463 73.1255
R11985 Vbias.n1928 Vbias.n1927 73.1255
R11986 Vbias.n1928 Vbias.n1526 73.1255
R11987 Vbias.n1926 Vbias.n1925 73.1255
R11988 Vbias.n1925 Vbias.n1921 73.1255
R11989 Vbias.n1942 Vbias.n1941 73.1255
R11990 Vbias.n1941 Vbias.n1922 73.1255
R11991 Vbias.n1934 Vbias.n1933 73.1255
R11992 Vbias.n1934 Vbias.n1464 73.1255
R11993 Vbias.n1860 Vbias.n1859 73.1255
R11994 Vbias.n1860 Vbias.n1527 73.1255
R11995 Vbias.n1858 Vbias.n1857 73.1255
R11996 Vbias.n1857 Vbias.n1853 73.1255
R11997 Vbias.n1866 Vbias.n1865 73.1255
R11998 Vbias.n1865 Vbias.n1854 73.1255
R11999 Vbias.n1868 Vbias.n1867 73.1255
R12000 Vbias.n1868 Vbias.n1465 73.1255
R12001 Vbias.n1807 Vbias.n1803 73.1255
R12002 Vbias.n1803 Vbias.n1531 73.1255
R12003 Vbias.n1802 Vbias.n1801 73.1255
R12004 Vbias.n1804 Vbias.n1802 73.1255
R12005 Vbias.n1766 Vbias.n1762 73.1255
R12006 Vbias.n1767 Vbias.n1766 73.1255
R12007 Vbias.n1758 Vbias.n1756 73.1255
R12008 Vbias.n1760 Vbias.n1758 73.1255
R12009 Vbias.n1805 Vbias.n1536 73.1255
R12010 Vbias.n1806 Vbias.n1805 73.1255
R12011 Vbias.n1768 Vbias.n1538 73.1255
R12012 Vbias.n1768 Vbias.n1765 73.1255
R12013 Vbias.n1770 Vbias.n1540 73.1255
R12014 Vbias.n1770 Vbias.n1759 73.1255
R12015 Vbias.n1774 Vbias.n1542 73.1255
R12016 Vbias.n1774 Vbias.n1466 73.1255
R12017 Vbias.n1634 Vbias.n1613 73.1255
R12018 Vbias.n5920 Vbias.n1634 73.1255
R12019 Vbias.n1632 Vbias.n1615 73.1255
R12020 Vbias.n1632 Vbias.n1630 73.1255
R12021 Vbias.n5928 Vbias.n1617 73.1255
R12022 Vbias.n5929 Vbias.n5928 73.1255
R12023 Vbias.n5931 Vbias.n1619 73.1255
R12024 Vbias.n5932 Vbias.n5931 73.1255
R12025 Vbias.n5934 Vbias.n1622 73.1255
R12026 Vbias.n5934 Vbias.n5933 73.1255
R12027 Vbias.n5939 Vbias.n1624 73.1255
R12028 Vbias.n5940 Vbias.n5939 73.1255
R12029 Vbias.n5943 Vbias.n5942 73.1255
R12030 Vbias.n5942 Vbias.n1532 73.1255
R12031 Vbias.n6099 Vbias.n6098 73.1255
R12032 Vbias.n6100 Vbias.n6099 73.1255
R12033 Vbias.n5279 Vbias.n5272 73.1255
R12034 Vbias.n5279 Vbias.n5278 73.1255
R12035 Vbias.n5411 Vbias.n5410 73.1255
R12036 Vbias.n5410 Vbias.n5409 73.1255
R12037 Vbias.n5401 Vbias.n5284 73.1255
R12038 Vbias.n5284 Vbias.n5282 73.1255
R12039 Vbias.n5403 Vbias.n5285 73.1255
R12040 Vbias.n5397 Vbias.n5285 73.1255
R12041 Vbias.n5395 Vbias.n5394 73.1255
R12042 Vbias.n5396 Vbias.n5395 73.1255
R12043 Vbias.n5391 Vbias.n5390 73.1255
R12044 Vbias.n5390 Vbias.n5389 73.1255
R12045 Vbias.n5386 Vbias.n5296 73.1255
R12046 Vbias.n5296 Vbias.n5294 73.1255
R12047 Vbias.n5308 Vbias.n5301 73.1255
R12048 Vbias.n5308 Vbias.n5307 73.1255
R12049 Vbias.n5380 Vbias.n5379 73.1255
R12050 Vbias.n5379 Vbias.n5378 73.1255
R12051 Vbias.n5370 Vbias.n5313 73.1255
R12052 Vbias.n5313 Vbias.n5311 73.1255
R12053 Vbias.n5372 Vbias.n5314 73.1255
R12054 Vbias.n5366 Vbias.n5314 73.1255
R12055 Vbias.n5364 Vbias.n5363 73.1255
R12056 Vbias.n5365 Vbias.n5364 73.1255
R12057 Vbias.n5325 Vbias.n5319 73.1255
R12058 Vbias.n5325 Vbias.n5323 73.1255
R12059 Vbias.n5330 Vbias.n5329 73.1255
R12060 Vbias.n5329 Vbias.n5324 73.1255
R12061 Vbias.n5337 Vbias.n5336 73.1255
R12062 Vbias.n5350 Vbias.n5337 73.1255
R12063 Vbias.n5348 Vbias.n5347 73.1255
R12064 Vbias.n5349 Vbias.n5348 73.1255
R12065 Vbias.n5345 Vbias.n5344 73.1255
R12066 Vbias.n5344 Vbias.n1639 73.1255
R12067 Vbias.n5483 Vbias.n5482 73.1255
R12068 Vbias.n5484 Vbias.n5483 73.1255
R12069 Vbias.n5427 Vbias.n5426 73.1255
R12070 Vbias.n5426 Vbias.n5425 73.1255
R12071 Vbias.n5434 Vbias.n5419 73.1255
R12072 Vbias.n5435 Vbias.n5434 73.1255
R12073 Vbias.n5475 Vbias.n5474 73.1255
R12074 Vbias.n5474 Vbias.n5473 73.1255
R12075 Vbias.n5471 Vbias.n5470 73.1255
R12076 Vbias.n5472 Vbias.n5471 73.1255
R12077 Vbias.n5449 Vbias.n5448 73.1255
R12078 Vbias.n5450 Vbias.n5449 73.1255
R12079 Vbias.n5465 Vbias.n5464 73.1255
R12080 Vbias.n5464 Vbias.n5463 73.1255
R12081 Vbias.n5461 Vbias.n5460 73.1255
R12082 Vbias.n5462 Vbias.n5461 73.1255
R12083 Vbias.n5456 Vbias.n5455 73.1255
R12084 Vbias.n5455 Vbias.n5454 73.1255
R12085 Vbias.n1671 Vbias.n1670 73.1255
R12086 Vbias.n1672 Vbias.n1671 73.1255
R12087 Vbias.n1669 Vbias.n1668 73.1255
R12088 Vbias.n1668 Vbias.n1664 73.1255
R12089 Vbias.n5885 Vbias.n5884 73.1255
R12090 Vbias.n5884 Vbias.n1665 73.1255
R12091 Vbias.n5896 Vbias.n5895 73.1255
R12092 Vbias.n5897 Vbias.n5896 73.1255
R12093 Vbias.n1655 Vbias.n1654 73.1255
R12094 Vbias.n5898 Vbias.n1655 73.1255
R12095 Vbias.n1653 Vbias.n1652 73.1255
R12096 Vbias.n1652 Vbias.n1648 73.1255
R12097 Vbias.n5905 Vbias.n5904 73.1255
R12098 Vbias.n5904 Vbias.n1649 73.1255
R12099 Vbias.n5916 Vbias.n5915 73.1255
R12100 Vbias.n5917 Vbias.n5916 73.1255
R12101 Vbias.n2369 Vbias.n2347 73.1255
R12102 Vbias.n2370 Vbias.n2369 73.1255
R12103 Vbias.n5188 Vbias.n5187 73.1255
R12104 Vbias.n5187 Vbias.n2345 73.1255
R12105 Vbias.n5195 Vbias.n5194 73.1255
R12106 Vbias.n5194 Vbias.n2340 73.1255
R12107 Vbias.n2339 Vbias.n2337 73.1255
R12108 Vbias.n2341 Vbias.n2339 73.1255
R12109 Vbias.n2334 Vbias.n2333 73.1255
R12110 Vbias.n2333 Vbias.n2331 73.1255
R12111 Vbias.n5210 Vbias.n5209 73.1255
R12112 Vbias.n5209 Vbias.n5208 73.1255
R12113 Vbias.n5214 Vbias.n5213 73.1255
R12114 Vbias.n5215 Vbias.n5214 73.1255
R12115 Vbias.n2323 Vbias.n2322 73.1255
R12116 Vbias.n5216 Vbias.n2323 73.1255
R12117 Vbias.n5219 Vbias.n5218 73.1255
R12118 Vbias.n5218 Vbias.n2318 73.1255
R12119 Vbias.n5233 Vbias.n5232 73.1255
R12120 Vbias.n5232 Vbias.n5231 73.1255
R12121 Vbias.n5237 Vbias.n5236 73.1255
R12122 Vbias.n5238 Vbias.n5237 73.1255
R12123 Vbias.n2310 Vbias.n2309 73.1255
R12124 Vbias.n5239 Vbias.n2310 73.1255
R12125 Vbias.n5242 Vbias.n5241 73.1255
R12126 Vbias.n5241 Vbias.n2305 73.1255
R12127 Vbias.n5256 Vbias.n5255 73.1255
R12128 Vbias.n5255 Vbias.n5254 73.1255
R12129 Vbias.n5260 Vbias.n5259 73.1255
R12130 Vbias.n5261 Vbias.n5260 73.1255
R12131 Vbias.n2296 Vbias.n2294 73.1255
R12132 Vbias.n5262 Vbias.n2296 73.1255
R12133 Vbias.n2297 Vbias.n2295 73.1255
R12134 Vbias.n5263 Vbias.n2297 73.1255
R12135 Vbias.n5124 Vbias.n2350 73.1255
R12136 Vbias.n5124 Vbias.n5123 73.1255
R12137 Vbias.n5128 Vbias.n2352 73.1255
R12138 Vbias.n5129 Vbias.n5128 73.1255
R12139 Vbias.n5131 Vbias.n2354 73.1255
R12140 Vbias.n5132 Vbias.n5131 73.1255
R12141 Vbias.n5138 Vbias.n2356 73.1255
R12142 Vbias.n5139 Vbias.n5138 73.1255
R12143 Vbias.n5141 Vbias.n2358 73.1255
R12144 Vbias.n5141 Vbias.n5140 73.1255
R12145 Vbias.n5147 Vbias.n2360 73.1255
R12146 Vbias.n5148 Vbias.n5147 73.1255
R12147 Vbias.n5170 Vbias.n5169 73.1255
R12148 Vbias.n5169 Vbias.n5168 73.1255
R12149 Vbias.n5166 Vbias.n5165 73.1255
R12150 Vbias.n5167 Vbias.n5166 73.1255
R12151 Vbias.n5160 Vbias.n5159 73.1255
R12152 Vbias.n5159 Vbias.n5158 73.1255
R12153 Vbias.n5156 Vbias.n5155 73.1255
R12154 Vbias.n5157 Vbias.n5156 73.1255
R12155 Vbias.n5507 Vbias.n5506 73.1255
R12156 Vbias.n5508 Vbias.n5507 73.1255
R12157 Vbias.n2263 Vbias.n2262 73.1255
R12158 Vbias.n2264 Vbias.n2263 73.1255
R12159 Vbias.n5500 Vbias.n5499 73.1255
R12160 Vbias.n5499 Vbias.n5498 73.1255
R12161 Vbias.n5496 Vbias.n5495 73.1255
R12162 Vbias.n5497 Vbias.n5496 73.1255
R12163 Vbias.n2279 Vbias.n2278 73.1255
R12164 Vbias.n2278 Vbias.n2277 73.1255
R12165 Vbias.n2286 Vbias.n2271 73.1255
R12166 Vbias.n2287 Vbias.n2286 73.1255
R12167 Vbias.n5488 Vbias.n5487 73.1255
R12168 Vbias.n5487 Vbias.n5486 73.1255
R12169 Vbias.n2447 Vbias.n2440 73.1255
R12170 Vbias.n2447 Vbias.n2446 73.1255
R12171 Vbias.n2579 Vbias.n2578 73.1255
R12172 Vbias.n2578 Vbias.n2577 73.1255
R12173 Vbias.n2569 Vbias.n2452 73.1255
R12174 Vbias.n2452 Vbias.n2450 73.1255
R12175 Vbias.n2571 Vbias.n2453 73.1255
R12176 Vbias.n2565 Vbias.n2453 73.1255
R12177 Vbias.n2563 Vbias.n2562 73.1255
R12178 Vbias.n2564 Vbias.n2563 73.1255
R12179 Vbias.n2559 Vbias.n2558 73.1255
R12180 Vbias.n2558 Vbias.n2557 73.1255
R12181 Vbias.n2554 Vbias.n2464 73.1255
R12182 Vbias.n2464 Vbias.n2462 73.1255
R12183 Vbias.n2476 Vbias.n2469 73.1255
R12184 Vbias.n2476 Vbias.n2475 73.1255
R12185 Vbias.n2548 Vbias.n2547 73.1255
R12186 Vbias.n2547 Vbias.n2546 73.1255
R12187 Vbias.n2538 Vbias.n2481 73.1255
R12188 Vbias.n2481 Vbias.n2479 73.1255
R12189 Vbias.n2540 Vbias.n2482 73.1255
R12190 Vbias.n2534 Vbias.n2482 73.1255
R12191 Vbias.n2532 Vbias.n2531 73.1255
R12192 Vbias.n2533 Vbias.n2532 73.1255
R12193 Vbias.n2493 Vbias.n2487 73.1255
R12194 Vbias.n2493 Vbias.n2491 73.1255
R12195 Vbias.n2498 Vbias.n2497 73.1255
R12196 Vbias.n2497 Vbias.n2492 73.1255
R12197 Vbias.n2505 Vbias.n2504 73.1255
R12198 Vbias.n2518 Vbias.n2505 73.1255
R12199 Vbias.n2516 Vbias.n2515 73.1255
R12200 Vbias.n2517 Vbias.n2516 73.1255
R12201 Vbias.n2513 Vbias.n2512 73.1255
R12202 Vbias.n2512 Vbias.n2371 73.1255
R12203 Vbias.n5059 Vbias.n2414 73.1255
R12204 Vbias.n5059 Vbias.n5058 73.1255
R12205 Vbias.n5064 Vbias.n5063 73.1255
R12206 Vbias.n5065 Vbias.n5064 73.1255
R12207 Vbias.n5070 Vbias.n5069 73.1255
R12208 Vbias.n5069 Vbias.n5068 73.1255
R12209 Vbias.n5066 Vbias.n2406 73.1255
R12210 Vbias.n5067 Vbias.n5066 73.1255
R12211 Vbias.n5078 Vbias.n5077 73.1255
R12212 Vbias.n5079 Vbias.n5078 73.1255
R12213 Vbias.n5081 Vbias.n2402 73.1255
R12214 Vbias.n5081 Vbias.n5080 73.1255
R12215 Vbias.n2401 Vbias.n2400 73.1255
R12216 Vbias.n2400 Vbias.n2396 73.1255
R12217 Vbias.n5088 Vbias.n5087 73.1255
R12218 Vbias.n5087 Vbias.n2397 73.1255
R12219 Vbias.n5099 Vbias.n5098 73.1255
R12220 Vbias.n5100 Vbias.n5099 73.1255
R12221 Vbias.n2387 Vbias.n2386 73.1255
R12222 Vbias.n5101 Vbias.n2387 73.1255
R12223 Vbias.n2385 Vbias.n2384 73.1255
R12224 Vbias.n2384 Vbias.n2380 73.1255
R12225 Vbias.n5108 Vbias.n5107 73.1255
R12226 Vbias.n5107 Vbias.n2381 73.1255
R12227 Vbias.n5119 Vbias.n5118 73.1255
R12228 Vbias.n5120 Vbias.n5119 73.1255
R12229 Vbias.n5056 Vbias.n5055 73.1255
R12230 Vbias.n5057 Vbias.n5056 73.1255
R12231 Vbias.n5045 Vbias.n5044 73.1255
R12232 Vbias.n5044 Vbias.n2426 73.1255
R12233 Vbias.n2430 Vbias.n2429 73.1255
R12234 Vbias.n2429 Vbias.n2425 73.1255
R12235 Vbias.n2432 Vbias.n2431 73.1255
R12236 Vbias.n5038 Vbias.n2432 73.1255
R12237 Vbias.n4105 Vbias.n4103 73.1255
R12238 Vbias.n4105 Vbias.n6 73.1255
R12239 Vbias.n4106 Vbias.n4104 73.1255
R12240 Vbias.n4107 Vbias.n4106 73.1255
R12241 Vbias.n4117 Vbias.n4116 73.1255
R12242 Vbias.n4116 Vbias.n3985 73.1255
R12243 Vbias.n4098 Vbias.n4097 73.1255
R12244 Vbias.n4097 Vbias.n3988 73.1255
R12245 Vbias.n4094 Vbias.n4093 73.1255
R12246 Vbias.n4093 Vbias.n3996 73.1255
R12247 Vbias.n4123 Vbias.n4005 73.1255
R12248 Vbias.n4235 Vbias.n4005 73.1255
R12249 Vbias.n4086 Vbias.n4006 73.1255
R12250 Vbias.n4234 Vbias.n4006 73.1255
R12251 Vbias.n4131 Vbias.n4085 73.1255
R12252 Vbias.n4131 Vbias.n4016 73.1255
R12253 Vbias.n4084 Vbias.n4083 73.1255
R12254 Vbias.n4083 Vbias.n4019 73.1255
R12255 Vbias.n4139 Vbias.n4031 73.1255
R12256 Vbias.n4219 Vbias.n4031 73.1255
R12257 Vbias.n4156 Vbias.n4146 73.1255
R12258 Vbias.n4156 Vbias.n4155 73.1255
R12259 Vbias.n4145 Vbias.n4044 73.1255
R12260 Vbias.n4207 Vbias.n4044 73.1255
R12261 Vbias.n4162 Vbias.n4047 73.1255
R12262 Vbias.n4201 Vbias.n4047 73.1255
R12263 Vbias.n4168 Vbias.n4048 73.1255
R12264 Vbias.n4200 Vbias.n4048 73.1255
R12265 Vbias.n4174 Vbias.n4167 73.1255
R12266 Vbias.n4174 Vbias.n4058 73.1255
R12267 Vbias.n4077 Vbias.n4076 73.1255
R12268 Vbias.n4076 Vbias.n4061 73.1255
R12269 Vbias.n4183 Vbias.n4073 73.1255
R12270 Vbias.n4073 Vbias.n2772 73.1255
R12271 Vbias.n3983 Vbias.n3981 73.1255
R12272 Vbias.n3985 Vbias.n3983 73.1255
R12273 Vbias.n3991 Vbias.n3990 73.1255
R12274 Vbias.n3990 Vbias.n3988 73.1255
R12275 Vbias.n3999 Vbias.n3998 73.1255
R12276 Vbias.n3998 Vbias.n3996 73.1255
R12277 Vbias.n4002 Vbias.n4001 73.1255
R12278 Vbias.n4235 Vbias.n4002 73.1255
R12279 Vbias.n4233 Vbias.n4232 73.1255
R12280 Vbias.n4234 Vbias.n4233 73.1255
R12281 Vbias.n4023 Vbias.n4022 73.1255
R12282 Vbias.n4022 Vbias.n4016 73.1255
R12283 Vbias.n4026 Vbias.n4025 73.1255
R12284 Vbias.n4025 Vbias.n4019 73.1255
R12285 Vbias.n4028 Vbias.n4027 73.1255
R12286 Vbias.n4219 Vbias.n4028 73.1255
R12287 Vbias.n4217 Vbias.n4216 73.1255
R12288 Vbias.n4218 Vbias.n4217 73.1255
R12289 Vbias.n4150 Vbias.n4035 73.1255
R12290 Vbias.n4151 Vbias.n4150 73.1255
R12291 Vbias.n4154 Vbias.n4038 73.1255
R12292 Vbias.n4155 Vbias.n4154 73.1255
R12293 Vbias.n4209 Vbias.n4208 73.1255
R12294 Vbias.n4208 Vbias.n4207 73.1255
R12295 Vbias.n4204 Vbias.n4203 73.1255
R12296 Vbias.n4203 Vbias.n4201 73.1255
R12297 Vbias.n4199 Vbias.n4198 73.1255
R12298 Vbias.n4200 Vbias.n4199 73.1255
R12299 Vbias.n4065 Vbias.n4064 73.1255
R12300 Vbias.n4064 Vbias.n4058 73.1255
R12301 Vbias.n4068 Vbias.n4067 73.1255
R12302 Vbias.n4067 Vbias.n4061 73.1255
R12303 Vbias.n4070 Vbias.n4069 73.1255
R12304 Vbias.n4070 Vbias.n2772 73.1255
R12305 Vbias.n3443 Vbias.n3441 73.1255
R12306 Vbias.n3443 Vbias.n7 73.1255
R12307 Vbias.n3444 Vbias.n3442 73.1255
R12308 Vbias.n3701 Vbias.n3444 73.1255
R12309 Vbias.n3449 Vbias.n3445 73.1255
R12310 Vbias.n3700 Vbias.n3445 73.1255
R12311 Vbias.n3669 Vbias.n3667 73.1255
R12312 Vbias.n3669 Vbias.n3459 73.1255
R12313 Vbias.n3679 Vbias.n3678 73.1255
R12314 Vbias.n3678 Vbias.n3461 73.1255
R12315 Vbias.n3683 Vbias.n3682 73.1255
R12316 Vbias.n3682 Vbias.n3663 73.1255
R12317 Vbias.n3478 Vbias.n3474 73.1255
R12318 Vbias.n3662 Vbias.n3474 73.1255
R12319 Vbias.n3631 Vbias.n3629 73.1255
R12320 Vbias.n3631 Vbias.n3488 73.1255
R12321 Vbias.n3641 Vbias.n3640 73.1255
R12322 Vbias.n3640 Vbias.n3490 73.1255
R12323 Vbias.n3645 Vbias.n3644 73.1255
R12324 Vbias.n3644 Vbias.n3625 73.1255
R12325 Vbias.n3599 Vbias.n3591 73.1255
R12326 Vbias.n3599 Vbias.n3598 73.1255
R12327 Vbias.n3590 Vbias.n3517 73.1255
R12328 Vbias.n3612 Vbias.n3517 73.1255
R12329 Vbias.n3606 Vbias.n3605 73.1255
R12330 Vbias.n3605 Vbias.n3587 73.1255
R12331 Vbias.n3525 Vbias.n3521 73.1255
R12332 Vbias.n3586 Vbias.n3521 73.1255
R12333 Vbias.n3555 Vbias.n3553 73.1255
R12334 Vbias.n3555 Vbias.n3535 73.1255
R12335 Vbias.n3565 Vbias.n3564 73.1255
R12336 Vbias.n3564 Vbias.n3537 73.1255
R12337 Vbias.n3569 Vbias.n3568 73.1255
R12338 Vbias.n3568 Vbias.n2773 73.1255
R12339 Vbias.n3699 Vbias.n3698 73.1255
R12340 Vbias.n3700 Vbias.n3699 73.1255
R12341 Vbias.n3466 Vbias.n3465 73.1255
R12342 Vbias.n3465 Vbias.n3459 73.1255
R12343 Vbias.n3469 Vbias.n3468 73.1255
R12344 Vbias.n3468 Vbias.n3461 73.1255
R12345 Vbias.n3471 Vbias.n3470 73.1255
R12346 Vbias.n3663 Vbias.n3471 73.1255
R12347 Vbias.n3661 Vbias.n3660 73.1255
R12348 Vbias.n3662 Vbias.n3661 73.1255
R12349 Vbias.n3495 Vbias.n3494 73.1255
R12350 Vbias.n3494 Vbias.n3488 73.1255
R12351 Vbias.n3498 Vbias.n3497 73.1255
R12352 Vbias.n3497 Vbias.n3490 73.1255
R12353 Vbias.n3500 Vbias.n3499 73.1255
R12354 Vbias.n3625 Vbias.n3500 73.1255
R12355 Vbias.n3623 Vbias.n3622 73.1255
R12356 Vbias.n3624 Vbias.n3623 73.1255
R12357 Vbias.n3592 Vbias.n3506 73.1255
R12358 Vbias.n3593 Vbias.n3592 73.1255
R12359 Vbias.n3597 Vbias.n3596 73.1255
R12360 Vbias.n3598 Vbias.n3597 73.1255
R12361 Vbias.n3614 Vbias.n3613 73.1255
R12362 Vbias.n3613 Vbias.n3612 73.1255
R12363 Vbias.n3609 Vbias.n3589 73.1255
R12364 Vbias.n3589 Vbias.n3587 73.1255
R12365 Vbias.n3585 Vbias.n3584 73.1255
R12366 Vbias.n3586 Vbias.n3585 73.1255
R12367 Vbias.n3542 Vbias.n3541 73.1255
R12368 Vbias.n3541 Vbias.n3535 73.1255
R12369 Vbias.n3545 Vbias.n3544 73.1255
R12370 Vbias.n3544 Vbias.n3537 73.1255
R12371 Vbias.n3547 Vbias.n3546 73.1255
R12372 Vbias.n3547 Vbias.n2773 73.1255
R12373 Vbias.n3174 Vbias.n3172 73.1255
R12374 Vbias.n3174 Vbias.n8 73.1255
R12375 Vbias.n3175 Vbias.n3173 73.1255
R12376 Vbias.n3432 Vbias.n3175 73.1255
R12377 Vbias.n3180 Vbias.n3176 73.1255
R12378 Vbias.n3431 Vbias.n3176 73.1255
R12379 Vbias.n3400 Vbias.n3398 73.1255
R12380 Vbias.n3400 Vbias.n3190 73.1255
R12381 Vbias.n3410 Vbias.n3409 73.1255
R12382 Vbias.n3409 Vbias.n3192 73.1255
R12383 Vbias.n3414 Vbias.n3413 73.1255
R12384 Vbias.n3413 Vbias.n3394 73.1255
R12385 Vbias.n3209 Vbias.n3205 73.1255
R12386 Vbias.n3393 Vbias.n3205 73.1255
R12387 Vbias.n3362 Vbias.n3360 73.1255
R12388 Vbias.n3362 Vbias.n3219 73.1255
R12389 Vbias.n3372 Vbias.n3371 73.1255
R12390 Vbias.n3371 Vbias.n3221 73.1255
R12391 Vbias.n3376 Vbias.n3375 73.1255
R12392 Vbias.n3375 Vbias.n3356 73.1255
R12393 Vbias.n3330 Vbias.n3322 73.1255
R12394 Vbias.n3330 Vbias.n3329 73.1255
R12395 Vbias.n3321 Vbias.n3248 73.1255
R12396 Vbias.n3343 Vbias.n3248 73.1255
R12397 Vbias.n3337 Vbias.n3336 73.1255
R12398 Vbias.n3336 Vbias.n3318 73.1255
R12399 Vbias.n3256 Vbias.n3252 73.1255
R12400 Vbias.n3317 Vbias.n3252 73.1255
R12401 Vbias.n3286 Vbias.n3284 73.1255
R12402 Vbias.n3286 Vbias.n3266 73.1255
R12403 Vbias.n3296 Vbias.n3295 73.1255
R12404 Vbias.n3295 Vbias.n3268 73.1255
R12405 Vbias.n3300 Vbias.n3299 73.1255
R12406 Vbias.n3299 Vbias.n2774 73.1255
R12407 Vbias.n3430 Vbias.n3429 73.1255
R12408 Vbias.n3431 Vbias.n3430 73.1255
R12409 Vbias.n3197 Vbias.n3196 73.1255
R12410 Vbias.n3196 Vbias.n3190 73.1255
R12411 Vbias.n3200 Vbias.n3199 73.1255
R12412 Vbias.n3199 Vbias.n3192 73.1255
R12413 Vbias.n3202 Vbias.n3201 73.1255
R12414 Vbias.n3394 Vbias.n3202 73.1255
R12415 Vbias.n3392 Vbias.n3391 73.1255
R12416 Vbias.n3393 Vbias.n3392 73.1255
R12417 Vbias.n3226 Vbias.n3225 73.1255
R12418 Vbias.n3225 Vbias.n3219 73.1255
R12419 Vbias.n3229 Vbias.n3228 73.1255
R12420 Vbias.n3228 Vbias.n3221 73.1255
R12421 Vbias.n3231 Vbias.n3230 73.1255
R12422 Vbias.n3356 Vbias.n3231 73.1255
R12423 Vbias.n3354 Vbias.n3353 73.1255
R12424 Vbias.n3355 Vbias.n3354 73.1255
R12425 Vbias.n3323 Vbias.n3237 73.1255
R12426 Vbias.n3324 Vbias.n3323 73.1255
R12427 Vbias.n3328 Vbias.n3327 73.1255
R12428 Vbias.n3329 Vbias.n3328 73.1255
R12429 Vbias.n3345 Vbias.n3344 73.1255
R12430 Vbias.n3344 Vbias.n3343 73.1255
R12431 Vbias.n3340 Vbias.n3320 73.1255
R12432 Vbias.n3320 Vbias.n3318 73.1255
R12433 Vbias.n3316 Vbias.n3315 73.1255
R12434 Vbias.n3317 Vbias.n3316 73.1255
R12435 Vbias.n3273 Vbias.n3272 73.1255
R12436 Vbias.n3272 Vbias.n3266 73.1255
R12437 Vbias.n3276 Vbias.n3275 73.1255
R12438 Vbias.n3275 Vbias.n3268 73.1255
R12439 Vbias.n3278 Vbias.n3277 73.1255
R12440 Vbias.n3278 Vbias.n2774 73.1255
R12441 Vbias.n3712 Vbias.n3710 73.1255
R12442 Vbias.n3712 Vbias.n9 73.1255
R12443 Vbias.n3713 Vbias.n3711 73.1255
R12444 Vbias.n3970 Vbias.n3713 73.1255
R12445 Vbias.n3718 Vbias.n3714 73.1255
R12446 Vbias.n3969 Vbias.n3714 73.1255
R12447 Vbias.n3938 Vbias.n3936 73.1255
R12448 Vbias.n3938 Vbias.n3728 73.1255
R12449 Vbias.n3948 Vbias.n3947 73.1255
R12450 Vbias.n3947 Vbias.n3730 73.1255
R12451 Vbias.n3952 Vbias.n3951 73.1255
R12452 Vbias.n3951 Vbias.n3932 73.1255
R12453 Vbias.n3747 Vbias.n3743 73.1255
R12454 Vbias.n3931 Vbias.n3743 73.1255
R12455 Vbias.n3900 Vbias.n3898 73.1255
R12456 Vbias.n3900 Vbias.n3757 73.1255
R12457 Vbias.n3910 Vbias.n3909 73.1255
R12458 Vbias.n3909 Vbias.n3759 73.1255
R12459 Vbias.n3914 Vbias.n3913 73.1255
R12460 Vbias.n3913 Vbias.n3894 73.1255
R12461 Vbias.n3868 Vbias.n3860 73.1255
R12462 Vbias.n3868 Vbias.n3867 73.1255
R12463 Vbias.n3859 Vbias.n3786 73.1255
R12464 Vbias.n3881 Vbias.n3786 73.1255
R12465 Vbias.n3875 Vbias.n3874 73.1255
R12466 Vbias.n3874 Vbias.n3856 73.1255
R12467 Vbias.n3794 Vbias.n3790 73.1255
R12468 Vbias.n3855 Vbias.n3790 73.1255
R12469 Vbias.n3824 Vbias.n3822 73.1255
R12470 Vbias.n3824 Vbias.n3804 73.1255
R12471 Vbias.n3834 Vbias.n3833 73.1255
R12472 Vbias.n3833 Vbias.n3806 73.1255
R12473 Vbias.n3838 Vbias.n3837 73.1255
R12474 Vbias.n3837 Vbias.n2775 73.1255
R12475 Vbias.n3968 Vbias.n3967 73.1255
R12476 Vbias.n3969 Vbias.n3968 73.1255
R12477 Vbias.n3735 Vbias.n3734 73.1255
R12478 Vbias.n3734 Vbias.n3728 73.1255
R12479 Vbias.n3738 Vbias.n3737 73.1255
R12480 Vbias.n3737 Vbias.n3730 73.1255
R12481 Vbias.n3740 Vbias.n3739 73.1255
R12482 Vbias.n3932 Vbias.n3740 73.1255
R12483 Vbias.n3930 Vbias.n3929 73.1255
R12484 Vbias.n3931 Vbias.n3930 73.1255
R12485 Vbias.n3764 Vbias.n3763 73.1255
R12486 Vbias.n3763 Vbias.n3757 73.1255
R12487 Vbias.n3767 Vbias.n3766 73.1255
R12488 Vbias.n3766 Vbias.n3759 73.1255
R12489 Vbias.n3769 Vbias.n3768 73.1255
R12490 Vbias.n3894 Vbias.n3769 73.1255
R12491 Vbias.n3892 Vbias.n3891 73.1255
R12492 Vbias.n3893 Vbias.n3892 73.1255
R12493 Vbias.n3861 Vbias.n3775 73.1255
R12494 Vbias.n3862 Vbias.n3861 73.1255
R12495 Vbias.n3866 Vbias.n3865 73.1255
R12496 Vbias.n3867 Vbias.n3866 73.1255
R12497 Vbias.n3883 Vbias.n3882 73.1255
R12498 Vbias.n3882 Vbias.n3881 73.1255
R12499 Vbias.n3878 Vbias.n3858 73.1255
R12500 Vbias.n3858 Vbias.n3856 73.1255
R12501 Vbias.n3854 Vbias.n3853 73.1255
R12502 Vbias.n3855 Vbias.n3854 73.1255
R12503 Vbias.n3811 Vbias.n3810 73.1255
R12504 Vbias.n3810 Vbias.n3804 73.1255
R12505 Vbias.n3814 Vbias.n3813 73.1255
R12506 Vbias.n3813 Vbias.n3806 73.1255
R12507 Vbias.n3816 Vbias.n3815 73.1255
R12508 Vbias.n3816 Vbias.n2775 73.1255
R12509 Vbias.n2903 Vbias.n2901 73.1255
R12510 Vbias.n2905 Vbias.n2903 73.1255
R12511 Vbias.n2904 Vbias.n2902 73.1255
R12512 Vbias.n3162 Vbias.n2904 73.1255
R12513 Vbias.n2910 Vbias.n2906 73.1255
R12514 Vbias.n3161 Vbias.n2906 73.1255
R12515 Vbias.n3130 Vbias.n3128 73.1255
R12516 Vbias.n3130 Vbias.n2920 73.1255
R12517 Vbias.n3140 Vbias.n3139 73.1255
R12518 Vbias.n3139 Vbias.n2922 73.1255
R12519 Vbias.n3144 Vbias.n3143 73.1255
R12520 Vbias.n3143 Vbias.n3124 73.1255
R12521 Vbias.n2939 Vbias.n2935 73.1255
R12522 Vbias.n3123 Vbias.n2935 73.1255
R12523 Vbias.n3092 Vbias.n3090 73.1255
R12524 Vbias.n3092 Vbias.n2949 73.1255
R12525 Vbias.n3102 Vbias.n3101 73.1255
R12526 Vbias.n3101 Vbias.n2951 73.1255
R12527 Vbias.n3106 Vbias.n3105 73.1255
R12528 Vbias.n3105 Vbias.n3086 73.1255
R12529 Vbias.n3060 Vbias.n3052 73.1255
R12530 Vbias.n3060 Vbias.n3059 73.1255
R12531 Vbias.n3051 Vbias.n2978 73.1255
R12532 Vbias.n3073 Vbias.n2978 73.1255
R12533 Vbias.n3067 Vbias.n3066 73.1255
R12534 Vbias.n3066 Vbias.n3048 73.1255
R12535 Vbias.n2986 Vbias.n2982 73.1255
R12536 Vbias.n3047 Vbias.n2982 73.1255
R12537 Vbias.n3016 Vbias.n3014 73.1255
R12538 Vbias.n3016 Vbias.n2996 73.1255
R12539 Vbias.n3026 Vbias.n3025 73.1255
R12540 Vbias.n3025 Vbias.n2998 73.1255
R12541 Vbias.n3030 Vbias.n3029 73.1255
R12542 Vbias.n3029 Vbias.n2776 73.1255
R12543 Vbias.n3160 Vbias.n3159 73.1255
R12544 Vbias.n3161 Vbias.n3160 73.1255
R12545 Vbias.n2927 Vbias.n2926 73.1255
R12546 Vbias.n2926 Vbias.n2920 73.1255
R12547 Vbias.n2930 Vbias.n2929 73.1255
R12548 Vbias.n2929 Vbias.n2922 73.1255
R12549 Vbias.n2932 Vbias.n2931 73.1255
R12550 Vbias.n3124 Vbias.n2932 73.1255
R12551 Vbias.n3122 Vbias.n3121 73.1255
R12552 Vbias.n3123 Vbias.n3122 73.1255
R12553 Vbias.n2956 Vbias.n2955 73.1255
R12554 Vbias.n2955 Vbias.n2949 73.1255
R12555 Vbias.n2959 Vbias.n2958 73.1255
R12556 Vbias.n2958 Vbias.n2951 73.1255
R12557 Vbias.n2961 Vbias.n2960 73.1255
R12558 Vbias.n3086 Vbias.n2961 73.1255
R12559 Vbias.n3084 Vbias.n3083 73.1255
R12560 Vbias.n3085 Vbias.n3084 73.1255
R12561 Vbias.n3053 Vbias.n2967 73.1255
R12562 Vbias.n3054 Vbias.n3053 73.1255
R12563 Vbias.n3058 Vbias.n3057 73.1255
R12564 Vbias.n3059 Vbias.n3058 73.1255
R12565 Vbias.n3075 Vbias.n3074 73.1255
R12566 Vbias.n3074 Vbias.n3073 73.1255
R12567 Vbias.n3070 Vbias.n3050 73.1255
R12568 Vbias.n3050 Vbias.n3048 73.1255
R12569 Vbias.n3046 Vbias.n3045 73.1255
R12570 Vbias.n3047 Vbias.n3046 73.1255
R12571 Vbias.n3003 Vbias.n3002 73.1255
R12572 Vbias.n3002 Vbias.n2996 73.1255
R12573 Vbias.n3006 Vbias.n3005 73.1255
R12574 Vbias.n3005 Vbias.n2998 73.1255
R12575 Vbias.n3008 Vbias.n3007 73.1255
R12576 Vbias.n3008 Vbias.n2776 73.1255
R12577 Vbias.n4843 Vbias.n4842 73.1255
R12578 Vbias.n4844 Vbias.n4843 73.1255
R12579 Vbias.n4840 Vbias.n4839 73.1255
R12580 Vbias.n4839 Vbias.n4838 73.1255
R12581 Vbias.n2671 Vbias.n2667 73.1255
R12582 Vbias.n4837 Vbias.n2667 73.1255
R12583 Vbias.n4806 Vbias.n4804 73.1255
R12584 Vbias.n4806 Vbias.n2681 73.1255
R12585 Vbias.n4816 Vbias.n4815 73.1255
R12586 Vbias.n4815 Vbias.n2683 73.1255
R12587 Vbias.n4820 Vbias.n4819 73.1255
R12588 Vbias.n4819 Vbias.n4800 73.1255
R12589 Vbias.n2700 Vbias.n2696 73.1255
R12590 Vbias.n4799 Vbias.n2696 73.1255
R12591 Vbias.n4768 Vbias.n4766 73.1255
R12592 Vbias.n4768 Vbias.n2710 73.1255
R12593 Vbias.n4778 Vbias.n4777 73.1255
R12594 Vbias.n4777 Vbias.n2712 73.1255
R12595 Vbias.n4782 Vbias.n4781 73.1255
R12596 Vbias.n4781 Vbias.n4762 73.1255
R12597 Vbias.n4736 Vbias.n4728 73.1255
R12598 Vbias.n4736 Vbias.n4735 73.1255
R12599 Vbias.n4727 Vbias.n2739 73.1255
R12600 Vbias.n4749 Vbias.n2739 73.1255
R12601 Vbias.n4743 Vbias.n4742 73.1255
R12602 Vbias.n4742 Vbias.n4724 73.1255
R12603 Vbias.n2747 Vbias.n2743 73.1255
R12604 Vbias.n4723 Vbias.n2743 73.1255
R12605 Vbias.n4692 Vbias.n4690 73.1255
R12606 Vbias.n4692 Vbias.n2757 73.1255
R12607 Vbias.n4702 Vbias.n4701 73.1255
R12608 Vbias.n4701 Vbias.n2759 73.1255
R12609 Vbias.n4706 Vbias.n4705 73.1255
R12610 Vbias.n4705 Vbias.n4686 73.1255
R12611 Vbias.n4836 Vbias.n4835 73.1255
R12612 Vbias.n4837 Vbias.n4836 73.1255
R12613 Vbias.n2688 Vbias.n2687 73.1255
R12614 Vbias.n2687 Vbias.n2681 73.1255
R12615 Vbias.n2691 Vbias.n2690 73.1255
R12616 Vbias.n2690 Vbias.n2683 73.1255
R12617 Vbias.n2693 Vbias.n2692 73.1255
R12618 Vbias.n4800 Vbias.n2693 73.1255
R12619 Vbias.n4798 Vbias.n4797 73.1255
R12620 Vbias.n4799 Vbias.n4798 73.1255
R12621 Vbias.n2717 Vbias.n2716 73.1255
R12622 Vbias.n2716 Vbias.n2710 73.1255
R12623 Vbias.n2720 Vbias.n2719 73.1255
R12624 Vbias.n2719 Vbias.n2712 73.1255
R12625 Vbias.n2722 Vbias.n2721 73.1255
R12626 Vbias.n4762 Vbias.n2722 73.1255
R12627 Vbias.n4760 Vbias.n4759 73.1255
R12628 Vbias.n4761 Vbias.n4760 73.1255
R12629 Vbias.n4729 Vbias.n2728 73.1255
R12630 Vbias.n4730 Vbias.n4729 73.1255
R12631 Vbias.n4734 Vbias.n4733 73.1255
R12632 Vbias.n4735 Vbias.n4734 73.1255
R12633 Vbias.n4751 Vbias.n4750 73.1255
R12634 Vbias.n4750 Vbias.n4749 73.1255
R12635 Vbias.n4746 Vbias.n4726 73.1255
R12636 Vbias.n4726 Vbias.n4724 73.1255
R12637 Vbias.n4722 Vbias.n4721 73.1255
R12638 Vbias.n4723 Vbias.n4722 73.1255
R12639 Vbias.n2764 Vbias.n2763 73.1255
R12640 Vbias.n2763 Vbias.n2757 73.1255
R12641 Vbias.n2767 Vbias.n2766 73.1255
R12642 Vbias.n2766 Vbias.n2759 73.1255
R12643 Vbias.n2769 Vbias.n2768 73.1255
R12644 Vbias.n4686 Vbias.n2769 73.1255
R12645 Vbias.n4906 Vbias.n4905 73.1255
R12646 Vbias.n4905 Vbias.n4904 73.1255
R12647 Vbias.n4909 Vbias.n4908 73.1255
R12648 Vbias.n4910 Vbias.n4909 73.1255
R12649 Vbias.n2659 Vbias.n2658 73.1255
R12650 Vbias.n4911 Vbias.n2659 73.1255
R12651 Vbias.n4914 Vbias.n4913 73.1255
R12652 Vbias.n4913 Vbias.n2653 73.1255
R12653 Vbias.n4927 Vbias.n4926 73.1255
R12654 Vbias.n4926 Vbias.n4925 73.1255
R12655 Vbias.n4931 Vbias.n4930 73.1255
R12656 Vbias.n4932 Vbias.n4931 73.1255
R12657 Vbias.n2645 Vbias.n2644 73.1255
R12658 Vbias.n4933 Vbias.n2645 73.1255
R12659 Vbias.n4936 Vbias.n4935 73.1255
R12660 Vbias.n4935 Vbias.n2639 73.1255
R12661 Vbias.n4950 Vbias.n4949 73.1255
R12662 Vbias.n4949 Vbias.n4948 73.1255
R12663 Vbias.n4954 Vbias.n4953 73.1255
R12664 Vbias.n4955 Vbias.n4954 73.1255
R12665 Vbias.n2631 Vbias.n2630 73.1255
R12666 Vbias.n4956 Vbias.n2631 73.1255
R12667 Vbias.n4962 Vbias.n4961 73.1255
R12668 Vbias.n4961 Vbias.n2623 73.1255
R12669 Vbias.n2622 Vbias.n2620 73.1255
R12670 Vbias.n2628 Vbias.n2622 73.1255
R12671 Vbias.n2626 Vbias.n2616 73.1255
R12672 Vbias.n2627 Vbias.n2626 73.1255
R12673 Vbias.n4973 Vbias.n4972 73.1255
R12674 Vbias.n4972 Vbias.n2614 73.1255
R12675 Vbias.n4980 Vbias.n4979 73.1255
R12676 Vbias.n4979 Vbias.n2609 73.1255
R12677 Vbias.n2608 Vbias.n2606 73.1255
R12678 Vbias.n2610 Vbias.n2608 73.1255
R12679 Vbias.n4549 Vbias.n4548 73.1255
R12680 Vbias.n4550 Vbias.n4549 73.1255
R12681 Vbias.n4416 Vbias.n4410 73.1255
R12682 Vbias.n4416 Vbias.n4414 73.1255
R12683 Vbias.n4421 Vbias.n4420 73.1255
R12684 Vbias.n4420 Vbias.n4415 73.1255
R12685 Vbias.n4425 Vbias.n4424 73.1255
R12686 Vbias.n4535 Vbias.n4425 73.1255
R12687 Vbias.n4533 Vbias.n4532 73.1255
R12688 Vbias.n4534 Vbias.n4533 73.1255
R12689 Vbias.n4435 Vbias.n4429 73.1255
R12690 Vbias.n4435 Vbias.n4433 73.1255
R12691 Vbias.n4432 Vbias.n4430 73.1255
R12692 Vbias.n4434 Vbias.n4432 73.1255
R12693 Vbias.n4451 Vbias.n4440 73.1255
R12694 Vbias.n4452 Vbias.n4451 73.1255
R12695 Vbias.n4448 Vbias.n4442 73.1255
R12696 Vbias.n4448 Vbias.n4446 73.1255
R12697 Vbias.n4457 Vbias.n4456 73.1255
R12698 Vbias.n4456 Vbias.n4447 73.1255
R12699 Vbias.n4459 Vbias.n4458 73.1255
R12700 Vbias.n4460 Vbias.n4459 73.1255
R12701 Vbias.n4473 Vbias.n4462 73.1255
R12702 Vbias.n4474 Vbias.n4473 73.1255
R12703 Vbias.n4470 Vbias.n4464 73.1255
R12704 Vbias.n4470 Vbias.n4468 73.1255
R12705 Vbias.n4479 Vbias.n4478 73.1255
R12706 Vbias.n4478 Vbias.n4469 73.1255
R12707 Vbias.n4481 Vbias.n4480 73.1255
R12708 Vbias.n4482 Vbias.n4481 73.1255
R12709 Vbias.n4489 Vbias.n4485 73.1255
R12710 Vbias.n4490 Vbias.n4489 73.1255
R12711 Vbias.n4493 Vbias.n4492 73.1255
R12712 Vbias.n4492 Vbias.n4491 73.1255
R12713 Vbias.n4669 Vbias.n4668 73.1255
R12714 Vbias.n4670 Vbias.n4669 73.1255
R12715 Vbias.n4587 Vbias.n4586 73.1255
R12716 Vbias.n4588 Vbias.n4587 73.1255
R12717 Vbias.n4663 Vbias.n4662 73.1255
R12718 Vbias.n4662 Vbias.n4661 73.1255
R12719 Vbias.n4659 Vbias.n4658 73.1255
R12720 Vbias.n4660 Vbias.n4659 73.1255
R12721 Vbias.n4616 Vbias.n4592 73.1255
R12722 Vbias.n4617 Vbias.n4616 73.1255
R12723 Vbias.n4619 Vbias.n4594 73.1255
R12724 Vbias.n4619 Vbias.n4618 73.1255
R12725 Vbias.n4615 Vbias.n4596 73.1255
R12726 Vbias.n4615 Vbias.n2592 73.1255
R12727 Vbias.n4624 Vbias.n4598 73.1255
R12728 Vbias.n4625 Vbias.n4624 73.1255
R12729 Vbias.n4631 Vbias.n4600 73.1255
R12730 Vbias.n4632 Vbias.n4631 73.1255
R12731 Vbias.n4611 Vbias.n4601 73.1255
R12732 Vbias.n4633 Vbias.n4611 73.1255
R12733 Vbias.n4608 Vbias.n4603 73.1255
R12734 Vbias.n4608 Vbias.n4606 73.1255
R12735 Vbias.n4638 Vbias.n4637 73.1255
R12736 Vbias.n4637 Vbias.n4607 73.1255
R12737 Vbias.n5035 Vbias.n5034 73.1255
R12738 Vbias.n5036 Vbias.n5035 73.1255
R12739 Vbias.n4673 Vbias.n4672 73.1255
R12740 Vbias.n4672 Vbias.n4671 73.1255
R12741 Vbias.n4572 Vbias.n4557 73.1255
R12742 Vbias.n4573 Vbias.n4572 73.1255
R12743 Vbias.n4565 Vbias.n4564 73.1255
R12744 Vbias.n4564 Vbias.n4563 73.1255
R12745 Vbias.n4680 Vbias.n4679 73.1255
R12746 Vbias.n4681 Vbias.n4680 73.1255
R12747 Vbias.n7327 Vbias.n7325 73.1255
R12748 Vbias.n7327 Vbias.n917 73.1255
R12749 Vbias.n7332 Vbias.n7331 73.1255
R12750 Vbias.n7331 Vbias.n7329 73.1255
R12751 Vbias.n7338 Vbias.n7337 73.1255
R12752 Vbias.n7337 Vbias.n7335 73.1255
R12753 Vbias.n7341 Vbias.n7340 73.1255
R12754 Vbias.n7450 Vbias.n7341 73.1255
R12755 Vbias.n7448 Vbias.n7447 73.1255
R12756 Vbias.n7449 Vbias.n7448 73.1255
R12757 Vbias.n7356 Vbias.n7355 73.1255
R12758 Vbias.n7355 Vbias.n7351 73.1255
R12759 Vbias.n7359 Vbias.n7358 73.1255
R12760 Vbias.n7358 Vbias.n7352 73.1255
R12761 Vbias.n7361 Vbias.n7360 73.1255
R12762 Vbias.n7434 Vbias.n7361 73.1255
R12763 Vbias.n7432 Vbias.n7431 73.1255
R12764 Vbias.n7433 Vbias.n7432 73.1255
R12765 Vbias.n7374 Vbias.n7365 73.1255
R12766 Vbias.n7375 Vbias.n7374 73.1255
R12767 Vbias.n7377 Vbias.n7368 73.1255
R12768 Vbias.n7377 Vbias.n7376 73.1255
R12769 Vbias.n7424 Vbias.n7423 73.1255
R12770 Vbias.n7423 Vbias.n7422 73.1255
R12771 Vbias.n7419 Vbias.n7418 73.1255
R12772 Vbias.n7418 Vbias.n7416 73.1255
R12773 Vbias.n7414 Vbias.n7413 73.1255
R12774 Vbias.n7415 Vbias.n7414 73.1255
R12775 Vbias.n7394 Vbias.n7393 73.1255
R12776 Vbias.n7393 Vbias.n7389 73.1255
R12777 Vbias.n7397 Vbias.n7396 73.1255
R12778 Vbias.n7396 Vbias.n7390 73.1255
R12779 Vbias.n7399 Vbias.n7398 73.1255
R12780 Vbias.n6503 Vbias.n860 73.1255
R12781 Vbias.n6504 Vbias.n6503 73.1255
R12782 Vbias.n6467 Vbias.n862 73.1255
R12783 Vbias.n6468 Vbias.n6467 73.1255
R12784 Vbias.n6496 Vbias.n864 73.1255
R12785 Vbias.n6497 Vbias.n6496 73.1255
R12786 Vbias.n6492 Vbias.n866 73.1255
R12787 Vbias.n6492 Vbias.n6491 73.1255
R12788 Vbias.n6489 Vbias.n868 73.1255
R12789 Vbias.n6490 Vbias.n6489 73.1255
R12790 Vbias.n6473 Vbias.n870 73.1255
R12791 Vbias.n6474 Vbias.n6473 73.1255
R12792 Vbias.n6482 Vbias.n872 73.1255
R12793 Vbias.n6483 Vbias.n6482 73.1255
R12794 Vbias.n6478 Vbias.n874 73.1255
R12795 Vbias.n6478 Vbias.n6477 73.1255
R12796 Vbias.n6475 Vbias.n875 73.1255
R12797 Vbias.n6476 Vbias.n6475 73.1255
R12798 Vbias.n7569 Vbias.n7568 73.1255
R12799 Vbias.n7568 Vbias.n7567 73.1255
R12800 Vbias.n7565 Vbias.n7564 73.1255
R12801 Vbias.n7566 Vbias.n7565 73.1255
R12802 Vbias.n891 Vbias.n890 73.1255
R12803 Vbias.n892 Vbias.n891 73.1255
R12804 Vbias.n7559 Vbias.n7558 73.1255
R12805 Vbias.n7558 Vbias.n7557 73.1255
R12806 Vbias.n7555 Vbias.n7554 73.1255
R12807 Vbias.n7556 Vbias.n7555 73.1255
R12808 Vbias.n908 Vbias.n907 73.1255
R12809 Vbias.n907 Vbias.n906 73.1255
R12810 Vbias.n915 Vbias.n900 73.1255
R12811 Vbias.n916 Vbias.n915 73.1255
R12812 Vbias.n7547 Vbias.n7546 73.1255
R12813 Vbias.n7546 Vbias.n7545 73.1255
R12814 Vbias.n6390 Vbias.n6365 73.1255
R12815 Vbias.n6390 Vbias.n6226 73.1255
R12816 Vbias.n6394 Vbias.n6367 73.1255
R12817 Vbias.n6395 Vbias.n6394 73.1255
R12818 Vbias.n6397 Vbias.n6369 73.1255
R12819 Vbias.n6398 Vbias.n6397 73.1255
R12820 Vbias.n6404 Vbias.n6371 73.1255
R12821 Vbias.n6405 Vbias.n6404 73.1255
R12822 Vbias.n6407 Vbias.n6373 73.1255
R12823 Vbias.n6407 Vbias.n6406 73.1255
R12824 Vbias.n6411 Vbias.n6375 73.1255
R12825 Vbias.n6412 Vbias.n6411 73.1255
R12826 Vbias.n6414 Vbias.n6377 73.1255
R12827 Vbias.n6415 Vbias.n6414 73.1255
R12828 Vbias.n6421 Vbias.n6379 73.1255
R12829 Vbias.n6422 Vbias.n6421 73.1255
R12830 Vbias.n6423 Vbias.n6380 73.1255
R12831 Vbias.n6424 Vbias.n6423 73.1255
R12832 Vbias.n6556 Vbias.n6555 73.1255
R12833 Vbias.n6555 Vbias.n6554 73.1255
R12834 Vbias.n6552 Vbias.n6551 73.1255
R12835 Vbias.n6553 Vbias.n6552 73.1255
R12836 Vbias.n6437 Vbias.n6436 73.1255
R12837 Vbias.n6438 Vbias.n6437 73.1255
R12838 Vbias.n6546 Vbias.n6545 73.1255
R12839 Vbias.n6545 Vbias.n6544 73.1255
R12840 Vbias.n6542 Vbias.n6541 73.1255
R12841 Vbias.n6543 Vbias.n6542 73.1255
R12842 Vbias.n6454 Vbias.n6453 73.1255
R12843 Vbias.n6453 Vbias.n6452 73.1255
R12844 Vbias.n6461 Vbias.n6446 73.1255
R12845 Vbias.n6462 Vbias.n6461 73.1255
R12846 Vbias.n6534 Vbias.n6533 73.1255
R12847 Vbias.n6533 Vbias.n6532 73.1255
R12848 Vbias.n6170 Vbias.n6155 73.1255
R12849 Vbias.n6170 Vbias.n6169 73.1255
R12850 Vbias.n6174 Vbias.n6157 73.1255
R12851 Vbias.n6175 Vbias.n6174 73.1255
R12852 Vbias.n6177 Vbias.n6159 73.1255
R12853 Vbias.n6178 Vbias.n6177 73.1255
R12854 Vbias.n6184 Vbias.n6161 73.1255
R12855 Vbias.n6185 Vbias.n6184 73.1255
R12856 Vbias.n6186 Vbias.n6162 73.1255
R12857 Vbias.n6187 Vbias.n6186 73.1255
R12858 Vbias.n6623 Vbias.n6622 73.1255
R12859 Vbias.n6622 Vbias.n6621 73.1255
R12860 Vbias.n6619 Vbias.n6618 73.1255
R12861 Vbias.n6620 Vbias.n6619 73.1255
R12862 Vbias.n6200 Vbias.n6199 73.1255
R12863 Vbias.n6201 Vbias.n6200 73.1255
R12864 Vbias.n6613 Vbias.n6612 73.1255
R12865 Vbias.n6612 Vbias.n6611 73.1255
R12866 Vbias.n6609 Vbias.n6608 73.1255
R12867 Vbias.n6610 Vbias.n6609 73.1255
R12868 Vbias.n6217 Vbias.n6216 73.1255
R12869 Vbias.n6216 Vbias.n6215 73.1255
R12870 Vbias.n6224 Vbias.n6209 73.1255
R12871 Vbias.n6225 Vbias.n6224 73.1255
R12872 Vbias.n6601 Vbias.n6600 73.1255
R12873 Vbias.n6600 Vbias.n6599 73.1255
R12874 Vbias.n6149 Vbias.n6148 73.1255
R12875 Vbias.n6150 Vbias.n6149 73.1255
R12876 Vbias.n6151 Vbias.n6147 73.1255
R12877 Vbias.n6151 Vbias.n6144 73.1255
R12878 Vbias.n6645 Vbias.n6644 73.1255
R12879 Vbias.n6644 Vbias.n6643 73.1255
R12880 Vbias.n6141 Vbias.n6135 73.1255
R12881 Vbias.n6141 Vbias.n755 73.1255
R12882 Vbias.n7734 Vbias.n7733 73.1255
R12883 Vbias.n7735 Vbias.n7734 73.1255
R12884 Vbias.n690 Vbias.n683 73.1255
R12885 Vbias.n690 Vbias.n688 73.1255
R12886 Vbias.n695 Vbias.n694 73.1255
R12887 Vbias.n694 Vbias.n689 73.1255
R12888 Vbias.n697 Vbias.n696 73.1255
R12889 Vbias.n698 Vbias.n697 73.1255
R12890 Vbias.n707 Vbias.n700 73.1255
R12891 Vbias.n707 Vbias.n706 73.1255
R12892 Vbias.n7716 Vbias.n7715 73.1255
R12893 Vbias.n7715 Vbias.n7714 73.1255
R12894 Vbias.n717 Vbias.n713 73.1255
R12895 Vbias.n717 Vbias.n710 73.1255
R12896 Vbias.n715 Vbias.n714 73.1255
R12897 Vbias.n716 Vbias.n715 73.1255
R12898 Vbias.n724 Vbias.n720 73.1255
R12899 Vbias.n725 Vbias.n724 73.1255
R12900 Vbias.n7702 Vbias.n7701 73.1255
R12901 Vbias.n7701 Vbias.n7700 73.1255
R12902 Vbias.n7698 Vbias.n7697 73.1255
R12903 Vbias.n7699 Vbias.n7698 73.1255
R12904 Vbias.n7688 Vbias.n7687 73.1255
R12905 Vbias.n7687 Vbias.n734 73.1255
R12906 Vbias.n733 Vbias.n731 73.1255
R12907 Vbias.n7685 Vbias.n733 73.1255
R12908 Vbias.n7683 Vbias.n7682 73.1255
R12909 Vbias.n7684 Vbias.n7683 73.1255
R12910 Vbias.n749 Vbias.n748 73.1255
R12911 Vbias.n748 Vbias.n744 73.1255
R12912 Vbias.n752 Vbias.n751 73.1255
R12913 Vbias.n751 Vbias.n745 73.1255
R12914 Vbias.n754 Vbias.n753 73.1255
R12915 Vbias.n7669 Vbias.n754 73.1255
R12916 Vbias.n6674 Vbias.n6673 73.1255
R12917 Vbias.n6675 Vbias.n6674 73.1255
R12918 Vbias.n1477 Vbias.n1471 73.1255
R12919 Vbias.n1477 Vbias.n1475 73.1255
R12920 Vbias.n1474 Vbias.n1472 73.1255
R12921 Vbias.n1476 Vbias.n1474 73.1255
R12922 Vbias.n1493 Vbias.n1482 73.1255
R12923 Vbias.n1493 Vbias.n1459 73.1255
R12924 Vbias.n1490 Vbias.n1484 73.1255
R12925 Vbias.n1490 Vbias.n1488 73.1255
R12926 Vbias.n1498 Vbias.n1497 73.1255
R12927 Vbias.n1497 Vbias.n1489 73.1255
R12928 Vbias.n1500 Vbias.n1499 73.1255
R12929 Vbias.n6132 Vbias.n1500 73.1255
R12930 Vbias.n6302 Vbias.n6298 73.1255
R12931 Vbias.n6303 Vbias.n6302 73.1255
R12932 Vbias.n6310 Vbias.n6309 73.1255
R12933 Vbias.n6309 Vbias.n6308 73.1255
R12934 Vbias.n6306 Vbias.n6295 73.1255
R12935 Vbias.n6307 Vbias.n6306 73.1255
R12936 Vbias.n6294 Vbias.n6293 73.1255
R12937 Vbias.n6293 Vbias.n6291 73.1255
R12938 Vbias.n6288 Vbias.n6287 73.1255
R12939 Vbias.n6287 Vbias.n6280 73.1255
R12940 Vbias.n6279 Vbias.n6277 73.1255
R12941 Vbias.n6285 Vbias.n6279 73.1255
R12942 Vbias.n6283 Vbias.n6273 73.1255
R12943 Vbias.n6284 Vbias.n6283 73.1255
R12944 Vbias.n6272 Vbias.n6271 73.1255
R12945 Vbias.n6271 Vbias.n6269 73.1255
R12946 Vbias.n6266 Vbias.n6265 73.1255
R12947 Vbias.n6265 Vbias.n6263 73.1255
R12948 Vbias.n6262 Vbias.n6259 73.1255
R12949 Vbias.n6262 Vbias.n6261 73.1255
R12950 Vbias.n6250 Vbias.n6249 73.1255
R12951 Vbias.n6252 Vbias.n6250 73.1255
R12952 Vbias.n6254 Vbias.n6248 73.1255
R12953 Vbias.n6254 Vbias.n6253 73.1255
R12954 Vbias.n6351 Vbias.n6350 73.1255
R12955 Vbias.n6352 Vbias.n6351 73.1255
R12956 Vbias.n6244 Vbias.n6243 73.1255
R12957 Vbias.n6353 Vbias.n6244 73.1255
R12958 Vbias.n6240 Vbias.n6239 73.1255
R12959 Vbias.n6239 Vbias.n6234 73.1255
R12960 Vbias.n6237 Vbias.n6230 73.1255
R12961 Vbias.n6237 Vbias.n6235 73.1255
R12962 Vbias.n6588 Vbias.n6587 73.1255
R12963 Vbias.n6589 Vbias.n6588 73.1255
R12964 Vbias.n7650 Vbias.n7649 73.1255
R12965 Vbias.n7651 Vbias.n7650 73.1255
R12966 Vbias.n7647 Vbias.n7646 73.1255
R12967 Vbias.n7646 Vbias.n7645 73.1255
R12968 Vbias.n7643 Vbias.n7642 73.1255
R12969 Vbias.n7644 Vbias.n7643 73.1255
R12970 Vbias.n790 Vbias.n784 73.1255
R12971 Vbias.n790 Vbias.n788 73.1255
R12972 Vbias.n796 Vbias.n795 73.1255
R12973 Vbias.n795 Vbias.n789 73.1255
R12974 Vbias.n799 Vbias.n798 73.1255
R12975 Vbias.n7630 Vbias.n799 73.1255
R12976 Vbias.n7628 Vbias.n7627 73.1255
R12977 Vbias.n7629 Vbias.n7628 73.1255
R12978 Vbias.n809 Vbias.n803 73.1255
R12979 Vbias.n809 Vbias.n807 73.1255
R12980 Vbias.n817 Vbias.n816 73.1255
R12981 Vbias.n816 Vbias.n808 73.1255
R12982 Vbias.n820 Vbias.n819 73.1255
R12983 Vbias.n7615 Vbias.n820 73.1255
R12984 Vbias.n7613 Vbias.n7612 73.1255
R12985 Vbias.n7614 Vbias.n7613 73.1255
R12986 Vbias.n831 Vbias.n825 73.1255
R12987 Vbias.n831 Vbias.n829 73.1255
R12988 Vbias.n828 Vbias.n826 73.1255
R12989 Vbias.n830 Vbias.n828 73.1255
R12990 Vbias.n848 Vbias.n837 73.1255
R12991 Vbias.n849 Vbias.n848 73.1255
R12992 Vbias.n845 Vbias.n839 73.1255
R12993 Vbias.n845 Vbias.n843 73.1255
R12994 Vbias.n854 Vbias.n853 73.1255
R12995 Vbias.n853 Vbias.n844 73.1255
R12996 Vbias.n856 Vbias.n855 73.1255
R12997 Vbias.n857 Vbias.n856 73.1255
R12998 Vbias.n7529 Vbias.n7528 73.1255
R12999 Vbias.n7530 Vbias.n7529 73.1255
R13000 Vbias.n7526 Vbias.n7525 73.1255
R13001 Vbias.n7525 Vbias.n7524 73.1255
R13002 Vbias.n7522 Vbias.n7521 73.1255
R13003 Vbias.n7523 Vbias.n7522 73.1255
R13004 Vbias.n941 Vbias.n935 73.1255
R13005 Vbias.n941 Vbias.n939 73.1255
R13006 Vbias.n951 Vbias.n950 73.1255
R13007 Vbias.n950 Vbias.n940 73.1255
R13008 Vbias.n954 Vbias.n953 73.1255
R13009 Vbias.n7509 Vbias.n954 73.1255
R13010 Vbias.n7507 Vbias.n7506 73.1255
R13011 Vbias.n7508 Vbias.n7507 73.1255
R13012 Vbias.n964 Vbias.n958 73.1255
R13013 Vbias.n964 Vbias.n962 73.1255
R13014 Vbias.n972 Vbias.n971 73.1255
R13015 Vbias.n971 Vbias.n963 73.1255
R13016 Vbias.n975 Vbias.n974 73.1255
R13017 Vbias.n7493 Vbias.n975 73.1255
R13018 Vbias.n7491 Vbias.n7490 73.1255
R13019 Vbias.n7492 Vbias.n7491 73.1255
R13020 Vbias.n986 Vbias.n980 73.1255
R13021 Vbias.n986 Vbias.n984 73.1255
R13022 Vbias.n983 Vbias.n981 73.1255
R13023 Vbias.n985 Vbias.n983 73.1255
R13024 Vbias.n1003 Vbias.n992 73.1255
R13025 Vbias.n1004 Vbias.n1003 73.1255
R13026 Vbias.n1000 Vbias.n994 73.1255
R13027 Vbias.n1000 Vbias.n998 73.1255
R13028 Vbias.n1009 Vbias.n1008 73.1255
R13029 Vbias.n1008 Vbias.n999 73.1255
R13030 Vbias.n1011 Vbias.n1010 73.1255
R13031 Vbias.n1018 Vbias.n1011 73.1255
R13032 Vbias.n1027 Vbias.n1019 73.1255
R13033 Vbias.n1028 Vbias.n1027 73.1255
R13034 Vbias.n7319 Vbias.n7318 73.1255
R13035 Vbias.n7318 Vbias.n7317 73.1255
R13036 Vbias.n7315 Vbias.n7314 73.1255
R13037 Vbias.n7316 Vbias.n7315 73.1255
R13038 Vbias.n1038 Vbias.n1032 73.1255
R13039 Vbias.n1038 Vbias.n1036 73.1255
R13040 Vbias.n1046 Vbias.n1045 73.1255
R13041 Vbias.n1045 Vbias.n1037 73.1255
R13042 Vbias.n1049 Vbias.n1048 73.1255
R13043 Vbias.n7302 Vbias.n1049 73.1255
R13044 Vbias.n7300 Vbias.n7299 73.1255
R13045 Vbias.n7301 Vbias.n7300 73.1255
R13046 Vbias.n1059 Vbias.n1053 73.1255
R13047 Vbias.n1059 Vbias.n1057 73.1255
R13048 Vbias.n1067 Vbias.n1066 73.1255
R13049 Vbias.n1066 Vbias.n1058 73.1255
R13050 Vbias.n1070 Vbias.n1069 73.1255
R13051 Vbias.n7287 Vbias.n1070 73.1255
R13052 Vbias.n7285 Vbias.n7284 73.1255
R13053 Vbias.n7286 Vbias.n7285 73.1255
R13054 Vbias.n7236 Vbias.n7230 73.1255
R13055 Vbias.n7236 Vbias.n7234 73.1255
R13056 Vbias.n7233 Vbias.n7231 73.1255
R13057 Vbias.n7235 Vbias.n7233 73.1255
R13058 Vbias.n7253 Vbias.n7242 73.1255
R13059 Vbias.n7254 Vbias.n7253 73.1255
R13060 Vbias.n7250 Vbias.n7244 73.1255
R13061 Vbias.n7250 Vbias.n7248 73.1255
R13062 Vbias.n7259 Vbias.n7258 73.1255
R13063 Vbias.n7258 Vbias.n7249 73.1255
R13064 Vbias.n7261 Vbias.n7260 73.1255
R13065 Vbias.n761 Vbias.n759 73.1255
R13066 Vbias.n759 Vbias.n756 73.1255
R13067 Vbias.n766 Vbias.n762 73.1255
R13068 Vbias.n766 Vbias.n757 73.1255
R13069 Vbias.n764 Vbias.n763 73.1255
R13070 Vbias.n765 Vbias.n764 73.1255
R13071 Vbias.n6591 Vbias.n772 73.1255
R13072 Vbias.n6591 Vbias.n6590 73.1255
R13073 Vbias.n6597 Vbias.n774 73.1255
R13074 Vbias.n6598 Vbias.n6597 73.1255
R13075 Vbias.n7654 Vbias.n7653 73.1255
R13076 Vbias.n7653 Vbias.n7652 73.1255
R13077 Vbias.n6510 Vbias.n6509 73.1255
R13078 Vbias.n6509 Vbias.n6508 73.1255
R13079 Vbias.n6516 Vbias.n6515 73.1255
R13080 Vbias.n6517 Vbias.n6516 73.1255
R13081 Vbias.n6524 Vbias.n6521 73.1255
R13082 Vbias.n6521 Vbias.n6518 73.1255
R13083 Vbias.n6527 Vbias.n6526 73.1255
R13084 Vbias.n6526 Vbias.n6519 73.1255
R13085 Vbias.n7533 Vbias.n7532 73.1255
R13086 Vbias.n7532 Vbias.n7531 73.1255
R13087 Vbias.n1016 Vbias.n1015 73.1255
R13088 Vbias.n1017 Vbias.n1016 73.1255
R13089 Vbias.n7543 Vbias.n7542 73.1255
R13090 Vbias.n7544 Vbias.n7543 73.1255
R13091 Vbias.n1025 Vbias.n923 73.1255
R13092 Vbias.n1026 Vbias.n1025 73.1255
R13093 Vbias.n1506 Vbias.n1505 73.1255
R13094 Vbias.n1505 Vbias.n1504 73.1255
R13095 Vbias.n6130 Vbias.n6129 73.1255
R13096 Vbias.n6131 Vbias.n6130 73.1255
R13097 Vbias.n347 Vbias.n346 73.1255
R13098 Vbias.n348 Vbias.n347 73.1255
R13099 Vbias.n344 Vbias.n343 73.1255
R13100 Vbias.n343 Vbias.n342 73.1255
R13101 Vbias.n340 Vbias.n339 73.1255
R13102 Vbias.n341 Vbias.n340 73.1255
R13103 Vbias.n334 Vbias.n333 73.1255
R13104 Vbias.n333 Vbias.n332 73.1255
R13105 Vbias.n7940 Vbias.n7939 73.1255
R13106 Vbias.n7939 Vbias.n7938 73.1255
R13107 Vbias.n5597 Vbias.n5596 73.1255
R13108 Vbias.n5596 Vbias.n174 73.1255
R13109 Vbias.n5600 Vbias.n5599 73.1255
R13110 Vbias.n5601 Vbias.n5600 73.1255
R13111 Vbias.n5589 Vbias.n5588 73.1255
R13112 Vbias.n5602 Vbias.n5589 73.1255
R13113 Vbias.n5585 Vbias.n5584 73.1255
R13114 Vbias.n5584 Vbias.n5579 73.1255
R13115 Vbias.n5582 Vbias.n5575 73.1255
R13116 Vbias.n5582 Vbias.n5580 73.1255
R13117 Vbias.n5618 Vbias.n5617 73.1255
R13118 Vbias.n5619 Vbias.n5618 73.1255
R13119 Vbias.n5571 Vbias.n5570 73.1255
R13120 Vbias.n5620 Vbias.n5571 73.1255
R13121 Vbias.n5567 Vbias.n5566 73.1255
R13122 Vbias.n5566 Vbias.n5561 73.1255
R13123 Vbias.n5564 Vbias.n5557 73.1255
R13124 Vbias.n5564 Vbias.n5562 73.1255
R13125 Vbias.n5637 Vbias.n5636 73.1255
R13126 Vbias.n5638 Vbias.n5637 73.1255
R13127 Vbias.n2227 Vbias.n2226 73.1255
R13128 Vbias.n5639 Vbias.n2227 73.1255
R13129 Vbias.n2225 Vbias.n2224 73.1255
R13130 Vbias.n2224 Vbias.n2217 73.1255
R13131 Vbias.n2216 Vbias.n2214 73.1255
R13132 Vbias.n2222 Vbias.n2216 73.1255
R13133 Vbias.n2220 Vbias.n2210 73.1255
R13134 Vbias.n2221 Vbias.n2220 73.1255
R13135 Vbias.n2209 Vbias.n2208 73.1255
R13136 Vbias.n2208 Vbias.n2206 73.1255
R13137 Vbias.n2203 Vbias.n2202 73.1255
R13138 Vbias.n2202 Vbias.n2200 73.1255
R13139 Vbias.n2199 Vbias.n2197 73.1255
R13140 Vbias.n2199 Vbias.n447 73.1255
R13141 Vbias.n7885 Vbias.n7884 73.1255
R13142 Vbias.n7886 Vbias.n7885 73.1255
R13143 Vbias.n7875 Vbias.n7874 73.1255
R13144 Vbias.n7874 Vbias.n456 73.1255
R13145 Vbias.n455 Vbias.n453 73.1255
R13146 Vbias.n7872 Vbias.n455 73.1255
R13147 Vbias.n5671 Vbias.n5670 73.1255
R13148 Vbias.n5670 Vbias.n457 73.1255
R13149 Vbias.n5674 Vbias.n5673 73.1255
R13150 Vbias.n5675 Vbias.n5674 73.1255
R13151 Vbias.n2192 Vbias.n2191 73.1255
R13152 Vbias.n5676 Vbias.n2192 73.1255
R13153 Vbias.n2188 Vbias.n2187 73.1255
R13154 Vbias.n2187 Vbias.n2182 73.1255
R13155 Vbias.n2185 Vbias.n2178 73.1255
R13156 Vbias.n2185 Vbias.n2183 73.1255
R13157 Vbias.n5692 Vbias.n5691 73.1255
R13158 Vbias.n5693 Vbias.n5692 73.1255
R13159 Vbias.n2174 Vbias.n2173 73.1255
R13160 Vbias.n5694 Vbias.n2174 73.1255
R13161 Vbias.n2170 Vbias.n2169 73.1255
R13162 Vbias.n2169 Vbias.n2164 73.1255
R13163 Vbias.n2167 Vbias.n2160 73.1255
R13164 Vbias.n2167 Vbias.n2165 73.1255
R13165 Vbias.n5711 Vbias.n5710 73.1255
R13166 Vbias.n5712 Vbias.n5711 73.1255
R13167 Vbias.n2156 Vbias.n2155 73.1255
R13168 Vbias.n5713 Vbias.n2156 73.1255
R13169 Vbias.n2154 Vbias.n2153 73.1255
R13170 Vbias.n2153 Vbias.n2146 73.1255
R13171 Vbias.n2145 Vbias.n2143 73.1255
R13172 Vbias.n2151 Vbias.n2145 73.1255
R13173 Vbias.n2149 Vbias.n2139 73.1255
R13174 Vbias.n2150 Vbias.n2149 73.1255
R13175 Vbias.n2138 Vbias.n2137 73.1255
R13176 Vbias.n2137 Vbias.n2135 73.1255
R13177 Vbias.n2132 Vbias.n2131 73.1255
R13178 Vbias.n2131 Vbias.n2129 73.1255
R13179 Vbias.n2128 Vbias.n2126 73.1255
R13180 Vbias.n2128 Vbias.n553 73.1255
R13181 Vbias.n7819 Vbias.n7818 73.1255
R13182 Vbias.n7820 Vbias.n7819 73.1255
R13183 Vbias.n565 Vbias.n557 73.1255
R13184 Vbias.n566 Vbias.n565 73.1255
R13185 Vbias.n568 Vbias.n559 73.1255
R13186 Vbias.n568 Vbias.n567 73.1255
R13187 Vbias.n7811 Vbias.n7810 73.1255
R13188 Vbias.n7810 Vbias.n7809 73.1255
R13189 Vbias.n7806 Vbias.n7805 73.1255
R13190 Vbias.n7805 Vbias.n7803 73.1255
R13191 Vbias.n5745 Vbias.n5742 73.1255
R13192 Vbias.n5745 Vbias.n571 73.1255
R13193 Vbias.n5753 Vbias.n5752 73.1255
R13194 Vbias.n5752 Vbias.n5751 73.1255
R13195 Vbias.n5749 Vbias.n2122 73.1255
R13196 Vbias.n5750 Vbias.n5749 73.1255
R13197 Vbias.n2121 Vbias.n2120 73.1255
R13198 Vbias.n2120 Vbias.n2118 73.1255
R13199 Vbias.n2115 Vbias.n2114 73.1255
R13200 Vbias.n2114 Vbias.n2107 73.1255
R13201 Vbias.n2106 Vbias.n2104 73.1255
R13202 Vbias.n2112 Vbias.n2106 73.1255
R13203 Vbias.n2110 Vbias.n2100 73.1255
R13204 Vbias.n2111 Vbias.n2110 73.1255
R13205 Vbias.n2099 Vbias.n2098 73.1255
R13206 Vbias.n2098 Vbias.n2094 73.1255
R13207 Vbias.n2095 Vbias.n2091 73.1255
R13208 Vbias.n2096 Vbias.n2095 73.1255
R13209 Vbias.n5781 Vbias.n2088 73.1255
R13210 Vbias.n5781 Vbias.n1674 73.1255
R13211 Vbias.n5801 Vbias.n5800 73.1255
R13212 Vbias.n5802 Vbias.n5801 73.1255
R13213 Vbias.n5799 Vbias.n5798 73.1255
R13214 Vbias.n5798 Vbias.n5791 73.1255
R13215 Vbias.n5790 Vbias.n5788 73.1255
R13216 Vbias.n5796 Vbias.n5790 73.1255
R13217 Vbias.n5794 Vbias.n2084 73.1255
R13218 Vbias.n5795 Vbias.n5794 73.1255
R13219 Vbias.n2083 Vbias.n2082 73.1255
R13220 Vbias.n2082 Vbias.n2080 73.1255
R13221 Vbias.n2077 Vbias.n2076 73.1255
R13222 Vbias.n2076 Vbias.n2074 73.1255
R13223 Vbias.n2073 Vbias.n2071 73.1255
R13224 Vbias.n2073 Vbias.n667 73.1255
R13225 Vbias.n7750 Vbias.n7749 73.1255
R13226 Vbias.n7751 Vbias.n7750 73.1255
R13227 Vbias.n7740 Vbias.n7739 73.1255
R13228 Vbias.n7739 Vbias.n677 73.1255
R13229 Vbias.n676 Vbias.n674 73.1255
R13230 Vbias.n7737 Vbias.n676 73.1255
R13231 Vbias.n5835 Vbias.n5832 73.1255
R13232 Vbias.n5835 Vbias.n678 73.1255
R13233 Vbias.n5839 Vbias.n5838 73.1255
R13234 Vbias.n5838 Vbias.n5837 73.1255
R13235 Vbias.n2065 Vbias.n2064 73.1255
R13236 Vbias.n2068 Vbias.n2065 73.1255
R13237 Vbias.n2066 Vbias.n2063 73.1255
R13238 Vbias.n2066 Vbias.n1693 73.1255
R13239 Vbias.n2061 Vbias.n1700 73.1255
R13240 Vbias.n2061 Vbias.n1694 73.1255
R13241 Vbias.n1703 Vbias.n1702 73.1255
R13242 Vbias.n2060 Vbias.n1703 73.1255
R13243 Vbias.n2058 Vbias.n2057 73.1255
R13244 Vbias.n2059 Vbias.n2058 73.1255
R13245 Vbias.n1711 Vbias.n1707 73.1255
R13246 Vbias.n1711 Vbias.n1530 73.1255
R13247 Vbias.n1722 Vbias.n1721 73.1255
R13248 Vbias.n1723 Vbias.n1722 73.1255
R13249 Vbias.n1720 Vbias.n1719 73.1255
R13250 Vbias.n1725 Vbias.n1720 73.1255
R13251 Vbias.n1739 Vbias.n1736 73.1255
R13252 Vbias.n1739 Vbias.n1529 73.1255
R13253 Vbias.n1740 Vbias.n1735 73.1255
R13254 Vbias.n1740 Vbias.n1724 73.1255
R13255 Vbias.n2041 Vbias.n2040 73.1255
R13256 Vbias.n2040 Vbias.n2039 73.1255
R13257 Vbias.n2037 Vbias.n2036 73.1255
R13258 Vbias.n2037 Vbias.n1467 73.1255
R13259 Vbias.n6748 Vbias.n6747 73.1255
R13260 Vbias.n6749 Vbias.n6748 73.1255
R13261 Vbias.n6725 Vbias.n1448 73.1255
R13262 Vbias.n6726 Vbias.n6725 73.1255
R13263 Vbias.n6728 Vbias.n6719 73.1255
R13264 Vbias.n6728 Vbias.n6727 73.1255
R13265 Vbias.n6734 Vbias.n6721 73.1255
R13266 Vbias.n6735 Vbias.n6734 73.1255
R13267 Vbias.n6739 Vbias.n6738 73.1255
R13268 Vbias.n6738 Vbias.n6737 73.1255
R13269 Vbias.n6702 Vbias.n6695 73.1255
R13270 Vbias.n6702 Vbias.n6701 73.1255
R13271 Vbias.n6708 Vbias.n6697 73.1255
R13272 Vbias.n6709 Vbias.n6708 73.1255
R13273 Vbias.n6712 Vbias.n6711 73.1255
R13274 Vbias.n6711 Vbias.n6710 73.1255
R13275 Vbias.n6689 Vbias.n6688 73.1255
R13276 Vbias.n6688 Vbias.n1443 73.1255
R13277 Vbias.n6685 Vbias.n6684 73.1255
R13278 Vbias.n6686 Vbias.n6685 73.1255
R13279 Vbias.n6680 Vbias.n1455 73.1255
R13280 Vbias.n6680 Vbias.n6679 73.1255
R13281 Vbias.n8074 Vbias.n8073 73.1255
R13282 Vbias.n8075 Vbias.n8074 73.1255
R13283 Vbias.n21 Vbias.n14 73.1255
R13284 Vbias.n21 Vbias.n19 73.1255
R13285 Vbias.n26 Vbias.n25 73.1255
R13286 Vbias.n25 Vbias.n20 73.1255
R13287 Vbias.n28 Vbias.n27 73.1255
R13288 Vbias.n29 Vbias.n28 73.1255
R13289 Vbias.n38 Vbias.n31 73.1255
R13290 Vbias.n38 Vbias.n37 73.1255
R13291 Vbias.n8056 Vbias.n8055 73.1255
R13292 Vbias.n8055 Vbias.n8054 73.1255
R13293 Vbias.n48 Vbias.n44 73.1255
R13294 Vbias.n48 Vbias.n41 73.1255
R13295 Vbias.n46 Vbias.n45 73.1255
R13296 Vbias.n47 Vbias.n46 73.1255
R13297 Vbias.n55 Vbias.n51 73.1255
R13298 Vbias.n56 Vbias.n55 73.1255
R13299 Vbias.n8042 Vbias.n8041 73.1255
R13300 Vbias.n8041 Vbias.n8040 73.1255
R13301 Vbias.n8038 Vbias.n8037 73.1255
R13302 Vbias.n8039 Vbias.n8038 73.1255
R13303 Vbias.n8028 Vbias.n8027 73.1255
R13304 Vbias.n8027 Vbias.n65 73.1255
R13305 Vbias.n64 Vbias.n62 73.1255
R13306 Vbias.n8025 Vbias.n64 73.1255
R13307 Vbias.n8023 Vbias.n8022 73.1255
R13308 Vbias.n8024 Vbias.n8023 73.1255
R13309 Vbias.n80 Vbias.n79 73.1255
R13310 Vbias.n79 Vbias.n75 73.1255
R13311 Vbias.n83 Vbias.n82 73.1255
R13312 Vbias.n82 Vbias.n76 73.1255
R13313 Vbias.n85 Vbias.n84 73.1255
R13314 Vbias.n8009 Vbias.n85 73.1255
R13315 Vbias.n8006 Vbias.n8005 73.1255
R13316 Vbias.n8007 Vbias.n8006 73.1255
R13317 Vbias.n8003 Vbias.n8002 73.1255
R13318 Vbias.n8002 Vbias.n8001 73.1255
R13319 Vbias.n7999 Vbias.n7998 73.1255
R13320 Vbias.n8000 Vbias.n7999 73.1255
R13321 Vbias.n99 Vbias.n93 73.1255
R13322 Vbias.n99 Vbias.n97 73.1255
R13323 Vbias.n105 Vbias.n104 73.1255
R13324 Vbias.n104 Vbias.n98 73.1255
R13325 Vbias.n108 Vbias.n107 73.1255
R13326 Vbias.n7986 Vbias.n108 73.1255
R13327 Vbias.n7984 Vbias.n7983 73.1255
R13328 Vbias.n7985 Vbias.n7984 73.1255
R13329 Vbias.n118 Vbias.n112 73.1255
R13330 Vbias.n118 Vbias.n116 73.1255
R13331 Vbias.n126 Vbias.n125 73.1255
R13332 Vbias.n125 Vbias.n117 73.1255
R13333 Vbias.n129 Vbias.n128 73.1255
R13334 Vbias.n7971 Vbias.n129 73.1255
R13335 Vbias.n7969 Vbias.n7968 73.1255
R13336 Vbias.n7970 Vbias.n7969 73.1255
R13337 Vbias.n139 Vbias.n133 73.1255
R13338 Vbias.n139 Vbias.n137 73.1255
R13339 Vbias.n136 Vbias.n134 73.1255
R13340 Vbias.n138 Vbias.n136 73.1255
R13341 Vbias.n156 Vbias.n145 73.1255
R13342 Vbias.n157 Vbias.n156 73.1255
R13343 Vbias.n153 Vbias.n147 73.1255
R13344 Vbias.n153 Vbias.n151 73.1255
R13345 Vbias.n162 Vbias.n161 73.1255
R13346 Vbias.n161 Vbias.n152 73.1255
R13347 Vbias.n164 Vbias.n163 73.1255
R13348 Vbias.n165 Vbias.n164 73.1255
R13349 Vbias.n4683 Vbias.n2603 73.1255
R13350 Vbias.n4684 Vbias.n4683 73.1255
R13351 Vbias.n4991 Vbias.n4990 73.1255
R13352 Vbias.n4992 Vbias.n4991 73.1255
R13353 Vbias.n2598 Vbias.n2597 73.1255
R13354 Vbias.n4993 Vbias.n2598 73.1255
R13355 Vbias.n4997 Vbias.n4996 73.1255
R13356 Vbias.n4996 Vbias.n4994 73.1255
R13357 Vbias.n5008 Vbias.n5007 73.1255
R13358 Vbias.n5009 Vbias.n5008 73.1255
R13359 Vbias.n5013 Vbias.n2586 73.1255
R13360 Vbias.n5013 Vbias.n5012 73.1255
R13361 Vbias.n5024 Vbias.n5023 73.1255
R13362 Vbias.n5023 Vbias.n5022 73.1255
R13363 Vbias.n5019 Vbias.n5018 73.1255
R13364 Vbias.n5018 Vbias.n5016 73.1255
R13365 Vbias.n5551 Vbias.n5550 73.1255
R13366 Vbias.n5552 Vbias.n5551 73.1255
R13367 Vbias.n2240 Vbias.n2232 73.1255
R13368 Vbias.n2241 Vbias.n2240 73.1255
R13369 Vbias.n2243 Vbias.n2234 73.1255
R13370 Vbias.n2243 Vbias.n2242 73.1255
R13371 Vbias.n5543 Vbias.n5542 73.1255
R13372 Vbias.n5542 Vbias.n5541 73.1255
R13373 Vbias.n5538 Vbias.n5537 73.1255
R13374 Vbias.n5537 Vbias.n5535 73.1255
R13375 Vbias.n5531 Vbias.n5530 73.1255
R13376 Vbias.n5532 Vbias.n5531 73.1255
R13377 Vbias.n5521 Vbias.n5520 73.1255
R13378 Vbias.n5520 Vbias.n5518 73.1255
R13379 Vbias.n5517 Vbias.n5515 73.1255
R13380 Vbias.n5517 Vbias.n1673 73.1255
R13381 Vbias.n5875 Vbias.n5874 73.1255
R13382 Vbias.n5876 Vbias.n5875 73.1255
R13383 Vbias.n1687 Vbias.n1678 73.1255
R13384 Vbias.n1688 Vbias.n1687 73.1255
R13385 Vbias.n1690 Vbias.n1681 73.1255
R13386 Vbias.n1690 Vbias.n1689 73.1255
R13387 Vbias.n5867 Vbias.n5866 73.1255
R13388 Vbias.n5866 Vbias.n5865 73.1255
R13389 Vbias.n5862 Vbias.n5861 73.1255
R13390 Vbias.n5861 Vbias.n5859 73.1255
R13391 Vbias.n4260 Vbias.n4256 73.1255
R13392 Vbias.n4261 Vbias.n4260 73.1255
R13393 Vbias.n4264 Vbias.n4263 73.1255
R13394 Vbias.n4263 Vbias.n4262 73.1255
R13395 Vbias.n2881 Vbias.n2880 73.1255
R13396 Vbias.n2883 Vbias.n2881 73.1255
R13397 Vbias.n2884 Vbias.n2879 73.1255
R13398 Vbias.n2884 Vbias.n2874 73.1255
R13399 Vbias.n4285 Vbias.n4284 73.1255
R13400 Vbias.n4284 Vbias.n2866 73.1255
R13401 Vbias.n4279 Vbias.n4278 73.1255
R13402 Vbias.n4278 Vbias.n2868 73.1255
R13403 Vbias.n2847 Vbias.n2846 73.1255
R13404 Vbias.n2849 Vbias.n2847 73.1255
R13405 Vbias.n2850 Vbias.n2845 73.1255
R13406 Vbias.n2850 Vbias.n2840 73.1255
R13407 Vbias.n4318 Vbias.n4317 73.1255
R13408 Vbias.n4317 Vbias.n2830 73.1255
R13409 Vbias.n4312 Vbias.n4311 73.1255
R13410 Vbias.n4311 Vbias.n2834 73.1255
R13411 Vbias.n4344 Vbias.n2819 73.1255
R13412 Vbias.n4344 Vbias.n4343 73.1255
R13413 Vbias.n4351 Vbias.n4350 73.1255
R13414 Vbias.n4352 Vbias.n4351 73.1255
R13415 Vbias.n2806 Vbias.n2802 73.1255
R13416 Vbias.n4364 Vbias.n2802 73.1255
R13417 Vbias.n2801 Vbias.n2800 73.1255
R13418 Vbias.n4365 Vbias.n2801 73.1255
R13419 Vbias.n4375 Vbias.n4374 73.1255
R13420 Vbias.n4374 Vbias.n2786 73.1255
R13421 Vbias.n4388 Vbias.n2783 73.1255
R13422 Vbias.n2790 Vbias.n2783 73.1255
R13423 Vbias.n4402 Vbias.n2777 73.1255
R13424 Vbias.n4406 Vbias.n2777 73.1255
R13425 Vbias.n4271 Vbias.n2888 73.1255
R13426 Vbias.n2888 Vbias.n2883 73.1255
R13427 Vbias.n2891 Vbias.n2890 73.1255
R13428 Vbias.n2890 Vbias.n2874 73.1255
R13429 Vbias.n2871 Vbias.n2870 73.1255
R13430 Vbias.n2870 Vbias.n2866 73.1255
R13431 Vbias.n4294 Vbias.n2865 73.1255
R13432 Vbias.n2868 Vbias.n2865 73.1255
R13433 Vbias.n4304 Vbias.n2854 73.1255
R13434 Vbias.n2854 Vbias.n2849 73.1255
R13435 Vbias.n2857 Vbias.n2856 73.1255
R13436 Vbias.n2856 Vbias.n2840 73.1255
R13437 Vbias.n2837 Vbias.n2836 73.1255
R13438 Vbias.n2836 Vbias.n2830 73.1255
R13439 Vbias.n4327 Vbias.n2829 73.1255
R13440 Vbias.n2834 Vbias.n2829 73.1255
R13441 Vbias.n2832 Vbias.n2823 73.1255
R13442 Vbias.n2833 Vbias.n2832 73.1255
R13443 Vbias.n4337 Vbias.n4336 73.1255
R13444 Vbias.n4338 Vbias.n4337 73.1255
R13445 Vbias.n4342 Vbias.n4341 73.1255
R13446 Vbias.n4343 Vbias.n4342 73.1255
R13447 Vbias.n4354 Vbias.n4353 73.1255
R13448 Vbias.n4353 Vbias.n4352 73.1255
R13449 Vbias.n4363 Vbias.n4362 73.1255
R13450 Vbias.n4364 Vbias.n4363 73.1255
R13451 Vbias.n4367 Vbias.n4366 73.1255
R13452 Vbias.n4366 Vbias.n4365 73.1255
R13453 Vbias.n4379 Vbias.n4378 73.1255
R13454 Vbias.n4378 Vbias.n2786 73.1255
R13455 Vbias.n4394 Vbias.n4393 73.1255
R13456 Vbias.n4393 Vbias.n2790 73.1255
R13457 Vbias.n4405 Vbias.n4404 73.1255
R13458 Vbias.n4406 Vbias.n4405 73.1255
R13459 Vbias.n6101 Vbias.n1529 71.34
R13460 Vbias.n6676 Vbias.n1467 71.34
R13461 Vbias.n2031 Vbias.t342 69.8913
R13462 Vbias.n2024 Vbias.t595 69.8913
R13463 Vbias.n2019 Vbias.t854 69.8913
R13464 Vbias.n1824 Vbias.t764 69.8913
R13465 Vbias.n1829 Vbias.t423 69.8913
R13466 Vbias.n1834 Vbias.t645 69.8913
R13467 Vbias.n1839 Vbias.t359 69.8913
R13468 Vbias.n1844 Vbias.t561 69.8913
R13469 Vbias.n1847 Vbias 68.0603
R13470 Vbias.n4891 Vbias.n4890 65.6517
R13471 Vbias.n6677 Vbias.t52 65.5144
R13472 Vbias.n6101 Vbias.n1530 65.3176
R13473 Vbias.n6101 Vbias.n1531 62.4595
R13474 Vbias.n4267 Vbias.t85 61.1579
R13475 Vbias.n4267 Vbias.t725 61.1579
R13476 Vbias.n4300 Vbias.t168 61.1579
R13477 Vbias.n4300 Vbias.t433 61.1579
R13478 Vbias.n4333 Vbias.t638 61.1579
R13479 Vbias.n2809 Vbias.t295 61.1579
R13480 Vbias.n2809 Vbias.t129 61.1579
R13481 Vbias.n2796 Vbias.t841 61.1579
R13482 Vbias.n2796 Vbias.t508 61.1579
R13483 Vbias.n4255 Vbias.t838 61.1579
R13484 Vbias.n5052 Vbias.t242 61.1579
R13485 Vbias.n5073 Vbias.t641 61.1579
R13486 Vbias.n5074 Vbias.t386 61.1579
R13487 Vbias.n5095 Vbias.t272 61.1579
R13488 Vbias.n5115 Vbias.t57 61.1579
R13489 Vbias.n5175 Vbias.t221 61.1579
R13490 Vbias.n5161 Vbias.t687 61.1579
R13491 Vbias.n5162 Vbias.t587 61.1579
R13492 Vbias.n2253 Vbias.t260 61.1579
R13493 Vbias.n2293 Vbias.t101 61.1579
R13494 Vbias.n5440 Vbias.t179 61.1579
R13495 Vbias.n5441 Vbias.t12 61.1579
R13496 Vbias.n5457 Vbias.t396 61.1579
R13497 Vbias.n5892 Vbias.t238 61.1579
R13498 Vbias.n5912 Vbias.t27 61.1579
R13499 Vbias.n5948 Vbias.t213 61.1579
R13500 Vbias.n1620 Vbias.t751 61.1579
R13501 Vbias.n6095 Vbias.t816 61.1579
R13502 Vbias.n6087 Vbias.t183 61.1579
R13503 Vbias.n6079 Vbias.t77 61.1579
R13504 Vbias.n6806 Vbias.t268 61.1579
R13505 Vbias.n1420 Vbias.t491 61.1579
R13506 Vbias.n6793 Vbias.t331 61.1579
R13507 Vbias.n6785 Vbias.t266 61.1579
R13508 Vbias.n7009 Vbias.t93 61.1579
R13509 Vbias.n7031 Vbias.t240 61.1579
R13510 Vbias.n7048 Vbias.t543 61.1579
R13511 Vbias.n7061 Vbias.t382 61.1579
R13512 Vbias.n7078 Vbias.t199 61.1579
R13513 Vbias.n7095 Vbias.t115 61.1579
R13514 Vbias.n7137 Vbias.t33 61.1579
R13515 Vbias.n7154 Vbias.t846 61.1579
R13516 Vbias.n7167 Vbias.t499 61.1579
R13517 Vbias.n7184 Vbias.t63 61.1579
R13518 Vbias.n7201 Vbias.t177 61.1579
R13519 Vbias.n7203 Vbias.t689 61.1579
R13520 Vbias.n7205 Vbias.t105 61.1579
R13521 Vbias.n1211 Vbias.t256 61.1579
R13522 Vbias.n1243 Vbias.t316 61.1579
R13523 Vbias.n1194 Vbias.t189 61.1579
R13524 Vbias.n7099 Vbias.t510 61.1579
R13525 Vbias.n7101 Vbias.t197 61.1579
R13526 Vbias.n6944 Vbias.t67 61.1579
R13527 Vbias.n6976 Vbias.t535 61.1579
R13528 Vbias.n6927 Vbias.t41 61.1579
R13529 Vbias.n6899 Vbias.t421 61.1579
R13530 Vbias.n6880 Vbias.t223 61.1579
R13531 Vbias.n6857 Vbias.t123 61.1579
R13532 Vbias.n6834 Vbias.t489 61.1579
R13533 Vbias.n6833 Vbias.t119 61.1579
R13534 Vbias.n6023 Vbias.t729 61.1579
R13535 Vbias.n6025 Vbias.t244 61.1579
R13536 Vbias.n5999 Vbias.t95 61.1579
R13537 Vbias.n5976 Vbias.t319 61.1579
R13538 Vbias.n5975 Vbias.t61 61.1579
R13539 Vbias.n5341 Vbias.t743 61.1579
R13540 Vbias.n5335 Vbias.t195 61.1579
R13541 Vbias.n5333 Vbias.t23 61.1579
R13542 Vbias.n5384 Vbias.t405 61.1579
R13543 Vbias.n5298 Vbias.t99 61.1579
R13544 Vbias.n5269 Vbias.t708 61.1579
R13545 Vbias.n5249 Vbias.t217 61.1579
R13546 Vbias.n5226 Vbias.t29 61.1579
R13547 Vbias.n5203 Vbias.t665 61.1579
R13548 Vbias.n5202 Vbias.t55 61.1579
R13549 Vbias.n2509 Vbias.t602 61.1579
R13550 Vbias.n2503 Vbias.t264 61.1579
R13551 Vbias.n2501 Vbias.t109 61.1579
R13552 Vbias.n2552 Vbias.t691 61.1579
R13553 Vbias.n2466 Vbias.t39 61.1579
R13554 Vbias.n4484 Vbias.t825 61.1579
R13555 Vbias.n4496 Vbias.t181 61.1579
R13556 Vbias.n4510 Vbias.t59 61.1579
R13557 Vbias.n4524 Vbias.t301 61.1579
R13558 Vbias.n4423 Vbias.t111 61.1579
R13559 Vbias.n3721 Vbias.t459 61.1579
R13560 Vbias.n3721 Vbias.t563 61.1579
R13561 Vbias.n3750 Vbias.t352 61.1579
R13562 Vbias.n3750 Vbias.t676 61.1579
R13563 Vbias.n3776 Vbias.t451 61.1579
R13564 Vbias.n3888 Vbias.t125 61.1579
R13565 Vbias.n3888 Vbias.t412 61.1579
R13566 Vbias.n3797 Vbias.t618 61.1579
R13567 Vbias.n3797 Vbias.t525 61.1579
R13568 Vbias.n3976 Vbias.t652 61.1579
R13569 Vbias.n3183 Vbias.t844 61.1579
R13570 Vbias.n3183 Vbias.t551 61.1579
R13571 Vbias.n3212 Vbias.t375 61.1579
R13572 Vbias.n3212 Vbias.t891 61.1579
R13573 Vbias.n3238 Vbias.t388 61.1579
R13574 Vbias.n3350 Vbias.t597 61.1579
R13575 Vbias.n3350 Vbias.t584 61.1579
R13576 Vbias.n3259 Vbias.t887 61.1579
R13577 Vbias.n3259 Vbias.t882 61.1579
R13578 Vbias.n3438 Vbias.t878 61.1579
R13579 Vbias.n3452 Vbias.t171 61.1579
R13580 Vbias.n3452 Vbias.t617 61.1579
R13581 Vbias.n3481 Vbias.t553 61.1579
R13582 Vbias.n3481 Vbias.t463 61.1579
R13583 Vbias.n3507 Vbias.t810 61.1579
R13584 Vbias.n3619 Vbias.t149 61.1579
R13585 Vbias.n3619 Vbias.t434 61.1579
R13586 Vbias.n3528 Vbias.t610 61.1579
R13587 Vbias.n3528 Vbias.t879 61.1579
R13588 Vbias.n3707 Vbias.t836 61.1579
R13589 Vbias.n4251 Vbias.t880 61.1579
R13590 Vbias.n4011 Vbias.t83 61.1579
R13591 Vbias.n4036 Vbias.t504 61.1579
R13592 Vbias.n4213 Vbias.t290 61.1579
R13593 Vbias.n4053 Vbias.t37 61.1579
R13594 Vbias.n4165 Vbias.t562 61.1579
R13595 Vbias.n4142 Vbias.t698 61.1579
R13596 Vbias.n4126 Vbias.t771 61.1579
R13597 Vbias.n4113 Vbias.t529 61.1579
R13598 Vbias.n4102 Vbias.t574 61.1579
R13599 Vbias.n2913 Vbias.t169 61.1579
R13600 Vbias.n2913 Vbias.t138 61.1579
R13601 Vbias.n2942 Vbias.t727 61.1579
R13602 Vbias.n2942 Vbias.t843 61.1579
R13603 Vbias.n2968 Vbias.t872 61.1579
R13604 Vbias.n3080 Vbias.t519 61.1579
R13605 Vbias.n3080 Vbias.t281 61.1579
R13606 Vbias.n2989 Vbias.t613 61.1579
R13607 Vbias.n2989 Vbias.t166 61.1579
R13608 Vbias.n3168 Vbias.t834 61.1579
R13609 Vbias.n2674 Vbias.t512 61.1579
R13610 Vbias.n2674 Vbias.t228 61.1579
R13611 Vbias.n2703 Vbias.t134 61.1579
R13612 Vbias.n2703 Vbias.t530 61.1579
R13613 Vbias.n2729 Vbias.t447 61.1579
R13614 Vbias.n4756 Vbias.t349 61.1579
R13615 Vbias.n4756 Vbias.t516 61.1579
R13616 Vbias.n2750 Vbias.t709 61.1579
R13617 Vbias.n2750 Vbias.t461 61.1579
R13618 Vbias.n2898 Vbias.t876 61.1579
R13619 Vbias.n4578 Vbias.t270 61.1579
R13620 Vbias.n4579 Vbias.t453 61.1579
R13621 Vbias.n4655 Vbias.t335 61.1579
R13622 Vbias.n4647 Vbias.t215 61.1579
R13623 Vbias.n5031 Vbias.t43 61.1579
R13624 Vbias.n7466 Vbias.t65 61.1579
R13625 Vbias.n7346 Vbias.t193 61.1579
R13626 Vbias.n7366 Vbias.t589 61.1579
R13627 Vbias.n7428 Vbias.t668 61.1579
R13628 Vbias.n7384 Vbias.t252 61.1579
R13629 Vbias.n6649 Vbias.t75 61.1579
R13630 Vbias.n6634 Vbias.t225 61.1579
R13631 Vbias.n6626 Vbias.t384 61.1579
R13632 Vbias.n6192 Vbias.t734 61.1579
R13633 Vbias.n6206 Vbias.t187 61.1579
R13634 Vbias.n6575 Vbias.t89 61.1579
R13635 Vbias.n6567 Vbias.t278 61.1579
R13636 Vbias.n6559 Vbias.t484 61.1579
R13637 Vbias.n6429 Vbias.t345 61.1579
R13638 Vbias.n6443 Vbias.t232 61.1579
R13639 Vbias.n7588 Vbias.t121 61.1579
R13640 Vbias.n7580 Vbias.t250 61.1579
R13641 Vbias.n7572 Vbias.t338 61.1579
R13642 Vbias.n883 Vbias.t808 61.1579
R13643 Vbias.n897 Vbias.t205 61.1579
R13644 Vbias.n7276 Vbias.t117 61.1579
R13645 Vbias.n7239 Vbias.t144 61.1579
R13646 Vbias.n1063 Vbias.t69 61.1579
R13647 Vbias.n1042 Vbias.t262 61.1579
R13648 Vbias.n7322 Vbias.t478 61.1579
R13649 Vbias.n7482 Vbias.t49 61.1579
R13650 Vbias.n989 Vbias.t572 61.1579
R13651 Vbias.n968 Vbias.t17 61.1579
R13652 Vbias.n947 Vbias.t209 61.1579
R13653 Vbias.n945 Vbias.t157 61.1579
R13654 Vbias.n7604 Vbias.t35 61.1579
R13655 Vbias.n834 Vbias.t565 61.1579
R13656 Vbias.n813 Vbias.t97 61.1579
R13657 Vbias.n6360 Vbias.t234 61.1579
R13658 Vbias.n6362 Vbias.t367 61.1579
R13659 Vbias.n6242 Vbias.t79 61.1579
R13660 Vbias.n6341 Vbias.t465 61.1579
R13661 Vbias.n6327 Vbias.t19 61.1579
R13662 Vbias.n6313 Vbias.t254 61.1579
R13663 Vbias.n6297 Vbias.t612 61.1579
R13664 Vbias.n6665 Vbias.t53 61.1579
R13665 Vbias.n1718 Vbias.t294 61.1579
R13666 Vbias.n1716 Vbias.t31 61.1579
R13667 Vbias.n5842 Vbias.t203 61.1579
R13668 Vbias.n5831 Vbias.t785 61.1579
R13669 Vbias.n5813 Vbias.t107 61.1579
R13670 Vbias.n5785 Vbias.t683 61.1579
R13671 Vbias.n5770 Vbias.t103 61.1579
R13672 Vbias.n5756 Vbias.t175 61.1579
R13673 Vbias.n5741 Vbias.t822 61.1579
R13674 Vbias.n5724 Vbias.t81 61.1579
R13675 Vbias.n5700 Vbias.t152 61.1579
R13676 Vbias.n2172 Vbias.t45 61.1579
R13677 Vbias.n2190 Vbias.t211 61.1579
R13678 Vbias.n5667 Vbias.t773 61.1579
R13679 Vbias.n5650 Vbias.t73 61.1579
R13680 Vbias.n5626 Vbias.t432 61.1579
R13681 Vbias.n5569 Vbias.t91 61.1579
R13682 Vbias.n5587 Vbias.t236 61.1579
R13683 Vbias.n5593 Vbias.t416 61.1579
R13684 Vbias.n7960 Vbias.t21 61.1579
R13685 Vbias.n142 Vbias.t357 61.1579
R13686 Vbias.n122 Vbias.t47 61.1579
R13687 Vbias.n250 Vbias.t258 61.1579
R13688 Vbias.n252 Vbias.t792 61.1579
R13689 Vbias.n256 Vbias.t71 61.1579
R13690 Vbias.n273 Vbias.t207 61.1579
R13691 Vbias.n292 Vbias.t864 61.1579
R13692 Vbias.n293 Vbias.t803 61.1579
R13693 Vbias.n312 Vbias.t248 61.1579
R13694 Vbias.n356 Vbias.t87 61.1579
R13695 Vbias.n380 Vbias.t173 61.1579
R13696 Vbias.n404 Vbias.t591 61.1579
R13697 Vbias.n7907 Vbias.t321 61.1579
R13698 Vbias.n427 Vbias.t191 61.1579
R13699 Vbias.n462 Vbias.t113 61.1579
R13700 Vbias.n486 Vbias.t219 61.1579
R13701 Vbias.n510 Vbias.t398 61.1579
R13702 Vbias.n7841 Vbias.t890 61.1579
R13703 Vbias.n533 Vbias.t185 61.1579
R13704 Vbias.n576 Vbias.t51 61.1579
R13705 Vbias.n600 Vbias.t276 61.1579
R13706 Vbias.n624 Vbias.t818 61.1579
R13707 Vbias.n7772 Vbias.t856 61.1579
R13708 Vbias.n647 Vbias.t274 61.1579
R13709 Vbias.n5827 Vbias.t25 61.1579
R13710 Vbias.n7720 Vbias.t246 61.1579
R13711 Vbias.n7705 Vbias.t333 61.1579
R13712 Vbias.n730 Vbias.t672 61.1579
R13713 Vbias.n739 Vbias.t201 61.1579
R13714 Vbias.n6126 Vbias.t616 61.1579
R13715 Vbias.n7659 Vbias.t482 61.1579
R13716 Vbias.n6511 Vbias.t15 61.1579
R13717 Vbias.n6512 Vbias.t369 61.1579
R13718 Vbias.n7536 Vbias.t329 61.1579
R13719 Vbias.n7538 Vbias.t718 61.1579
R13720 Vbias.n169 Vbias.t812 61.1579
R13721 Vbias.n452 Vbias.t768 61.1579
R13722 Vbias.n7815 Vbias.t629 61.1579
R13723 Vbias.n672 Vbias.t486 61.1579
R13724 Vbias.n673 Vbias.t714 61.1579
R13725 Vbias.n327 Vbias.t622 61.1579
R13726 Vbias.n2584 Vbias.t830 61.1579
R13727 Vbias.n5547 Vbias.t656 61.1579
R13728 Vbias.n5513 Vbias.t720 61.1579
R13729 Vbias.n5514 Vbias.t136 61.1579
R13730 Vbias.n5871 Vbias.t371 61.1579
R13731 Vbias.n1679 Vbias.t8 61.1579
R13732 Vbias.n6692 Vbias.t724 61.1579
R13733 Vbias.n6744 Vbias.t761 61.1579
R13734 Vbias.n6717 Vbias.t738 61.1579
R13735 Vbias.n6693 Vbias.t678 61.1579
R13736 Vbias.n4987 Vbias.t740 61.1579
R13737 Vbias.n5004 Vbias.t701 61.1579
R13738 Vbias.n4969 Vbias.t827 61.1579
R13739 Vbias.n4943 Vbias.t425 61.1579
R13740 Vbias.n2643 Vbias.t832 61.1579
R13741 Vbias.n2657 Vbias.t527 61.1579
R13742 Vbias.n2895 Vbias.t840 61.1579
R13743 Vbias.n3171 Vbias.t159 61.1579
R13744 Vbias.n8060 Vbias.t675 61.1579
R13745 Vbias.n8045 Vbias.t324 61.1579
R13746 Vbias.n61 Vbias.t419 61.1579
R13747 Vbias.n70 Vbias.t523 61.1579
R13748 Vbias Vbias.t428 61.1525
R13749 Vbias Vbias.t794 61.1525
R13750 Vbias.n1734 Vbias.t558 61.1525
R13751 Vbias Vbias.t141 61.1525
R13752 Vbias Vbias.t663 61.1525
R13753 Vbias Vbias.t747 61.1525
R13754 Vbias Vbias.t869 61.1525
R13755 Vbias Vbias.t759 61.1525
R13756 Vbias.n7266 Vbias.n7265 59.792
R13757 Vbias.n349 Vbias.n348 59.5094
R13758 Vbias.n7938 Vbias.n7937 59.5094
R13759 Vbias.n7887 Vbias.n7886 59.5094
R13760 Vbias.n7872 Vbias.n7871 59.5094
R13761 Vbias.n7821 Vbias.n7820 59.5094
R13762 Vbias.n7803 Vbias.n7802 59.5094
R13763 Vbias.n7752 Vbias.n7751 59.5094
R13764 Vbias.n7737 Vbias.n7736 59.5094
R13765 Vbias.n1881 Vbias 58.3538
R13766 Vbias.n6751 Vbias.n6750 54.9156
R13767 Vbias.n6736 Vbias.n1305 54.9156
R13768 Vbias.n5553 Vbias.n2228 54.9156
R13769 Vbias.n5534 Vbias.n5533 54.9156
R13770 Vbias.n5878 Vbias.n5877 54.9156
R13771 Vbias.n8010 Vbias.n72 52.5417
R13772 Vbias.n8018 Vbias.n72 52.5417
R13773 Vbias.n8018 Vbias.n69 52.5417
R13774 Vbias.n8021 Vbias.n69 52.5417
R13775 Vbias.n8033 Vbias.n60 52.5417
R13776 Vbias.n8036 Vbias.n60 52.5417
R13777 Vbias.n8047 Vbias.n50 52.5417
R13778 Vbias.n50 Vbias.n33 52.5417
R13779 Vbias.n8057 Vbias.n33 52.5417
R13780 Vbias.n8058 Vbias.n8057 52.5417
R13781 Vbias.n5006 Vbias.n2596 52.5417
R13782 Vbias.n5002 Vbias.n2596 52.5417
R13783 Vbias.n6714 Vbias.n6713 52.5417
R13784 Vbias.n6715 Vbias.n6714 52.5417
R13785 Vbias.n6741 Vbias.n6740 52.5417
R13786 Vbias.n6742 Vbias.n6741 52.5417
R13787 Vbias.n7745 Vbias.n671 52.5417
R13788 Vbias.n7748 Vbias.n671 52.5417
R13789 Vbias.n7812 Vbias.n561 52.5417
R13790 Vbias.n7813 Vbias.n7812 52.5417
R13791 Vbias.n7880 Vbias.n451 52.5417
R13792 Vbias.n7883 Vbias.n451 52.5417
R13793 Vbias.n338 Vbias.n170 52.5417
R13794 Vbias.n7941 Vbias.n170 52.5417
R13795 Vbias.n7541 Vbias.n7540 52.5417
R13796 Vbias.n7541 Vbias.n921 52.5417
R13797 Vbias.n7534 Vbias.n925 52.5417
R13798 Vbias.n6523 Vbias.n925 52.5417
R13799 Vbias.n7656 Vbias.n7655 52.5417
R13800 Vbias.n7657 Vbias.n7656 52.5417
R13801 Vbias.n7661 Vbias.n768 52.5417
R13802 Vbias.n769 Vbias.n768 52.5417
R13803 Vbias.n7670 Vbias.n741 52.5417
R13804 Vbias.n7678 Vbias.n741 52.5417
R13805 Vbias.n7678 Vbias.n738 52.5417
R13806 Vbias.n7681 Vbias.n738 52.5417
R13807 Vbias.n7693 Vbias.n729 52.5417
R13808 Vbias.n7696 Vbias.n729 52.5417
R13809 Vbias.n7707 Vbias.n719 52.5417
R13810 Vbias.n719 Vbias.n702 52.5417
R13811 Vbias.n7717 Vbias.n702 52.5417
R13812 Vbias.n7718 Vbias.n7717 52.5417
R13813 Vbias.n7757 Vbias.n7756 52.5417
R13814 Vbias.n7758 Vbias.n7757 52.5417
R13815 Vbias.n7758 Vbias.n646 52.5417
R13816 Vbias.n7761 Vbias.n646 52.5417
R13817 Vbias.n7769 Vbias.n7768 52.5417
R13818 Vbias.n7770 Vbias.n7769 52.5417
R13819 Vbias.n7782 Vbias.n7781 52.5417
R13820 Vbias.n7783 Vbias.n7782 52.5417
R13821 Vbias.n7783 Vbias.n599 52.5417
R13822 Vbias.n7786 Vbias.n599 52.5417
R13823 Vbias.n7794 Vbias.n7793 52.5417
R13824 Vbias.n7795 Vbias.n7794 52.5417
R13825 Vbias.n7795 Vbias.n575 52.5417
R13826 Vbias.n7798 Vbias.n575 52.5417
R13827 Vbias.n7826 Vbias.n7825 52.5417
R13828 Vbias.n7827 Vbias.n7826 52.5417
R13829 Vbias.n7827 Vbias.n532 52.5417
R13830 Vbias.n7830 Vbias.n532 52.5417
R13831 Vbias.n7838 Vbias.n7837 52.5417
R13832 Vbias.n7839 Vbias.n7838 52.5417
R13833 Vbias.n7851 Vbias.n7850 52.5417
R13834 Vbias.n7852 Vbias.n7851 52.5417
R13835 Vbias.n7852 Vbias.n485 52.5417
R13836 Vbias.n7855 Vbias.n485 52.5417
R13837 Vbias.n7863 Vbias.n7862 52.5417
R13838 Vbias.n7864 Vbias.n7863 52.5417
R13839 Vbias.n7864 Vbias.n461 52.5417
R13840 Vbias.n7867 Vbias.n461 52.5417
R13841 Vbias.n7892 Vbias.n7891 52.5417
R13842 Vbias.n7893 Vbias.n7892 52.5417
R13843 Vbias.n7893 Vbias.n426 52.5417
R13844 Vbias.n7896 Vbias.n426 52.5417
R13845 Vbias.n7904 Vbias.n7903 52.5417
R13846 Vbias.n7905 Vbias.n7904 52.5417
R13847 Vbias.n7917 Vbias.n7916 52.5417
R13848 Vbias.n7918 Vbias.n7917 52.5417
R13849 Vbias.n7918 Vbias.n379 52.5417
R13850 Vbias.n7921 Vbias.n379 52.5417
R13851 Vbias.n7929 Vbias.n7928 52.5417
R13852 Vbias.n7930 Vbias.n7929 52.5417
R13853 Vbias.n7930 Vbias.n178 52.5417
R13854 Vbias.n7933 Vbias.n178 52.5417
R13855 Vbias.n353 Vbias.n180 52.5417
R13856 Vbias.n196 Vbias.n180 52.5417
R13857 Vbias.n197 Vbias.n196 52.5417
R13858 Vbias.n314 Vbias.n197 52.5417
R13859 Vbias.n310 Vbias.n199 52.5417
R13860 Vbias.n206 Vbias.n199 52.5417
R13861 Vbias.n290 Vbias.n213 52.5417
R13862 Vbias.n229 Vbias.n213 52.5417
R13863 Vbias.n230 Vbias.n229 52.5417
R13864 Vbias.n275 Vbias.n230 52.5417
R13865 Vbias.n271 Vbias.n232 52.5417
R13866 Vbias.n246 Vbias.n232 52.5417
R13867 Vbias.n248 Vbias.n246 52.5417
R13868 Vbias.n258 Vbias.n248 52.5417
R13869 Vbias.n7958 Vbias.n7957 52.5417
R13870 Vbias.n7957 Vbias.n7956 52.5417
R13871 Vbias.n7956 Vbias.n148 52.5417
R13872 Vbias.n7948 Vbias.n148 52.5417
R13873 Vbias.n141 Vbias.n132 52.5417
R13874 Vbias.n7962 Vbias.n141 52.5417
R13875 Vbias.n121 Vbias.n111 52.5417
R13876 Vbias.n7977 Vbias.n121 52.5417
R13877 Vbias.n7977 Vbias.n7976 52.5417
R13878 Vbias.n7976 Vbias.n7975 52.5417
R13879 Vbias.n102 Vbias.n92 52.5417
R13880 Vbias.n7992 Vbias.n102 52.5417
R13881 Vbias.n7992 Vbias.n7991 52.5417
R13882 Vbias.n7991 Vbias.n7990 52.5417
R13883 Vbias.n5033 Vbias.n2437 52.5417
R13884 Vbias.n4643 Vbias.n2437 52.5417
R13885 Vbias.n4644 Vbias.n4643 52.5417
R13886 Vbias.n4645 Vbias.n4644 52.5417
R13887 Vbias.n4650 Vbias.n4649 52.5417
R13888 Vbias.n4651 Vbias.n4650 52.5417
R13889 Vbias.n4652 Vbias.n4651 52.5417
R13890 Vbias.n4653 Vbias.n4652 52.5417
R13891 Vbias.n4664 Vbias.n4577 52.5417
R13892 Vbias.n4667 Vbias.n4577 52.5417
R13893 Vbias.n4508 Vbias.n4507 52.5417
R13894 Vbias.n4507 Vbias.n4506 52.5417
R13895 Vbias.n4506 Vbias.n4465 52.5417
R13896 Vbias.n4498 Vbias.n4465 52.5417
R13897 Vbias.n4522 Vbias.n4521 52.5417
R13898 Vbias.n4521 Vbias.n4520 52.5417
R13899 Vbias.n4520 Vbias.n4443 52.5417
R13900 Vbias.n4512 Vbias.n4443 52.5417
R13901 Vbias.n4437 Vbias.n4428 52.5417
R13902 Vbias.n4526 Vbias.n4437 52.5417
R13903 Vbias.n4542 Vbias.n4419 52.5417
R13904 Vbias.n4542 Vbias.n4422 52.5417
R13905 Vbias.n5117 Vbias.n2375 52.5417
R13906 Vbias.n5113 Vbias.n2375 52.5417
R13907 Vbias.n5113 Vbias.n2377 52.5417
R13908 Vbias.n5102 Vbias.n2377 52.5417
R13909 Vbias.n5097 Vbias.n2391 52.5417
R13910 Vbias.n5093 Vbias.n2391 52.5417
R13911 Vbias.n5093 Vbias.n2393 52.5417
R13912 Vbias.n5082 Vbias.n2393 52.5417
R13913 Vbias.n5071 Vbias.n2408 52.5417
R13914 Vbias.n2415 Vbias.n2408 52.5417
R13915 Vbias.n5490 Vbias.n5489 52.5417
R13916 Vbias.n5491 Vbias.n5490 52.5417
R13917 Vbias.n5491 Vbias.n2268 52.5417
R13918 Vbias.n5494 Vbias.n2268 52.5417
R13919 Vbias.n5501 Vbias.n2251 52.5417
R13920 Vbias.n5504 Vbias.n2251 52.5417
R13921 Vbias.n5505 Vbias.n5504 52.5417
R13922 Vbias.n5505 Vbias.n2249 52.5417
R13923 Vbias.n5172 Vbias.n5171 52.5417
R13924 Vbias.n5173 Vbias.n5172 52.5417
R13925 Vbias.n5178 Vbias.n5177 52.5417
R13926 Vbias.n5179 Vbias.n5178 52.5417
R13927 Vbias.n5180 Vbias.n5179 52.5417
R13928 Vbias.n5181 Vbias.n5180 52.5417
R13929 Vbias.n5914 Vbias.n1643 52.5417
R13930 Vbias.n5910 Vbias.n1643 52.5417
R13931 Vbias.n5910 Vbias.n1645 52.5417
R13932 Vbias.n5899 Vbias.n1645 52.5417
R13933 Vbias.n5894 Vbias.n1659 52.5417
R13934 Vbias.n5890 Vbias.n1659 52.5417
R13935 Vbias.n5890 Vbias.n1661 52.5417
R13936 Vbias.n5879 Vbias.n1661 52.5417
R13937 Vbias.n5466 Vbias.n5439 52.5417
R13938 Vbias.n5469 Vbias.n5439 52.5417
R13939 Vbias.n5477 Vbias.n5476 52.5417
R13940 Vbias.n5478 Vbias.n5477 52.5417
R13941 Vbias.n5478 Vbias.n2292 52.5417
R13942 Vbias.n5481 Vbias.n2292 52.5417
R13943 Vbias.n5945 Vbias.n5944 52.5417
R13944 Vbias.n5946 Vbias.n5945 52.5417
R13945 Vbias.n5951 Vbias.n5950 52.5417
R13946 Vbias.n5952 Vbias.n5951 52.5417
R13947 Vbias.n5953 Vbias.n5952 52.5417
R13948 Vbias.n5954 Vbias.n5953 52.5417
R13949 Vbias.n1884 Vbias.n1882 52.5417
R13950 Vbias.n1897 Vbias.n1882 52.5417
R13951 Vbias.n6121 Vbias.n1511 52.5417
R13952 Vbias.n6121 Vbias.n1512 52.5417
R13953 Vbias.n1511 Vbias.n1510 52.5417
R13954 Vbias.n6111 Vbias.n1512 52.5417
R13955 Vbias.n2000 Vbias.n1998 52.5417
R13956 Vbias.n1998 Vbias.n1985 52.5417
R13957 Vbias.n2001 Vbias.n2000 52.5417
R13958 Vbias.n2014 Vbias.n1985 52.5417
R13959 Vbias.n1981 Vbias.n1951 52.5417
R13960 Vbias.n1981 Vbias.n1952 52.5417
R13961 Vbias.n1951 Vbias.n1950 52.5417
R13962 Vbias.n1971 Vbias.n1952 52.5417
R13963 Vbias.n1947 Vbias.n1917 52.5417
R13964 Vbias.n1947 Vbias.n1918 52.5417
R13965 Vbias.n1917 Vbias.n1916 52.5417
R13966 Vbias.n1937 Vbias.n1918 52.5417
R13967 Vbias.n1800 Vbias.n1754 52.5417
R13968 Vbias.n1800 Vbias.n1753 52.5417
R13969 Vbias.n1755 Vbias.n1753 52.5417
R13970 Vbias.n1819 Vbias.n1755 52.5417
R13971 Vbias.n1849 Vbias.n1848 52.5417
R13972 Vbias.n1879 Vbias.n1849 52.5417
R13973 Vbias.n1879 Vbias.n1850 52.5417
R13974 Vbias.n1871 Vbias.n1850 52.5417
R13975 Vbias.n1745 Vbias.n1744 52.5417
R13976 Vbias.n1745 Vbias.n1731 52.5417
R13977 Vbias.n1744 Vbias.n1743 52.5417
R13978 Vbias.n2035 Vbias.n1731 52.5417
R13979 Vbias.n1913 Vbias.n1884 52.5417
R13980 Vbias.n1900 Vbias.n1897 52.5417
R13981 Vbias.n6082 Vbias.n6081 52.5417
R13982 Vbias.n6083 Vbias.n6082 52.5417
R13983 Vbias.n6084 Vbias.n6083 52.5417
R13984 Vbias.n6085 Vbias.n6084 52.5417
R13985 Vbias.n6090 Vbias.n6089 52.5417
R13986 Vbias.n6091 Vbias.n6090 52.5417
R13987 Vbias.n6092 Vbias.n6091 52.5417
R13988 Vbias.n6093 Vbias.n6092 52.5417
R13989 Vbias.n7011 Vbias.n1344 52.5417
R13990 Vbias.n6781 Vbias.n1344 52.5417
R13991 Vbias.n6782 Vbias.n6781 52.5417
R13992 Vbias.n6783 Vbias.n6782 52.5417
R13993 Vbias.n6788 Vbias.n6787 52.5417
R13994 Vbias.n6789 Vbias.n6788 52.5417
R13995 Vbias.n6790 Vbias.n6789 52.5417
R13996 Vbias.n6791 Vbias.n6790 52.5417
R13997 Vbias.n6803 Vbias.n6802 52.5417
R13998 Vbias.n6804 Vbias.n6803 52.5417
R13999 Vbias.n6809 Vbias.n6808 52.5417
R14000 Vbias.n6810 Vbias.n6809 52.5417
R14001 Vbias.n6811 Vbias.n6810 52.5417
R14002 Vbias.n6812 Vbias.n6811 52.5417
R14003 Vbias.n7093 Vbias.n1275 52.5417
R14004 Vbias.n1290 Vbias.n1275 52.5417
R14005 Vbias.n1291 Vbias.n1290 52.5417
R14006 Vbias.n7080 Vbias.n1291 52.5417
R14007 Vbias.n7076 Vbias.n1293 52.5417
R14008 Vbias.n1310 Vbias.n1293 52.5417
R14009 Vbias.n1311 Vbias.n1310 52.5417
R14010 Vbias.n7063 Vbias.n1311 52.5417
R14011 Vbias.n7050 Vbias.n1319 52.5417
R14012 Vbias.n7046 Vbias.n1319 52.5417
R14013 Vbias.n7033 Vbias.n1326 52.5417
R14014 Vbias.n7029 Vbias.n1326 52.5417
R14015 Vbias.n7029 Vbias.n1328 52.5417
R14016 Vbias.n7018 Vbias.n1328 52.5417
R14017 Vbias.n7199 Vbias.n1088 52.5417
R14018 Vbias.n1103 Vbias.n1088 52.5417
R14019 Vbias.n1104 Vbias.n1103 52.5417
R14020 Vbias.n7186 Vbias.n1104 52.5417
R14021 Vbias.n7182 Vbias.n1106 52.5417
R14022 Vbias.n1122 Vbias.n1106 52.5417
R14023 Vbias.n1123 Vbias.n1122 52.5417
R14024 Vbias.n7169 Vbias.n1123 52.5417
R14025 Vbias.n7156 Vbias.n1131 52.5417
R14026 Vbias.n7152 Vbias.n1131 52.5417
R14027 Vbias.n7139 Vbias.n1138 52.5417
R14028 Vbias.n7135 Vbias.n1138 52.5417
R14029 Vbias.n7135 Vbias.n1140 52.5417
R14030 Vbias.n7124 Vbias.n1140 52.5417
R14031 Vbias.n7208 Vbias.n1085 52.5417
R14032 Vbias.n7208 Vbias.n1079 52.5417
R14033 Vbias.n1216 Vbias.n1085 52.5417
R14034 Vbias.n1079 Vbias.n1077 52.5417
R14035 Vbias.n1240 Vbias.n1199 52.5417
R14036 Vbias.n1228 Vbias.n1199 52.5417
R14037 Vbias.n1241 Vbias.n1240 52.5417
R14038 Vbias.n1228 Vbias.n1213 52.5417
R14039 Vbias.n1187 Vbias.n1185 52.5417
R14040 Vbias.n1246 Vbias.n1187 52.5417
R14041 Vbias.n1271 Vbias.n1171 52.5417
R14042 Vbias.n1259 Vbias.n1171 52.5417
R14043 Vbias.n1272 Vbias.n1271 52.5417
R14044 Vbias.n1259 Vbias.n1182 52.5417
R14045 Vbias.n7104 Vbias.n1166 52.5417
R14046 Vbias.n7104 Vbias.n1160 52.5417
R14047 Vbias.n6949 Vbias.n1166 52.5417
R14048 Vbias.n1160 Vbias.n1158 52.5417
R14049 Vbias.n6973 Vbias.n6932 52.5417
R14050 Vbias.n6961 Vbias.n6932 52.5417
R14051 Vbias.n6974 Vbias.n6973 52.5417
R14052 Vbias.n6961 Vbias.n6946 52.5417
R14053 Vbias.n6920 Vbias.n6918 52.5417
R14054 Vbias.n6979 Vbias.n6920 52.5417
R14055 Vbias.n7004 Vbias.n6904 52.5417
R14056 Vbias.n6992 Vbias.n6904 52.5417
R14057 Vbias.n7005 Vbias.n7004 52.5417
R14058 Vbias.n6992 Vbias.n6915 52.5417
R14059 Vbias.n6883 Vbias.n1360 52.5417
R14060 Vbias.n6883 Vbias.n1354 52.5417
R14061 Vbias.n6878 Vbias.n1360 52.5417
R14062 Vbias.n1354 Vbias.n1352 52.5417
R14063 Vbias.n6860 Vbias.n1373 52.5417
R14064 Vbias.n6860 Vbias.n1367 52.5417
R14065 Vbias.n6855 Vbias.n1373 52.5417
R14066 Vbias.n1367 Vbias.n1365 52.5417
R14067 Vbias.n6837 Vbias.n1380 52.5417
R14068 Vbias.n1380 Vbias.n1378 52.5417
R14069 Vbias.n6821 Vbias.n6820 52.5417
R14070 Vbias.n6821 Vbias.n1388 52.5417
R14071 Vbias.n6820 Vbias.n6817 52.5417
R14072 Vbias.n6831 Vbias.n1388 52.5417
R14073 Vbias.n6028 Vbias.n1571 52.5417
R14074 Vbias.n6028 Vbias.n1565 52.5417
R14075 Vbias.n6020 Vbias.n1571 52.5417
R14076 Vbias.n1565 Vbias.n1563 52.5417
R14077 Vbias.n6002 Vbias.n1584 52.5417
R14078 Vbias.n6002 Vbias.n1578 52.5417
R14079 Vbias.n5997 Vbias.n1584 52.5417
R14080 Vbias.n1578 Vbias.n1576 52.5417
R14081 Vbias.n5979 Vbias.n1591 52.5417
R14082 Vbias.n1591 Vbias.n1589 52.5417
R14083 Vbias.n5963 Vbias.n5962 52.5417
R14084 Vbias.n5963 Vbias.n1599 52.5417
R14085 Vbias.n5962 Vbias.n5959 52.5417
R14086 Vbias.n5973 Vbias.n1599 52.5417
R14087 Vbias.n5357 Vbias.n5328 52.5417
R14088 Vbias.n5357 Vbias.n5331 52.5417
R14089 Vbias.n5328 Vbias.n5318 52.5417
R14090 Vbias.n5354 Vbias.n5331 52.5417
R14091 Vbias.n5381 Vbias.n5303 52.5417
R14092 Vbias.n5369 Vbias.n5303 52.5417
R14093 Vbias.n5382 Vbias.n5381 52.5417
R14094 Vbias.n5369 Vbias.n5315 52.5417
R14095 Vbias.n5291 Vbias.n5289 52.5417
R14096 Vbias.n5387 Vbias.n5291 52.5417
R14097 Vbias.n5412 Vbias.n5274 52.5417
R14098 Vbias.n5400 Vbias.n5274 52.5417
R14099 Vbias.n5413 Vbias.n5412 52.5417
R14100 Vbias.n5400 Vbias.n5286 52.5417
R14101 Vbias.n5252 Vbias.n2308 52.5417
R14102 Vbias.n5252 Vbias.n2302 52.5417
R14103 Vbias.n5247 Vbias.n2308 52.5417
R14104 Vbias.n2302 Vbias.n2300 52.5417
R14105 Vbias.n5229 Vbias.n2321 52.5417
R14106 Vbias.n5229 Vbias.n2315 52.5417
R14107 Vbias.n5224 Vbias.n2321 52.5417
R14108 Vbias.n2315 Vbias.n2313 52.5417
R14109 Vbias.n5206 Vbias.n2328 52.5417
R14110 Vbias.n2328 Vbias.n2326 52.5417
R14111 Vbias.n5190 Vbias.n5189 52.5417
R14112 Vbias.n5190 Vbias.n2336 52.5417
R14113 Vbias.n5189 Vbias.n5186 52.5417
R14114 Vbias.n5200 Vbias.n2336 52.5417
R14115 Vbias.n2525 Vbias.n2496 52.5417
R14116 Vbias.n2525 Vbias.n2499 52.5417
R14117 Vbias.n2496 Vbias.n2486 52.5417
R14118 Vbias.n2522 Vbias.n2499 52.5417
R14119 Vbias.n2549 Vbias.n2471 52.5417
R14120 Vbias.n2537 Vbias.n2471 52.5417
R14121 Vbias.n2550 Vbias.n2549 52.5417
R14122 Vbias.n2537 Vbias.n2483 52.5417
R14123 Vbias.n2459 Vbias.n2457 52.5417
R14124 Vbias.n2555 Vbias.n2459 52.5417
R14125 Vbias.n2580 Vbias.n2442 52.5417
R14126 Vbias.n2568 Vbias.n2442 52.5417
R14127 Vbias.n2581 Vbias.n2580 52.5417
R14128 Vbias.n2568 Vbias.n2454 52.5417
R14129 Vbias.n5054 Vbias.n2420 52.5417
R14130 Vbias.n5050 Vbias.n2420 52.5417
R14131 Vbias.n5050 Vbias.n2422 52.5417
R14132 Vbias.n5039 Vbias.n2422 52.5417
R14133 Vbias.n4419 Vbias.n4409 52.5417
R14134 Vbias.n4539 Vbias.n4422 52.5417
R14135 Vbias.n4186 Vbias.n4055 52.5417
R14136 Vbias.n4194 Vbias.n4055 52.5417
R14137 Vbias.n4194 Vbias.n4052 52.5417
R14138 Vbias.n4197 Vbias.n4052 52.5417
R14139 Vbias.n4210 Vbias.n4040 52.5417
R14140 Vbias.n4211 Vbias.n4210 52.5417
R14141 Vbias.n4220 Vbias.n4013 52.5417
R14142 Vbias.n4228 Vbias.n4013 52.5417
R14143 Vbias.n4228 Vbias.n4010 52.5417
R14144 Vbias.n4231 Vbias.n4010 52.5417
R14145 Vbias.n4240 Vbias.n4239 52.5417
R14146 Vbias.n4241 Vbias.n4240 52.5417
R14147 Vbias.n4241 Vbias.n3982 52.5417
R14148 Vbias.n4249 Vbias.n3982 52.5417
R14149 Vbias.n4178 Vbias.n4177 52.5417
R14150 Vbias.n4179 Vbias.n4178 52.5417
R14151 Vbias.n4179 Vbias.n4078 52.5417
R14152 Vbias.n4182 Vbias.n4078 52.5417
R14153 Vbias.n4148 Vbias.n4144 52.5417
R14154 Vbias.n4163 Vbias.n4144 52.5417
R14155 Vbias.n4128 Vbias.n4088 52.5417
R14156 Vbias.n4088 Vbias.n4087 52.5417
R14157 Vbias.n4087 Vbias.n4080 52.5417
R14158 Vbias.n4140 Vbias.n4080 52.5417
R14159 Vbias.n4115 Vbias.n4100 52.5417
R14160 Vbias.n4100 Vbias.n4099 52.5417
R14161 Vbias.n4099 Vbias.n4090 52.5417
R14162 Vbias.n4124 Vbias.n4090 52.5417
R14163 Vbias.n4975 Vbias.n4974 52.5417
R14164 Vbias.n4975 Vbias.n2605 52.5417
R14165 Vbias.n4974 Vbias.n4971 52.5417
R14166 Vbias.n4985 Vbias.n2605 52.5417
R14167 Vbias.n4957 Vbias.n2619 52.5417
R14168 Vbias.n4967 Vbias.n2619 52.5417
R14169 Vbias.n4946 Vbias.n2642 52.5417
R14170 Vbias.n4946 Vbias.n2636 52.5417
R14171 Vbias.n4941 Vbias.n2642 52.5417
R14172 Vbias.n2636 Vbias.n2634 52.5417
R14173 Vbias.n4923 Vbias.n2656 52.5417
R14174 Vbias.n4923 Vbias.n2650 52.5417
R14175 Vbias.n4919 Vbias.n2656 52.5417
R14176 Vbias.n2650 Vbias.n2648 52.5417
R14177 Vbias.n4675 Vbias.n4674 52.5417
R14178 Vbias.n4676 Vbias.n4675 52.5417
R14179 Vbias.n4676 Vbias.n4554 52.5417
R14180 Vbias.n4678 Vbias.n4554 52.5417
R14181 Vbias.n5653 Vbias.n5652 52.5417
R14182 Vbias.n5654 Vbias.n5653 52.5417
R14183 Vbias.n5654 Vbias.n2196 52.5417
R14184 Vbias.n5662 Vbias.n2196 52.5417
R14185 Vbias.n5640 Vbias.n2213 52.5417
R14186 Vbias.n5648 Vbias.n2213 52.5417
R14187 Vbias.n5624 Vbias.n5568 52.5417
R14188 Vbias.n5630 Vbias.n5568 52.5417
R14189 Vbias.n5630 Vbias.n5629 52.5417
R14190 Vbias.n5629 Vbias.n5556 52.5417
R14191 Vbias.n5606 Vbias.n5586 52.5417
R14192 Vbias.n5611 Vbias.n5586 52.5417
R14193 Vbias.n5611 Vbias.n5610 52.5417
R14194 Vbias.n5610 Vbias.n5574 52.5417
R14195 Vbias.n5727 Vbias.n5726 52.5417
R14196 Vbias.n5728 Vbias.n5727 52.5417
R14197 Vbias.n5728 Vbias.n2125 52.5417
R14198 Vbias.n5736 Vbias.n2125 52.5417
R14199 Vbias.n5714 Vbias.n2142 52.5417
R14200 Vbias.n5722 Vbias.n2142 52.5417
R14201 Vbias.n5698 Vbias.n2171 52.5417
R14202 Vbias.n5704 Vbias.n2171 52.5417
R14203 Vbias.n5704 Vbias.n5703 52.5417
R14204 Vbias.n5703 Vbias.n2159 52.5417
R14205 Vbias.n5680 Vbias.n2189 52.5417
R14206 Vbias.n5685 Vbias.n2189 52.5417
R14207 Vbias.n5685 Vbias.n5684 52.5417
R14208 Vbias.n5684 Vbias.n2177 52.5417
R14209 Vbias.n5816 Vbias.n5815 52.5417
R14210 Vbias.n5817 Vbias.n5816 52.5417
R14211 Vbias.n5817 Vbias.n2070 52.5417
R14212 Vbias.n5825 Vbias.n2070 52.5417
R14213 Vbias.n5803 Vbias.n5787 52.5417
R14214 Vbias.n5811 Vbias.n5787 52.5417
R14215 Vbias.n5773 Vbias.n5772 52.5417
R14216 Vbias.n5774 Vbias.n5773 52.5417
R14217 Vbias.n5774 Vbias.n2087 52.5417
R14218 Vbias.n5783 Vbias.n2087 52.5417
R14219 Vbias.n5759 Vbias.n5758 52.5417
R14220 Vbias.n5760 Vbias.n5759 52.5417
R14221 Vbias.n5760 Vbias.n2103 52.5417
R14222 Vbias.n5768 Vbias.n2103 52.5417
R14223 Vbias.n6663 Vbias.n6662 52.5417
R14224 Vbias.n6662 Vbias.n6661 52.5417
R14225 Vbias.n6661 Vbias.n1485 52.5417
R14226 Vbias.n6653 Vbias.n1485 52.5417
R14227 Vbias.n1479 Vbias.n1470 52.5417
R14228 Vbias.n6667 Vbias.n1479 52.5417
R14229 Vbias.n2051 Vbias.n1714 52.5417
R14230 Vbias.n2051 Vbias.n1715 52.5417
R14231 Vbias.n5844 Vbias.n1698 52.5417
R14232 Vbias.n5856 Vbias.n1698 52.5417
R14233 Vbias.n5856 Vbias.n5855 52.5417
R14234 Vbias.n5855 Vbias.n5854 52.5417
R14235 Vbias.n6357 Vbias.n6241 52.5417
R14236 Vbias.n6581 Vbias.n6241 52.5417
R14237 Vbias.n6581 Vbias.n6580 52.5417
R14238 Vbias.n6580 Vbias.n6229 52.5417
R14239 Vbias.n6344 Vbias.n6256 52.5417
R14240 Vbias.n6256 Vbias.n6247 52.5417
R14241 Vbias.n6330 Vbias.n6329 52.5417
R14242 Vbias.n6331 Vbias.n6330 52.5417
R14243 Vbias.n6331 Vbias.n6258 52.5417
R14244 Vbias.n6339 Vbias.n6258 52.5417
R14245 Vbias.n6316 Vbias.n6315 52.5417
R14246 Vbias.n6317 Vbias.n6316 52.5417
R14247 Vbias.n6317 Vbias.n6276 52.5417
R14248 Vbias.n6325 Vbias.n6276 52.5417
R14249 Vbias.n7602 Vbias.n7601 52.5417
R14250 Vbias.n7601 Vbias.n7600 52.5417
R14251 Vbias.n7600 Vbias.n840 52.5417
R14252 Vbias.n7592 Vbias.n840 52.5417
R14253 Vbias.n833 Vbias.n824 52.5417
R14254 Vbias.n7606 Vbias.n833 52.5417
R14255 Vbias.n812 Vbias.n802 52.5417
R14256 Vbias.n7621 Vbias.n812 52.5417
R14257 Vbias.n7621 Vbias.n7620 52.5417
R14258 Vbias.n7620 Vbias.n7619 52.5417
R14259 Vbias.n793 Vbias.n783 52.5417
R14260 Vbias.n7636 Vbias.n793 52.5417
R14261 Vbias.n7636 Vbias.n7635 52.5417
R14262 Vbias.n7635 Vbias.n7634 52.5417
R14263 Vbias.n7480 Vbias.n7479 52.5417
R14264 Vbias.n7479 Vbias.n7478 52.5417
R14265 Vbias.n7478 Vbias.n995 52.5417
R14266 Vbias.n7470 Vbias.n995 52.5417
R14267 Vbias.n988 Vbias.n979 52.5417
R14268 Vbias.n7484 Vbias.n988 52.5417
R14269 Vbias.n967 Vbias.n957 52.5417
R14270 Vbias.n7500 Vbias.n967 52.5417
R14271 Vbias.n7500 Vbias.n7499 52.5417
R14272 Vbias.n7499 Vbias.n7498 52.5417
R14273 Vbias.n944 Vbias.n934 52.5417
R14274 Vbias.n7515 Vbias.n944 52.5417
R14275 Vbias.n7515 Vbias.n7514 52.5417
R14276 Vbias.n7514 Vbias.n7513 52.5417
R14277 Vbias.n6603 Vbias.n6602 52.5417
R14278 Vbias.n6604 Vbias.n6603 52.5417
R14279 Vbias.n6604 Vbias.n6205 52.5417
R14280 Vbias.n6607 Vbias.n6205 52.5417
R14281 Vbias.n6614 Vbias.n6191 52.5417
R14282 Vbias.n6617 Vbias.n6191 52.5417
R14283 Vbias.n6629 Vbias.n6628 52.5417
R14284 Vbias.n6630 Vbias.n6629 52.5417
R14285 Vbias.n6631 Vbias.n6630 52.5417
R14286 Vbias.n6632 Vbias.n6631 52.5417
R14287 Vbias.n6536 Vbias.n6535 52.5417
R14288 Vbias.n6537 Vbias.n6536 52.5417
R14289 Vbias.n6537 Vbias.n6442 52.5417
R14290 Vbias.n6540 Vbias.n6442 52.5417
R14291 Vbias.n6547 Vbias.n6428 52.5417
R14292 Vbias.n6550 Vbias.n6428 52.5417
R14293 Vbias.n6562 Vbias.n6561 52.5417
R14294 Vbias.n6563 Vbias.n6562 52.5417
R14295 Vbias.n6564 Vbias.n6563 52.5417
R14296 Vbias.n6565 Vbias.n6564 52.5417
R14297 Vbias.n6570 Vbias.n6569 52.5417
R14298 Vbias.n6571 Vbias.n6570 52.5417
R14299 Vbias.n6572 Vbias.n6571 52.5417
R14300 Vbias.n6573 Vbias.n6572 52.5417
R14301 Vbias.n7549 Vbias.n7548 52.5417
R14302 Vbias.n7550 Vbias.n7549 52.5417
R14303 Vbias.n7550 Vbias.n896 52.5417
R14304 Vbias.n7553 Vbias.n896 52.5417
R14305 Vbias.n7560 Vbias.n882 52.5417
R14306 Vbias.n7563 Vbias.n882 52.5417
R14307 Vbias.n7575 Vbias.n7574 52.5417
R14308 Vbias.n7576 Vbias.n7575 52.5417
R14309 Vbias.n7577 Vbias.n7576 52.5417
R14310 Vbias.n7578 Vbias.n7577 52.5417
R14311 Vbias.n7583 Vbias.n7582 52.5417
R14312 Vbias.n7584 Vbias.n7583 52.5417
R14313 Vbias.n7585 Vbias.n7584 52.5417
R14314 Vbias.n7586 Vbias.n7585 52.5417
R14315 Vbias.n7400 Vbias.n7386 52.5417
R14316 Vbias.n7409 Vbias.n7386 52.5417
R14317 Vbias.n7409 Vbias.n7383 52.5417
R14318 Vbias.n7412 Vbias.n7383 52.5417
R14319 Vbias.n7425 Vbias.n7370 52.5417
R14320 Vbias.n7426 Vbias.n7425 52.5417
R14321 Vbias.n7435 Vbias.n7348 52.5417
R14322 Vbias.n7443 Vbias.n7348 52.5417
R14323 Vbias.n7443 Vbias.n7345 52.5417
R14324 Vbias.n7446 Vbias.n7345 52.5417
R14325 Vbias.n7455 Vbias.n7454 52.5417
R14326 Vbias.n7456 Vbias.n7455 52.5417
R14327 Vbias.n7456 Vbias.n7326 52.5417
R14328 Vbias.n7464 Vbias.n7326 52.5417
R14329 Vbias.n6636 Vbias.n6153 52.5417
R14330 Vbias.n6153 Vbias.n6137 52.5417
R14331 Vbias.n6646 Vbias.n6137 52.5417
R14332 Vbias.n6647 Vbias.n6646 52.5417
R14333 Vbias.n7274 Vbias.n7273 52.5417
R14334 Vbias.n7273 Vbias.n7272 52.5417
R14335 Vbias.n7272 Vbias.n7245 52.5417
R14336 Vbias.n7263 Vbias.n7245 52.5417
R14337 Vbias.n7238 Vbias.n7229 52.5417
R14338 Vbias.n7278 Vbias.n7238 52.5417
R14339 Vbias.n1062 Vbias.n1052 52.5417
R14340 Vbias.n7293 Vbias.n1062 52.5417
R14341 Vbias.n7293 Vbias.n7292 52.5417
R14342 Vbias.n7292 Vbias.n7291 52.5417
R14343 Vbias.n1041 Vbias.n1031 52.5417
R14344 Vbias.n7308 Vbias.n1041 52.5417
R14345 Vbias.n7308 Vbias.n7307 52.5417
R14346 Vbias.n7307 Vbias.n7306 52.5417
R14347 Vbias.n7722 Vbias.n685 52.5417
R14348 Vbias.n7730 Vbias.n685 52.5417
R14349 Vbias.n7731 Vbias.n7730 52.5417
R14350 Vbias.n7732 Vbias.n7731 52.5417
R14351 Vbias.n1714 Vbias.n1706 52.5417
R14352 Vbias.n2048 Vbias.n1715 52.5417
R14353 Vbias.n6690 Vbias.n1450 52.5417
R14354 Vbias.n1456 Vbias.n1450 52.5417
R14355 Vbias.n5868 Vbias.n1683 52.5417
R14356 Vbias.n5869 Vbias.n5868 52.5417
R14357 Vbias.n5526 Vbias.n5512 52.5417
R14358 Vbias.n5529 Vbias.n5512 52.5417
R14359 Vbias.n5544 Vbias.n2236 52.5417
R14360 Vbias.n5545 Vbias.n5544 52.5417
R14361 Vbias.n5025 Vbias.n2588 52.5417
R14362 Vbias.n5026 Vbias.n5025 52.5417
R14363 Vbias.n8062 Vbias.n16 52.5417
R14364 Vbias.n8070 Vbias.n16 52.5417
R14365 Vbias.n8071 Vbias.n8070 52.5417
R14366 Vbias.n8072 Vbias.n8071 52.5417
R14367 Vbias.n4685 Vbias.n4684 52.3938
R14368 Vbias.n4870 Vbias.t468 51.5416
R14369 Vbias.n8078 Vbias.t468 51.5416
R14370 Vbias.n1915 Vbias 48.6472
R14371 Vbias.n7402 Vbias.n7401 46.247
R14372 Vbias.n6101 Vbias.n1524 45.6728
R14373 Vbias.n6676 Vbias.n1461 45.6728
R14374 Vbias.n6679 Vbias.t744 45.3202
R14375 Vbias.n6686 Vbias.t744 45.3202
R14376 Vbias.t723 Vbias.n6686 45.3202
R14377 Vbias.t723 Vbias.n1443 45.3202
R14378 Vbias.n6749 Vbias.t760 45.3202
R14379 Vbias.n6726 Vbias.t760 45.3202
R14380 Vbias.n6727 Vbias.t407 45.3202
R14381 Vbias.n6735 Vbias.t407 45.3202
R14382 Vbias.t737 Vbias.n6735 45.3202
R14383 Vbias.n6737 Vbias.t737 45.3202
R14384 Vbias.n6701 Vbias.t229 45.3202
R14385 Vbias.n6709 Vbias.t229 45.3202
R14386 Vbias.t677 Vbias.n6709 45.3202
R14387 Vbias.n6710 Vbias.t677 45.3202
R14388 Vbias.n4684 Vbias.t739 45.3202
R14389 Vbias.n4992 Vbias.t739 45.3202
R14390 Vbias.t410 Vbias.n4993 45.3202
R14391 Vbias.t410 Vbias.n4994 45.3202
R14392 Vbias.n4994 Vbias.t700 45.3202
R14393 Vbias.n5009 Vbias.t700 45.3202
R14394 Vbias.t787 Vbias.n5012 45.3202
R14395 Vbias.n5022 Vbias.t787 45.3202
R14396 Vbias.n5022 Vbias.t829 45.3202
R14397 Vbias.t829 Vbias.n5016 45.3202
R14398 Vbias.n5552 Vbias.t655 45.3202
R14399 Vbias.n2241 Vbias.t655 45.3202
R14400 Vbias.t862 Vbias.n2242 45.3202
R14401 Vbias.n5541 Vbias.t862 45.3202
R14402 Vbias.n5541 Vbias.t719 45.3202
R14403 Vbias.t719 Vbias.n5535 45.3202
R14404 Vbias.n5532 Vbias.t604 45.3202
R14405 Vbias.n5518 Vbias.t604 45.3202
R14406 Vbias.t135 Vbias.n5518 45.3202
R14407 Vbias.t135 Vbias.n1673 45.3202
R14408 Vbias.n5876 Vbias.t370 45.3202
R14409 Vbias.n1688 Vbias.t370 45.3202
R14410 Vbias.t409 Vbias.n1689 45.3202
R14411 Vbias.n5865 Vbias.t409 45.3202
R14412 Vbias.n5865 Vbias.t7 45.3202
R14413 Vbias.t7 Vbias.n5859 45.3202
R14414 Vbias.n6678 Vbias.n1458 44.1007
R14415 Vbias.n4685 Vbias.n2610 43.0923
R14416 Vbias.n6676 Vbias.n1466 42.2805
R14417 Vbias.t299 Vbias.n7402 35.4181
R14418 Vbias.n7945 Vbias.n167 33.6641
R14419 Vbias.n4894 Vbias.n4846 32.5005
R14420 Vbias.n4897 Vbias.n4893 32.5005
R14421 Vbias.n4893 Vbias.n4892 32.4429
R14422 Vbias.n4381 Vbias.n4376 29.7417
R14423 Vbias.n4376 Vbias.n2795 29.7417
R14424 Vbias.n4389 Vbias.n4387 29.7417
R14425 Vbias.n4390 Vbias.n4389 29.7417
R14426 Vbias.n4391 Vbias.n4387 29.7417
R14427 Vbias.n4391 Vbias.n4390 29.7417
R14428 Vbias.n4381 Vbias.n4380 29.7417
R14429 Vbias.n4380 Vbias.n2795 29.7417
R14430 Vbias.n4356 Vbias.n2813 29.7417
R14431 Vbias.n2813 Vbias.n2807 29.7417
R14432 Vbias.n4356 Vbias.n4355 29.7417
R14433 Vbias.n4355 Vbias.n2807 29.7417
R14434 Vbias.n2859 Vbias.n2855 29.7417
R14435 Vbias.n2855 Vbias.n2844 29.7417
R14436 Vbias.n4321 Vbias.n4319 29.7417
R14437 Vbias.n4319 Vbias.n2825 29.7417
R14438 Vbias.n4321 Vbias.n4320 29.7417
R14439 Vbias.n4320 Vbias.n2825 29.7417
R14440 Vbias.n2859 Vbias.n2858 29.7417
R14441 Vbias.n2858 Vbias.n2844 29.7417
R14442 Vbias.n2893 Vbias.n2889 29.7417
R14443 Vbias.n2889 Vbias.n2878 29.7417
R14444 Vbias.n4288 Vbias.n4286 29.7417
R14445 Vbias.n4286 Vbias.n2861 29.7417
R14446 Vbias.n4288 Vbias.n4287 29.7417
R14447 Vbias.n4287 Vbias.n2861 29.7417
R14448 Vbias.n2893 Vbias.n2892 29.7417
R14449 Vbias.n2892 Vbias.n2878 29.7417
R14450 Vbias.n3821 Vbias.n3796 29.7417
R14451 Vbias.n3821 Vbias.n3799 29.7417
R14452 Vbias.n3830 Vbias.n3801 29.7417
R14453 Vbias.n3830 Vbias.n3820 29.7417
R14454 Vbias.n3819 Vbias.n3801 29.7417
R14455 Vbias.n3820 Vbias.n3819 29.7417
R14456 Vbias.n3809 Vbias.n3796 29.7417
R14457 Vbias.n3809 Vbias.n3799 29.7417
R14458 Vbias.n3885 Vbias.n3781 29.7417
R14459 Vbias.n3782 Vbias.n3781 29.7417
R14460 Vbias.n3885 Vbias.n3884 29.7417
R14461 Vbias.n3884 Vbias.n3782 29.7417
R14462 Vbias.n3897 Vbias.n3749 29.7417
R14463 Vbias.n3897 Vbias.n3752 29.7417
R14464 Vbias.n3906 Vbias.n3754 29.7417
R14465 Vbias.n3906 Vbias.n3896 29.7417
R14466 Vbias.n3895 Vbias.n3754 29.7417
R14467 Vbias.n3896 Vbias.n3895 29.7417
R14468 Vbias.n3762 Vbias.n3749 29.7417
R14469 Vbias.n3762 Vbias.n3752 29.7417
R14470 Vbias.n3935 Vbias.n3720 29.7417
R14471 Vbias.n3935 Vbias.n3723 29.7417
R14472 Vbias.n3944 Vbias.n3725 29.7417
R14473 Vbias.n3944 Vbias.n3934 29.7417
R14474 Vbias.n3933 Vbias.n3725 29.7417
R14475 Vbias.n3934 Vbias.n3933 29.7417
R14476 Vbias.n3733 Vbias.n3720 29.7417
R14477 Vbias.n3733 Vbias.n3723 29.7417
R14478 Vbias.n3283 Vbias.n3258 29.7417
R14479 Vbias.n3283 Vbias.n3261 29.7417
R14480 Vbias.n3292 Vbias.n3263 29.7417
R14481 Vbias.n3292 Vbias.n3282 29.7417
R14482 Vbias.n3281 Vbias.n3263 29.7417
R14483 Vbias.n3282 Vbias.n3281 29.7417
R14484 Vbias.n3271 Vbias.n3258 29.7417
R14485 Vbias.n3271 Vbias.n3261 29.7417
R14486 Vbias.n3347 Vbias.n3243 29.7417
R14487 Vbias.n3244 Vbias.n3243 29.7417
R14488 Vbias.n3347 Vbias.n3346 29.7417
R14489 Vbias.n3346 Vbias.n3244 29.7417
R14490 Vbias.n3359 Vbias.n3211 29.7417
R14491 Vbias.n3359 Vbias.n3214 29.7417
R14492 Vbias.n3368 Vbias.n3216 29.7417
R14493 Vbias.n3368 Vbias.n3358 29.7417
R14494 Vbias.n3357 Vbias.n3216 29.7417
R14495 Vbias.n3358 Vbias.n3357 29.7417
R14496 Vbias.n3224 Vbias.n3211 29.7417
R14497 Vbias.n3224 Vbias.n3214 29.7417
R14498 Vbias.n3397 Vbias.n3182 29.7417
R14499 Vbias.n3397 Vbias.n3185 29.7417
R14500 Vbias.n3406 Vbias.n3187 29.7417
R14501 Vbias.n3406 Vbias.n3396 29.7417
R14502 Vbias.n3395 Vbias.n3187 29.7417
R14503 Vbias.n3396 Vbias.n3395 29.7417
R14504 Vbias.n3195 Vbias.n3182 29.7417
R14505 Vbias.n3195 Vbias.n3185 29.7417
R14506 Vbias.n3552 Vbias.n3527 29.7417
R14507 Vbias.n3552 Vbias.n3530 29.7417
R14508 Vbias.n3561 Vbias.n3532 29.7417
R14509 Vbias.n3561 Vbias.n3551 29.7417
R14510 Vbias.n3550 Vbias.n3532 29.7417
R14511 Vbias.n3551 Vbias.n3550 29.7417
R14512 Vbias.n3540 Vbias.n3527 29.7417
R14513 Vbias.n3540 Vbias.n3530 29.7417
R14514 Vbias.n3616 Vbias.n3512 29.7417
R14515 Vbias.n3513 Vbias.n3512 29.7417
R14516 Vbias.n3616 Vbias.n3615 29.7417
R14517 Vbias.n3615 Vbias.n3513 29.7417
R14518 Vbias.n3628 Vbias.n3480 29.7417
R14519 Vbias.n3628 Vbias.n3483 29.7417
R14520 Vbias.n3637 Vbias.n3485 29.7417
R14521 Vbias.n3637 Vbias.n3627 29.7417
R14522 Vbias.n3626 Vbias.n3485 29.7417
R14523 Vbias.n3627 Vbias.n3626 29.7417
R14524 Vbias.n3493 Vbias.n3480 29.7417
R14525 Vbias.n3493 Vbias.n3483 29.7417
R14526 Vbias.n3666 Vbias.n3451 29.7417
R14527 Vbias.n3666 Vbias.n3454 29.7417
R14528 Vbias.n3675 Vbias.n3456 29.7417
R14529 Vbias.n3675 Vbias.n3665 29.7417
R14530 Vbias.n3664 Vbias.n3456 29.7417
R14531 Vbias.n3665 Vbias.n3664 29.7417
R14532 Vbias.n3464 Vbias.n3451 29.7417
R14533 Vbias.n3464 Vbias.n3454 29.7417
R14534 Vbias.n3013 Vbias.n2988 29.7417
R14535 Vbias.n3013 Vbias.n2991 29.7417
R14536 Vbias.n3022 Vbias.n2993 29.7417
R14537 Vbias.n3022 Vbias.n3012 29.7417
R14538 Vbias.n3011 Vbias.n2993 29.7417
R14539 Vbias.n3012 Vbias.n3011 29.7417
R14540 Vbias.n3001 Vbias.n2988 29.7417
R14541 Vbias.n3001 Vbias.n2991 29.7417
R14542 Vbias.n3077 Vbias.n2973 29.7417
R14543 Vbias.n2974 Vbias.n2973 29.7417
R14544 Vbias.n3077 Vbias.n3076 29.7417
R14545 Vbias.n3076 Vbias.n2974 29.7417
R14546 Vbias.n3089 Vbias.n2941 29.7417
R14547 Vbias.n3089 Vbias.n2944 29.7417
R14548 Vbias.n3098 Vbias.n2946 29.7417
R14549 Vbias.n3098 Vbias.n3088 29.7417
R14550 Vbias.n3087 Vbias.n2946 29.7417
R14551 Vbias.n3088 Vbias.n3087 29.7417
R14552 Vbias.n2954 Vbias.n2941 29.7417
R14553 Vbias.n2954 Vbias.n2944 29.7417
R14554 Vbias.n3127 Vbias.n2912 29.7417
R14555 Vbias.n3127 Vbias.n2915 29.7417
R14556 Vbias.n3136 Vbias.n2917 29.7417
R14557 Vbias.n3136 Vbias.n3126 29.7417
R14558 Vbias.n3125 Vbias.n2917 29.7417
R14559 Vbias.n3126 Vbias.n3125 29.7417
R14560 Vbias.n2925 Vbias.n2912 29.7417
R14561 Vbias.n2925 Vbias.n2915 29.7417
R14562 Vbias.n4689 Vbias.n2749 29.7417
R14563 Vbias.n4689 Vbias.n2752 29.7417
R14564 Vbias.n4698 Vbias.n2754 29.7417
R14565 Vbias.n4698 Vbias.n4688 29.7417
R14566 Vbias.n4687 Vbias.n2754 29.7417
R14567 Vbias.n4688 Vbias.n4687 29.7417
R14568 Vbias.n2762 Vbias.n2749 29.7417
R14569 Vbias.n2762 Vbias.n2752 29.7417
R14570 Vbias.n4753 Vbias.n2734 29.7417
R14571 Vbias.n2735 Vbias.n2734 29.7417
R14572 Vbias.n4753 Vbias.n4752 29.7417
R14573 Vbias.n4752 Vbias.n2735 29.7417
R14574 Vbias.n4765 Vbias.n2702 29.7417
R14575 Vbias.n4765 Vbias.n2705 29.7417
R14576 Vbias.n4774 Vbias.n2707 29.7417
R14577 Vbias.n4774 Vbias.n4764 29.7417
R14578 Vbias.n4763 Vbias.n2707 29.7417
R14579 Vbias.n4764 Vbias.n4763 29.7417
R14580 Vbias.n2715 Vbias.n2702 29.7417
R14581 Vbias.n2715 Vbias.n2705 29.7417
R14582 Vbias.n4803 Vbias.n2673 29.7417
R14583 Vbias.n4803 Vbias.n2676 29.7417
R14584 Vbias.n4812 Vbias.n2678 29.7417
R14585 Vbias.n4812 Vbias.n4802 29.7417
R14586 Vbias.n4801 Vbias.n2678 29.7417
R14587 Vbias.n4802 Vbias.n4801 29.7417
R14588 Vbias.n2686 Vbias.n2673 29.7417
R14589 Vbias.n2686 Vbias.n2676 29.7417
R14590 Vbias.n1949 Vbias 29.2342
R14591 Vbias.n6678 Vbias.n6677 27.4581
R14592 Vbias.n5858 Vbias.n1528 27.4581
R14593 Vbias Vbias.n7658 26.3103
R14594 Vbias.n6513 Vbias 26.3103
R14595 Vbias.n7537 Vbias 26.3103
R14596 Vbias.n7882 Vbias 26.3103
R14597 Vbias.n7816 Vbias 26.3103
R14598 Vbias.n7747 Vbias 26.3103
R14599 Vbias.n5548 Vbias 26.3103
R14600 Vbias.n5528 Vbias 26.3103
R14601 Vbias.n5872 Vbias 26.3103
R14602 Vbias Vbias.n1449 26.3103
R14603 Vbias.n6745 Vbias 26.3103
R14604 Vbias Vbias.n6716 26.3103
R14605 Vbias.n4887 Vbias.n4886 26.3005
R14606 Vbias.n4886 Vbias.n4885 26.3005
R14607 Vbias.n4890 Vbias.n4847 26.261
R14608 Vbias.t893 Vbias.t472 26.261
R14609 Vbias.n4878 Vbias.n4855 26.261
R14610 Vbias.t470 Vbias.t548 26.261
R14611 Vbias.n4871 Vbias.n4868 26.261
R14612 Vbias.t472 Vbias.n4847 25.2811
R14613 Vbias.n4878 Vbias.t893 25.2811
R14614 Vbias.t470 Vbias.n4855 25.2811
R14615 Vbias.n4868 Vbias.t548 25.2811
R14616 Vbias.n5028 Vbias 24.2016
R14617 Vbias.n7265 Vbias.t566 21.3141
R14618 Vbias.n1804 Vbias.n1765 20.1796
R14619 Vbias.t795 Vbias.t317 20.1796
R14620 Vbias.n1767 Vbias.n1759 20.1796
R14621 Vbias.t560 Vbias.t414 20.1796
R14622 Vbias.n1760 Vbias.n1466 20.1796
R14623 Vbias.n1983 Vbias 19.5277
R14624 Vbias.n1949 Vbias 19.2885
R14625 Vbias.n6727 Vbias.n6726 19.1913
R14626 Vbias.n4993 Vbias.n4992 19.1913
R14627 Vbias.n2242 Vbias.n2241 19.1913
R14628 Vbias.n1689 Vbias.n1688 19.1913
R14629 Vbias.n7097 Vbias.n7096 18.6076
R14630 Vbias.n7008 Vbias.n7007 18.6076
R14631 Vbias.n6815 Vbias.n6814 18.6076
R14632 Vbias.n5957 Vbias.n5956 18.6076
R14633 Vbias.n5416 Vbias.n5415 18.6076
R14634 Vbias.n5184 Vbias.n5183 18.6076
R14635 Vbias.n7468 Vbias.n7467 18.6076
R14636 Vbias.n7590 Vbias.n7589 18.6076
R14637 Vbias.n6577 Vbias.n6576 18.6076
R14638 Vbias.n6651 Vbias.n6650 18.6076
R14639 Vbias.n355 Vbias.n166 18.6076
R14640 Vbias.n5665 Vbias.n5664 18.6076
R14641 Vbias.n5739 Vbias.n5738 18.6076
R14642 Vbias.n5829 Vbias.n5828 18.6076
R14643 Vbias.n4869 Vbias.n1 17.7278
R14644 Vbias.n4870 Vbias.n4869 17.7278
R14645 Vbias.n8080 Vbias.n8079 17.7278
R14646 Vbias.n8079 Vbias.n8078 17.7278
R14647 Vbias.n6125 Vbias.n6124 17.3253
R14648 Vbias.n4254 Vbias 17.1782
R14649 Vbias.n3977 Vbias 17.1782
R14650 Vbias.n3439 Vbias 17.1782
R14651 Vbias.n3708 Vbias 17.1782
R14652 Vbias.n4101 Vbias 17.1782
R14653 Vbias.n3169 Vbias 17.1782
R14654 Vbias.n2899 Vbias 17.1782
R14655 Vbias.n7323 Vbias 17.1782
R14656 Vbias.n858 Vbias 17.1782
R14657 Vbias.n6363 Vbias 17.1782
R14658 Vbias.n6133 Vbias 17.1782
R14659 Vbias.n5830 Vbias 17.1782
R14660 Vbias.n5740 Vbias 17.1782
R14661 Vbias.n5666 Vbias 17.1782
R14662 Vbias.n5592 Vbias 17.1782
R14663 Vbias.n253 Vbias 17.1782
R14664 Vbias.n2896 Vbias 17.1782
R14665 Vbias.n8084 Vbias.t469 16.8637
R14666 Vbias.n6127 Vbias.n6125 15.8782
R14667 Vbias.n8085 Vbias.t471 14.02
R14668 Vbias.n8086 Vbias.t473 14.02
R14669 Vbias.n4390 Vbias.n2781 13.8976
R14670 Vbias.n4403 Vbias.n2781 13.8976
R14671 Vbias.n4386 Vbias.n2795 13.8976
R14672 Vbias.n4387 Vbias.n4386 13.8976
R14673 Vbias.n4382 Vbias.n2797 13.8976
R14674 Vbias.n4382 Vbias.n4381 13.8976
R14675 Vbias.n4360 Vbias.n2807 13.8976
R14676 Vbias.n4361 Vbias.n4360 13.8976
R14677 Vbias.n4357 Vbias.n2810 13.8976
R14678 Vbias.n4357 Vbias.n4356 13.8976
R14679 Vbias.n4331 Vbias.n2825 13.8976
R14680 Vbias.n4331 Vbias.n2827 13.8976
R14681 Vbias.n4322 Vbias.n2844 13.8976
R14682 Vbias.n4322 Vbias.n4321 13.8976
R14683 Vbias.n4303 Vbias.n4302 13.8976
R14684 Vbias.n4302 Vbias.n2859 13.8976
R14685 Vbias.n4298 Vbias.n2861 13.8976
R14686 Vbias.n4298 Vbias.n2863 13.8976
R14687 Vbias.n4289 Vbias.n2878 13.8976
R14688 Vbias.n4289 Vbias.n4288 13.8976
R14689 Vbias.n4270 Vbias.n4269 13.8976
R14690 Vbias.n4269 Vbias.n2893 13.8976
R14691 Vbias.n3840 Vbias.n3820 13.8976
R14692 Vbias.n3840 Vbias.n3839 13.8976
R14693 Vbias.n3848 Vbias.n3799 13.8976
R14694 Vbias.n3848 Vbias.n3801 13.8976
R14695 Vbias.n3852 Vbias.n3851 13.8976
R14696 Vbias.n3851 Vbias.n3796 13.8976
R14697 Vbias.n3876 Vbias.n3782 13.8976
R14698 Vbias.n3877 Vbias.n3876 13.8976
R14699 Vbias.n3886 Vbias.n3778 13.8976
R14700 Vbias.n3886 Vbias.n3885 13.8976
R14701 Vbias.n3916 Vbias.n3896 13.8976
R14702 Vbias.n3916 Vbias.n3915 13.8976
R14703 Vbias.n3924 Vbias.n3752 13.8976
R14704 Vbias.n3924 Vbias.n3754 13.8976
R14705 Vbias.n3928 Vbias.n3927 13.8976
R14706 Vbias.n3927 Vbias.n3749 13.8976
R14707 Vbias.n3954 Vbias.n3934 13.8976
R14708 Vbias.n3954 Vbias.n3953 13.8976
R14709 Vbias.n3962 Vbias.n3723 13.8976
R14710 Vbias.n3962 Vbias.n3725 13.8976
R14711 Vbias.n3966 Vbias.n3965 13.8976
R14712 Vbias.n3965 Vbias.n3720 13.8976
R14713 Vbias.n3302 Vbias.n3282 13.8976
R14714 Vbias.n3302 Vbias.n3301 13.8976
R14715 Vbias.n3310 Vbias.n3261 13.8976
R14716 Vbias.n3310 Vbias.n3263 13.8976
R14717 Vbias.n3314 Vbias.n3313 13.8976
R14718 Vbias.n3313 Vbias.n3258 13.8976
R14719 Vbias.n3338 Vbias.n3244 13.8976
R14720 Vbias.n3339 Vbias.n3338 13.8976
R14721 Vbias.n3348 Vbias.n3240 13.8976
R14722 Vbias.n3348 Vbias.n3347 13.8976
R14723 Vbias.n3378 Vbias.n3358 13.8976
R14724 Vbias.n3378 Vbias.n3377 13.8976
R14725 Vbias.n3386 Vbias.n3214 13.8976
R14726 Vbias.n3386 Vbias.n3216 13.8976
R14727 Vbias.n3390 Vbias.n3389 13.8976
R14728 Vbias.n3389 Vbias.n3211 13.8976
R14729 Vbias.n3416 Vbias.n3396 13.8976
R14730 Vbias.n3416 Vbias.n3415 13.8976
R14731 Vbias.n3424 Vbias.n3185 13.8976
R14732 Vbias.n3424 Vbias.n3187 13.8976
R14733 Vbias.n3428 Vbias.n3427 13.8976
R14734 Vbias.n3427 Vbias.n3182 13.8976
R14735 Vbias.n3571 Vbias.n3551 13.8976
R14736 Vbias.n3571 Vbias.n3570 13.8976
R14737 Vbias.n3579 Vbias.n3530 13.8976
R14738 Vbias.n3579 Vbias.n3532 13.8976
R14739 Vbias.n3583 Vbias.n3582 13.8976
R14740 Vbias.n3582 Vbias.n3527 13.8976
R14741 Vbias.n3607 Vbias.n3513 13.8976
R14742 Vbias.n3608 Vbias.n3607 13.8976
R14743 Vbias.n3617 Vbias.n3509 13.8976
R14744 Vbias.n3617 Vbias.n3616 13.8976
R14745 Vbias.n3647 Vbias.n3627 13.8976
R14746 Vbias.n3647 Vbias.n3646 13.8976
R14747 Vbias.n3655 Vbias.n3483 13.8976
R14748 Vbias.n3655 Vbias.n3485 13.8976
R14749 Vbias.n3659 Vbias.n3658 13.8976
R14750 Vbias.n3658 Vbias.n3480 13.8976
R14751 Vbias.n3685 Vbias.n3665 13.8976
R14752 Vbias.n3685 Vbias.n3684 13.8976
R14753 Vbias.n3693 Vbias.n3454 13.8976
R14754 Vbias.n3693 Vbias.n3456 13.8976
R14755 Vbias.n3697 Vbias.n3696 13.8976
R14756 Vbias.n3696 Vbias.n3451 13.8976
R14757 Vbias.n3032 Vbias.n3012 13.8976
R14758 Vbias.n3032 Vbias.n3031 13.8976
R14759 Vbias.n3040 Vbias.n2991 13.8976
R14760 Vbias.n3040 Vbias.n2993 13.8976
R14761 Vbias.n3044 Vbias.n3043 13.8976
R14762 Vbias.n3043 Vbias.n2988 13.8976
R14763 Vbias.n3068 Vbias.n2974 13.8976
R14764 Vbias.n3069 Vbias.n3068 13.8976
R14765 Vbias.n3078 Vbias.n2970 13.8976
R14766 Vbias.n3078 Vbias.n3077 13.8976
R14767 Vbias.n3108 Vbias.n3088 13.8976
R14768 Vbias.n3108 Vbias.n3107 13.8976
R14769 Vbias.n3116 Vbias.n2944 13.8976
R14770 Vbias.n3116 Vbias.n2946 13.8976
R14771 Vbias.n3120 Vbias.n3119 13.8976
R14772 Vbias.n3119 Vbias.n2941 13.8976
R14773 Vbias.n3146 Vbias.n3126 13.8976
R14774 Vbias.n3146 Vbias.n3145 13.8976
R14775 Vbias.n3154 Vbias.n2915 13.8976
R14776 Vbias.n3154 Vbias.n2917 13.8976
R14777 Vbias.n3158 Vbias.n3157 13.8976
R14778 Vbias.n3157 Vbias.n2912 13.8976
R14779 Vbias.n4708 Vbias.n4688 13.8976
R14780 Vbias.n4708 Vbias.n4707 13.8976
R14781 Vbias.n4716 Vbias.n2752 13.8976
R14782 Vbias.n4716 Vbias.n2754 13.8976
R14783 Vbias.n4720 Vbias.n4719 13.8976
R14784 Vbias.n4719 Vbias.n2749 13.8976
R14785 Vbias.n4744 Vbias.n2735 13.8976
R14786 Vbias.n4745 Vbias.n4744 13.8976
R14787 Vbias.n4754 Vbias.n2731 13.8976
R14788 Vbias.n4754 Vbias.n4753 13.8976
R14789 Vbias.n4784 Vbias.n4764 13.8976
R14790 Vbias.n4784 Vbias.n4783 13.8976
R14791 Vbias.n4792 Vbias.n2705 13.8976
R14792 Vbias.n4792 Vbias.n2707 13.8976
R14793 Vbias.n4796 Vbias.n4795 13.8976
R14794 Vbias.n4795 Vbias.n2702 13.8976
R14795 Vbias.n4822 Vbias.n4802 13.8976
R14796 Vbias.n4822 Vbias.n4821 13.8976
R14797 Vbias.n4830 Vbias.n2676 13.8976
R14798 Vbias.n4830 Vbias.n2678 13.8976
R14799 Vbias.n4834 Vbias.n4833 13.8976
R14800 Vbias.n4833 Vbias.n2673 13.8976
R14801 Vbias.n3440 Vbias.n3171 13.2764
R14802 Vbias.n4859 Vbias.n4857 12.4473
R14803 Vbias.n4857 Vbias.n4847 12.4473
R14804 Vbias.n4862 Vbias.n4860 12.4473
R14805 Vbias.n4862 Vbias.n4855 12.4473
R14806 Vbias.n4872 Vbias.n4861 12.4473
R14807 Vbias.n4872 Vbias.n4871 12.4473
R14808 Vbias.n8087 Vbias.n8086 11.5578
R14809 Vbias.n2900 Vbias.n2896 10.7601
R14810 Vbias.n5029 Vbias.n2583 10.6976
R14811 Vbias.n256 GND 10.5092
R14812 Vbias.n4252 Vbias.n4251 10.4893
R14813 Vbias.n6125 Vbias 10.3837
R14814 Vbias.n1509 Vbias 9.81028
R14815 Vbias.n8083 Vbias.t567 9.78785
R14816 Vbias.n5029 Vbias.n5028 9.62522
R14817 Vbias Vbias.n1509 9.59289
R14818 Vbias.n1881 Vbias 9.58202
R14819 Vbias.n1983 Vbias 9.58202
R14820 Vbias.n1915 Vbias 9.58202
R14821 Vbias.n6123 Vbias 9.53583
R14822 Vbias.n4889 Vbias.n4888 9.43598
R14823 Vbias.n4890 Vbias.n4889 9.43598
R14824 Vbias.n4879 Vbias.n4851 9.43598
R14825 Vbias.n4879 Vbias.n4878 9.43598
R14826 Vbias.n4854 Vbias.n4852 9.43598
R14827 Vbias.n4868 Vbias.n4854 9.43598
R14828 Vbias.n1847 Vbias 8.38365
R14829 Vbias.n1845 Vbias.n1844 8.32958
R14830 Vbias.n2032 Vbias.n2031 8.32958
R14831 Vbias.n7946 Vbias.n7945 8.16273
R14832 Vbias.n8083 Vbias.n8082 8.14785
R14833 Vbias.n254 Vbias.n253 7.9965
R14834 Vbias.n4254 Vbias.n4253 7.973
R14835 Vbias.n3978 Vbias.n3977 7.973
R14836 Vbias.n3440 Vbias.n3439 7.973
R14837 Vbias.n3709 Vbias.n3708 7.973
R14838 Vbias.n4101 Vbias.n3979 7.973
R14839 Vbias.n3170 Vbias.n3169 7.973
R14840 Vbias.n2900 Vbias.n2899 7.973
R14841 Vbias.n2023 Vbias.n1508 7.9105
R14842 Vbias.n2018 Vbias.n2017 7.9105
R14843 Vbias.n1825 Vbias.n1749 7.9105
R14844 Vbias.n1830 Vbias.n1750 7.9105
R14845 Vbias.n1835 Vbias.n1751 7.9105
R14846 Vbias.n1840 Vbias.n1752 7.9105
R14847 Vbias.n5030 Vbias.n5029 7.9105
R14848 Vbias.n7945 Vbias.n7944 7.9105
R14849 Vbias.n5183 Vbias.n5182 7.0005
R14850 Vbias.n5480 Vbias.n5416 7.0005
R14851 Vbias.n5956 Vbias.n5955 7.0005
R14852 Vbias.n6814 Vbias.n6813 7.0005
R14853 Vbias.n7008 Vbias.n1327 7.0005
R14854 Vbias.n7096 Vbias.n1139 7.0005
R14855 Vbias.n7097 Vbias.n1273 7.0005
R14856 Vbias.n7007 Vbias.n7006 7.0005
R14857 Vbias.n6816 Vbias.n6815 7.0005
R14858 Vbias.n5958 Vbias.n5957 7.0005
R14859 Vbias.n5415 Vbias.n5414 7.0005
R14860 Vbias.n5185 Vbias.n5184 7.0005
R14861 Vbias.n2583 Vbias.n2582 7.0005
R14862 Vbias.n6650 Vbias 5.98963
R14863 Vbias.n6576 Vbias 5.98963
R14864 Vbias.n7589 Vbias 5.98963
R14865 Vbias.n7467 Vbias 5.98963
R14866 Vbias Vbias.n7468 5.98963
R14867 Vbias Vbias.n7590 5.98963
R14868 Vbias Vbias.n6577 5.98963
R14869 Vbias Vbias.n6651 5.98963
R14870 Vbias.n5829 Vbias 5.98963
R14871 Vbias.n5739 Vbias 5.98963
R14872 Vbias.n5665 Vbias 5.98963
R14873 Vbias.n355 Vbias 5.98963
R14874 Vbias.n5664 Vbias 5.98963
R14875 Vbias.n5738 Vbias 5.98963
R14876 Vbias.n5828 Vbias 5.98963
R14877 Vbias.n4897 Vbias 4.71008
R14878 Vbias.n1826 Vbias.n1825 4.47177
R14879 Vbias Vbias.n7946 4.35376
R14880 Vbias.n5030 Vbias.n167 4.15267
R14881 Vbias.n8084 Vbias.n8083 3.4105
R14882 Vbias.n4541 Vbias.n4409 3.21898
R14883 Vbias.n4678 Vbias.n4677 3.21898
R14884 Vbias Vbias.n1242 3.03311
R14885 Vbias Vbias.n6975 3.03311
R14886 Vbias.n6856 Vbias 3.03311
R14887 Vbias.n5998 Vbias 3.03311
R14888 Vbias Vbias.n5383 3.03311
R14889 Vbias.n5225 Vbias 3.03311
R14890 Vbias Vbias.n2551 3.03311
R14891 Vbias Vbias.n4523 3.03311
R14892 Vbias.n8082 Vbias.n8081 2.92115
R14893 Vbias.n2421 Vbias.n167 2.79941
R14894 Vbias.n3170 Vbias.n2900 2.7876
R14895 Vbias.n4253 Vbias.n3170 2.7876
R14896 Vbias.n4253 Vbias.n4252 2.7876
R14897 Vbias.n3979 Vbias.n3978 2.7876
R14898 Vbias.n3978 Vbias.n3709 2.7876
R14899 Vbias.n3709 Vbias.n3440 2.7876
R14900 Vbias.n255 Vbias.n254 2.7406
R14901 Vbias.n7467 Vbias.n7466 2.5793
R14902 Vbias.n6650 Vbias.n6649 2.5793
R14903 Vbias.n6576 Vbias.n6575 2.5793
R14904 Vbias.n7589 Vbias.n7588 2.5793
R14905 Vbias.n356 Vbias.n355 2.5793
R14906 Vbias.n5664 Vbias.n462 2.5793
R14907 Vbias.n5738 Vbias.n576 2.5793
R14908 Vbias.n5828 Vbias.n5827 2.5793
R14909 Vbias.n254 GND 2.49506
R14910 Vbias.n8082 Vbias.n0 2.47333
R14911 Vbias.n4142 Vbias 2.42713
R14912 Vbias.n7239 Vbias 2.42713
R14913 Vbias.n989 Vbias 2.42713
R14914 Vbias.n834 Vbias 2.42713
R14915 Vbias.n6341 Vbias 2.42713
R14916 Vbias Vbias.n1718 2.42713
R14917 Vbias.n5785 Vbias 2.42713
R14918 Vbias Vbias.n5700 2.42713
R14919 Vbias Vbias.n5626 2.42713
R14920 Vbias.n142 Vbias 2.42713
R14921 Vbias Vbias.n4943 2.42713
R14922 Vbias.n1747 Vbias 2.32659
R14923 Vbias.n5183 Vbias 2.17441
R14924 Vbias.n5416 Vbias 2.17441
R14925 Vbias.n5956 Vbias 2.17441
R14926 Vbias.n6814 Vbias 2.17441
R14927 Vbias Vbias.n7008 2.17441
R14928 Vbias.n7096 Vbias 2.17441
R14929 Vbias Vbias.n5030 2.17441
R14930 Vbias.n345 Vbias.n327 2.15648
R14931 Vbias.n5028 Vbias.n5027 2.06028
R14932 Vbias.n4988 Vbias 1.74454
R14933 Vbias.n2023 Vbias.n2022 1.67683
R14934 Vbias.n1831 Vbias.n1830 1.6737
R14935 Vbias.n2018 Vbias.n1748 1.6737
R14936 Vbias.n1836 Vbias.n1835 1.67363
R14937 Vbias.n4268 Vbias.n2860 1.66898
R14938 Vbias.n4299 Vbias.n2860 1.66898
R14939 Vbias.n4301 Vbias.n2824 1.66898
R14940 Vbias.n4332 Vbias.n2824 1.66898
R14941 Vbias.n4359 Vbias.n4358 1.66898
R14942 Vbias.n4385 Vbias.n4383 1.66898
R14943 Vbias.n4385 Vbias.n4384 1.66898
R14944 Vbias.n5051 Vbias.n2421 1.66898
R14945 Vbias.n5053 Vbias.n5051 1.66898
R14946 Vbias.n5072 Vbias.n2407 1.66898
R14947 Vbias.n5094 Vbias.n2392 1.66898
R14948 Vbias.n5096 Vbias.n5094 1.66898
R14949 Vbias.n5114 Vbias.n2376 1.66898
R14950 Vbias.n5116 Vbias.n5114 1.66898
R14951 Vbias.n5182 Vbias.n2349 1.66898
R14952 Vbias.n5176 Vbias.n2349 1.66898
R14953 Vbias.n5174 Vbias.n2357 1.66898
R14954 Vbias.n5503 Vbias.n2252 1.66898
R14955 Vbias.n5503 Vbias.n5502 1.66898
R14956 Vbias.n5493 Vbias.n5492 1.66898
R14957 Vbias.n5492 Vbias.n2269 1.66898
R14958 Vbias.n5480 Vbias.n5479 1.66898
R14959 Vbias.n5479 Vbias.n5417 1.66898
R14960 Vbias.n5468 Vbias.n5467 1.66898
R14961 Vbias.n5891 Vbias.n1660 1.66898
R14962 Vbias.n5893 Vbias.n5891 1.66898
R14963 Vbias.n5911 Vbias.n1644 1.66898
R14964 Vbias.n5913 Vbias.n5911 1.66898
R14965 Vbias.n5955 Vbias.n1612 1.66898
R14966 Vbias.n5949 Vbias.n1612 1.66898
R14967 Vbias.n5947 Vbias.n1621 1.66898
R14968 Vbias.n6094 Vbias.n1537 1.66898
R14969 Vbias.n6088 Vbias.n1537 1.66898
R14970 Vbias.n6086 Vbias.n1545 1.66898
R14971 Vbias.n6080 Vbias.n1545 1.66898
R14972 Vbias.n6813 Vbias.n1401 1.66898
R14973 Vbias.n6807 Vbias.n1401 1.66898
R14974 Vbias.n6805 Vbias.n1409 1.66898
R14975 Vbias.n6792 Vbias.n1421 1.66898
R14976 Vbias.n6786 Vbias.n1421 1.66898
R14977 Vbias.n6784 Vbias.n1345 1.66898
R14978 Vbias.n7010 Vbias.n1345 1.66898
R14979 Vbias.n7030 Vbias.n1327 1.66898
R14980 Vbias.n7032 Vbias.n7030 1.66898
R14981 Vbias.n7049 Vbias.n7047 1.66898
R14982 Vbias.n7062 Vbias.n1292 1.66898
R14983 Vbias.n7077 Vbias.n1292 1.66898
R14984 Vbias.n7079 Vbias.n1274 1.66898
R14985 Vbias.n7094 Vbias.n1274 1.66898
R14986 Vbias.n7136 Vbias.n1139 1.66898
R14987 Vbias.n7138 Vbias.n7136 1.66898
R14988 Vbias.n7155 Vbias.n7153 1.66898
R14989 Vbias.n7168 Vbias.n1105 1.66898
R14990 Vbias.n7183 Vbias.n1105 1.66898
R14991 Vbias.n7185 Vbias.n1087 1.66898
R14992 Vbias.n7200 Vbias.n1087 1.66898
R14993 Vbias.n1273 Vbias.n1168 1.66898
R14994 Vbias.n1193 Vbias.n1168 1.66898
R14995 Vbias.n1244 Vbias.n1195 1.66898
R14996 Vbias.n1242 Vbias.n1196 1.66898
R14997 Vbias.n1212 Vbias.n1196 1.66898
R14998 Vbias.n7207 Vbias.n1086 1.66898
R14999 Vbias.n7207 Vbias.n7206 1.66898
R15000 Vbias.n7006 Vbias.n6901 1.66898
R15001 Vbias.n6926 Vbias.n6901 1.66898
R15002 Vbias.n6977 Vbias.n6928 1.66898
R15003 Vbias.n6975 Vbias.n6929 1.66898
R15004 Vbias.n6945 Vbias.n6929 1.66898
R15005 Vbias.n7103 Vbias.n1167 1.66898
R15006 Vbias.n7103 Vbias.n7102 1.66898
R15007 Vbias.n6816 Vbias.n1387 1.66898
R15008 Vbias.n6832 Vbias.n1387 1.66898
R15009 Vbias.n6836 Vbias.n6835 1.66898
R15010 Vbias.n6859 Vbias.n6856 1.66898
R15011 Vbias.n6859 Vbias.n6858 1.66898
R15012 Vbias.n6882 Vbias.n6879 1.66898
R15013 Vbias.n6882 Vbias.n6881 1.66898
R15014 Vbias.n5958 Vbias.n1598 1.66898
R15015 Vbias.n5974 Vbias.n1598 1.66898
R15016 Vbias.n5978 Vbias.n5977 1.66898
R15017 Vbias.n6001 Vbias.n5998 1.66898
R15018 Vbias.n6001 Vbias.n6000 1.66898
R15019 Vbias.n6027 Vbias.n6021 1.66898
R15020 Vbias.n6027 Vbias.n6026 1.66898
R15021 Vbias.n5414 Vbias.n5271 1.66898
R15022 Vbias.n5297 Vbias.n5271 1.66898
R15023 Vbias.n5385 Vbias.n5299 1.66898
R15024 Vbias.n5383 Vbias.n5300 1.66898
R15025 Vbias.n5332 Vbias.n5300 1.66898
R15026 Vbias.n5356 Vbias.n5334 1.66898
R15027 Vbias.n5356 Vbias.n5355 1.66898
R15028 Vbias.n5185 Vbias.n2335 1.66898
R15029 Vbias.n5201 Vbias.n2335 1.66898
R15030 Vbias.n5205 Vbias.n5204 1.66898
R15031 Vbias.n5228 Vbias.n5225 1.66898
R15032 Vbias.n5228 Vbias.n5227 1.66898
R15033 Vbias.n5251 Vbias.n5248 1.66898
R15034 Vbias.n5251 Vbias.n5250 1.66898
R15035 Vbias.n2582 Vbias.n2439 1.66898
R15036 Vbias.n2465 Vbias.n2439 1.66898
R15037 Vbias.n2553 Vbias.n2467 1.66898
R15038 Vbias.n2551 Vbias.n2468 1.66898
R15039 Vbias.n2500 Vbias.n2468 1.66898
R15040 Vbias.n2524 Vbias.n2502 1.66898
R15041 Vbias.n2524 Vbias.n2523 1.66898
R15042 Vbias.n4541 Vbias.n4540 1.66898
R15043 Vbias.n4525 Vbias.n4438 1.66898
R15044 Vbias.n4523 Vbias.n4439 1.66898
R15045 Vbias.n4511 Vbias.n4439 1.66898
R15046 Vbias.n4509 Vbias.n4461 1.66898
R15047 Vbias.n4497 Vbias.n4461 1.66898
R15048 Vbias.n3964 Vbias.n3963 1.66898
R15049 Vbias.n3963 Vbias.n3722 1.66898
R15050 Vbias.n3926 Vbias.n3925 1.66898
R15051 Vbias.n3925 Vbias.n3751 1.66898
R15052 Vbias.n3887 Vbias.n3777 1.66898
R15053 Vbias.n3850 Vbias.n3849 1.66898
R15054 Vbias.n3849 Vbias.n3798 1.66898
R15055 Vbias.n3426 Vbias.n3425 1.66898
R15056 Vbias.n3425 Vbias.n3184 1.66898
R15057 Vbias.n3388 Vbias.n3387 1.66898
R15058 Vbias.n3387 Vbias.n3213 1.66898
R15059 Vbias.n3349 Vbias.n3239 1.66898
R15060 Vbias.n3312 Vbias.n3311 1.66898
R15061 Vbias.n3311 Vbias.n3260 1.66898
R15062 Vbias.n3695 Vbias.n3694 1.66898
R15063 Vbias.n3694 Vbias.n3453 1.66898
R15064 Vbias.n3657 Vbias.n3656 1.66898
R15065 Vbias.n3656 Vbias.n3482 1.66898
R15066 Vbias.n3618 Vbias.n3508 1.66898
R15067 Vbias.n3581 Vbias.n3580 1.66898
R15068 Vbias.n3580 Vbias.n3529 1.66898
R15069 Vbias.n4250 Vbias.n3980 1.66898
R15070 Vbias.n4000 Vbias.n3980 1.66898
R15071 Vbias.n4230 Vbias.n4229 1.66898
R15072 Vbias.n4229 Vbias.n4012 1.66898
R15073 Vbias.n4212 Vbias.n4037 1.66898
R15074 Vbias.n4196 Vbias.n4195 1.66898
R15075 Vbias.n4195 Vbias.n4054 1.66898
R15076 Vbias.n4114 Vbias.n4089 1.66898
R15077 Vbias.n4125 Vbias.n4089 1.66898
R15078 Vbias.n4127 Vbias.n4079 1.66898
R15079 Vbias.n4141 Vbias.n4079 1.66898
R15080 Vbias.n4164 Vbias.n4143 1.66898
R15081 Vbias.n4180 Vbias.n4166 1.66898
R15082 Vbias.n4181 Vbias.n4180 1.66898
R15083 Vbias.n3156 Vbias.n3155 1.66898
R15084 Vbias.n3155 Vbias.n2914 1.66898
R15085 Vbias.n3118 Vbias.n3117 1.66898
R15086 Vbias.n3117 Vbias.n2943 1.66898
R15087 Vbias.n3079 Vbias.n2969 1.66898
R15088 Vbias.n3042 Vbias.n3041 1.66898
R15089 Vbias.n3041 Vbias.n2990 1.66898
R15090 Vbias.n4832 Vbias.n4831 1.66898
R15091 Vbias.n4831 Vbias.n2675 1.66898
R15092 Vbias.n4794 Vbias.n4793 1.66898
R15093 Vbias.n4793 Vbias.n2704 1.66898
R15094 Vbias.n4755 Vbias.n2730 1.66898
R15095 Vbias.n4718 Vbias.n4717 1.66898
R15096 Vbias.n4717 Vbias.n2751 1.66898
R15097 Vbias.n4677 Vbias.n4555 1.66898
R15098 Vbias.n4666 Vbias.n4665 1.66898
R15099 Vbias.n4654 Vbias.n4593 1.66898
R15100 Vbias.n4648 Vbias.n4593 1.66898
R15101 Vbias.n4646 Vbias.n2438 1.66898
R15102 Vbias.n5032 Vbias.n2438 1.66898
R15103 Vbias.n7465 Vbias.n7324 1.66898
R15104 Vbias.n7339 Vbias.n7324 1.66898
R15105 Vbias.n7445 Vbias.n7444 1.66898
R15106 Vbias.n7444 Vbias.n7347 1.66898
R15107 Vbias.n7427 Vbias.n7367 1.66898
R15108 Vbias.n7411 Vbias.n7410 1.66898
R15109 Vbias.n7410 Vbias.n7385 1.66898
R15110 Vbias.n6648 Vbias.n6134 1.66898
R15111 Vbias.n6635 Vbias.n6134 1.66898
R15112 Vbias.n6633 Vbias.n6154 1.66898
R15113 Vbias.n6627 Vbias.n6154 1.66898
R15114 Vbias.n6616 Vbias.n6615 1.66898
R15115 Vbias.n6606 Vbias.n6605 1.66898
R15116 Vbias.n6605 Vbias.n6207 1.66898
R15117 Vbias.n6574 Vbias.n6364 1.66898
R15118 Vbias.n6568 Vbias.n6364 1.66898
R15119 Vbias.n6566 Vbias.n6372 1.66898
R15120 Vbias.n6560 Vbias.n6372 1.66898
R15121 Vbias.n6549 Vbias.n6548 1.66898
R15122 Vbias.n6539 Vbias.n6538 1.66898
R15123 Vbias.n6538 Vbias.n6444 1.66898
R15124 Vbias.n7587 Vbias.n859 1.66898
R15125 Vbias.n7581 Vbias.n859 1.66898
R15126 Vbias.n7579 Vbias.n867 1.66898
R15127 Vbias.n7573 Vbias.n867 1.66898
R15128 Vbias.n7562 Vbias.n7561 1.66898
R15129 Vbias.n7552 Vbias.n7551 1.66898
R15130 Vbias.n7551 Vbias.n898 1.66898
R15131 Vbias.n1044 Vbias.n1043 1.66898
R15132 Vbias.n1047 Vbias.n1044 1.66898
R15133 Vbias.n1065 Vbias.n1064 1.66898
R15134 Vbias.n1068 Vbias.n1065 1.66898
R15135 Vbias.n7277 Vbias.n7240 1.66898
R15136 Vbias.n7275 Vbias.n7241 1.66898
R15137 Vbias.n7262 Vbias.n7241 1.66898
R15138 Vbias.n949 Vbias.n948 1.66898
R15139 Vbias.n952 Vbias.n949 1.66898
R15140 Vbias.n970 Vbias.n969 1.66898
R15141 Vbias.n973 Vbias.n970 1.66898
R15142 Vbias.n7483 Vbias.n990 1.66898
R15143 Vbias.n7481 Vbias.n991 1.66898
R15144 Vbias.n7469 Vbias.n991 1.66898
R15145 Vbias.n6359 Vbias.n794 1.66898
R15146 Vbias.n797 Vbias.n794 1.66898
R15147 Vbias.n815 Vbias.n814 1.66898
R15148 Vbias.n818 Vbias.n815 1.66898
R15149 Vbias.n7605 Vbias.n835 1.66898
R15150 Vbias.n7603 Vbias.n836 1.66898
R15151 Vbias.n7591 Vbias.n836 1.66898
R15152 Vbias.n6314 Vbias.n6275 1.66898
R15153 Vbias.n6326 Vbias.n6275 1.66898
R15154 Vbias.n6328 Vbias.n6257 1.66898
R15155 Vbias.n6340 Vbias.n6257 1.66898
R15156 Vbias.n6343 Vbias.n6342 1.66898
R15157 Vbias.n6579 Vbias.n6358 1.66898
R15158 Vbias.n6579 Vbias.n6578 1.66898
R15159 Vbias.n5843 Vbias.n1699 1.66898
R15160 Vbias.n1701 Vbias.n1699 1.66898
R15161 Vbias.n2050 Vbias.n1717 1.66898
R15162 Vbias.n2050 Vbias.n2049 1.66898
R15163 Vbias.n6666 Vbias.n1480 1.66898
R15164 Vbias.n6664 Vbias.n1481 1.66898
R15165 Vbias.n6652 Vbias.n1481 1.66898
R15166 Vbias.n5757 Vbias.n2102 1.66898
R15167 Vbias.n5769 Vbias.n2102 1.66898
R15168 Vbias.n5771 Vbias.n2086 1.66898
R15169 Vbias.n5784 Vbias.n2086 1.66898
R15170 Vbias.n5812 Vbias.n5786 1.66898
R15171 Vbias.n5814 Vbias.n2069 1.66898
R15172 Vbias.n5826 Vbias.n2069 1.66898
R15173 Vbias.n5683 Vbias.n5681 1.66898
R15174 Vbias.n5683 Vbias.n5682 1.66898
R15175 Vbias.n5702 Vbias.n5699 1.66898
R15176 Vbias.n5702 Vbias.n5701 1.66898
R15177 Vbias.n5723 Vbias.n2141 1.66898
R15178 Vbias.n5725 Vbias.n2124 1.66898
R15179 Vbias.n5737 Vbias.n2124 1.66898
R15180 Vbias.n5609 Vbias.n5607 1.66898
R15181 Vbias.n5609 Vbias.n5608 1.66898
R15182 Vbias.n5628 Vbias.n5625 1.66898
R15183 Vbias.n5628 Vbias.n5627 1.66898
R15184 Vbias.n5649 Vbias.n2212 1.66898
R15185 Vbias.n5651 Vbias.n2195 1.66898
R15186 Vbias.n5663 Vbias.n2195 1.66898
R15187 Vbias.n249 Vbias.n103 1.66898
R15188 Vbias.n106 Vbias.n103 1.66898
R15189 Vbias.n124 Vbias.n123 1.66898
R15190 Vbias.n127 Vbias.n124 1.66898
R15191 Vbias.n7961 Vbias.n143 1.66898
R15192 Vbias.n7959 Vbias.n144 1.66898
R15193 Vbias.n7947 Vbias.n144 1.66898
R15194 Vbias.n257 Vbias.n231 1.66898
R15195 Vbias.n272 Vbias.n231 1.66898
R15196 Vbias.n274 Vbias.n212 1.66898
R15197 Vbias.n291 Vbias.n212 1.66898
R15198 Vbias.n311 Vbias.n198 1.66898
R15199 Vbias.n313 Vbias.n179 1.66898
R15200 Vbias.n354 Vbias.n179 1.66898
R15201 Vbias.n7932 Vbias.n7931 1.66898
R15202 Vbias.n7931 Vbias.n357 1.66898
R15203 Vbias.n7920 Vbias.n7919 1.66898
R15204 Vbias.n7919 Vbias.n381 1.66898
R15205 Vbias.n7906 Vbias.n405 1.66898
R15206 Vbias.n7895 Vbias.n7894 1.66898
R15207 Vbias.n7894 Vbias.n428 1.66898
R15208 Vbias.n7866 Vbias.n7865 1.66898
R15209 Vbias.n7865 Vbias.n463 1.66898
R15210 Vbias.n7854 Vbias.n7853 1.66898
R15211 Vbias.n7853 Vbias.n487 1.66898
R15212 Vbias.n7840 Vbias.n511 1.66898
R15213 Vbias.n7829 Vbias.n7828 1.66898
R15214 Vbias.n7828 Vbias.n534 1.66898
R15215 Vbias.n7797 Vbias.n7796 1.66898
R15216 Vbias.n7796 Vbias.n577 1.66898
R15217 Vbias.n7785 Vbias.n7784 1.66898
R15218 Vbias.n7784 Vbias.n601 1.66898
R15219 Vbias.n7771 Vbias.n625 1.66898
R15220 Vbias.n7760 Vbias.n7759 1.66898
R15221 Vbias.n7759 Vbias.n648 1.66898
R15222 Vbias.n684 Vbias.n682 1.66898
R15223 Vbias.n7721 Vbias.n684 1.66898
R15224 Vbias.n7719 Vbias.n699 1.66898
R15225 Vbias.n7706 Vbias.n699 1.66898
R15226 Vbias.n7695 Vbias.n7694 1.66898
R15227 Vbias.n7680 Vbias.n7679 1.66898
R15228 Vbias.n7679 Vbias.n740 1.66898
R15229 Vbias.n7660 Vbias.n770 1.66898
R15230 Vbias.n7658 Vbias.n771 1.66898
R15231 Vbias.n7535 Vbias.n924 1.66898
R15232 Vbias.n7539 Vbias.n7537 1.66898
R15233 Vbias.n7882 Vbias.n7881 1.66898
R15234 Vbias.n7814 Vbias.n558 1.66898
R15235 Vbias.n7747 Vbias.n7746 1.66898
R15236 Vbias.n5027 Vbias.n2585 1.66898
R15237 Vbias.n5546 Vbias.n2233 1.66898
R15238 Vbias.n5528 Vbias.n5527 1.66898
R15239 Vbias.n5870 Vbias.n1680 1.66898
R15240 Vbias.n6691 Vbias.n1449 1.66898
R15241 Vbias.n6743 Vbias.n6718 1.66898
R15242 Vbias.n6716 Vbias.n6694 1.66898
R15243 Vbias.n5005 Vbias.n5003 1.66898
R15244 Vbias.n4922 Vbias.n4920 1.66898
R15245 Vbias.n4922 Vbias.n4921 1.66898
R15246 Vbias.n4945 Vbias.n4942 1.66898
R15247 Vbias.n4945 Vbias.n4944 1.66898
R15248 Vbias.n4968 Vbias.n2618 1.66898
R15249 Vbias.n4970 Vbias.n2604 1.66898
R15250 Vbias.n4986 Vbias.n2604 1.66898
R15251 Vbias.n15 Vbias.n13 1.66898
R15252 Vbias.n8061 Vbias.n15 1.66898
R15253 Vbias.n8059 Vbias.n30 1.66898
R15254 Vbias.n8046 Vbias.n30 1.66898
R15255 Vbias.n8035 Vbias.n8034 1.66898
R15256 Vbias.n8020 Vbias.n8019 1.66898
R15257 Vbias.n8019 Vbias.n71 1.66898
R15258 Vbias.n168 Vbias 1.66083
R15259 Vbias.n4252 Vbias.n3979 1.65255
R15260 Vbias.n7946 Vbias.n166 1.58746
R15261 Vbias.n4266 Vbias.n4265 1.5505
R15262 Vbias.n4269 Vbias.n4268 1.5505
R15263 Vbias.n4289 Vbias.n2860 1.5505
R15264 Vbias.n4299 Vbias.n4298 1.5505
R15265 Vbias.n4302 Vbias.n4301 1.5505
R15266 Vbias.n4322 Vbias.n2824 1.5505
R15267 Vbias.n4332 Vbias.n4331 1.5505
R15268 Vbias.n4335 Vbias.n4334 1.5505
R15269 Vbias.n4358 Vbias.n4357 1.5505
R15270 Vbias.n4360 Vbias.n4359 1.5505
R15271 Vbias.n4383 Vbias.n4382 1.5505
R15272 Vbias.n4386 Vbias.n4385 1.5505
R15273 Vbias.n4384 Vbias.n2781 1.5505
R15274 Vbias.n6111 Vbias.n6110 1.5505
R15275 Vbias.n2015 Vbias.n2014 1.5505
R15276 Vbias.n1971 Vbias.n1970 1.5505
R15277 Vbias.n1937 Vbias.n1936 1.5505
R15278 Vbias.n1820 Vbias.n1819 1.5505
R15279 Vbias.n1871 Vbias.n1870 1.5505
R15280 Vbias.n1880 Vbias.n1848 1.5505
R15281 Vbias.n1880 Vbias.n1879 1.5505
R15282 Vbias.n1846 Vbias.n1754 1.5505
R15283 Vbias.n1846 Vbias.n1753 1.5505
R15284 Vbias.n2035 Vbias.n2034 1.5505
R15285 Vbias.n1743 Vbias.n1507 1.5505
R15286 Vbias.n1746 Vbias.n1745 1.5505
R15287 Vbias.n6122 Vbias.n1510 1.5505
R15288 Vbias.n6122 Vbias.n6121 1.5505
R15289 Vbias.n2001 Vbias.n1984 1.5505
R15290 Vbias.n1998 Vbias.n1984 1.5505
R15291 Vbias.n1982 Vbias.n1950 1.5505
R15292 Vbias.n1982 Vbias.n1981 1.5505
R15293 Vbias.n1948 Vbias.n1916 1.5505
R15294 Vbias.n1948 Vbias.n1947 1.5505
R15295 Vbias.n1914 Vbias.n1882 1.5505
R15296 Vbias.n1914 Vbias.n1913 1.5505
R15297 Vbias.n1900 Vbias.n1899 1.5505
R15298 Vbias.n5039 Vbias.n2421 1.5505
R15299 Vbias.n5051 Vbias.n5050 1.5505
R15300 Vbias.n5054 Vbias.n5053 1.5505
R15301 Vbias.n2415 Vbias.n2407 1.5505
R15302 Vbias.n5072 Vbias.n5071 1.5505
R15303 Vbias.n5076 Vbias.n5075 1.5505
R15304 Vbias.n5082 Vbias.n2392 1.5505
R15305 Vbias.n5094 Vbias.n5093 1.5505
R15306 Vbias.n5097 Vbias.n5096 1.5505
R15307 Vbias.n5102 Vbias.n2376 1.5505
R15308 Vbias.n5114 Vbias.n5113 1.5505
R15309 Vbias.n5117 Vbias.n5116 1.5505
R15310 Vbias.n5182 Vbias.n5181 1.5505
R15311 Vbias.n5179 Vbias.n2349 1.5505
R15312 Vbias.n5177 Vbias.n5176 1.5505
R15313 Vbias.n5174 Vbias.n5173 1.5505
R15314 Vbias.n5171 Vbias.n2357 1.5505
R15315 Vbias.n5164 Vbias.n5163 1.5505
R15316 Vbias.n2252 Vbias.n2249 1.5505
R15317 Vbias.n5504 Vbias.n5503 1.5505
R15318 Vbias.n5502 Vbias.n5501 1.5505
R15319 Vbias.n5494 Vbias.n5493 1.5505
R15320 Vbias.n5492 Vbias.n5491 1.5505
R15321 Vbias.n5489 Vbias.n2269 1.5505
R15322 Vbias.n5481 Vbias.n5480 1.5505
R15323 Vbias.n5479 Vbias.n5478 1.5505
R15324 Vbias.n5476 Vbias.n5417 1.5505
R15325 Vbias.n5469 Vbias.n5468 1.5505
R15326 Vbias.n5467 Vbias.n5466 1.5505
R15327 Vbias.n5459 Vbias.n5458 1.5505
R15328 Vbias.n5879 Vbias.n1660 1.5505
R15329 Vbias.n5891 Vbias.n5890 1.5505
R15330 Vbias.n5894 Vbias.n5893 1.5505
R15331 Vbias.n5899 Vbias.n1644 1.5505
R15332 Vbias.n5911 Vbias.n5910 1.5505
R15333 Vbias.n5914 Vbias.n5913 1.5505
R15334 Vbias.n5955 Vbias.n5954 1.5505
R15335 Vbias.n5952 Vbias.n1612 1.5505
R15336 Vbias.n5950 Vbias.n5949 1.5505
R15337 Vbias.n5947 Vbias.n5946 1.5505
R15338 Vbias.n5944 Vbias.n1621 1.5505
R15339 Vbias.n6097 Vbias.n6096 1.5505
R15340 Vbias.n6094 Vbias.n6093 1.5505
R15341 Vbias.n6091 Vbias.n1537 1.5505
R15342 Vbias.n6089 Vbias.n6088 1.5505
R15343 Vbias.n6086 Vbias.n6085 1.5505
R15344 Vbias.n6083 Vbias.n1545 1.5505
R15345 Vbias.n6081 Vbias.n6080 1.5505
R15346 Vbias.n6813 Vbias.n6812 1.5505
R15347 Vbias.n6810 Vbias.n1401 1.5505
R15348 Vbias.n6808 Vbias.n6807 1.5505
R15349 Vbias.n6805 Vbias.n6804 1.5505
R15350 Vbias.n6802 Vbias.n1409 1.5505
R15351 Vbias.n6795 Vbias.n6794 1.5505
R15352 Vbias.n6792 Vbias.n6791 1.5505
R15353 Vbias.n6789 Vbias.n1421 1.5505
R15354 Vbias.n6787 Vbias.n6786 1.5505
R15355 Vbias.n6784 Vbias.n6783 1.5505
R15356 Vbias.n6781 Vbias.n1345 1.5505
R15357 Vbias.n7011 Vbias.n7010 1.5505
R15358 Vbias.n7018 Vbias.n1327 1.5505
R15359 Vbias.n7030 Vbias.n7029 1.5505
R15360 Vbias.n7033 Vbias.n7032 1.5505
R15361 Vbias.n7047 Vbias.n7046 1.5505
R15362 Vbias.n7050 Vbias.n7049 1.5505
R15363 Vbias.n7060 Vbias.n7059 1.5505
R15364 Vbias.n7063 Vbias.n7062 1.5505
R15365 Vbias.n1310 Vbias.n1292 1.5505
R15366 Vbias.n7077 Vbias.n7076 1.5505
R15367 Vbias.n7080 Vbias.n7079 1.5505
R15368 Vbias.n1290 Vbias.n1274 1.5505
R15369 Vbias.n7094 Vbias.n7093 1.5505
R15370 Vbias.n7124 Vbias.n1139 1.5505
R15371 Vbias.n7136 Vbias.n7135 1.5505
R15372 Vbias.n7139 Vbias.n7138 1.5505
R15373 Vbias.n7153 Vbias.n7152 1.5505
R15374 Vbias.n7156 Vbias.n7155 1.5505
R15375 Vbias.n7166 Vbias.n7165 1.5505
R15376 Vbias.n7169 Vbias.n7168 1.5505
R15377 Vbias.n1122 Vbias.n1105 1.5505
R15378 Vbias.n7183 Vbias.n7182 1.5505
R15379 Vbias.n7186 Vbias.n7185 1.5505
R15380 Vbias.n1103 Vbias.n1087 1.5505
R15381 Vbias.n7200 Vbias.n7199 1.5505
R15382 Vbias.n1273 Vbias.n1272 1.5505
R15383 Vbias.n1171 Vbias.n1168 1.5505
R15384 Vbias.n1193 Vbias.n1182 1.5505
R15385 Vbias.n1195 Vbias.n1185 1.5505
R15386 Vbias.n1246 Vbias.n1244 1.5505
R15387 Vbias.n1242 Vbias.n1241 1.5505
R15388 Vbias.n1199 Vbias.n1196 1.5505
R15389 Vbias.n1213 Vbias.n1212 1.5505
R15390 Vbias.n1216 Vbias.n1086 1.5505
R15391 Vbias.n7208 Vbias.n7207 1.5505
R15392 Vbias.n7206 Vbias.n1077 1.5505
R15393 Vbias.n7204 Vbias.n1074 1.5505
R15394 Vbias.n7006 Vbias.n7005 1.5505
R15395 Vbias.n6904 Vbias.n6901 1.5505
R15396 Vbias.n6926 Vbias.n6915 1.5505
R15397 Vbias.n6928 Vbias.n6918 1.5505
R15398 Vbias.n6979 Vbias.n6977 1.5505
R15399 Vbias.n6975 Vbias.n6974 1.5505
R15400 Vbias.n6932 Vbias.n6929 1.5505
R15401 Vbias.n6946 Vbias.n6945 1.5505
R15402 Vbias.n6949 Vbias.n1167 1.5505
R15403 Vbias.n7104 Vbias.n7103 1.5505
R15404 Vbias.n7102 Vbias.n1158 1.5505
R15405 Vbias.n7100 Vbias.n1155 1.5505
R15406 Vbias.n6817 Vbias.n6816 1.5505
R15407 Vbias.n6821 Vbias.n1387 1.5505
R15408 Vbias.n6832 Vbias.n6831 1.5505
R15409 Vbias.n6837 Vbias.n6836 1.5505
R15410 Vbias.n6835 Vbias.n1378 1.5505
R15411 Vbias.n6856 Vbias.n6855 1.5505
R15412 Vbias.n6860 Vbias.n6859 1.5505
R15413 Vbias.n6858 Vbias.n1365 1.5505
R15414 Vbias.n6879 Vbias.n6878 1.5505
R15415 Vbias.n6883 Vbias.n6882 1.5505
R15416 Vbias.n6881 Vbias.n1352 1.5505
R15417 Vbias.n6898 Vbias.n6897 1.5505
R15418 Vbias.n5959 Vbias.n5958 1.5505
R15419 Vbias.n5963 Vbias.n1598 1.5505
R15420 Vbias.n5974 Vbias.n5973 1.5505
R15421 Vbias.n5979 Vbias.n5978 1.5505
R15422 Vbias.n5977 Vbias.n1589 1.5505
R15423 Vbias.n5998 Vbias.n5997 1.5505
R15424 Vbias.n6002 Vbias.n6001 1.5505
R15425 Vbias.n6000 Vbias.n1576 1.5505
R15426 Vbias.n6021 Vbias.n6020 1.5505
R15427 Vbias.n6028 Vbias.n6027 1.5505
R15428 Vbias.n6026 Vbias.n1563 1.5505
R15429 Vbias.n6024 Vbias.n1560 1.5505
R15430 Vbias.n5414 Vbias.n5413 1.5505
R15431 Vbias.n5274 Vbias.n5271 1.5505
R15432 Vbias.n5297 Vbias.n5286 1.5505
R15433 Vbias.n5299 Vbias.n5289 1.5505
R15434 Vbias.n5387 Vbias.n5385 1.5505
R15435 Vbias.n5383 Vbias.n5382 1.5505
R15436 Vbias.n5303 Vbias.n5300 1.5505
R15437 Vbias.n5332 Vbias.n5315 1.5505
R15438 Vbias.n5334 Vbias.n5318 1.5505
R15439 Vbias.n5357 Vbias.n5356 1.5505
R15440 Vbias.n5355 Vbias.n5354 1.5505
R15441 Vbias.n5343 Vbias.n5342 1.5505
R15442 Vbias.n5186 Vbias.n5185 1.5505
R15443 Vbias.n5190 Vbias.n2335 1.5505
R15444 Vbias.n5201 Vbias.n5200 1.5505
R15445 Vbias.n5206 Vbias.n5205 1.5505
R15446 Vbias.n5204 Vbias.n2326 1.5505
R15447 Vbias.n5225 Vbias.n5224 1.5505
R15448 Vbias.n5229 Vbias.n5228 1.5505
R15449 Vbias.n5227 Vbias.n2313 1.5505
R15450 Vbias.n5248 Vbias.n5247 1.5505
R15451 Vbias.n5252 Vbias.n5251 1.5505
R15452 Vbias.n5250 Vbias.n2300 1.5505
R15453 Vbias.n5268 Vbias.n5267 1.5505
R15454 Vbias.n2582 Vbias.n2581 1.5505
R15455 Vbias.n2442 Vbias.n2439 1.5505
R15456 Vbias.n2465 Vbias.n2454 1.5505
R15457 Vbias.n2467 Vbias.n2457 1.5505
R15458 Vbias.n2555 Vbias.n2553 1.5505
R15459 Vbias.n2551 Vbias.n2550 1.5505
R15460 Vbias.n2471 Vbias.n2468 1.5505
R15461 Vbias.n2500 Vbias.n2483 1.5505
R15462 Vbias.n2502 Vbias.n2486 1.5505
R15463 Vbias.n2525 Vbias.n2524 1.5505
R15464 Vbias.n2523 Vbias.n2522 1.5505
R15465 Vbias.n2511 Vbias.n2510 1.5505
R15466 Vbias.n4542 Vbias.n4541 1.5505
R15467 Vbias.n4438 Vbias.n4428 1.5505
R15468 Vbias.n4526 Vbias.n4525 1.5505
R15469 Vbias.n4523 Vbias.n4522 1.5505
R15470 Vbias.n4520 Vbias.n4439 1.5505
R15471 Vbias.n4512 Vbias.n4511 1.5505
R15472 Vbias.n4509 Vbias.n4508 1.5505
R15473 Vbias.n4506 Vbias.n4461 1.5505
R15474 Vbias.n4498 Vbias.n4497 1.5505
R15475 Vbias.n4495 Vbias.n4494 1.5505
R15476 Vbias.n4540 Vbias.n4539 1.5505
R15477 Vbias.n3965 Vbias.n3964 1.5505
R15478 Vbias.n3963 Vbias.n3962 1.5505
R15479 Vbias.n3954 Vbias.n3722 1.5505
R15480 Vbias.n3927 Vbias.n3926 1.5505
R15481 Vbias.n3925 Vbias.n3924 1.5505
R15482 Vbias.n3916 Vbias.n3751 1.5505
R15483 Vbias.n3890 Vbias.n3889 1.5505
R15484 Vbias.n3887 Vbias.n3886 1.5505
R15485 Vbias.n3876 Vbias.n3777 1.5505
R15486 Vbias.n3851 Vbias.n3850 1.5505
R15487 Vbias.n3849 Vbias.n3848 1.5505
R15488 Vbias.n3840 Vbias.n3798 1.5505
R15489 Vbias.n3975 Vbias.n3974 1.5505
R15490 Vbias.n3427 Vbias.n3426 1.5505
R15491 Vbias.n3425 Vbias.n3424 1.5505
R15492 Vbias.n3416 Vbias.n3184 1.5505
R15493 Vbias.n3389 Vbias.n3388 1.5505
R15494 Vbias.n3387 Vbias.n3386 1.5505
R15495 Vbias.n3378 Vbias.n3213 1.5505
R15496 Vbias.n3352 Vbias.n3351 1.5505
R15497 Vbias.n3349 Vbias.n3348 1.5505
R15498 Vbias.n3338 Vbias.n3239 1.5505
R15499 Vbias.n3313 Vbias.n3312 1.5505
R15500 Vbias.n3311 Vbias.n3310 1.5505
R15501 Vbias.n3302 Vbias.n3260 1.5505
R15502 Vbias.n3437 Vbias.n3436 1.5505
R15503 Vbias.n3696 Vbias.n3695 1.5505
R15504 Vbias.n3694 Vbias.n3693 1.5505
R15505 Vbias.n3685 Vbias.n3453 1.5505
R15506 Vbias.n3658 Vbias.n3657 1.5505
R15507 Vbias.n3656 Vbias.n3655 1.5505
R15508 Vbias.n3647 Vbias.n3482 1.5505
R15509 Vbias.n3621 Vbias.n3620 1.5505
R15510 Vbias.n3618 Vbias.n3617 1.5505
R15511 Vbias.n3607 Vbias.n3508 1.5505
R15512 Vbias.n3582 Vbias.n3581 1.5505
R15513 Vbias.n3580 Vbias.n3579 1.5505
R15514 Vbias.n3571 Vbias.n3529 1.5505
R15515 Vbias.n3706 Vbias.n3705 1.5505
R15516 Vbias.n4231 Vbias.n4230 1.5505
R15517 Vbias.n4229 Vbias.n4228 1.5505
R15518 Vbias.n4220 Vbias.n4012 1.5505
R15519 Vbias.n4215 Vbias.n4214 1.5505
R15520 Vbias.n4212 Vbias.n4211 1.5505
R15521 Vbias.n4040 Vbias.n4037 1.5505
R15522 Vbias.n4197 Vbias.n4196 1.5505
R15523 Vbias.n4195 Vbias.n4194 1.5505
R15524 Vbias.n4186 Vbias.n4054 1.5505
R15525 Vbias.n4239 Vbias.n4000 1.5505
R15526 Vbias.n4241 Vbias.n3980 1.5505
R15527 Vbias.n4250 Vbias.n4249 1.5505
R15528 Vbias.n4115 Vbias.n4114 1.5505
R15529 Vbias.n4099 Vbias.n4089 1.5505
R15530 Vbias.n4125 Vbias.n4124 1.5505
R15531 Vbias.n4128 Vbias.n4127 1.5505
R15532 Vbias.n4087 Vbias.n4079 1.5505
R15533 Vbias.n4141 Vbias.n4140 1.5505
R15534 Vbias.n4148 Vbias.n4143 1.5505
R15535 Vbias.n4164 Vbias.n4163 1.5505
R15536 Vbias.n4177 Vbias.n4166 1.5505
R15537 Vbias.n4180 Vbias.n4179 1.5505
R15538 Vbias.n4182 Vbias.n4181 1.5505
R15539 Vbias.n4112 Vbias.n4111 1.5505
R15540 Vbias.n3157 Vbias.n3156 1.5505
R15541 Vbias.n3155 Vbias.n3154 1.5505
R15542 Vbias.n3146 Vbias.n2914 1.5505
R15543 Vbias.n3119 Vbias.n3118 1.5505
R15544 Vbias.n3117 Vbias.n3116 1.5505
R15545 Vbias.n3108 Vbias.n2943 1.5505
R15546 Vbias.n3082 Vbias.n3081 1.5505
R15547 Vbias.n3079 Vbias.n3078 1.5505
R15548 Vbias.n3068 Vbias.n2969 1.5505
R15549 Vbias.n3043 Vbias.n3042 1.5505
R15550 Vbias.n3041 Vbias.n3040 1.5505
R15551 Vbias.n3032 Vbias.n2990 1.5505
R15552 Vbias.n3167 Vbias.n3166 1.5505
R15553 Vbias.n4833 Vbias.n4832 1.5505
R15554 Vbias.n4831 Vbias.n4830 1.5505
R15555 Vbias.n4822 Vbias.n2675 1.5505
R15556 Vbias.n4795 Vbias.n4794 1.5505
R15557 Vbias.n4793 Vbias.n4792 1.5505
R15558 Vbias.n4784 Vbias.n2704 1.5505
R15559 Vbias.n4758 Vbias.n4757 1.5505
R15560 Vbias.n4755 Vbias.n4754 1.5505
R15561 Vbias.n4744 Vbias.n2730 1.5505
R15562 Vbias.n4719 Vbias.n4718 1.5505
R15563 Vbias.n4717 Vbias.n4716 1.5505
R15564 Vbias.n4708 Vbias.n2751 1.5505
R15565 Vbias.n2897 Vbias.n2666 1.5505
R15566 Vbias.n4677 Vbias.n4676 1.5505
R15567 Vbias.n4674 Vbias.n4555 1.5505
R15568 Vbias.n4667 Vbias.n4666 1.5505
R15569 Vbias.n4665 Vbias.n4664 1.5505
R15570 Vbias.n4657 Vbias.n4656 1.5505
R15571 Vbias.n4654 Vbias.n4653 1.5505
R15572 Vbias.n4651 Vbias.n4593 1.5505
R15573 Vbias.n4649 Vbias.n4648 1.5505
R15574 Vbias.n4646 Vbias.n4645 1.5505
R15575 Vbias.n4643 Vbias.n2438 1.5505
R15576 Vbias.n5033 Vbias.n5032 1.5505
R15577 Vbias.n7446 Vbias.n7445 1.5505
R15578 Vbias.n7444 Vbias.n7443 1.5505
R15579 Vbias.n7435 Vbias.n7347 1.5505
R15580 Vbias.n7430 Vbias.n7429 1.5505
R15581 Vbias.n7427 Vbias.n7426 1.5505
R15582 Vbias.n7370 Vbias.n7367 1.5505
R15583 Vbias.n7412 Vbias.n7411 1.5505
R15584 Vbias.n7410 Vbias.n7409 1.5505
R15585 Vbias.n7400 Vbias.n7385 1.5505
R15586 Vbias.n7454 Vbias.n7339 1.5505
R15587 Vbias.n7456 Vbias.n7324 1.5505
R15588 Vbias.n7465 Vbias.n7464 1.5505
R15589 Vbias.n6648 Vbias.n6647 1.5505
R15590 Vbias.n6137 Vbias.n6134 1.5505
R15591 Vbias.n6636 Vbias.n6635 1.5505
R15592 Vbias.n6633 Vbias.n6632 1.5505
R15593 Vbias.n6630 Vbias.n6154 1.5505
R15594 Vbias.n6628 Vbias.n6627 1.5505
R15595 Vbias.n6625 Vbias.n6624 1.5505
R15596 Vbias.n6617 Vbias.n6616 1.5505
R15597 Vbias.n6615 Vbias.n6614 1.5505
R15598 Vbias.n6607 Vbias.n6606 1.5505
R15599 Vbias.n6605 Vbias.n6604 1.5505
R15600 Vbias.n6602 Vbias.n6207 1.5505
R15601 Vbias.n6574 Vbias.n6573 1.5505
R15602 Vbias.n6571 Vbias.n6364 1.5505
R15603 Vbias.n6569 Vbias.n6568 1.5505
R15604 Vbias.n6566 Vbias.n6565 1.5505
R15605 Vbias.n6563 Vbias.n6372 1.5505
R15606 Vbias.n6561 Vbias.n6560 1.5505
R15607 Vbias.n6558 Vbias.n6557 1.5505
R15608 Vbias.n6550 Vbias.n6549 1.5505
R15609 Vbias.n6548 Vbias.n6547 1.5505
R15610 Vbias.n6540 Vbias.n6539 1.5505
R15611 Vbias.n6538 Vbias.n6537 1.5505
R15612 Vbias.n6535 Vbias.n6444 1.5505
R15613 Vbias.n7587 Vbias.n7586 1.5505
R15614 Vbias.n7584 Vbias.n859 1.5505
R15615 Vbias.n7582 Vbias.n7581 1.5505
R15616 Vbias.n7579 Vbias.n7578 1.5505
R15617 Vbias.n7576 Vbias.n867 1.5505
R15618 Vbias.n7574 Vbias.n7573 1.5505
R15619 Vbias.n7571 Vbias.n7570 1.5505
R15620 Vbias.n7563 Vbias.n7562 1.5505
R15621 Vbias.n7561 Vbias.n7560 1.5505
R15622 Vbias.n7553 Vbias.n7552 1.5505
R15623 Vbias.n7551 Vbias.n7550 1.5505
R15624 Vbias.n7548 Vbias.n898 1.5505
R15625 Vbias.n7321 Vbias.n7320 1.5505
R15626 Vbias.n1043 Vbias.n1031 1.5505
R15627 Vbias.n7308 Vbias.n1044 1.5505
R15628 Vbias.n7306 Vbias.n1047 1.5505
R15629 Vbias.n1064 Vbias.n1052 1.5505
R15630 Vbias.n7293 Vbias.n1065 1.5505
R15631 Vbias.n7291 Vbias.n1068 1.5505
R15632 Vbias.n7240 Vbias.n7229 1.5505
R15633 Vbias.n7278 Vbias.n7277 1.5505
R15634 Vbias.n7275 Vbias.n7274 1.5505
R15635 Vbias.n7272 Vbias.n7241 1.5505
R15636 Vbias.n7263 Vbias.n7262 1.5505
R15637 Vbias.n946 Vbias.n931 1.5505
R15638 Vbias.n948 Vbias.n934 1.5505
R15639 Vbias.n7515 Vbias.n949 1.5505
R15640 Vbias.n7513 Vbias.n952 1.5505
R15641 Vbias.n969 Vbias.n957 1.5505
R15642 Vbias.n7500 Vbias.n970 1.5505
R15643 Vbias.n7498 Vbias.n973 1.5505
R15644 Vbias.n990 Vbias.n979 1.5505
R15645 Vbias.n7484 Vbias.n7483 1.5505
R15646 Vbias.n7481 Vbias.n7480 1.5505
R15647 Vbias.n7478 Vbias.n991 1.5505
R15648 Vbias.n7470 Vbias.n7469 1.5505
R15649 Vbias.n6361 Vbias.n780 1.5505
R15650 Vbias.n6359 Vbias.n783 1.5505
R15651 Vbias.n7636 Vbias.n794 1.5505
R15652 Vbias.n7634 Vbias.n797 1.5505
R15653 Vbias.n814 Vbias.n802 1.5505
R15654 Vbias.n7621 Vbias.n815 1.5505
R15655 Vbias.n7619 Vbias.n818 1.5505
R15656 Vbias.n835 Vbias.n824 1.5505
R15657 Vbias.n7606 Vbias.n7605 1.5505
R15658 Vbias.n7603 Vbias.n7602 1.5505
R15659 Vbias.n7600 Vbias.n836 1.5505
R15660 Vbias.n7592 Vbias.n7591 1.5505
R15661 Vbias.n6312 Vbias.n6311 1.5505
R15662 Vbias.n6315 Vbias.n6314 1.5505
R15663 Vbias.n6317 Vbias.n6275 1.5505
R15664 Vbias.n6326 Vbias.n6325 1.5505
R15665 Vbias.n6329 Vbias.n6328 1.5505
R15666 Vbias.n6331 Vbias.n6257 1.5505
R15667 Vbias.n6340 Vbias.n6339 1.5505
R15668 Vbias.n6344 Vbias.n6343 1.5505
R15669 Vbias.n6342 Vbias.n6247 1.5505
R15670 Vbias.n6358 Vbias.n6357 1.5505
R15671 Vbias.n6581 Vbias.n6579 1.5505
R15672 Vbias.n6578 Vbias.n6229 1.5505
R15673 Vbias.n5841 Vbias.n5840 1.5505
R15674 Vbias.n5844 Vbias.n5843 1.5505
R15675 Vbias.n5856 Vbias.n1699 1.5505
R15676 Vbias.n5854 Vbias.n1701 1.5505
R15677 Vbias.n2051 Vbias.n2050 1.5505
R15678 Vbias.n1480 Vbias.n1470 1.5505
R15679 Vbias.n6667 Vbias.n6666 1.5505
R15680 Vbias.n6664 Vbias.n6663 1.5505
R15681 Vbias.n6661 Vbias.n1481 1.5505
R15682 Vbias.n6653 Vbias.n6652 1.5505
R15683 Vbias.n5755 Vbias.n5754 1.5505
R15684 Vbias.n5758 Vbias.n5757 1.5505
R15685 Vbias.n5760 Vbias.n2102 1.5505
R15686 Vbias.n5769 Vbias.n5768 1.5505
R15687 Vbias.n5772 Vbias.n5771 1.5505
R15688 Vbias.n5774 Vbias.n2086 1.5505
R15689 Vbias.n5784 Vbias.n5783 1.5505
R15690 Vbias.n5803 Vbias.n5786 1.5505
R15691 Vbias.n5812 Vbias.n5811 1.5505
R15692 Vbias.n5815 Vbias.n5814 1.5505
R15693 Vbias.n5817 Vbias.n2069 1.5505
R15694 Vbias.n5826 Vbias.n5825 1.5505
R15695 Vbias.n5669 Vbias.n5668 1.5505
R15696 Vbias.n5681 Vbias.n5680 1.5505
R15697 Vbias.n5685 Vbias.n5683 1.5505
R15698 Vbias.n5682 Vbias.n2177 1.5505
R15699 Vbias.n5699 Vbias.n5698 1.5505
R15700 Vbias.n5704 Vbias.n5702 1.5505
R15701 Vbias.n5701 Vbias.n2159 1.5505
R15702 Vbias.n5714 Vbias.n2141 1.5505
R15703 Vbias.n5723 Vbias.n5722 1.5505
R15704 Vbias.n5726 Vbias.n5725 1.5505
R15705 Vbias.n5728 Vbias.n2124 1.5505
R15706 Vbias.n5737 Vbias.n5736 1.5505
R15707 Vbias.n5595 Vbias.n5594 1.5505
R15708 Vbias.n5607 Vbias.n5606 1.5505
R15709 Vbias.n5611 Vbias.n5609 1.5505
R15710 Vbias.n5608 Vbias.n5574 1.5505
R15711 Vbias.n5625 Vbias.n5624 1.5505
R15712 Vbias.n5630 Vbias.n5628 1.5505
R15713 Vbias.n5627 Vbias.n5556 1.5505
R15714 Vbias.n5640 Vbias.n2212 1.5505
R15715 Vbias.n5649 Vbias.n5648 1.5505
R15716 Vbias.n5652 Vbias.n5651 1.5505
R15717 Vbias.n5654 Vbias.n2195 1.5505
R15718 Vbias.n5663 Vbias.n5662 1.5505
R15719 Vbias.n251 Vbias.n89 1.5505
R15720 Vbias.n249 Vbias.n92 1.5505
R15721 Vbias.n7992 Vbias.n103 1.5505
R15722 Vbias.n7990 Vbias.n106 1.5505
R15723 Vbias.n123 Vbias.n111 1.5505
R15724 Vbias.n7977 Vbias.n124 1.5505
R15725 Vbias.n7975 Vbias.n127 1.5505
R15726 Vbias.n143 Vbias.n132 1.5505
R15727 Vbias.n7962 Vbias.n7961 1.5505
R15728 Vbias.n7959 Vbias.n7958 1.5505
R15729 Vbias.n7956 Vbias.n144 1.5505
R15730 Vbias.n7948 Vbias.n7947 1.5505
R15731 Vbias.n258 Vbias.n257 1.5505
R15732 Vbias.n246 Vbias.n231 1.5505
R15733 Vbias.n272 Vbias.n271 1.5505
R15734 Vbias.n275 Vbias.n274 1.5505
R15735 Vbias.n229 Vbias.n212 1.5505
R15736 Vbias.n291 Vbias.n290 1.5505
R15737 Vbias.n295 Vbias.n294 1.5505
R15738 Vbias.n206 Vbias.n198 1.5505
R15739 Vbias.n311 Vbias.n310 1.5505
R15740 Vbias.n314 Vbias.n313 1.5505
R15741 Vbias.n196 Vbias.n179 1.5505
R15742 Vbias.n354 Vbias.n353 1.5505
R15743 Vbias.n7933 Vbias.n7932 1.5505
R15744 Vbias.n7931 Vbias.n7930 1.5505
R15745 Vbias.n7928 Vbias.n357 1.5505
R15746 Vbias.n7921 Vbias.n7920 1.5505
R15747 Vbias.n7919 Vbias.n7918 1.5505
R15748 Vbias.n7916 Vbias.n381 1.5505
R15749 Vbias.n7909 Vbias.n7908 1.5505
R15750 Vbias.n7906 Vbias.n7905 1.5505
R15751 Vbias.n7903 Vbias.n405 1.5505
R15752 Vbias.n7896 Vbias.n7895 1.5505
R15753 Vbias.n7894 Vbias.n7893 1.5505
R15754 Vbias.n7891 Vbias.n428 1.5505
R15755 Vbias.n7867 Vbias.n7866 1.5505
R15756 Vbias.n7865 Vbias.n7864 1.5505
R15757 Vbias.n7862 Vbias.n463 1.5505
R15758 Vbias.n7855 Vbias.n7854 1.5505
R15759 Vbias.n7853 Vbias.n7852 1.5505
R15760 Vbias.n7850 Vbias.n487 1.5505
R15761 Vbias.n7843 Vbias.n7842 1.5505
R15762 Vbias.n7840 Vbias.n7839 1.5505
R15763 Vbias.n7837 Vbias.n511 1.5505
R15764 Vbias.n7830 Vbias.n7829 1.5505
R15765 Vbias.n7828 Vbias.n7827 1.5505
R15766 Vbias.n7825 Vbias.n534 1.5505
R15767 Vbias.n7798 Vbias.n7797 1.5505
R15768 Vbias.n7796 Vbias.n7795 1.5505
R15769 Vbias.n7793 Vbias.n577 1.5505
R15770 Vbias.n7786 Vbias.n7785 1.5505
R15771 Vbias.n7784 Vbias.n7783 1.5505
R15772 Vbias.n7781 Vbias.n601 1.5505
R15773 Vbias.n7774 Vbias.n7773 1.5505
R15774 Vbias.n7771 Vbias.n7770 1.5505
R15775 Vbias.n7768 Vbias.n625 1.5505
R15776 Vbias.n7761 Vbias.n7760 1.5505
R15777 Vbias.n7759 Vbias.n7758 1.5505
R15778 Vbias.n7756 Vbias.n648 1.5505
R15779 Vbias.n7719 Vbias.n7718 1.5505
R15780 Vbias.n702 Vbias.n699 1.5505
R15781 Vbias.n7707 Vbias.n7706 1.5505
R15782 Vbias.n7704 Vbias.n7703 1.5505
R15783 Vbias.n7696 Vbias.n7695 1.5505
R15784 Vbias.n7694 Vbias.n7693 1.5505
R15785 Vbias.n7681 Vbias.n7680 1.5505
R15786 Vbias.n7679 Vbias.n7678 1.5505
R15787 Vbias.n7670 Vbias.n740 1.5505
R15788 Vbias.n7722 Vbias.n7721 1.5505
R15789 Vbias.n7730 Vbias.n684 1.5505
R15790 Vbias.n7732 Vbias.n682 1.5505
R15791 Vbias.n6128 Vbias.n6127 1.5505
R15792 Vbias.n770 Vbias.n769 1.5505
R15793 Vbias.n7661 Vbias.n7660 1.5505
R15794 Vbias.n7658 Vbias.n7657 1.5505
R15795 Vbias.n7655 Vbias.n771 1.5505
R15796 Vbias.n6514 Vbias.n6513 1.5505
R15797 Vbias.n6523 Vbias.n924 1.5505
R15798 Vbias.n7535 Vbias.n7534 1.5505
R15799 Vbias.n7537 Vbias.n921 1.5505
R15800 Vbias.n7540 Vbias.n7539 1.5505
R15801 Vbias.n7942 Vbias.n7941 1.5505
R15802 Vbias.n7883 Vbias.n7882 1.5505
R15803 Vbias.n7881 Vbias.n7880 1.5505
R15804 Vbias.n7817 Vbias.n7816 1.5505
R15805 Vbias.n7814 Vbias.n7813 1.5505
R15806 Vbias.n561 Vbias.n558 1.5505
R15807 Vbias.n7748 Vbias.n7747 1.5505
R15808 Vbias.n7746 Vbias.n7745 1.5505
R15809 Vbias.n338 Vbias.n337 1.5505
R15810 Vbias.n1717 Vbias.n1706 1.5505
R15811 Vbias.n2049 Vbias.n2048 1.5505
R15812 Vbias.n5027 Vbias.n5026 1.5505
R15813 Vbias.n2588 Vbias.n2585 1.5505
R15814 Vbias.n5549 Vbias.n5548 1.5505
R15815 Vbias.n5546 Vbias.n5545 1.5505
R15816 Vbias.n2236 Vbias.n2233 1.5505
R15817 Vbias.n5529 Vbias.n5528 1.5505
R15818 Vbias.n5527 Vbias.n5526 1.5505
R15819 Vbias.n5873 Vbias.n5872 1.5505
R15820 Vbias.n5870 Vbias.n5869 1.5505
R15821 Vbias.n1683 Vbias.n1680 1.5505
R15822 Vbias.n1456 Vbias.n1449 1.5505
R15823 Vbias.n6691 Vbias.n6690 1.5505
R15824 Vbias.n6746 Vbias.n6745 1.5505
R15825 Vbias.n6743 Vbias.n6742 1.5505
R15826 Vbias.n6740 Vbias.n6718 1.5505
R15827 Vbias.n6716 Vbias.n6715 1.5505
R15828 Vbias.n6713 Vbias.n6694 1.5505
R15829 Vbias.n4989 Vbias.n4988 1.5505
R15830 Vbias.n5003 Vbias.n5002 1.5505
R15831 Vbias.n5006 Vbias.n5005 1.5505
R15832 Vbias.n2894 Vbias.n2662 1.5505
R15833 Vbias.n4920 Vbias.n4919 1.5505
R15834 Vbias.n4923 Vbias.n4922 1.5505
R15835 Vbias.n4921 Vbias.n2648 1.5505
R15836 Vbias.n4942 Vbias.n4941 1.5505
R15837 Vbias.n4946 Vbias.n4945 1.5505
R15838 Vbias.n4944 Vbias.n2634 1.5505
R15839 Vbias.n4957 Vbias.n2618 1.5505
R15840 Vbias.n4968 Vbias.n4967 1.5505
R15841 Vbias.n4971 Vbias.n4970 1.5505
R15842 Vbias.n4975 Vbias.n2604 1.5505
R15843 Vbias.n4986 Vbias.n4985 1.5505
R15844 Vbias.n8059 Vbias.n8058 1.5505
R15845 Vbias.n33 Vbias.n30 1.5505
R15846 Vbias.n8047 Vbias.n8046 1.5505
R15847 Vbias.n8044 Vbias.n8043 1.5505
R15848 Vbias.n8036 Vbias.n8035 1.5505
R15849 Vbias.n8034 Vbias.n8033 1.5505
R15850 Vbias.n8021 Vbias.n8020 1.5505
R15851 Vbias.n8019 Vbias.n8018 1.5505
R15852 Vbias.n8010 Vbias.n71 1.5505
R15853 Vbias.n8062 Vbias.n8061 1.5505
R15854 Vbias.n8070 Vbias.n15 1.5505
R15855 Vbias.n8072 Vbias.n13 1.5505
R15856 Vbias.n6109 Vbias 1.54738
R15857 Vbias.n2016 Vbias 1.54738
R15858 Vbias.n1969 Vbias 1.54738
R15859 Vbias.n1935 Vbias 1.54738
R15860 Vbias.n1898 Vbias 1.54738
R15861 Vbias.n1869 Vbias 1.54738
R15862 Vbias.n1821 Vbias 1.54738
R15863 Vbias.n2033 Vbias 1.54738
R15864 Vbias.n8085 Vbias.n8084 1.37007
R15865 Vbias.n8086 Vbias.n8085 1.36735
R15866 Vbias.n1841 Vbias.n1840 1.32825
R15867 Vbias.n4899 Vbias.n4898 1.28905
R15868 Vbias.n4900 Vbias.n4899 1.28905
R15869 Vbias.n4896 Vbias.n4895 1.28905
R15870 Vbias.n6110 Vbias.n6109 1.1418
R15871 Vbias.n2016 Vbias.n2015 1.1418
R15872 Vbias.n1970 Vbias.n1969 1.1418
R15873 Vbias.n1936 Vbias.n1935 1.1418
R15874 Vbias.n1899 Vbias.n1898 1.1418
R15875 Vbias.n1821 Vbias.n1820 1.1418
R15876 Vbias.n1870 Vbias.n1869 1.1418
R15877 Vbias.n2034 Vbias.n2033 1.1418
R15878 Vbias.n6124 Vbias.n1507 1.11191
R15879 Vbias.n7943 Vbias 1.06886
R15880 Vbias.n1746 Vbias.n1734 1.06843
R15881 Vbias.n337 Vbias.n168 1.01952
R15882 Vbias Vbias.n4266 1.01137
R15883 Vbias Vbias.n4299 1.01137
R15884 Vbias Vbias.n4332 1.01137
R15885 Vbias.n4334 Vbias 1.01137
R15886 Vbias.n4359 Vbias 1.01137
R15887 Vbias.n4384 Vbias 1.01137
R15888 Vbias.n6110 Vbias 1.01137
R15889 Vbias.n2015 Vbias 1.01137
R15890 Vbias.n1970 Vbias 1.01137
R15891 Vbias.n1936 Vbias 1.01137
R15892 Vbias.n1899 Vbias 1.01137
R15893 Vbias.n1820 Vbias 1.01137
R15894 Vbias.n1870 Vbias 1.01137
R15895 Vbias.n2034 Vbias 1.01137
R15896 Vbias Vbias.n2407 1.01137
R15897 Vbias.n5075 Vbias 1.01137
R15898 Vbias Vbias.n2392 1.01137
R15899 Vbias Vbias.n2376 1.01137
R15900 Vbias Vbias.n5174 1.01137
R15901 Vbias.n5163 Vbias 1.01137
R15902 Vbias Vbias.n2252 1.01137
R15903 Vbias.n5493 Vbias 1.01137
R15904 Vbias.n5468 Vbias 1.01137
R15905 Vbias.n5458 Vbias 1.01137
R15906 Vbias Vbias.n1660 1.01137
R15907 Vbias Vbias.n1644 1.01137
R15908 Vbias Vbias.n5947 1.01137
R15909 Vbias.n6096 Vbias 1.01137
R15910 Vbias Vbias.n6094 1.01137
R15911 Vbias Vbias.n6086 1.01137
R15912 Vbias Vbias.n6805 1.01137
R15913 Vbias.n6794 Vbias 1.01137
R15914 Vbias Vbias.n6792 1.01137
R15915 Vbias Vbias.n6784 1.01137
R15916 Vbias.n7047 Vbias 1.01137
R15917 Vbias.n7060 Vbias 1.01137
R15918 Vbias.n7062 Vbias 1.01137
R15919 Vbias.n7079 Vbias 1.01137
R15920 Vbias.n7153 Vbias 1.01137
R15921 Vbias.n7166 Vbias 1.01137
R15922 Vbias.n7168 Vbias 1.01137
R15923 Vbias.n7185 Vbias 1.01137
R15924 Vbias.n1195 Vbias 1.01137
R15925 Vbias Vbias.n1086 1.01137
R15926 Vbias Vbias.n7204 1.01137
R15927 Vbias.n6928 Vbias 1.01137
R15928 Vbias Vbias.n1167 1.01137
R15929 Vbias Vbias.n7100 1.01137
R15930 Vbias.n6836 Vbias 1.01137
R15931 Vbias.n6879 Vbias 1.01137
R15932 Vbias.n6898 Vbias 1.01137
R15933 Vbias.n5978 Vbias 1.01137
R15934 Vbias.n6021 Vbias 1.01137
R15935 Vbias Vbias.n6024 1.01137
R15936 Vbias.n5299 Vbias 1.01137
R15937 Vbias.n5334 Vbias 1.01137
R15938 Vbias.n5342 Vbias 1.01137
R15939 Vbias.n5205 Vbias 1.01137
R15940 Vbias.n5248 Vbias 1.01137
R15941 Vbias.n5268 Vbias 1.01137
R15942 Vbias.n2467 Vbias 1.01137
R15943 Vbias.n2502 Vbias 1.01137
R15944 Vbias.n2510 Vbias 1.01137
R15945 Vbias.n4438 Vbias 1.01137
R15946 Vbias Vbias.n4509 1.01137
R15947 Vbias Vbias.n4495 1.01137
R15948 Vbias.n3975 Vbias 1.01137
R15949 Vbias Vbias.n3722 1.01137
R15950 Vbias Vbias.n3751 1.01137
R15951 Vbias.n3889 Vbias 1.01137
R15952 Vbias Vbias.n3777 1.01137
R15953 Vbias.n3798 Vbias 1.01137
R15954 Vbias.n3437 Vbias 1.01137
R15955 Vbias Vbias.n3184 1.01137
R15956 Vbias Vbias.n3213 1.01137
R15957 Vbias.n3351 Vbias 1.01137
R15958 Vbias Vbias.n3239 1.01137
R15959 Vbias.n3260 Vbias 1.01137
R15960 Vbias.n3706 Vbias 1.01137
R15961 Vbias Vbias.n3453 1.01137
R15962 Vbias Vbias.n3482 1.01137
R15963 Vbias.n3620 Vbias 1.01137
R15964 Vbias Vbias.n3508 1.01137
R15965 Vbias.n3529 Vbias 1.01137
R15966 Vbias Vbias.n4000 1.01137
R15967 Vbias Vbias.n4012 1.01137
R15968 Vbias.n4214 Vbias 1.01137
R15969 Vbias Vbias.n4037 1.01137
R15970 Vbias.n4054 Vbias 1.01137
R15971 Vbias Vbias.n4112 1.01137
R15972 Vbias Vbias.n4125 1.01137
R15973 Vbias Vbias.n4141 1.01137
R15974 Vbias Vbias.n4164 1.01137
R15975 Vbias.n4181 Vbias 1.01137
R15976 Vbias.n3167 Vbias 1.01137
R15977 Vbias Vbias.n2914 1.01137
R15978 Vbias Vbias.n2943 1.01137
R15979 Vbias.n3081 Vbias 1.01137
R15980 Vbias Vbias.n2969 1.01137
R15981 Vbias.n2990 Vbias 1.01137
R15982 Vbias.n2897 Vbias 1.01137
R15983 Vbias Vbias.n2675 1.01137
R15984 Vbias Vbias.n2704 1.01137
R15985 Vbias.n4757 Vbias 1.01137
R15986 Vbias Vbias.n2730 1.01137
R15987 Vbias.n2751 Vbias 1.01137
R15988 Vbias.n4666 Vbias 1.01137
R15989 Vbias.n4656 Vbias 1.01137
R15990 Vbias Vbias.n4654 1.01137
R15991 Vbias Vbias.n4646 1.01137
R15992 Vbias Vbias.n7339 1.01137
R15993 Vbias Vbias.n7347 1.01137
R15994 Vbias.n7429 Vbias 1.01137
R15995 Vbias Vbias.n7367 1.01137
R15996 Vbias.n7385 Vbias 1.01137
R15997 Vbias.n6635 Vbias 1.01137
R15998 Vbias.n6627 Vbias 1.01137
R15999 Vbias.n6625 Vbias 1.01137
R16000 Vbias.n6615 Vbias 1.01137
R16001 Vbias Vbias.n6207 1.01137
R16002 Vbias.n6568 Vbias 1.01137
R16003 Vbias.n6560 Vbias 1.01137
R16004 Vbias.n6558 Vbias 1.01137
R16005 Vbias.n6548 Vbias 1.01137
R16006 Vbias.n6444 Vbias 1.01137
R16007 Vbias.n7581 Vbias 1.01137
R16008 Vbias.n7573 Vbias 1.01137
R16009 Vbias.n7571 Vbias 1.01137
R16010 Vbias.n7561 Vbias 1.01137
R16011 Vbias Vbias.n898 1.01137
R16012 Vbias.n7321 Vbias 1.01137
R16013 Vbias Vbias.n1047 1.01137
R16014 Vbias Vbias.n1068 1.01137
R16015 Vbias.n7277 Vbias 1.01137
R16016 Vbias.n7262 Vbias 1.01137
R16017 Vbias Vbias.n946 1.01137
R16018 Vbias Vbias.n952 1.01137
R16019 Vbias Vbias.n973 1.01137
R16020 Vbias.n7483 Vbias 1.01137
R16021 Vbias.n7469 Vbias 1.01137
R16022 Vbias.n6361 Vbias 1.01137
R16023 Vbias Vbias.n797 1.01137
R16024 Vbias Vbias.n818 1.01137
R16025 Vbias.n7605 Vbias 1.01137
R16026 Vbias.n7591 Vbias 1.01137
R16027 Vbias Vbias.n6312 1.01137
R16028 Vbias Vbias.n6326 1.01137
R16029 Vbias Vbias.n6340 1.01137
R16030 Vbias.n6342 Vbias 1.01137
R16031 Vbias.n6578 Vbias 1.01137
R16032 Vbias Vbias.n5841 1.01137
R16033 Vbias Vbias.n1701 1.01137
R16034 Vbias.n2049 Vbias 1.01137
R16035 Vbias.n6666 Vbias 1.01137
R16036 Vbias.n6652 Vbias 1.01137
R16037 Vbias Vbias.n5755 1.01137
R16038 Vbias Vbias.n5769 1.01137
R16039 Vbias Vbias.n5784 1.01137
R16040 Vbias Vbias.n5812 1.01137
R16041 Vbias Vbias.n5826 1.01137
R16042 Vbias.n5668 Vbias 1.01137
R16043 Vbias.n5682 Vbias 1.01137
R16044 Vbias.n5701 Vbias 1.01137
R16045 Vbias Vbias.n5723 1.01137
R16046 Vbias Vbias.n5737 1.01137
R16047 Vbias.n5594 Vbias 1.01137
R16048 Vbias.n5608 Vbias 1.01137
R16049 Vbias.n5627 Vbias 1.01137
R16050 Vbias Vbias.n5649 1.01137
R16051 Vbias Vbias.n5663 1.01137
R16052 Vbias.n251 Vbias 1.01137
R16053 Vbias Vbias.n106 1.01137
R16054 Vbias Vbias.n127 1.01137
R16055 Vbias.n7961 Vbias 1.01137
R16056 Vbias.n7947 Vbias 1.01137
R16057 Vbias Vbias.n272 1.01137
R16058 Vbias Vbias.n291 1.01137
R16059 Vbias.n294 Vbias 1.01137
R16060 Vbias Vbias.n311 1.01137
R16061 Vbias Vbias.n354 1.01137
R16062 Vbias Vbias.n357 1.01137
R16063 Vbias Vbias.n381 1.01137
R16064 Vbias.n7908 Vbias 1.01137
R16065 Vbias Vbias.n405 1.01137
R16066 Vbias Vbias.n428 1.01137
R16067 Vbias Vbias.n463 1.01137
R16068 Vbias Vbias.n487 1.01137
R16069 Vbias.n7842 Vbias 1.01137
R16070 Vbias Vbias.n511 1.01137
R16071 Vbias Vbias.n534 1.01137
R16072 Vbias Vbias.n577 1.01137
R16073 Vbias Vbias.n601 1.01137
R16074 Vbias.n7773 Vbias 1.01137
R16075 Vbias Vbias.n625 1.01137
R16076 Vbias Vbias.n648 1.01137
R16077 Vbias.n7721 Vbias 1.01137
R16078 Vbias.n7706 Vbias 1.01137
R16079 Vbias.n7704 Vbias 1.01137
R16080 Vbias.n7694 Vbias 1.01137
R16081 Vbias Vbias.n740 1.01137
R16082 Vbias Vbias.n770 1.01137
R16083 Vbias Vbias.n924 1.01137
R16084 Vbias Vbias.n7814 1.01137
R16085 Vbias.n337 Vbias 1.01137
R16086 Vbias Vbias.n5546 1.01137
R16087 Vbias Vbias.n5870 1.01137
R16088 Vbias Vbias.n6743 1.01137
R16089 Vbias.n5003 Vbias 1.01137
R16090 Vbias.n2894 Vbias 1.01137
R16091 Vbias.n4921 Vbias 1.01137
R16092 Vbias.n4944 Vbias 1.01137
R16093 Vbias Vbias.n4968 1.01137
R16094 Vbias Vbias.n4986 1.01137
R16095 Vbias.n8061 Vbias 1.01137
R16096 Vbias.n8046 Vbias 1.01137
R16097 Vbias.n8044 Vbias 1.01137
R16098 Vbias.n8034 Vbias 1.01137
R16099 Vbias.n71 Vbias 1.01137
R16100 Vbias.n1843 Vbias.n1842 0.645183
R16101 Vbias.n1838 Vbias.n1837 0.645183
R16102 Vbias.n1833 Vbias.n1832 0.645183
R16103 Vbias.n1828 Vbias.n1827 0.645183
R16104 Vbias.n1823 Vbias.n1822 0.645183
R16105 Vbias.n2021 Vbias.n2020 0.645183
R16106 Vbias.n2026 Vbias.n2025 0.645183
R16107 Vbias.n2030 Vbias.n2029 0.645183
R16108 Vbias.n4886 Vbias.n0 0.6205
R16109 Vbias.n4266 Vbias.n4255 0.606478
R16110 Vbias.n4268 Vbias.n4267 0.606478
R16111 Vbias.n4301 Vbias.n4300 0.606478
R16112 Vbias.n4334 Vbias.n4333 0.606478
R16113 Vbias.n4358 Vbias.n2809 0.606478
R16114 Vbias.n4383 Vbias.n2796 0.606478
R16115 Vbias.n5053 Vbias.n5052 0.606478
R16116 Vbias.n5073 Vbias.n5072 0.606478
R16117 Vbias.n5075 Vbias.n5074 0.606478
R16118 Vbias.n5096 Vbias.n5095 0.606478
R16119 Vbias.n5116 Vbias.n5115 0.606478
R16120 Vbias.n5176 Vbias.n5175 0.606478
R16121 Vbias.n5161 Vbias.n2357 0.606478
R16122 Vbias.n5163 Vbias.n5162 0.606478
R16123 Vbias.n5502 Vbias.n2253 0.606478
R16124 Vbias.n2293 Vbias.n2269 0.606478
R16125 Vbias.n5440 Vbias.n5417 0.606478
R16126 Vbias.n5467 Vbias.n5441 0.606478
R16127 Vbias.n5458 Vbias.n5457 0.606478
R16128 Vbias.n5893 Vbias.n5892 0.606478
R16129 Vbias.n5913 Vbias.n5912 0.606478
R16130 Vbias.n5949 Vbias.n5948 0.606478
R16131 Vbias.n1621 Vbias.n1620 0.606478
R16132 Vbias.n6096 Vbias.n6095 0.606478
R16133 Vbias.n6088 Vbias.n6087 0.606478
R16134 Vbias.n6080 Vbias.n6079 0.606478
R16135 Vbias.n6807 Vbias.n6806 0.606478
R16136 Vbias.n1420 Vbias.n1409 0.606478
R16137 Vbias.n6794 Vbias.n6793 0.606478
R16138 Vbias.n6786 Vbias.n6785 0.606478
R16139 Vbias.n7010 Vbias.n7009 0.606478
R16140 Vbias.n7032 Vbias.n7031 0.606478
R16141 Vbias.n7049 Vbias.n7048 0.606478
R16142 Vbias.n7061 Vbias.n7060 0.606478
R16143 Vbias.n7078 Vbias.n7077 0.606478
R16144 Vbias.n7095 Vbias.n7094 0.606478
R16145 Vbias.n7138 Vbias.n7137 0.606478
R16146 Vbias.n7155 Vbias.n7154 0.606478
R16147 Vbias.n7167 Vbias.n7166 0.606478
R16148 Vbias.n7184 Vbias.n7183 0.606478
R16149 Vbias.n7201 Vbias.n7200 0.606478
R16150 Vbias.n1194 Vbias.n1193 0.606478
R16151 Vbias.n1244 Vbias.n1243 0.606478
R16152 Vbias.n1212 Vbias.n1211 0.606478
R16153 Vbias.n7206 Vbias.n7205 0.606478
R16154 Vbias.n7204 Vbias.n7203 0.606478
R16155 Vbias.n6927 Vbias.n6926 0.606478
R16156 Vbias.n6977 Vbias.n6976 0.606478
R16157 Vbias.n6945 Vbias.n6944 0.606478
R16158 Vbias.n7102 Vbias.n7101 0.606478
R16159 Vbias.n7100 Vbias.n7099 0.606478
R16160 Vbias.n6833 Vbias.n6832 0.606478
R16161 Vbias.n6835 Vbias.n6834 0.606478
R16162 Vbias.n6858 Vbias.n6857 0.606478
R16163 Vbias.n6881 Vbias.n6880 0.606478
R16164 Vbias.n6899 Vbias.n6898 0.606478
R16165 Vbias.n5975 Vbias.n5974 0.606478
R16166 Vbias.n5977 Vbias.n5976 0.606478
R16167 Vbias.n6000 Vbias.n5999 0.606478
R16168 Vbias.n6026 Vbias.n6025 0.606478
R16169 Vbias.n6024 Vbias.n6023 0.606478
R16170 Vbias.n5298 Vbias.n5297 0.606478
R16171 Vbias.n5385 Vbias.n5384 0.606478
R16172 Vbias.n5333 Vbias.n5332 0.606478
R16173 Vbias.n5355 Vbias.n5335 0.606478
R16174 Vbias.n5342 Vbias.n5341 0.606478
R16175 Vbias.n5202 Vbias.n5201 0.606478
R16176 Vbias.n5204 Vbias.n5203 0.606478
R16177 Vbias.n5227 Vbias.n5226 0.606478
R16178 Vbias.n5250 Vbias.n5249 0.606478
R16179 Vbias.n5269 Vbias.n5268 0.606478
R16180 Vbias.n2466 Vbias.n2465 0.606478
R16181 Vbias.n2553 Vbias.n2552 0.606478
R16182 Vbias.n2501 Vbias.n2500 0.606478
R16183 Vbias.n2523 Vbias.n2503 0.606478
R16184 Vbias.n2510 Vbias.n2509 0.606478
R16185 Vbias.n4540 Vbias.n4423 0.606478
R16186 Vbias.n4525 Vbias.n4524 0.606478
R16187 Vbias.n4511 Vbias.n4510 0.606478
R16188 Vbias.n4497 Vbias.n4496 0.606478
R16189 Vbias.n4495 Vbias.n4484 0.606478
R16190 Vbias.n3976 Vbias.n3975 0.606478
R16191 Vbias.n3964 Vbias.n3721 0.606478
R16192 Vbias.n3926 Vbias.n3750 0.606478
R16193 Vbias.n3889 Vbias.n3776 0.606478
R16194 Vbias.n3888 Vbias.n3887 0.606478
R16195 Vbias.n3850 Vbias.n3797 0.606478
R16196 Vbias.n3438 Vbias.n3437 0.606478
R16197 Vbias.n3426 Vbias.n3183 0.606478
R16198 Vbias.n3388 Vbias.n3212 0.606478
R16199 Vbias.n3351 Vbias.n3238 0.606478
R16200 Vbias.n3350 Vbias.n3349 0.606478
R16201 Vbias.n3312 Vbias.n3259 0.606478
R16202 Vbias.n3707 Vbias.n3706 0.606478
R16203 Vbias.n3695 Vbias.n3452 0.606478
R16204 Vbias.n3657 Vbias.n3481 0.606478
R16205 Vbias.n3620 Vbias.n3507 0.606478
R16206 Vbias.n3619 Vbias.n3618 0.606478
R16207 Vbias.n3581 Vbias.n3528 0.606478
R16208 Vbias.n4251 Vbias.n4250 0.606478
R16209 Vbias.n4230 Vbias.n4011 0.606478
R16210 Vbias.n4214 Vbias.n4036 0.606478
R16211 Vbias.n4213 Vbias.n4212 0.606478
R16212 Vbias.n4196 Vbias.n4053 0.606478
R16213 Vbias.n4112 Vbias.n4102 0.606478
R16214 Vbias.n4114 Vbias.n4113 0.606478
R16215 Vbias.n4127 Vbias.n4126 0.606478
R16216 Vbias.n4143 Vbias.n4142 0.606478
R16217 Vbias.n4166 Vbias.n4165 0.606478
R16218 Vbias.n3168 Vbias.n3167 0.606478
R16219 Vbias.n3156 Vbias.n2913 0.606478
R16220 Vbias.n3118 Vbias.n2942 0.606478
R16221 Vbias.n3081 Vbias.n2968 0.606478
R16222 Vbias.n3080 Vbias.n3079 0.606478
R16223 Vbias.n3042 Vbias.n2989 0.606478
R16224 Vbias.n2898 Vbias.n2897 0.606478
R16225 Vbias.n4832 Vbias.n2674 0.606478
R16226 Vbias.n4794 Vbias.n2703 0.606478
R16227 Vbias.n4757 Vbias.n2729 0.606478
R16228 Vbias.n4756 Vbias.n4755 0.606478
R16229 Vbias.n4718 Vbias.n2750 0.606478
R16230 Vbias.n4578 Vbias.n4555 0.606478
R16231 Vbias.n4665 Vbias.n4579 0.606478
R16232 Vbias.n4656 Vbias.n4655 0.606478
R16233 Vbias.n4648 Vbias.n4647 0.606478
R16234 Vbias.n5032 Vbias.n5031 0.606478
R16235 Vbias.n7466 Vbias.n7465 0.606478
R16236 Vbias.n7445 Vbias.n7346 0.606478
R16237 Vbias.n7429 Vbias.n7366 0.606478
R16238 Vbias.n7428 Vbias.n7427 0.606478
R16239 Vbias.n7411 Vbias.n7384 0.606478
R16240 Vbias.n6649 Vbias.n6648 0.606478
R16241 Vbias.n6634 Vbias.n6633 0.606478
R16242 Vbias.n6626 Vbias.n6625 0.606478
R16243 Vbias.n6616 Vbias.n6192 0.606478
R16244 Vbias.n6606 Vbias.n6206 0.606478
R16245 Vbias.n6575 Vbias.n6574 0.606478
R16246 Vbias.n6567 Vbias.n6566 0.606478
R16247 Vbias.n6559 Vbias.n6558 0.606478
R16248 Vbias.n6549 Vbias.n6429 0.606478
R16249 Vbias.n6539 Vbias.n6443 0.606478
R16250 Vbias.n7588 Vbias.n7587 0.606478
R16251 Vbias.n7580 Vbias.n7579 0.606478
R16252 Vbias.n7572 Vbias.n7571 0.606478
R16253 Vbias.n7562 Vbias.n883 0.606478
R16254 Vbias.n7552 Vbias.n897 0.606478
R16255 Vbias.n7322 Vbias.n7321 0.606478
R16256 Vbias.n1043 Vbias.n1042 0.606478
R16257 Vbias.n1064 Vbias.n1063 0.606478
R16258 Vbias.n7240 Vbias.n7239 0.606478
R16259 Vbias.n7276 Vbias.n7275 0.606478
R16260 Vbias.n946 Vbias.n945 0.606478
R16261 Vbias.n948 Vbias.n947 0.606478
R16262 Vbias.n969 Vbias.n968 0.606478
R16263 Vbias.n990 Vbias.n989 0.606478
R16264 Vbias.n7482 Vbias.n7481 0.606478
R16265 Vbias.n6362 Vbias.n6361 0.606478
R16266 Vbias.n6360 Vbias.n6359 0.606478
R16267 Vbias.n814 Vbias.n813 0.606478
R16268 Vbias.n835 Vbias.n834 0.606478
R16269 Vbias.n7604 Vbias.n7603 0.606478
R16270 Vbias.n6312 Vbias.n6297 0.606478
R16271 Vbias.n6314 Vbias.n6313 0.606478
R16272 Vbias.n6328 Vbias.n6327 0.606478
R16273 Vbias.n6343 Vbias.n6341 0.606478
R16274 Vbias.n6358 Vbias.n6242 0.606478
R16275 Vbias.n5841 Vbias.n5831 0.606478
R16276 Vbias.n5843 Vbias.n5842 0.606478
R16277 Vbias.n1717 Vbias.n1716 0.606478
R16278 Vbias.n1718 Vbias.n1480 0.606478
R16279 Vbias.n6665 Vbias.n6664 0.606478
R16280 Vbias.n5755 Vbias.n5741 0.606478
R16281 Vbias.n5757 Vbias.n5756 0.606478
R16282 Vbias.n5771 Vbias.n5770 0.606478
R16283 Vbias.n5786 Vbias.n5785 0.606478
R16284 Vbias.n5814 Vbias.n5813 0.606478
R16285 Vbias.n5668 Vbias.n5667 0.606478
R16286 Vbias.n5681 Vbias.n2190 0.606478
R16287 Vbias.n5699 Vbias.n2172 0.606478
R16288 Vbias.n5700 Vbias.n2141 0.606478
R16289 Vbias.n5725 Vbias.n5724 0.606478
R16290 Vbias.n5594 Vbias.n5593 0.606478
R16291 Vbias.n5607 Vbias.n5587 0.606478
R16292 Vbias.n5625 Vbias.n5569 0.606478
R16293 Vbias.n5626 Vbias.n2212 0.606478
R16294 Vbias.n5651 Vbias.n5650 0.606478
R16295 Vbias.n252 Vbias.n251 0.606478
R16296 Vbias.n250 Vbias.n249 0.606478
R16297 Vbias.n123 Vbias.n122 0.606478
R16298 Vbias.n143 Vbias.n142 0.606478
R16299 Vbias.n7960 Vbias.n7959 0.606478
R16300 Vbias.n257 Vbias.n256 0.606478
R16301 Vbias.n274 Vbias.n273 0.606478
R16302 Vbias.n294 Vbias.n292 0.606478
R16303 Vbias.n293 Vbias.n198 0.606478
R16304 Vbias.n313 Vbias.n312 0.606478
R16305 Vbias.n7932 Vbias.n356 0.606478
R16306 Vbias.n7920 Vbias.n380 0.606478
R16307 Vbias.n7908 Vbias.n404 0.606478
R16308 Vbias.n7907 Vbias.n7906 0.606478
R16309 Vbias.n7895 Vbias.n427 0.606478
R16310 Vbias.n7866 Vbias.n462 0.606478
R16311 Vbias.n7854 Vbias.n486 0.606478
R16312 Vbias.n7842 Vbias.n510 0.606478
R16313 Vbias.n7841 Vbias.n7840 0.606478
R16314 Vbias.n7829 Vbias.n533 0.606478
R16315 Vbias.n7797 Vbias.n576 0.606478
R16316 Vbias.n7785 Vbias.n600 0.606478
R16317 Vbias.n7773 Vbias.n624 0.606478
R16318 Vbias.n7772 Vbias.n7771 0.606478
R16319 Vbias.n7760 Vbias.n647 0.606478
R16320 Vbias.n5827 Vbias.n682 0.606478
R16321 Vbias.n7720 Vbias.n7719 0.606478
R16322 Vbias.n7705 Vbias.n7704 0.606478
R16323 Vbias.n7695 Vbias.n730 0.606478
R16324 Vbias.n7680 Vbias.n739 0.606478
R16325 Vbias.n6127 Vbias.n6126 0.606478
R16326 Vbias.n7660 Vbias.n7659 0.606478
R16327 Vbias.n6511 Vbias.n771 0.606478
R16328 Vbias.n6513 Vbias.n6512 0.606478
R16329 Vbias.n7536 Vbias.n7535 0.606478
R16330 Vbias.n7539 Vbias.n7538 0.606478
R16331 Vbias.n7942 Vbias.n169 0.606478
R16332 Vbias.n7881 Vbias.n452 0.606478
R16333 Vbias.n7816 Vbias.n7815 0.606478
R16334 Vbias.n672 Vbias.n558 0.606478
R16335 Vbias.n7746 Vbias.n673 0.606478
R16336 Vbias.n2585 Vbias.n2584 0.606478
R16337 Vbias.n5548 Vbias.n5547 0.606478
R16338 Vbias.n5513 Vbias.n2233 0.606478
R16339 Vbias.n5527 Vbias.n5514 0.606478
R16340 Vbias.n5872 Vbias.n5871 0.606478
R16341 Vbias.n1680 Vbias.n1679 0.606478
R16342 Vbias.n6692 Vbias.n6691 0.606478
R16343 Vbias.n6745 Vbias.n6744 0.606478
R16344 Vbias.n6718 Vbias.n6717 0.606478
R16345 Vbias.n6694 Vbias.n6693 0.606478
R16346 Vbias.n4988 Vbias.n4987 0.606478
R16347 Vbias.n5005 Vbias.n5004 0.606478
R16348 Vbias.n2895 Vbias.n2894 0.606478
R16349 Vbias.n4920 Vbias.n2657 0.606478
R16350 Vbias.n4942 Vbias.n2643 0.606478
R16351 Vbias.n4943 Vbias.n2618 0.606478
R16352 Vbias.n4970 Vbias.n4969 0.606478
R16353 Vbias.n3171 Vbias.n13 0.606478
R16354 Vbias.n8060 Vbias.n8059 0.606478
R16355 Vbias.n8045 Vbias.n8044 0.606478
R16356 Vbias.n8035 Vbias.n61 0.606478
R16357 Vbias.n8020 Vbias.n70 0.606478
R16358 Vbias.n1734 Vbias.n1507 0.601043
R16359 Vbias.n1843 Vbias 0.590136
R16360 Vbias.n1838 Vbias 0.590136
R16361 Vbias.n1833 Vbias 0.590136
R16362 Vbias.n1828 Vbias 0.590136
R16363 Vbias.n1823 Vbias 0.590136
R16364 Vbias.n2020 Vbias 0.590136
R16365 Vbias.n2025 Vbias 0.590136
R16366 Vbias.n2029 Vbias 0.590136
R16367 Vbias.n2028 Vbias.n2027 0.547267
R16368 Vbias.n4255 Vbias.n4254 0.495065
R16369 Vbias.n3977 Vbias.n3976 0.495065
R16370 Vbias.n3439 Vbias.n3438 0.495065
R16371 Vbias.n3708 Vbias.n3707 0.495065
R16372 Vbias.n4102 Vbias.n4101 0.495065
R16373 Vbias.n3169 Vbias.n3168 0.495065
R16374 Vbias.n2899 Vbias.n2898 0.495065
R16375 Vbias.n7323 Vbias.n7322 0.495065
R16376 Vbias.n945 Vbias.n858 0.495065
R16377 Vbias.n6363 Vbias.n6362 0.495065
R16378 Vbias.n6297 Vbias.n6133 0.495065
R16379 Vbias.n5831 Vbias.n5830 0.495065
R16380 Vbias.n5741 Vbias.n5740 0.495065
R16381 Vbias.n5667 Vbias.n5666 0.495065
R16382 Vbias.n5593 Vbias.n5592 0.495065
R16383 Vbias.n253 Vbias.n252 0.495065
R16384 Vbias.n2896 Vbias.n2895 0.495065
R16385 Vbias.n7943 Vbias.n7942 0.476043
R16386 Vbias.n1840 Vbias.n1839 0.419583
R16387 Vbias.n1835 Vbias.n1834 0.419583
R16388 Vbias.n1830 Vbias.n1829 0.419583
R16389 Vbias.n1825 Vbias.n1824 0.419583
R16390 Vbias.n2019 Vbias.n2018 0.419583
R16391 Vbias.n2024 Vbias.n2023 0.419583
R16392 Vbias.n4267 Vbias 0.405391
R16393 Vbias.n4300 Vbias 0.405391
R16394 Vbias.n4333 Vbias 0.405391
R16395 Vbias Vbias.n2809 0.405391
R16396 Vbias Vbias.n2796 0.405391
R16397 Vbias.n5052 Vbias 0.405391
R16398 Vbias Vbias.n5073 0.405391
R16399 Vbias.n5074 Vbias 0.405391
R16400 Vbias.n5095 Vbias 0.405391
R16401 Vbias.n5115 Vbias 0.405391
R16402 Vbias.n5175 Vbias 0.405391
R16403 Vbias Vbias.n5161 0.405391
R16404 Vbias.n5162 Vbias 0.405391
R16405 Vbias Vbias.n2253 0.405391
R16406 Vbias Vbias.n2293 0.405391
R16407 Vbias Vbias.n5440 0.405391
R16408 Vbias Vbias.n5441 0.405391
R16409 Vbias.n5457 Vbias 0.405391
R16410 Vbias.n5892 Vbias 0.405391
R16411 Vbias.n5912 Vbias 0.405391
R16412 Vbias.n5948 Vbias 0.405391
R16413 Vbias.n1620 Vbias 0.405391
R16414 Vbias.n6095 Vbias 0.405391
R16415 Vbias.n6087 Vbias 0.405391
R16416 Vbias.n6079 Vbias 0.405391
R16417 Vbias.n6806 Vbias 0.405391
R16418 Vbias Vbias.n1420 0.405391
R16419 Vbias.n6793 Vbias 0.405391
R16420 Vbias.n6785 Vbias 0.405391
R16421 Vbias.n7009 Vbias 0.405391
R16422 Vbias.n7031 Vbias 0.405391
R16423 Vbias.n7048 Vbias 0.405391
R16424 Vbias Vbias.n7061 0.405391
R16425 Vbias Vbias.n7078 0.405391
R16426 Vbias Vbias.n7095 0.405391
R16427 Vbias.n7137 Vbias 0.405391
R16428 Vbias.n7154 Vbias 0.405391
R16429 Vbias Vbias.n7167 0.405391
R16430 Vbias Vbias.n7184 0.405391
R16431 Vbias Vbias.n7201 0.405391
R16432 Vbias Vbias.n1194 0.405391
R16433 Vbias.n1243 Vbias 0.405391
R16434 Vbias.n1211 Vbias 0.405391
R16435 Vbias.n7205 Vbias 0.405391
R16436 Vbias.n7203 Vbias 0.405391
R16437 Vbias Vbias.n6927 0.405391
R16438 Vbias.n6976 Vbias 0.405391
R16439 Vbias.n6944 Vbias 0.405391
R16440 Vbias.n7101 Vbias 0.405391
R16441 Vbias.n7099 Vbias 0.405391
R16442 Vbias Vbias.n6833 0.405391
R16443 Vbias.n6834 Vbias 0.405391
R16444 Vbias.n6857 Vbias 0.405391
R16445 Vbias.n6880 Vbias 0.405391
R16446 Vbias Vbias.n6899 0.405391
R16447 Vbias Vbias.n5975 0.405391
R16448 Vbias.n5976 Vbias 0.405391
R16449 Vbias.n5999 Vbias 0.405391
R16450 Vbias.n6025 Vbias 0.405391
R16451 Vbias.n6023 Vbias 0.405391
R16452 Vbias Vbias.n5298 0.405391
R16453 Vbias.n5384 Vbias 0.405391
R16454 Vbias Vbias.n5333 0.405391
R16455 Vbias Vbias.n5335 0.405391
R16456 Vbias.n5341 Vbias 0.405391
R16457 Vbias Vbias.n5202 0.405391
R16458 Vbias.n5203 Vbias 0.405391
R16459 Vbias.n5226 Vbias 0.405391
R16460 Vbias.n5249 Vbias 0.405391
R16461 Vbias Vbias.n5269 0.405391
R16462 Vbias Vbias.n2466 0.405391
R16463 Vbias.n2552 Vbias 0.405391
R16464 Vbias Vbias.n2501 0.405391
R16465 Vbias Vbias.n2503 0.405391
R16466 Vbias.n2509 Vbias 0.405391
R16467 Vbias Vbias.n4423 0.405391
R16468 Vbias.n4524 Vbias 0.405391
R16469 Vbias.n4510 Vbias 0.405391
R16470 Vbias.n4496 Vbias 0.405391
R16471 Vbias.n4484 Vbias 0.405391
R16472 Vbias.n3721 Vbias 0.405391
R16473 Vbias.n3750 Vbias 0.405391
R16474 Vbias.n3776 Vbias 0.405391
R16475 Vbias Vbias.n3888 0.405391
R16476 Vbias.n3797 Vbias 0.405391
R16477 Vbias.n3183 Vbias 0.405391
R16478 Vbias.n3212 Vbias 0.405391
R16479 Vbias.n3238 Vbias 0.405391
R16480 Vbias Vbias.n3350 0.405391
R16481 Vbias.n3259 Vbias 0.405391
R16482 Vbias.n3452 Vbias 0.405391
R16483 Vbias.n3481 Vbias 0.405391
R16484 Vbias.n3507 Vbias 0.405391
R16485 Vbias Vbias.n3619 0.405391
R16486 Vbias.n3528 Vbias 0.405391
R16487 Vbias.n4011 Vbias 0.405391
R16488 Vbias.n4036 Vbias 0.405391
R16489 Vbias Vbias.n4213 0.405391
R16490 Vbias.n4053 Vbias 0.405391
R16491 Vbias.n4113 Vbias 0.405391
R16492 Vbias.n4126 Vbias 0.405391
R16493 Vbias.n4165 Vbias 0.405391
R16494 Vbias.n2913 Vbias 0.405391
R16495 Vbias.n2942 Vbias 0.405391
R16496 Vbias.n2968 Vbias 0.405391
R16497 Vbias Vbias.n3080 0.405391
R16498 Vbias.n2989 Vbias 0.405391
R16499 Vbias Vbias.n2674 0.405391
R16500 Vbias.n2703 Vbias 0.405391
R16501 Vbias.n2729 Vbias 0.405391
R16502 Vbias Vbias.n4756 0.405391
R16503 Vbias.n2750 Vbias 0.405391
R16504 Vbias Vbias.n4578 0.405391
R16505 Vbias Vbias.n4579 0.405391
R16506 Vbias.n4655 Vbias 0.405391
R16507 Vbias.n4647 Vbias 0.405391
R16508 Vbias.n5031 Vbias 0.405391
R16509 Vbias.n7346 Vbias 0.405391
R16510 Vbias.n7366 Vbias 0.405391
R16511 Vbias Vbias.n7428 0.405391
R16512 Vbias.n7384 Vbias 0.405391
R16513 Vbias Vbias.n6634 0.405391
R16514 Vbias Vbias.n6626 0.405391
R16515 Vbias.n6192 Vbias 0.405391
R16516 Vbias.n6206 Vbias 0.405391
R16517 Vbias Vbias.n6567 0.405391
R16518 Vbias Vbias.n6559 0.405391
R16519 Vbias.n6429 Vbias 0.405391
R16520 Vbias.n6443 Vbias 0.405391
R16521 Vbias Vbias.n7580 0.405391
R16522 Vbias Vbias.n7572 0.405391
R16523 Vbias.n883 Vbias 0.405391
R16524 Vbias.n897 Vbias 0.405391
R16525 Vbias.n1042 Vbias 0.405391
R16526 Vbias.n1063 Vbias 0.405391
R16527 Vbias Vbias.n7276 0.405391
R16528 Vbias.n947 Vbias 0.405391
R16529 Vbias.n968 Vbias 0.405391
R16530 Vbias Vbias.n7482 0.405391
R16531 Vbias Vbias.n6360 0.405391
R16532 Vbias.n813 Vbias 0.405391
R16533 Vbias Vbias.n7604 0.405391
R16534 Vbias.n6313 Vbias 0.405391
R16535 Vbias.n6327 Vbias 0.405391
R16536 Vbias Vbias.n6242 0.405391
R16537 Vbias.n5842 Vbias 0.405391
R16538 Vbias.n1716 Vbias 0.405391
R16539 Vbias Vbias.n6665 0.405391
R16540 Vbias.n5756 Vbias 0.405391
R16541 Vbias.n5770 Vbias 0.405391
R16542 Vbias.n5813 Vbias 0.405391
R16543 Vbias Vbias.n2190 0.405391
R16544 Vbias Vbias.n2172 0.405391
R16545 Vbias.n5724 Vbias 0.405391
R16546 Vbias Vbias.n5587 0.405391
R16547 Vbias Vbias.n5569 0.405391
R16548 Vbias.n5650 Vbias 0.405391
R16549 Vbias Vbias.n250 0.405391
R16550 Vbias.n122 Vbias 0.405391
R16551 Vbias Vbias.n7960 0.405391
R16552 Vbias.n273 Vbias 0.405391
R16553 Vbias.n292 Vbias 0.405391
R16554 Vbias Vbias.n293 0.405391
R16555 Vbias.n312 Vbias 0.405391
R16556 Vbias.n380 Vbias 0.405391
R16557 Vbias.n404 Vbias 0.405391
R16558 Vbias Vbias.n7907 0.405391
R16559 Vbias.n427 Vbias 0.405391
R16560 Vbias.n486 Vbias 0.405391
R16561 Vbias.n510 Vbias 0.405391
R16562 Vbias Vbias.n7841 0.405391
R16563 Vbias.n533 Vbias 0.405391
R16564 Vbias.n600 Vbias 0.405391
R16565 Vbias.n624 Vbias 0.405391
R16566 Vbias Vbias.n7772 0.405391
R16567 Vbias.n647 Vbias 0.405391
R16568 Vbias Vbias.n7720 0.405391
R16569 Vbias Vbias.n7705 0.405391
R16570 Vbias.n730 Vbias 0.405391
R16571 Vbias.n739 Vbias 0.405391
R16572 Vbias.n6126 Vbias 0.405391
R16573 Vbias.n7659 Vbias 0.405391
R16574 Vbias Vbias.n6511 0.405391
R16575 Vbias.n6512 Vbias 0.405391
R16576 Vbias Vbias.n7536 0.405391
R16577 Vbias.n7538 Vbias 0.405391
R16578 Vbias Vbias.n169 0.405391
R16579 Vbias Vbias.n452 0.405391
R16580 Vbias.n7815 Vbias 0.405391
R16581 Vbias Vbias.n672 0.405391
R16582 Vbias Vbias.n673 0.405391
R16583 Vbias Vbias.n327 0.405391
R16584 Vbias.n2584 Vbias 0.405391
R16585 Vbias.n5547 Vbias 0.405391
R16586 Vbias Vbias.n5513 0.405391
R16587 Vbias.n5514 Vbias 0.405391
R16588 Vbias.n5871 Vbias 0.405391
R16589 Vbias.n1679 Vbias 0.405391
R16590 Vbias Vbias.n6692 0.405391
R16591 Vbias.n6744 Vbias 0.405391
R16592 Vbias.n6717 Vbias 0.405391
R16593 Vbias.n6693 Vbias 0.405391
R16594 Vbias.n4987 Vbias 0.405391
R16595 Vbias.n5004 Vbias 0.405391
R16596 Vbias Vbias.n2657 0.405391
R16597 Vbias Vbias.n2643 0.405391
R16598 Vbias.n4969 Vbias 0.405391
R16599 Vbias Vbias.n8060 0.405391
R16600 Vbias Vbias.n8045 0.405391
R16601 Vbias.n61 Vbias 0.405391
R16602 Vbias.n70 Vbias 0.405391
R16603 Vbias.n1747 Vbias.n1746 0.353761
R16604 Vbias.n8087 Vbias.n0 0.340174
R16605 Vbias.n6123 Vbias 0.149957
R16606 Vbias Vbias.n7202 0.0901739
R16607 Vbias Vbias.n7098 0.0901739
R16608 Vbias.n6900 Vbias 0.0901739
R16609 Vbias Vbias.n6022 0.0901739
R16610 Vbias Vbias.n5340 0.0901739
R16611 Vbias.n5270 Vbias 0.0901739
R16612 Vbias Vbias.n2508 0.0901739
R16613 Vbias Vbias.n4483 0.0901739
R16614 Vbias.n6122 Vbias.n1508 0.063
R16615 Vbias.n6109 Vbias.n1508 0.063
R16616 Vbias.n2017 Vbias.n1984 0.063
R16617 Vbias.n2017 Vbias.n2016 0.063
R16618 Vbias.n1982 Vbias.n1749 0.063
R16619 Vbias.n1969 Vbias.n1749 0.063
R16620 Vbias.n1948 Vbias.n1750 0.063
R16621 Vbias.n1935 Vbias.n1750 0.063
R16622 Vbias.n1914 Vbias.n1751 0.063
R16623 Vbias.n1898 Vbias.n1751 0.063
R16624 Vbias.n1880 Vbias.n1752 0.063
R16625 Vbias.n1869 Vbias.n1752 0.063
R16626 Vbias.n1846 Vbias.n1845 0.063
R16627 Vbias.n1845 Vbias.n1821 0.063
R16628 Vbias.n2032 Vbias.n1747 0.063
R16629 Vbias.n2033 Vbias.n2032 0.063
R16630 Vbias.n6124 Vbias.n6123 0.063
R16631 Vbias.n7468 Vbias.n7323 0.063
R16632 Vbias.n7590 Vbias.n858 0.063
R16633 Vbias.n6577 Vbias.n6363 0.063
R16634 Vbias.n6651 Vbias.n6133 0.063
R16635 Vbias.n5830 Vbias.n5829 0.063
R16636 Vbias.n5740 Vbias.n5739 0.063
R16637 Vbias.n5666 Vbias.n5665 0.063
R16638 Vbias.n5592 Vbias.n166 0.063
R16639 Vbias.n7944 Vbias.n168 0.063
R16640 Vbias.n7944 Vbias.n7943 0.063
R16641 Vbias Vbias.n8087 0.0512812
R16642 Vbias.t702 Vbias.n4892 0.047916
R16643 Vbias.n6124 Vbias 0.0454219
R16644 Vbias Vbias.n7097 0.0454219
R16645 Vbias.n7007 Vbias 0.0454219
R16646 Vbias.n6815 Vbias 0.0454219
R16647 Vbias.n5957 Vbias 0.0454219
R16648 Vbias.n5415 Vbias 0.0454219
R16649 Vbias.n5184 Vbias 0.0454219
R16650 Vbias Vbias.n2583 0.0454219
R16651 Vbias.n7202 Vbias 0.0249565
R16652 Vbias.n7098 Vbias 0.0249565
R16653 Vbias.n6900 Vbias 0.0249565
R16654 Vbias.n6022 Vbias 0.0249565
R16655 Vbias.n5340 Vbias 0.0249565
R16656 Vbias.n5270 Vbias 0.0249565
R16657 Vbias.n2508 Vbias 0.0249565
R16658 Vbias.n4483 Vbias 0.0249565
R16659 Vbias.n1844 Vbias.n1843 0.024
R16660 Vbias.n1839 Vbias.n1838 0.024
R16661 Vbias.n1834 Vbias.n1833 0.024
R16662 Vbias.n1829 Vbias.n1828 0.024
R16663 Vbias.n1824 Vbias.n1823 0.024
R16664 Vbias.n2020 Vbias.n2019 0.024
R16665 Vbias.n2025 Vbias.n2024 0.024
R16666 Vbias.n2029 Vbias.n2028 0.024
R16667 Vbias Vbias.n1841 0.0204394
R16668 Vbias Vbias.n1836 0.0204394
R16669 Vbias Vbias.n1831 0.0204394
R16670 Vbias Vbias.n1826 0.0204394
R16671 Vbias Vbias.n1748 0.0204394
R16672 Vbias.n2022 Vbias 0.0204394
R16673 Vbias.n2027 Vbias 0.0204394
R16674 Vbias.n2031 Vbias 0.0204394
R16675 Vbias.n7202 Vbias 0.0180781
R16676 Vbias.n7098 Vbias 0.0180781
R16677 Vbias Vbias.n6900 0.0180781
R16678 Vbias.n6022 Vbias 0.0180781
R16679 Vbias.n5340 Vbias 0.0180781
R16680 Vbias Vbias.n5270 0.0180781
R16681 Vbias.n2508 Vbias 0.0180781
R16682 Vbias.n4483 Vbias 0.0180781
R16683 Vbias.n1842 Vbias 0.00441667
R16684 Vbias.n1837 Vbias 0.00441667
R16685 Vbias.n1832 Vbias 0.00441667
R16686 Vbias.n1827 Vbias 0.00441667
R16687 Vbias.n1822 Vbias 0.00441667
R16688 Vbias.n2021 Vbias 0.00441667
R16689 Vbias.n2026 Vbias 0.00441667
R16690 Vbias.n2030 Vbias 0.00441667
R16691 Vbias.n255 GND 0.00441667
R16692 Vbias.n1842 Vbias 0.00406061
R16693 Vbias.n1837 Vbias 0.00406061
R16694 Vbias.n1832 Vbias 0.00406061
R16695 Vbias.n1827 Vbias 0.00406061
R16696 Vbias.n1822 Vbias 0.00406061
R16697 Vbias Vbias.n2021 0.00406061
R16698 Vbias Vbias.n2026 0.00406061
R16699 Vbias Vbias.n2030 0.00406061
R16700 GND Vbias.n255 0.00406061
R16701 Vbias.n1880 Vbias.n1847 0.00287997
R16702 Vbias Vbias.n1880 0.00287997
R16703 Vbias Vbias.n1846 0.00287997
R16704 Vbias.n6122 Vbias.n1509 0.00287997
R16705 Vbias Vbias.n6122 0.00287997
R16706 Vbias.n1984 Vbias.n1983 0.00287997
R16707 Vbias.n1984 Vbias 0.00287997
R16708 Vbias.n1982 Vbias.n1949 0.00287997
R16709 Vbias Vbias.n1982 0.00287997
R16710 Vbias.n1948 Vbias.n1915 0.00287997
R16711 Vbias Vbias.n1948 0.00287997
R16712 Vbias.n1914 Vbias.n1881 0.00287997
R16713 Vbias Vbias.n1914 0.00287997
R16714 CLK.n244 CLK.t23 158.207
R16715 CLK.n231 CLK.t8 158.207
R16716 CLK.n218 CLK.t59 158.207
R16717 CLK.n205 CLK.t2 158.207
R16718 CLK.n192 CLK.t93 158.207
R16719 CLK.n179 CLK.t22 158.207
R16720 CLK.n166 CLK.t5 158.207
R16721 CLK.n154 CLK.t102 158.207
R16722 CLK.n104 CLK.t13 158.207
R16723 CLK.n91 CLK.t80 158.207
R16724 CLK.n78 CLK.t51 158.207
R16725 CLK.n65 CLK.t114 158.207
R16726 CLK.n52 CLK.t84 158.207
R16727 CLK.n39 CLK.t54 158.207
R16728 CLK.n27 CLK.t117 158.207
R16729 CLK.n15 CLK.t27 158.207
R16730 CLK.n3 CLK.t95 158.207
R16731 CLK CLK.t100 158.202
R16732 CLK CLK.t72 158.202
R16733 CLK CLK.t15 158.202
R16734 CLK CLK.t62 158.202
R16735 CLK CLK.t37 158.202
R16736 CLK CLK.t97 158.202
R16737 CLK CLK.t69 158.202
R16738 CLK CLK.t45 158.202
R16739 CLK CLK.t83 158.202
R16740 CLK CLK.t30 158.202
R16741 CLK CLK.t16 158.202
R16742 CLK CLK.t63 158.202
R16743 CLK CLK.t38 158.202
R16744 CLK CLK.t19 158.202
R16745 CLK CLK.t70 158.202
R16746 CLK CLK.t113 158.202
R16747 CLK CLK.t42 158.202
R16748 CLK.n246 CLK.t39 150.293
R16749 CLK.t100 CLK.n249 150.293
R16750 CLK.n233 CLK.t26 150.293
R16751 CLK.t72 CLK.n236 150.293
R16752 CLK.n220 CLK.t108 150.293
R16753 CLK.t15 CLK.n223 150.293
R16754 CLK.n207 CLK.t75 150.293
R16755 CLK.t62 CLK.n210 150.293
R16756 CLK.n194 CLK.t47 150.293
R16757 CLK.t37 CLK.n197 150.293
R16758 CLK.n181 CLK.t111 150.293
R16759 CLK.t97 CLK.n184 150.293
R16760 CLK.n168 CLK.t78 150.293
R16761 CLK.t69 CLK.n171 150.293
R16762 CLK.n156 CLK.t17 150.293
R16763 CLK.t45 CLK.n159 150.293
R16764 CLK.n128 CLK.t44 150.293
R16765 CLK.n131 CLK.t87 150.293
R16766 CLK.n134 CLK.t34 150.293
R16767 CLK.n125 CLK.t18 150.293
R16768 CLK.n106 CLK.t31 150.293
R16769 CLK.t83 CLK.n109 150.293
R16770 CLK.n93 CLK.t52 150.293
R16771 CLK.t30 CLK.n96 150.293
R16772 CLK.n80 CLK.t25 150.293
R16773 CLK.t16 CLK.n83 150.293
R16774 CLK.n67 CLK.t11 150.293
R16775 CLK.t63 CLK.n70 150.293
R16776 CLK.n54 CLK.t55 150.293
R16777 CLK.t38 CLK.n57 150.293
R16778 CLK.n41 CLK.t28 150.293
R16779 CLK.t19 CLK.n44 150.293
R16780 CLK.n29 CLK.t88 150.293
R16781 CLK.t70 CLK.n32 150.293
R16782 CLK.n17 CLK.t57 150.293
R16783 CLK.t113 CLK.n20 150.293
R16784 CLK.n5 CLK.t33 150.293
R16785 CLK.t42 CLK.n8 150.293
R16786 CLK.t23 CLK.n243 150.273
R16787 CLK.t8 CLK.n230 150.273
R16788 CLK.t59 CLK.n217 150.273
R16789 CLK.t2 CLK.n204 150.273
R16790 CLK.t93 CLK.n191 150.273
R16791 CLK.t22 CLK.n178 150.273
R16792 CLK.t5 CLK.n165 150.273
R16793 CLK.t102 CLK.n153 150.273
R16794 CLK.n123 CLK.t105 150.273
R16795 CLK.n119 CLK.t77 150.273
R16796 CLK.n141 CLK.t74 150.273
R16797 CLK.n146 CLK.t110 150.273
R16798 CLK.t13 CLK.n103 150.273
R16799 CLK.t80 CLK.n90 150.273
R16800 CLK.t51 CLK.n77 150.273
R16801 CLK.t114 CLK.n64 150.273
R16802 CLK.t84 CLK.n51 150.273
R16803 CLK.t54 CLK.n38 150.273
R16804 CLK.t117 CLK.n26 150.273
R16805 CLK.t27 CLK.n14 150.273
R16806 CLK.t95 CLK.n2 150.273
R16807 CLK.n241 CLK.t40 73.6406
R16808 CLK.n228 CLK.t98 73.6406
R16809 CLK.n215 CLK.t29 73.6406
R16810 CLK.n202 CLK.t89 73.6406
R16811 CLK.n189 CLK.t60 73.6406
R16812 CLK.n176 CLK.t35 73.6406
R16813 CLK.n163 CLK.t96 73.6406
R16814 CLK.n151 CLK.t68 73.6406
R16815 CLK.n101 CLK.t20 73.6406
R16816 CLK.n88 CLK.t91 73.6406
R16817 CLK.n75 CLK.t65 73.6406
R16818 CLK.n62 CLK.t41 73.6406
R16819 CLK.n49 CLK.t99 73.6406
R16820 CLK.n36 CLK.t71 73.6406
R16821 CLK.n24 CLK.t9 73.6406
R16822 CLK.n12 CLK.t46 73.6406
R16823 CLK.n0 CLK.t64 73.6406
R16824 CLK.n248 CLK.t58 73.6304
R16825 CLK.n247 CLK.t107 73.6304
R16826 CLK.n235 CLK.t1 73.6304
R16827 CLK.n234 CLK.t94 73.6304
R16828 CLK.n222 CLK.t53 73.6304
R16829 CLK.n221 CLK.t67 73.6304
R16830 CLK.n209 CLK.t116 73.6304
R16831 CLK.n208 CLK.t6 73.6304
R16832 CLK.n196 CLK.t85 73.6304
R16833 CLK.n195 CLK.t103 73.6304
R16834 CLK.n183 CLK.t56 73.6304
R16835 CLK.n182 CLK.t24 73.6304
R16836 CLK.n170 CLK.t0 73.6304
R16837 CLK.n169 CLK.t10 73.6304
R16838 CLK.n158 CLK.t90 73.6304
R16839 CLK.n157 CLK.t106 73.6304
R16840 CLK.n129 CLK.t81 73.6304
R16841 CLK.n132 CLK.t48 73.6304
R16842 CLK.n120 CLK.t21 73.6304
R16843 CLK.n116 CLK.t3 73.6304
R16844 CLK.n138 CLK.t115 73.6304
R16845 CLK.n143 CLK.t61 73.6304
R16846 CLK.n135 CLK.t43 73.6304
R16847 CLK.n126 CLK.t49 73.6304
R16848 CLK.n108 CLK.t50 73.6304
R16849 CLK.n107 CLK.t104 73.6304
R16850 CLK.n95 CLK.t12 73.6304
R16851 CLK.n94 CLK.t32 73.6304
R16852 CLK.n82 CLK.t109 73.6304
R16853 CLK.n81 CLK.t92 73.6304
R16854 CLK.n69 CLK.t76 73.6304
R16855 CLK.n68 CLK.t66 73.6304
R16856 CLK.n56 CLK.t14 73.6304
R16857 CLK.n55 CLK.t4 73.6304
R16858 CLK.n43 CLK.t112 73.6304
R16859 CLK.n42 CLK.t101 73.6304
R16860 CLK.n31 CLK.t36 73.6304
R16861 CLK.n30 CLK.t73 73.6304
R16862 CLK.n19 CLK.t79 73.6304
R16863 CLK.n18 CLK.t7 73.6304
R16864 CLK.n7 CLK.t86 73.6304
R16865 CLK.n6 CLK.t82 73.6304
R16866 CLK.n124 CLK.n119 64.4516
R16867 CLK.n147 CLK.n142 59.9516
R16868 CLK.n133 CLK.n130 59.9516
R16869 CLK.n136 CLK.n135 54.8429
R16870 CLK.n142 CLK.n137 37.8646
R16871 CLK.n127 CLK.n126 34.5521
R16872 CLK.n137 CLK.n136 30.474
R16873 CLK.n130 CLK.n127 29.8239
R16874 CLK.n148 CLK.n115 23.654
R16875 CLK.n137 CLK.n124 22.0114
R16876 CLK.n248 CLK.n247 16.332
R16877 CLK.n235 CLK.n234 16.332
R16878 CLK.n222 CLK.n221 16.332
R16879 CLK.n209 CLK.n208 16.332
R16880 CLK.n196 CLK.n195 16.332
R16881 CLK.n183 CLK.n182 16.332
R16882 CLK.n170 CLK.n169 16.332
R16883 CLK.n158 CLK.n157 16.332
R16884 CLK.n108 CLK.n107 16.332
R16885 CLK.n95 CLK.n94 16.332
R16886 CLK.n82 CLK.n81 16.332
R16887 CLK.n69 CLK.n68 16.332
R16888 CLK.n56 CLK.n55 16.332
R16889 CLK.n43 CLK.n42 16.332
R16890 CLK.n31 CLK.n30 16.332
R16891 CLK.n19 CLK.n18 16.332
R16892 CLK.n7 CLK.n6 16.332
R16893 CLK.n175 CLK.n162 12.0538
R16894 CLK.n48 CLK.n35 12.0538
R16895 CLK.n136 CLK.n133 9.53311
R16896 CLK.n149 CLK.n11 9.40927
R16897 CLK.n188 CLK.n175 8.6438
R16898 CLK.n201 CLK.n188 8.6438
R16899 CLK.n214 CLK.n201 8.6438
R16900 CLK.n227 CLK.n214 8.6438
R16901 CLK.n240 CLK.n227 8.6438
R16902 CLK.n253 CLK.n240 8.6438
R16903 CLK.n61 CLK.n48 8.6438
R16904 CLK.n74 CLK.n61 8.6438
R16905 CLK.n87 CLK.n74 8.6438
R16906 CLK.n100 CLK.n87 8.6438
R16907 CLK.n113 CLK.n100 8.6438
R16908 CLK.n114 CLK.n23 6.21797
R16909 CLK.n115 CLK.n114 6.0284
R16910 CLK.n149 CLK.n148 5.92422
R16911 CLK.n114 CLK.n113 5.83163
R16912 CLK.n148 CLK.n147 4.90235
R16913 CLK.n124 CLK.n123 4.5005
R16914 CLK.n147 CLK.n146 4.5005
R16915 CLK.n142 CLK.n141 4.5005
R16916 CLK.n133 CLK.n132 4.5005
R16917 CLK.n130 CLK.n129 4.5005
R16918 CLK.n175 CLK.n174 3.4105
R16919 CLK.n188 CLK.n187 3.4105
R16920 CLK.n201 CLK.n200 3.4105
R16921 CLK.n214 CLK.n213 3.4105
R16922 CLK.n227 CLK.n226 3.4105
R16923 CLK.n240 CLK.n239 3.4105
R16924 CLK.n48 CLK.n47 3.4105
R16925 CLK.n61 CLK.n60 3.4105
R16926 CLK.n74 CLK.n73 3.4105
R16927 CLK.n87 CLK.n86 3.4105
R16928 CLK.n100 CLK.n99 3.4105
R16929 CLK.n113 CLK.n112 3.4105
R16930 CLK.n127 CLK.n115 3.4105
R16931 CLK.n253 CLK.n252 3.4105
R16932 CLK.n254 CLK.n150 2.59333
R16933 CLK.n150 CLK 2.35833
R16934 CLK.n242 CLK.n241 1.19615
R16935 CLK.n229 CLK.n228 1.19615
R16936 CLK.n216 CLK.n215 1.19615
R16937 CLK.n203 CLK.n202 1.19615
R16938 CLK.n190 CLK.n189 1.19615
R16939 CLK.n177 CLK.n176 1.19615
R16940 CLK.n164 CLK.n163 1.19615
R16941 CLK.n152 CLK.n151 1.19615
R16942 CLK.n102 CLK.n101 1.19615
R16943 CLK.n89 CLK.n88 1.19615
R16944 CLK.n76 CLK.n75 1.19615
R16945 CLK.n63 CLK.n62 1.19615
R16946 CLK.n50 CLK.n49 1.19615
R16947 CLK.n37 CLK.n36 1.19615
R16948 CLK.n25 CLK.n24 1.19615
R16949 CLK.n13 CLK.n12 1.19615
R16950 CLK.n1 CLK.n0 1.19615
R16951 CLK.n247 CLK.n246 1.1717
R16952 CLK.n249 CLK.n248 1.1717
R16953 CLK.n234 CLK.n233 1.1717
R16954 CLK.n236 CLK.n235 1.1717
R16955 CLK.n221 CLK.n220 1.1717
R16956 CLK.n223 CLK.n222 1.1717
R16957 CLK.n208 CLK.n207 1.1717
R16958 CLK.n210 CLK.n209 1.1717
R16959 CLK.n195 CLK.n194 1.1717
R16960 CLK.n197 CLK.n196 1.1717
R16961 CLK.n182 CLK.n181 1.1717
R16962 CLK.n184 CLK.n183 1.1717
R16963 CLK.n169 CLK.n168 1.1717
R16964 CLK.n171 CLK.n170 1.1717
R16965 CLK.n157 CLK.n156 1.1717
R16966 CLK.n159 CLK.n158 1.1717
R16967 CLK.n129 CLK.n128 1.1717
R16968 CLK.n132 CLK.n131 1.1717
R16969 CLK.n122 CLK.n121 1.1717
R16970 CLK.n118 CLK.n117 1.1717
R16971 CLK.n140 CLK.n139 1.1717
R16972 CLK.n145 CLK.n144 1.1717
R16973 CLK.n135 CLK.n134 1.1717
R16974 CLK.n126 CLK.n125 1.1717
R16975 CLK.n107 CLK.n106 1.1717
R16976 CLK.n109 CLK.n108 1.1717
R16977 CLK.n94 CLK.n93 1.1717
R16978 CLK.n96 CLK.n95 1.1717
R16979 CLK.n81 CLK.n80 1.1717
R16980 CLK.n83 CLK.n82 1.1717
R16981 CLK.n68 CLK.n67 1.1717
R16982 CLK.n70 CLK.n69 1.1717
R16983 CLK.n55 CLK.n54 1.1717
R16984 CLK.n57 CLK.n56 1.1717
R16985 CLK.n42 CLK.n41 1.1717
R16986 CLK.n44 CLK.n43 1.1717
R16987 CLK.n30 CLK.n29 1.1717
R16988 CLK.n32 CLK.n31 1.1717
R16989 CLK.n18 CLK.n17 1.1717
R16990 CLK.n20 CLK.n19 1.1717
R16991 CLK.n6 CLK.n5 1.1717
R16992 CLK.n8 CLK.n7 1.1717
R16993 CLK.n122 CLK 0.932141
R16994 CLK.n118 CLK 0.932141
R16995 CLK.n140 CLK 0.932141
R16996 CLK.n145 CLK 0.932141
R16997 CLK.n249 CLK 0.447191
R16998 CLK.n236 CLK 0.447191
R16999 CLK.n223 CLK 0.447191
R17000 CLK.n210 CLK 0.447191
R17001 CLK.n197 CLK 0.447191
R17002 CLK.n184 CLK 0.447191
R17003 CLK.n171 CLK 0.447191
R17004 CLK.n159 CLK 0.447191
R17005 CLK.n128 CLK 0.447191
R17006 CLK.n131 CLK 0.447191
R17007 CLK.n134 CLK 0.447191
R17008 CLK.n125 CLK 0.447191
R17009 CLK.n109 CLK 0.447191
R17010 CLK.n96 CLK 0.447191
R17011 CLK.n83 CLK 0.447191
R17012 CLK.n70 CLK 0.447191
R17013 CLK.n57 CLK 0.447191
R17014 CLK.n44 CLK 0.447191
R17015 CLK.n32 CLK 0.447191
R17016 CLK.n20 CLK 0.447191
R17017 CLK.n8 CLK 0.447191
R17018 CLK.n246 CLK 0.436162
R17019 CLK.n233 CLK 0.436162
R17020 CLK.n220 CLK 0.436162
R17021 CLK.n207 CLK 0.436162
R17022 CLK.n194 CLK 0.436162
R17023 CLK.n181 CLK 0.436162
R17024 CLK.n168 CLK 0.436162
R17025 CLK.n156 CLK 0.436162
R17026 CLK.n106 CLK 0.436162
R17027 CLK.n93 CLK 0.436162
R17028 CLK.n80 CLK 0.436162
R17029 CLK.n67 CLK 0.436162
R17030 CLK.n54 CLK 0.436162
R17031 CLK.n41 CLK 0.436162
R17032 CLK.n29 CLK 0.436162
R17033 CLK.n17 CLK 0.436162
R17034 CLK.n5 CLK 0.436162
R17035 CLK.n244 CLK 0.321667
R17036 CLK.n231 CLK 0.321667
R17037 CLK.n218 CLK 0.321667
R17038 CLK.n205 CLK 0.321667
R17039 CLK.n192 CLK 0.321667
R17040 CLK.n179 CLK 0.321667
R17041 CLK.n166 CLK 0.321667
R17042 CLK.n154 CLK 0.321667
R17043 CLK.n104 CLK 0.321667
R17044 CLK.n91 CLK 0.321667
R17045 CLK.n78 CLK 0.321667
R17046 CLK.n65 CLK 0.321667
R17047 CLK.n52 CLK 0.321667
R17048 CLK.n39 CLK 0.321667
R17049 CLK.n27 CLK 0.321667
R17050 CLK.n15 CLK 0.321667
R17051 CLK.n3 CLK 0.321667
R17052 CLK.n241 CLK 0.217464
R17053 CLK.n228 CLK 0.217464
R17054 CLK.n215 CLK 0.217464
R17055 CLK.n202 CLK 0.217464
R17056 CLK.n189 CLK 0.217464
R17057 CLK.n176 CLK 0.217464
R17058 CLK.n163 CLK 0.217464
R17059 CLK.n151 CLK 0.217464
R17060 CLK.n101 CLK 0.217464
R17061 CLK.n88 CLK 0.217464
R17062 CLK.n75 CLK 0.217464
R17063 CLK.n62 CLK 0.217464
R17064 CLK.n49 CLK 0.217464
R17065 CLK.n36 CLK 0.217464
R17066 CLK.n24 CLK 0.217464
R17067 CLK.n12 CLK 0.217464
R17068 CLK.n0 CLK 0.217464
R17069 CLK.n245 CLK 0.208867
R17070 CLK.n232 CLK 0.208867
R17071 CLK.n219 CLK 0.208867
R17072 CLK.n206 CLK 0.208867
R17073 CLK.n193 CLK 0.208867
R17074 CLK.n180 CLK 0.208867
R17075 CLK.n167 CLK 0.208867
R17076 CLK.n155 CLK 0.208867
R17077 CLK.n105 CLK 0.208867
R17078 CLK.n92 CLK 0.208867
R17079 CLK.n79 CLK 0.208867
R17080 CLK.n66 CLK 0.208867
R17081 CLK.n53 CLK 0.208867
R17082 CLK.n40 CLK 0.208867
R17083 CLK.n28 CLK 0.208867
R17084 CLK.n16 CLK 0.208867
R17085 CLK.n4 CLK 0.208867
R17086 CLK.n248 CLK 0.149957
R17087 CLK.n235 CLK 0.149957
R17088 CLK.n222 CLK 0.149957
R17089 CLK.n209 CLK 0.149957
R17090 CLK.n196 CLK 0.149957
R17091 CLK.n183 CLK 0.149957
R17092 CLK.n170 CLK 0.149957
R17093 CLK.n158 CLK 0.149957
R17094 CLK.n129 CLK 0.149957
R17095 CLK.n132 CLK 0.149957
R17096 CLK.n135 CLK 0.149957
R17097 CLK.n126 CLK 0.149957
R17098 CLK.n108 CLK 0.149957
R17099 CLK.n95 CLK 0.149957
R17100 CLK.n82 CLK 0.149957
R17101 CLK.n69 CLK 0.149957
R17102 CLK.n56 CLK 0.149957
R17103 CLK.n43 CLK 0.149957
R17104 CLK.n31 CLK 0.149957
R17105 CLK.n19 CLK 0.149957
R17106 CLK.n7 CLK 0.149957
R17107 CLK.n245 CLK.n244 0.145417
R17108 CLK.n251 CLK.n250 0.145417
R17109 CLK.n232 CLK.n231 0.145417
R17110 CLK.n238 CLK.n237 0.145417
R17111 CLK.n219 CLK.n218 0.145417
R17112 CLK.n225 CLK.n224 0.145417
R17113 CLK.n206 CLK.n205 0.145417
R17114 CLK.n212 CLK.n211 0.145417
R17115 CLK.n193 CLK.n192 0.145417
R17116 CLK.n199 CLK.n198 0.145417
R17117 CLK.n180 CLK.n179 0.145417
R17118 CLK.n186 CLK.n185 0.145417
R17119 CLK.n167 CLK.n166 0.145417
R17120 CLK.n173 CLK.n172 0.145417
R17121 CLK.n155 CLK.n154 0.145417
R17122 CLK.n161 CLK.n160 0.145417
R17123 CLK.n105 CLK.n104 0.145417
R17124 CLK.n111 CLK.n110 0.145417
R17125 CLK.n92 CLK.n91 0.145417
R17126 CLK.n98 CLK.n97 0.145417
R17127 CLK.n79 CLK.n78 0.145417
R17128 CLK.n85 CLK.n84 0.145417
R17129 CLK.n66 CLK.n65 0.145417
R17130 CLK.n72 CLK.n71 0.145417
R17131 CLK.n53 CLK.n52 0.145417
R17132 CLK.n59 CLK.n58 0.145417
R17133 CLK.n40 CLK.n39 0.145417
R17134 CLK.n46 CLK.n45 0.145417
R17135 CLK.n28 CLK.n27 0.145417
R17136 CLK.n34 CLK.n33 0.145417
R17137 CLK.n16 CLK.n15 0.145417
R17138 CLK.n22 CLK.n21 0.145417
R17139 CLK.n4 CLK.n3 0.145417
R17140 CLK.n10 CLK.n9 0.145417
R17141 CLK.n242 CLK 0.1255
R17142 CLK.n229 CLK 0.1255
R17143 CLK.n216 CLK 0.1255
R17144 CLK.n203 CLK 0.1255
R17145 CLK.n190 CLK 0.1255
R17146 CLK.n177 CLK 0.1255
R17147 CLK.n164 CLK 0.1255
R17148 CLK.n152 CLK 0.1255
R17149 CLK.n121 CLK 0.1255
R17150 CLK.n117 CLK 0.1255
R17151 CLK.n139 CLK 0.1255
R17152 CLK.n144 CLK 0.1255
R17153 CLK.n102 CLK 0.1255
R17154 CLK.n89 CLK 0.1255
R17155 CLK.n76 CLK 0.1255
R17156 CLK.n63 CLK 0.1255
R17157 CLK.n50 CLK 0.1255
R17158 CLK.n37 CLK 0.1255
R17159 CLK.n25 CLK 0.1255
R17160 CLK.n13 CLK 0.1255
R17161 CLK.n1 CLK 0.1255
R17162 CLK.n251 CLK 0.118
R17163 CLK.n238 CLK 0.118
R17164 CLK.n225 CLK 0.118
R17165 CLK.n212 CLK 0.118
R17166 CLK.n199 CLK 0.118
R17167 CLK.n186 CLK 0.118
R17168 CLK.n173 CLK 0.118
R17169 CLK.n161 CLK 0.118
R17170 CLK.n111 CLK 0.118
R17171 CLK.n98 CLK 0.118
R17172 CLK.n85 CLK 0.118
R17173 CLK.n72 CLK 0.118
R17174 CLK.n59 CLK 0.118
R17175 CLK.n46 CLK 0.118
R17176 CLK.n34 CLK 0.118
R17177 CLK.n22 CLK 0.118
R17178 CLK.n10 CLK 0.118
R17179 CLK.n247 CLK 0.117348
R17180 CLK.n234 CLK 0.117348
R17181 CLK.n221 CLK 0.117348
R17182 CLK.n208 CLK 0.117348
R17183 CLK.n195 CLK 0.117348
R17184 CLK.n182 CLK 0.117348
R17185 CLK.n169 CLK 0.117348
R17186 CLK.n157 CLK 0.117348
R17187 CLK.n107 CLK 0.117348
R17188 CLK.n94 CLK 0.117348
R17189 CLK.n81 CLK 0.117348
R17190 CLK.n68 CLK 0.117348
R17191 CLK.n55 CLK 0.117348
R17192 CLK.n42 CLK 0.117348
R17193 CLK.n30 CLK 0.117348
R17194 CLK.n18 CLK 0.117348
R17195 CLK.n6 CLK 0.117348
R17196 CLK.n123 CLK.n122 0.063
R17197 CLK.n119 CLK.n118 0.063
R17198 CLK.n141 CLK.n140 0.063
R17199 CLK.n146 CLK.n145 0.063
R17200 CLK.n247 CLK 0.0454219
R17201 CLK.n248 CLK 0.0454219
R17202 CLK.n234 CLK 0.0454219
R17203 CLK.n235 CLK 0.0454219
R17204 CLK.n221 CLK 0.0454219
R17205 CLK.n222 CLK 0.0454219
R17206 CLK.n208 CLK 0.0454219
R17207 CLK.n209 CLK 0.0454219
R17208 CLK.n195 CLK 0.0454219
R17209 CLK.n196 CLK 0.0454219
R17210 CLK.n182 CLK 0.0454219
R17211 CLK.n183 CLK 0.0454219
R17212 CLK.n169 CLK 0.0454219
R17213 CLK.n170 CLK 0.0454219
R17214 CLK.n157 CLK 0.0454219
R17215 CLK.n158 CLK 0.0454219
R17216 CLK.n129 CLK 0.0454219
R17217 CLK.n132 CLK 0.0454219
R17218 CLK.n135 CLK 0.0454219
R17219 CLK.n126 CLK 0.0454219
R17220 CLK.n107 CLK 0.0454219
R17221 CLK.n108 CLK 0.0454219
R17222 CLK.n94 CLK 0.0454219
R17223 CLK.n95 CLK 0.0454219
R17224 CLK.n81 CLK 0.0454219
R17225 CLK.n82 CLK 0.0454219
R17226 CLK.n68 CLK 0.0454219
R17227 CLK.n69 CLK 0.0454219
R17228 CLK.n55 CLK 0.0454219
R17229 CLK.n56 CLK 0.0454219
R17230 CLK.n42 CLK 0.0454219
R17231 CLK.n43 CLK 0.0454219
R17232 CLK.n30 CLK 0.0454219
R17233 CLK.n31 CLK 0.0454219
R17234 CLK.n18 CLK 0.0454219
R17235 CLK.n19 CLK 0.0454219
R17236 CLK.n6 CLK 0.0454219
R17237 CLK.n7 CLK 0.0454219
R17238 CLK.n252 CLK.n245 0.024
R17239 CLK.n252 CLK.n251 0.024
R17240 CLK.n239 CLK.n232 0.024
R17241 CLK.n239 CLK.n238 0.024
R17242 CLK.n226 CLK.n219 0.024
R17243 CLK.n226 CLK.n225 0.024
R17244 CLK.n213 CLK.n206 0.024
R17245 CLK.n213 CLK.n212 0.024
R17246 CLK.n200 CLK.n193 0.024
R17247 CLK.n200 CLK.n199 0.024
R17248 CLK.n187 CLK.n180 0.024
R17249 CLK.n187 CLK.n186 0.024
R17250 CLK.n174 CLK.n167 0.024
R17251 CLK.n174 CLK.n173 0.024
R17252 CLK.n162 CLK.n155 0.024
R17253 CLK.n162 CLK.n161 0.024
R17254 CLK.n112 CLK.n105 0.024
R17255 CLK.n112 CLK.n111 0.024
R17256 CLK.n99 CLK.n92 0.024
R17257 CLK.n99 CLK.n98 0.024
R17258 CLK.n86 CLK.n79 0.024
R17259 CLK.n86 CLK.n85 0.024
R17260 CLK.n73 CLK.n66 0.024
R17261 CLK.n73 CLK.n72 0.024
R17262 CLK.n60 CLK.n53 0.024
R17263 CLK.n60 CLK.n59 0.024
R17264 CLK.n47 CLK.n40 0.024
R17265 CLK.n47 CLK.n46 0.024
R17266 CLK.n35 CLK.n28 0.024
R17267 CLK.n35 CLK.n34 0.024
R17268 CLK.n23 CLK.n16 0.024
R17269 CLK.n23 CLK.n22 0.024
R17270 CLK.n11 CLK.n4 0.024
R17271 CLK.n11 CLK.n10 0.024
R17272 CLK.n150 CLK.n149 0.024
R17273 CLK CLK.n253 0.0232879
R17274 CLK.n243 CLK.n242 0.0216397
R17275 CLK.n243 CLK 0.0216397
R17276 CLK.n230 CLK.n229 0.0216397
R17277 CLK.n230 CLK 0.0216397
R17278 CLK.n217 CLK.n216 0.0216397
R17279 CLK.n217 CLK 0.0216397
R17280 CLK.n204 CLK.n203 0.0216397
R17281 CLK.n204 CLK 0.0216397
R17282 CLK.n191 CLK.n190 0.0216397
R17283 CLK.n191 CLK 0.0216397
R17284 CLK.n178 CLK.n177 0.0216397
R17285 CLK.n178 CLK 0.0216397
R17286 CLK.n165 CLK.n164 0.0216397
R17287 CLK.n165 CLK 0.0216397
R17288 CLK.n153 CLK.n152 0.0216397
R17289 CLK.n153 CLK 0.0216397
R17290 CLK.n103 CLK.n102 0.0216397
R17291 CLK.n103 CLK 0.0216397
R17292 CLK.n90 CLK.n89 0.0216397
R17293 CLK.n90 CLK 0.0216397
R17294 CLK.n77 CLK.n76 0.0216397
R17295 CLK.n77 CLK 0.0216397
R17296 CLK.n64 CLK.n63 0.0216397
R17297 CLK.n64 CLK 0.0216397
R17298 CLK.n51 CLK.n50 0.0216397
R17299 CLK.n51 CLK 0.0216397
R17300 CLK.n38 CLK.n37 0.0216397
R17301 CLK.n38 CLK 0.0216397
R17302 CLK.n26 CLK.n25 0.0216397
R17303 CLK.n26 CLK 0.0216397
R17304 CLK.n14 CLK.n13 0.0216397
R17305 CLK.n14 CLK 0.0216397
R17306 CLK.n2 CLK.n1 0.0216397
R17307 CLK.n2 CLK 0.0216397
R17308 CLK.n121 CLK.n120 0.0107679
R17309 CLK.n120 CLK 0.0107679
R17310 CLK.n117 CLK.n116 0.0107679
R17311 CLK.n116 CLK 0.0107679
R17312 CLK.n139 CLK.n138 0.0107679
R17313 CLK.n138 CLK 0.0107679
R17314 CLK.n144 CLK.n143 0.0107679
R17315 CLK.n143 CLK 0.0107679
R17316 CLK.n250 CLK 0.00441667
R17317 CLK.n237 CLK 0.00441667
R17318 CLK.n224 CLK 0.00441667
R17319 CLK.n211 CLK 0.00441667
R17320 CLK.n198 CLK 0.00441667
R17321 CLK.n185 CLK 0.00441667
R17322 CLK.n172 CLK 0.00441667
R17323 CLK.n160 CLK 0.00441667
R17324 CLK.n110 CLK 0.00441667
R17325 CLK.n97 CLK 0.00441667
R17326 CLK.n84 CLK 0.00441667
R17327 CLK.n71 CLK 0.00441667
R17328 CLK.n58 CLK 0.00441667
R17329 CLK.n45 CLK 0.00441667
R17330 CLK.n33 CLK 0.00441667
R17331 CLK.n21 CLK 0.00441667
R17332 CLK.n9 CLK 0.00441667
R17333 CLK.n250 CLK 0.00406061
R17334 CLK.n237 CLK 0.00406061
R17335 CLK.n224 CLK 0.00406061
R17336 CLK.n211 CLK 0.00406061
R17337 CLK.n198 CLK 0.00406061
R17338 CLK.n185 CLK 0.00406061
R17339 CLK.n172 CLK 0.00406061
R17340 CLK.n160 CLK 0.00406061
R17341 CLK.n110 CLK 0.00406061
R17342 CLK.n97 CLK 0.00406061
R17343 CLK.n84 CLK 0.00406061
R17344 CLK.n71 CLK 0.00406061
R17345 CLK.n58 CLK 0.00406061
R17346 CLK.n45 CLK 0.00406061
R17347 CLK.n33 CLK 0.00406061
R17348 CLK.n21 CLK 0.00406061
R17349 CLK.n9 CLK 0.00406061
R17350 CLK.n254 CLK 0.00128333
R17351 CLK.n254 CLK 0.00121212
R17352 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 169.46
R17353 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 168.089
R17354 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 167.809
R17355 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 150.293
R17356 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 73.6304
R17357 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 60.4568
R17358 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 12.0358
R17359 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 11.4489
R17360 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.981478
R17361 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 0.788543
R17362 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.769522
R17363 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 0.720633
R17364 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 0.682565
R17365 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.580578
R17366 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 0.55213
R17367 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 0.470609
R17368 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.447191
R17369 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.428234
R17370 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.1255
R17371 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.1255
R17372 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 0.063
R17373 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 0.063
R17374 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.063
R17375 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 0.063
R17376 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 0.063
R17377 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 0.0435206
R17378 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 0.0107679
R17379 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.0107679
R17380 Nand_Gate_4.A.n33 Nand_Gate_4.A.t0 169.46
R17381 Nand_Gate_4.A.n33 Nand_Gate_4.A.t3 167.809
R17382 Nand_Gate_4.A.n35 Nand_Gate_4.A.t2 167.809
R17383 Nand_Gate_4.A Nand_Gate_4.A.t4 158.585
R17384 Nand_Gate_4.A.n21 Nand_Gate_4.A.t8 150.293
R17385 Nand_Gate_4.A.t4 Nand_Gate_4.A.n2 150.293
R17386 Nand_Gate_4.A.n14 Nand_Gate_4.A.t7 150.273
R17387 Nand_Gate_4.A.n8 Nand_Gate_4.A.t11 150.273
R17388 Nand_Gate_4.A.n12 Nand_Gate_4.A.t9 73.6406
R17389 Nand_Gate_4.A.n6 Nand_Gate_4.A.t5 73.6406
R17390 Nand_Gate_4.A.n23 Nand_Gate_4.A.t6 73.6304
R17391 Nand_Gate_4.A.n0 Nand_Gate_4.A.t10 73.6304
R17392 Nand_Gate_4.A.n4 Nand_Gate_4.A.t1 60.3809
R17393 Nand_Gate_4.A.n27 Nand_Gate_4.A.n26 14.3097
R17394 Nand_Gate_4.A.n34 Nand_Gate_4.A.n33 11.4489
R17395 Nand_Gate_4.A.n36 Nand_Gate_4.A.n35 8.21389
R17396 Nand_Gate_4.A.n18 Nand_Gate_4.A.n11 8.1418
R17397 Nand_Gate_4.A.n29 Nand_Gate_4.A.n28 5.61191
R17398 Nand_Gate_4.A.n29 Nand_Gate_4.A 5.35402
R17399 Nand_Gate_4.A.n30 Nand_Gate_4.A.n29 4.563
R17400 Nand_Gate_4.A.n18 Nand_Gate_4.A.n17 4.5005
R17401 Nand_Gate_4.A.n28 Nand_Gate_4.A 1.83746
R17402 Nand_Gate_4.A.n20 Nand_Gate_4.A.n19 1.62007
R17403 Nand_Gate_4.A.n2 Nand_Gate_4.A.n1 1.19615
R17404 Nand_Gate_4.A.n5 Nand_Gate_4.A 1.08746
R17405 Nand_Gate_4.A.n20 Nand_Gate_4.A 1.01739
R17406 Nand_Gate_4.A.n13 Nand_Gate_4.A 0.851043
R17407 Nand_Gate_4.A.n7 Nand_Gate_4.A 0.851043
R17408 Nand_Gate_4.A.n4 Nand_Gate_4.A 0.848156
R17409 Nand_Gate_4.A.n32 Nand_Gate_4.A.n31 0.788543
R17410 Nand_Gate_4.A.n22 Nand_Gate_4.A 0.769522
R17411 Nand_Gate_4.A.n5 Nand_Gate_4.A.n4 0.682565
R17412 Nand_Gate_4.A.n31 Nand_Gate_4.A 0.65675
R17413 Nand_Gate_4.A.n22 Nand_Gate_4.A.n21 0.55213
R17414 Nand_Gate_4.A.n16 Nand_Gate_4.A.n15 0.55213
R17415 Nand_Gate_4.A.n10 Nand_Gate_4.A.n9 0.55213
R17416 Nand_Gate_4.A.n16 Nand_Gate_4.A 0.486828
R17417 Nand_Gate_4.A.n10 Nand_Gate_4.A 0.486828
R17418 Nand_Gate_4.A.n25 Nand_Gate_4.A.n24 0.470609
R17419 Nand_Gate_4.A.n13 Nand_Gate_4.A.n12 0.470609
R17420 Nand_Gate_4.A.n7 Nand_Gate_4.A.n6 0.470609
R17421 Nand_Gate_4.A.n21 Nand_Gate_4.A 0.447191
R17422 Nand_Gate_4.A.n2 Nand_Gate_4.A 0.447191
R17423 Nand_Gate_4.A.n25 Nand_Gate_4.A 0.428234
R17424 Nand_Gate_4.A.n36 Nand_Gate_4.A.n3 0.425067
R17425 Nand_Gate_4.A Nand_Gate_4.A.n36 0.39003
R17426 Nand_Gate_4.A.n35 Nand_Gate_4.A.n34 0.280391
R17427 Nand_Gate_4.A.n34 Nand_Gate_4.A.n32 0.262643
R17428 Nand_Gate_4.A.n12 Nand_Gate_4.A 0.217464
R17429 Nand_Gate_4.A.n6 Nand_Gate_4.A 0.217464
R17430 Nand_Gate_4.A.n24 Nand_Gate_4.A 0.1255
R17431 Nand_Gate_4.A.n15 Nand_Gate_4.A 0.1255
R17432 Nand_Gate_4.A.n9 Nand_Gate_4.A 0.1255
R17433 Nand_Gate_4.A.n32 Nand_Gate_4.A 0.1255
R17434 Nand_Gate_4.A.n1 Nand_Gate_4.A 0.1255
R17435 Nand_Gate_4.A.n26 Nand_Gate_4.A.n22 0.063
R17436 Nand_Gate_4.A.n26 Nand_Gate_4.A.n25 0.063
R17437 Nand_Gate_4.A.n17 Nand_Gate_4.A.n13 0.063
R17438 Nand_Gate_4.A.n17 Nand_Gate_4.A.n16 0.063
R17439 Nand_Gate_4.A.n11 Nand_Gate_4.A.n7 0.063
R17440 Nand_Gate_4.A.n11 Nand_Gate_4.A.n10 0.063
R17441 Nand_Gate_4.A.n28 Nand_Gate_4.A.n27 0.063
R17442 Nand_Gate_4.A.n27 Nand_Gate_4.A.n20 0.063
R17443 Nand_Gate_4.A.n30 Nand_Gate_4.A.n5 0.063
R17444 Nand_Gate_4.A.n31 Nand_Gate_4.A.n30 0.063
R17445 Nand_Gate_4.A.n32 Nand_Gate_4.A 0.063
R17446 Nand_Gate_4.A Nand_Gate_4.A.n18 0.0512812
R17447 Nand_Gate_4.A.n15 Nand_Gate_4.A.n14 0.0216397
R17448 Nand_Gate_4.A.n14 Nand_Gate_4.A 0.0216397
R17449 Nand_Gate_4.A.n9 Nand_Gate_4.A.n8 0.0216397
R17450 Nand_Gate_4.A.n8 Nand_Gate_4.A 0.0216397
R17451 Nand_Gate_4.A.n19 Nand_Gate_4.A 0.0168043
R17452 Nand_Gate_4.A.n19 Nand_Gate_4.A 0.0122188
R17453 Nand_Gate_4.A.n24 Nand_Gate_4.A.n23 0.0107679
R17454 Nand_Gate_4.A.n23 Nand_Gate_4.A 0.0107679
R17455 Nand_Gate_4.A.n1 Nand_Gate_4.A.n0 0.0107679
R17456 Nand_Gate_4.A.n0 Nand_Gate_4.A 0.0107679
R17457 Nand_Gate_4.A.n3 Nand_Gate_4.A 0.00441667
R17458 Nand_Gate_4.A.n3 Nand_Gate_4.A 0.00406061
R17459 VDD.n275 VDD.n269 12650.1
R17460 VDD.n273 VDD.n272 12650.1
R17461 VDD.n257 VDD.n254 10684.6
R17462 VDD.n263 VDD.n249 10684.6
R17463 VDD.n251 VDD.n248 10167.6
R17464 VDD.n252 VDD.n251 10167.6
R17465 VDD.n276 VDD.n270 2427.48
R17466 VDD.n270 VDD.n268 2427.48
R17467 VDD.n277 VDD.n276 2349.78
R17468 VDD.n277 VDD.n268 2349.78
R17469 VDD.n260 VDD.n247 2051.01
R17470 VDD.n258 VDD.n253 2051.01
R17471 VDD.n264 VDD.n247 1973.31
R17472 VDD.n253 VDD.n246 1973.31
R17473 VDD.n265 VDD.n245 1952
R17474 VDD.n259 VDD.n245 1952
R17475 VDD.n7601 VDD.n7588 1084.97
R17476 VDD.n7601 VDD.n7589 1084.97
R17477 VDD.n7608 VDD.n7589 1084.97
R17478 VDD.n7608 VDD.n7588 1084.97
R17479 VDD.n7611 VDD.n7578 1084.97
R17480 VDD.n7611 VDD.n7579 1084.97
R17481 VDD.n7618 VDD.n7579 1084.97
R17482 VDD.n7618 VDD.n7578 1084.97
R17483 VDD.n7621 VDD.n7567 1084.97
R17484 VDD.n7621 VDD.n7568 1084.97
R17485 VDD.n7628 VDD.n7568 1084.97
R17486 VDD.n7628 VDD.n7567 1084.97
R17487 VDD.n7631 VDD.n7554 1084.97
R17488 VDD.n7631 VDD.n7555 1084.97
R17489 VDD.n7638 VDD.n7555 1084.97
R17490 VDD.n7638 VDD.n7554 1084.97
R17491 VDD.n7641 VDD.n7542 1084.97
R17492 VDD.n7641 VDD.n7543 1084.97
R17493 VDD.n7648 VDD.n7543 1084.97
R17494 VDD.n7648 VDD.n7542 1084.97
R17495 VDD.n7658 VDD.n7526 1084.97
R17496 VDD.n7658 VDD.n7527 1084.97
R17497 VDD.n7665 VDD.n7527 1084.97
R17498 VDD.n7665 VDD.n7526 1084.97
R17499 VDD.n7668 VDD.n7516 1084.97
R17500 VDD.n7668 VDD.n7517 1084.97
R17501 VDD.n7675 VDD.n7517 1084.97
R17502 VDD.n7675 VDD.n7516 1084.97
R17503 VDD.n7678 VDD.n7505 1084.97
R17504 VDD.n7678 VDD.n7506 1084.97
R17505 VDD.n7685 VDD.n7506 1084.97
R17506 VDD.n7685 VDD.n7505 1084.97
R17507 VDD.n7688 VDD.n7492 1084.97
R17508 VDD.n7688 VDD.n7493 1084.97
R17509 VDD.n7695 VDD.n7493 1084.97
R17510 VDD.n7695 VDD.n7492 1084.97
R17511 VDD.n7698 VDD.n7483 1084.97
R17512 VDD.n7698 VDD.n7484 1084.97
R17513 VDD.n7705 VDD.n7484 1084.97
R17514 VDD.n7705 VDD.n7483 1084.97
R17515 VDD.n7713 VDD.n7709 1084.97
R17516 VDD.n7709 VDD.n7463 1084.97
R17517 VDD.n7708 VDD.n7463 1084.97
R17518 VDD.n7713 VDD.n7708 1084.97
R17519 VDD.n7604 VDD.n7603 1084.97
R17520 VDD.n7603 VDD.n7597 1084.97
R17521 VDD.n7597 VDD.n7587 1084.97
R17522 VDD.n7604 VDD.n7587 1084.97
R17523 VDD.n7614 VDD.n7613 1084.97
R17524 VDD.n7613 VDD.n7584 1084.97
R17525 VDD.n7584 VDD.n7577 1084.97
R17526 VDD.n7614 VDD.n7577 1084.97
R17527 VDD.n7624 VDD.n7623 1084.97
R17528 VDD.n7623 VDD.n7574 1084.97
R17529 VDD.n7574 VDD.n7566 1084.97
R17530 VDD.n7624 VDD.n7566 1084.97
R17531 VDD.n7634 VDD.n7633 1084.97
R17532 VDD.n7633 VDD.n7563 1084.97
R17533 VDD.n7563 VDD.n7553 1084.97
R17534 VDD.n7634 VDD.n7553 1084.97
R17535 VDD.n7644 VDD.n7643 1084.97
R17536 VDD.n7643 VDD.n7550 1084.97
R17537 VDD.n7550 VDD.n7541 1084.97
R17538 VDD.n7644 VDD.n7541 1084.97
R17539 VDD.n7651 VDD.n7538 1084.97
R17540 VDD.n7651 VDD.n7539 1084.97
R17541 VDD.n7655 VDD.n7539 1084.97
R17542 VDD.n7655 VDD.n7538 1084.97
R17543 VDD.n7661 VDD.n7660 1084.97
R17544 VDD.n7660 VDD.n7535 1084.97
R17545 VDD.n7535 VDD.n7525 1084.97
R17546 VDD.n7661 VDD.n7525 1084.97
R17547 VDD.n7671 VDD.n7670 1084.97
R17548 VDD.n7670 VDD.n7522 1084.97
R17549 VDD.n7522 VDD.n7515 1084.97
R17550 VDD.n7671 VDD.n7515 1084.97
R17551 VDD.n7681 VDD.n7680 1084.97
R17552 VDD.n7680 VDD.n7512 1084.97
R17553 VDD.n7512 VDD.n7504 1084.97
R17554 VDD.n7681 VDD.n7504 1084.97
R17555 VDD.n7691 VDD.n7690 1084.97
R17556 VDD.n7690 VDD.n7501 1084.97
R17557 VDD.n7501 VDD.n7491 1084.97
R17558 VDD.n7691 VDD.n7491 1084.97
R17559 VDD.n7701 VDD.n7700 1084.97
R17560 VDD.n7700 VDD.n7488 1084.97
R17561 VDD.n7488 VDD.n7482 1084.97
R17562 VDD.n7701 VDD.n7482 1084.97
R17563 VDD.n7714 VDD.n7466 1084.97
R17564 VDD.n7481 VDD.n7466 1084.97
R17565 VDD.n7481 VDD.n7465 1084.97
R17566 VDD.n7714 VDD.n7465 1084.97
R17567 VDD.n7471 VDD.n7467 1084.97
R17568 VDD.n7475 VDD.n7467 1084.97
R17569 VDD.n7475 VDD.n7468 1084.97
R17570 VDD.n1719 VDD.n1706 1084.97
R17571 VDD.n1719 VDD.n1707 1084.97
R17572 VDD.n1726 VDD.n1707 1084.97
R17573 VDD.n1726 VDD.n1706 1084.97
R17574 VDD.n1729 VDD.n1696 1084.97
R17575 VDD.n1729 VDD.n1697 1084.97
R17576 VDD.n1736 VDD.n1697 1084.97
R17577 VDD.n1736 VDD.n1696 1084.97
R17578 VDD.n1739 VDD.n1685 1084.97
R17579 VDD.n1739 VDD.n1686 1084.97
R17580 VDD.n1746 VDD.n1686 1084.97
R17581 VDD.n1746 VDD.n1685 1084.97
R17582 VDD.n1749 VDD.n1672 1084.97
R17583 VDD.n1749 VDD.n1673 1084.97
R17584 VDD.n1756 VDD.n1673 1084.97
R17585 VDD.n1756 VDD.n1672 1084.97
R17586 VDD.n1759 VDD.n1660 1084.97
R17587 VDD.n1759 VDD.n1661 1084.97
R17588 VDD.n1766 VDD.n1661 1084.97
R17589 VDD.n1766 VDD.n1660 1084.97
R17590 VDD.n1776 VDD.n1644 1084.97
R17591 VDD.n1776 VDD.n1645 1084.97
R17592 VDD.n1783 VDD.n1645 1084.97
R17593 VDD.n1783 VDD.n1644 1084.97
R17594 VDD.n1786 VDD.n1634 1084.97
R17595 VDD.n1786 VDD.n1635 1084.97
R17596 VDD.n1793 VDD.n1635 1084.97
R17597 VDD.n1793 VDD.n1634 1084.97
R17598 VDD.n1796 VDD.n1623 1084.97
R17599 VDD.n1796 VDD.n1624 1084.97
R17600 VDD.n1803 VDD.n1624 1084.97
R17601 VDD.n1803 VDD.n1623 1084.97
R17602 VDD.n1806 VDD.n1610 1084.97
R17603 VDD.n1806 VDD.n1611 1084.97
R17604 VDD.n1813 VDD.n1611 1084.97
R17605 VDD.n1813 VDD.n1610 1084.97
R17606 VDD.n1816 VDD.n1600 1084.97
R17607 VDD.n1816 VDD.n1601 1084.97
R17608 VDD.n1823 VDD.n1601 1084.97
R17609 VDD.n1823 VDD.n1600 1084.97
R17610 VDD.n1826 VDD.n1589 1084.97
R17611 VDD.n1826 VDD.n1590 1084.97
R17612 VDD.n1833 VDD.n1590 1084.97
R17613 VDD.n1833 VDD.n1589 1084.97
R17614 VDD.n1722 VDD.n1721 1084.97
R17615 VDD.n1721 VDD.n1715 1084.97
R17616 VDD.n1715 VDD.n1705 1084.97
R17617 VDD.n1722 VDD.n1705 1084.97
R17618 VDD.n1732 VDD.n1731 1084.97
R17619 VDD.n1731 VDD.n1702 1084.97
R17620 VDD.n1702 VDD.n1695 1084.97
R17621 VDD.n1732 VDD.n1695 1084.97
R17622 VDD.n1742 VDD.n1741 1084.97
R17623 VDD.n1741 VDD.n1692 1084.97
R17624 VDD.n1692 VDD.n1684 1084.97
R17625 VDD.n1742 VDD.n1684 1084.97
R17626 VDD.n1752 VDD.n1751 1084.97
R17627 VDD.n1751 VDD.n1681 1084.97
R17628 VDD.n1681 VDD.n1671 1084.97
R17629 VDD.n1752 VDD.n1671 1084.97
R17630 VDD.n1762 VDD.n1761 1084.97
R17631 VDD.n1761 VDD.n1668 1084.97
R17632 VDD.n1668 VDD.n1659 1084.97
R17633 VDD.n1762 VDD.n1659 1084.97
R17634 VDD.n1769 VDD.n1656 1084.97
R17635 VDD.n1769 VDD.n1657 1084.97
R17636 VDD.n1773 VDD.n1657 1084.97
R17637 VDD.n1773 VDD.n1656 1084.97
R17638 VDD.n1779 VDD.n1778 1084.97
R17639 VDD.n1778 VDD.n1653 1084.97
R17640 VDD.n1653 VDD.n1643 1084.97
R17641 VDD.n1779 VDD.n1643 1084.97
R17642 VDD.n1789 VDD.n1788 1084.97
R17643 VDD.n1788 VDD.n1640 1084.97
R17644 VDD.n1640 VDD.n1633 1084.97
R17645 VDD.n1789 VDD.n1633 1084.97
R17646 VDD.n1799 VDD.n1798 1084.97
R17647 VDD.n1798 VDD.n1630 1084.97
R17648 VDD.n1630 VDD.n1622 1084.97
R17649 VDD.n1799 VDD.n1622 1084.97
R17650 VDD.n1809 VDD.n1808 1084.97
R17651 VDD.n1808 VDD.n1619 1084.97
R17652 VDD.n1619 VDD.n1609 1084.97
R17653 VDD.n1809 VDD.n1609 1084.97
R17654 VDD.n1819 VDD.n1818 1084.97
R17655 VDD.n1818 VDD.n1606 1084.97
R17656 VDD.n1606 VDD.n1599 1084.97
R17657 VDD.n1819 VDD.n1599 1084.97
R17658 VDD.n1829 VDD.n1828 1084.97
R17659 VDD.n1828 VDD.n1596 1084.97
R17660 VDD.n1596 VDD.n1588 1084.97
R17661 VDD.n1829 VDD.n1588 1084.97
R17662 VDD.n1586 VDD.n1585 1084.97
R17663 VDD.n1836 VDD.n1585 1084.97
R17664 VDD.n1836 VDD.n1583 1084.97
R17665 VDD.n1459 VDD.n1446 1084.97
R17666 VDD.n1459 VDD.n1447 1084.97
R17667 VDD.n1466 VDD.n1447 1084.97
R17668 VDD.n1466 VDD.n1446 1084.97
R17669 VDD.n1469 VDD.n1436 1084.97
R17670 VDD.n1469 VDD.n1437 1084.97
R17671 VDD.n1476 VDD.n1437 1084.97
R17672 VDD.n1476 VDD.n1436 1084.97
R17673 VDD.n1479 VDD.n1425 1084.97
R17674 VDD.n1479 VDD.n1426 1084.97
R17675 VDD.n1486 VDD.n1426 1084.97
R17676 VDD.n1486 VDD.n1425 1084.97
R17677 VDD.n1489 VDD.n1412 1084.97
R17678 VDD.n1489 VDD.n1413 1084.97
R17679 VDD.n1496 VDD.n1413 1084.97
R17680 VDD.n1496 VDD.n1412 1084.97
R17681 VDD.n1499 VDD.n1400 1084.97
R17682 VDD.n1499 VDD.n1401 1084.97
R17683 VDD.n1506 VDD.n1401 1084.97
R17684 VDD.n1506 VDD.n1400 1084.97
R17685 VDD.n1516 VDD.n1384 1084.97
R17686 VDD.n1516 VDD.n1385 1084.97
R17687 VDD.n1523 VDD.n1385 1084.97
R17688 VDD.n1523 VDD.n1384 1084.97
R17689 VDD.n1526 VDD.n1374 1084.97
R17690 VDD.n1526 VDD.n1375 1084.97
R17691 VDD.n1533 VDD.n1375 1084.97
R17692 VDD.n1533 VDD.n1374 1084.97
R17693 VDD.n1536 VDD.n1363 1084.97
R17694 VDD.n1536 VDD.n1364 1084.97
R17695 VDD.n1543 VDD.n1364 1084.97
R17696 VDD.n1543 VDD.n1363 1084.97
R17697 VDD.n1546 VDD.n1350 1084.97
R17698 VDD.n1546 VDD.n1351 1084.97
R17699 VDD.n1553 VDD.n1351 1084.97
R17700 VDD.n1553 VDD.n1350 1084.97
R17701 VDD.n1556 VDD.n1340 1084.97
R17702 VDD.n1556 VDD.n1341 1084.97
R17703 VDD.n1563 VDD.n1341 1084.97
R17704 VDD.n1563 VDD.n1340 1084.97
R17705 VDD.n1566 VDD.n1329 1084.97
R17706 VDD.n1566 VDD.n1330 1084.97
R17707 VDD.n1573 VDD.n1330 1084.97
R17708 VDD.n1573 VDD.n1329 1084.97
R17709 VDD.n1462 VDD.n1461 1084.97
R17710 VDD.n1461 VDD.n1455 1084.97
R17711 VDD.n1455 VDD.n1445 1084.97
R17712 VDD.n1462 VDD.n1445 1084.97
R17713 VDD.n1472 VDD.n1471 1084.97
R17714 VDD.n1471 VDD.n1442 1084.97
R17715 VDD.n1442 VDD.n1435 1084.97
R17716 VDD.n1472 VDD.n1435 1084.97
R17717 VDD.n1482 VDD.n1481 1084.97
R17718 VDD.n1481 VDD.n1432 1084.97
R17719 VDD.n1432 VDD.n1424 1084.97
R17720 VDD.n1482 VDD.n1424 1084.97
R17721 VDD.n1492 VDD.n1491 1084.97
R17722 VDD.n1491 VDD.n1421 1084.97
R17723 VDD.n1421 VDD.n1411 1084.97
R17724 VDD.n1492 VDD.n1411 1084.97
R17725 VDD.n1502 VDD.n1501 1084.97
R17726 VDD.n1501 VDD.n1408 1084.97
R17727 VDD.n1408 VDD.n1399 1084.97
R17728 VDD.n1502 VDD.n1399 1084.97
R17729 VDD.n1509 VDD.n1396 1084.97
R17730 VDD.n1509 VDD.n1397 1084.97
R17731 VDD.n1513 VDD.n1397 1084.97
R17732 VDD.n1513 VDD.n1396 1084.97
R17733 VDD.n1519 VDD.n1518 1084.97
R17734 VDD.n1518 VDD.n1393 1084.97
R17735 VDD.n1393 VDD.n1383 1084.97
R17736 VDD.n1519 VDD.n1383 1084.97
R17737 VDD.n1529 VDD.n1528 1084.97
R17738 VDD.n1528 VDD.n1380 1084.97
R17739 VDD.n1380 VDD.n1373 1084.97
R17740 VDD.n1529 VDD.n1373 1084.97
R17741 VDD.n1539 VDD.n1538 1084.97
R17742 VDD.n1538 VDD.n1370 1084.97
R17743 VDD.n1370 VDD.n1362 1084.97
R17744 VDD.n1539 VDD.n1362 1084.97
R17745 VDD.n1549 VDD.n1548 1084.97
R17746 VDD.n1548 VDD.n1359 1084.97
R17747 VDD.n1359 VDD.n1349 1084.97
R17748 VDD.n1549 VDD.n1349 1084.97
R17749 VDD.n1559 VDD.n1558 1084.97
R17750 VDD.n1558 VDD.n1346 1084.97
R17751 VDD.n1346 VDD.n1339 1084.97
R17752 VDD.n1559 VDD.n1339 1084.97
R17753 VDD.n1569 VDD.n1568 1084.97
R17754 VDD.n1568 VDD.n1336 1084.97
R17755 VDD.n1336 VDD.n1328 1084.97
R17756 VDD.n1569 VDD.n1328 1084.97
R17757 VDD.n1326 VDD.n1325 1084.97
R17758 VDD.n1576 VDD.n1325 1084.97
R17759 VDD.n1576 VDD.n1323 1084.97
R17760 VDD.n1199 VDD.n1186 1084.97
R17761 VDD.n1199 VDD.n1187 1084.97
R17762 VDD.n1206 VDD.n1187 1084.97
R17763 VDD.n1206 VDD.n1186 1084.97
R17764 VDD.n1209 VDD.n1176 1084.97
R17765 VDD.n1209 VDD.n1177 1084.97
R17766 VDD.n1216 VDD.n1177 1084.97
R17767 VDD.n1216 VDD.n1176 1084.97
R17768 VDD.n1219 VDD.n1165 1084.97
R17769 VDD.n1219 VDD.n1166 1084.97
R17770 VDD.n1226 VDD.n1166 1084.97
R17771 VDD.n1226 VDD.n1165 1084.97
R17772 VDD.n1229 VDD.n1152 1084.97
R17773 VDD.n1229 VDD.n1153 1084.97
R17774 VDD.n1236 VDD.n1153 1084.97
R17775 VDD.n1236 VDD.n1152 1084.97
R17776 VDD.n1239 VDD.n1140 1084.97
R17777 VDD.n1239 VDD.n1141 1084.97
R17778 VDD.n1246 VDD.n1141 1084.97
R17779 VDD.n1246 VDD.n1140 1084.97
R17780 VDD.n1256 VDD.n1124 1084.97
R17781 VDD.n1256 VDD.n1125 1084.97
R17782 VDD.n1263 VDD.n1125 1084.97
R17783 VDD.n1263 VDD.n1124 1084.97
R17784 VDD.n1266 VDD.n1114 1084.97
R17785 VDD.n1266 VDD.n1115 1084.97
R17786 VDD.n1273 VDD.n1115 1084.97
R17787 VDD.n1273 VDD.n1114 1084.97
R17788 VDD.n1276 VDD.n1103 1084.97
R17789 VDD.n1276 VDD.n1104 1084.97
R17790 VDD.n1283 VDD.n1104 1084.97
R17791 VDD.n1283 VDD.n1103 1084.97
R17792 VDD.n1286 VDD.n1090 1084.97
R17793 VDD.n1286 VDD.n1091 1084.97
R17794 VDD.n1293 VDD.n1091 1084.97
R17795 VDD.n1293 VDD.n1090 1084.97
R17796 VDD.n1296 VDD.n1080 1084.97
R17797 VDD.n1296 VDD.n1081 1084.97
R17798 VDD.n1303 VDD.n1081 1084.97
R17799 VDD.n1303 VDD.n1080 1084.97
R17800 VDD.n1306 VDD.n1069 1084.97
R17801 VDD.n1306 VDD.n1070 1084.97
R17802 VDD.n1313 VDD.n1070 1084.97
R17803 VDD.n1313 VDD.n1069 1084.97
R17804 VDD.n1202 VDD.n1201 1084.97
R17805 VDD.n1201 VDD.n1195 1084.97
R17806 VDD.n1195 VDD.n1185 1084.97
R17807 VDD.n1202 VDD.n1185 1084.97
R17808 VDD.n1212 VDD.n1211 1084.97
R17809 VDD.n1211 VDD.n1182 1084.97
R17810 VDD.n1182 VDD.n1175 1084.97
R17811 VDD.n1212 VDD.n1175 1084.97
R17812 VDD.n1222 VDD.n1221 1084.97
R17813 VDD.n1221 VDD.n1172 1084.97
R17814 VDD.n1172 VDD.n1164 1084.97
R17815 VDD.n1222 VDD.n1164 1084.97
R17816 VDD.n1232 VDD.n1231 1084.97
R17817 VDD.n1231 VDD.n1161 1084.97
R17818 VDD.n1161 VDD.n1151 1084.97
R17819 VDD.n1232 VDD.n1151 1084.97
R17820 VDD.n1242 VDD.n1241 1084.97
R17821 VDD.n1241 VDD.n1148 1084.97
R17822 VDD.n1148 VDD.n1139 1084.97
R17823 VDD.n1242 VDD.n1139 1084.97
R17824 VDD.n1249 VDD.n1136 1084.97
R17825 VDD.n1249 VDD.n1137 1084.97
R17826 VDD.n1253 VDD.n1137 1084.97
R17827 VDD.n1253 VDD.n1136 1084.97
R17828 VDD.n1259 VDD.n1258 1084.97
R17829 VDD.n1258 VDD.n1133 1084.97
R17830 VDD.n1133 VDD.n1123 1084.97
R17831 VDD.n1259 VDD.n1123 1084.97
R17832 VDD.n1269 VDD.n1268 1084.97
R17833 VDD.n1268 VDD.n1120 1084.97
R17834 VDD.n1120 VDD.n1113 1084.97
R17835 VDD.n1269 VDD.n1113 1084.97
R17836 VDD.n1279 VDD.n1278 1084.97
R17837 VDD.n1278 VDD.n1110 1084.97
R17838 VDD.n1110 VDD.n1102 1084.97
R17839 VDD.n1279 VDD.n1102 1084.97
R17840 VDD.n1289 VDD.n1288 1084.97
R17841 VDD.n1288 VDD.n1099 1084.97
R17842 VDD.n1099 VDD.n1089 1084.97
R17843 VDD.n1289 VDD.n1089 1084.97
R17844 VDD.n1299 VDD.n1298 1084.97
R17845 VDD.n1298 VDD.n1086 1084.97
R17846 VDD.n1086 VDD.n1079 1084.97
R17847 VDD.n1299 VDD.n1079 1084.97
R17848 VDD.n1309 VDD.n1308 1084.97
R17849 VDD.n1308 VDD.n1076 1084.97
R17850 VDD.n1076 VDD.n1068 1084.97
R17851 VDD.n1309 VDD.n1068 1084.97
R17852 VDD.n1066 VDD.n1065 1084.97
R17853 VDD.n1316 VDD.n1065 1084.97
R17854 VDD.n1316 VDD.n1063 1084.97
R17855 VDD.n939 VDD.n926 1084.97
R17856 VDD.n939 VDD.n927 1084.97
R17857 VDD.n946 VDD.n927 1084.97
R17858 VDD.n946 VDD.n926 1084.97
R17859 VDD.n949 VDD.n916 1084.97
R17860 VDD.n949 VDD.n917 1084.97
R17861 VDD.n956 VDD.n917 1084.97
R17862 VDD.n956 VDD.n916 1084.97
R17863 VDD.n959 VDD.n905 1084.97
R17864 VDD.n959 VDD.n906 1084.97
R17865 VDD.n966 VDD.n906 1084.97
R17866 VDD.n966 VDD.n905 1084.97
R17867 VDD.n969 VDD.n892 1084.97
R17868 VDD.n969 VDD.n893 1084.97
R17869 VDD.n976 VDD.n893 1084.97
R17870 VDD.n976 VDD.n892 1084.97
R17871 VDD.n979 VDD.n880 1084.97
R17872 VDD.n979 VDD.n881 1084.97
R17873 VDD.n986 VDD.n881 1084.97
R17874 VDD.n986 VDD.n880 1084.97
R17875 VDD.n996 VDD.n864 1084.97
R17876 VDD.n996 VDD.n865 1084.97
R17877 VDD.n1003 VDD.n865 1084.97
R17878 VDD.n1003 VDD.n864 1084.97
R17879 VDD.n1006 VDD.n854 1084.97
R17880 VDD.n1006 VDD.n855 1084.97
R17881 VDD.n1013 VDD.n855 1084.97
R17882 VDD.n1013 VDD.n854 1084.97
R17883 VDD.n1016 VDD.n843 1084.97
R17884 VDD.n1016 VDD.n844 1084.97
R17885 VDD.n1023 VDD.n844 1084.97
R17886 VDD.n1023 VDD.n843 1084.97
R17887 VDD.n1026 VDD.n830 1084.97
R17888 VDD.n1026 VDD.n831 1084.97
R17889 VDD.n1033 VDD.n831 1084.97
R17890 VDD.n1033 VDD.n830 1084.97
R17891 VDD.n1036 VDD.n820 1084.97
R17892 VDD.n1036 VDD.n821 1084.97
R17893 VDD.n1043 VDD.n821 1084.97
R17894 VDD.n1043 VDD.n820 1084.97
R17895 VDD.n1046 VDD.n809 1084.97
R17896 VDD.n1046 VDD.n810 1084.97
R17897 VDD.n1053 VDD.n810 1084.97
R17898 VDD.n1053 VDD.n809 1084.97
R17899 VDD.n942 VDD.n941 1084.97
R17900 VDD.n941 VDD.n935 1084.97
R17901 VDD.n935 VDD.n925 1084.97
R17902 VDD.n942 VDD.n925 1084.97
R17903 VDD.n952 VDD.n951 1084.97
R17904 VDD.n951 VDD.n922 1084.97
R17905 VDD.n922 VDD.n915 1084.97
R17906 VDD.n952 VDD.n915 1084.97
R17907 VDD.n962 VDD.n961 1084.97
R17908 VDD.n961 VDD.n912 1084.97
R17909 VDD.n912 VDD.n904 1084.97
R17910 VDD.n962 VDD.n904 1084.97
R17911 VDD.n972 VDD.n971 1084.97
R17912 VDD.n971 VDD.n901 1084.97
R17913 VDD.n901 VDD.n891 1084.97
R17914 VDD.n972 VDD.n891 1084.97
R17915 VDD.n982 VDD.n981 1084.97
R17916 VDD.n981 VDD.n888 1084.97
R17917 VDD.n888 VDD.n879 1084.97
R17918 VDD.n982 VDD.n879 1084.97
R17919 VDD.n989 VDD.n876 1084.97
R17920 VDD.n989 VDD.n877 1084.97
R17921 VDD.n993 VDD.n877 1084.97
R17922 VDD.n993 VDD.n876 1084.97
R17923 VDD.n999 VDD.n998 1084.97
R17924 VDD.n998 VDD.n873 1084.97
R17925 VDD.n873 VDD.n863 1084.97
R17926 VDD.n999 VDD.n863 1084.97
R17927 VDD.n1009 VDD.n1008 1084.97
R17928 VDD.n1008 VDD.n860 1084.97
R17929 VDD.n860 VDD.n853 1084.97
R17930 VDD.n1009 VDD.n853 1084.97
R17931 VDD.n1019 VDD.n1018 1084.97
R17932 VDD.n1018 VDD.n850 1084.97
R17933 VDD.n850 VDD.n842 1084.97
R17934 VDD.n1019 VDD.n842 1084.97
R17935 VDD.n1029 VDD.n1028 1084.97
R17936 VDD.n1028 VDD.n839 1084.97
R17937 VDD.n839 VDD.n829 1084.97
R17938 VDD.n1029 VDD.n829 1084.97
R17939 VDD.n1039 VDD.n1038 1084.97
R17940 VDD.n1038 VDD.n826 1084.97
R17941 VDD.n826 VDD.n819 1084.97
R17942 VDD.n1039 VDD.n819 1084.97
R17943 VDD.n1049 VDD.n1048 1084.97
R17944 VDD.n1048 VDD.n816 1084.97
R17945 VDD.n816 VDD.n808 1084.97
R17946 VDD.n1049 VDD.n808 1084.97
R17947 VDD.n806 VDD.n805 1084.97
R17948 VDD.n1056 VDD.n805 1084.97
R17949 VDD.n1056 VDD.n803 1084.97
R17950 VDD.n679 VDD.n666 1084.97
R17951 VDD.n679 VDD.n667 1084.97
R17952 VDD.n686 VDD.n667 1084.97
R17953 VDD.n686 VDD.n666 1084.97
R17954 VDD.n689 VDD.n656 1084.97
R17955 VDD.n689 VDD.n657 1084.97
R17956 VDD.n696 VDD.n657 1084.97
R17957 VDD.n696 VDD.n656 1084.97
R17958 VDD.n699 VDD.n645 1084.97
R17959 VDD.n699 VDD.n646 1084.97
R17960 VDD.n706 VDD.n646 1084.97
R17961 VDD.n706 VDD.n645 1084.97
R17962 VDD.n709 VDD.n632 1084.97
R17963 VDD.n709 VDD.n633 1084.97
R17964 VDD.n716 VDD.n633 1084.97
R17965 VDD.n716 VDD.n632 1084.97
R17966 VDD.n719 VDD.n620 1084.97
R17967 VDD.n719 VDD.n621 1084.97
R17968 VDD.n726 VDD.n621 1084.97
R17969 VDD.n726 VDD.n620 1084.97
R17970 VDD.n736 VDD.n604 1084.97
R17971 VDD.n736 VDD.n605 1084.97
R17972 VDD.n743 VDD.n605 1084.97
R17973 VDD.n743 VDD.n604 1084.97
R17974 VDD.n746 VDD.n594 1084.97
R17975 VDD.n746 VDD.n595 1084.97
R17976 VDD.n753 VDD.n595 1084.97
R17977 VDD.n753 VDD.n594 1084.97
R17978 VDD.n756 VDD.n583 1084.97
R17979 VDD.n756 VDD.n584 1084.97
R17980 VDD.n763 VDD.n584 1084.97
R17981 VDD.n763 VDD.n583 1084.97
R17982 VDD.n766 VDD.n570 1084.97
R17983 VDD.n766 VDD.n571 1084.97
R17984 VDD.n773 VDD.n571 1084.97
R17985 VDD.n773 VDD.n570 1084.97
R17986 VDD.n776 VDD.n560 1084.97
R17987 VDD.n776 VDD.n561 1084.97
R17988 VDD.n783 VDD.n561 1084.97
R17989 VDD.n783 VDD.n560 1084.97
R17990 VDD.n786 VDD.n549 1084.97
R17991 VDD.n786 VDD.n550 1084.97
R17992 VDD.n793 VDD.n550 1084.97
R17993 VDD.n793 VDD.n549 1084.97
R17994 VDD.n682 VDD.n681 1084.97
R17995 VDD.n681 VDD.n675 1084.97
R17996 VDD.n675 VDD.n665 1084.97
R17997 VDD.n682 VDD.n665 1084.97
R17998 VDD.n692 VDD.n691 1084.97
R17999 VDD.n691 VDD.n662 1084.97
R18000 VDD.n662 VDD.n655 1084.97
R18001 VDD.n692 VDD.n655 1084.97
R18002 VDD.n702 VDD.n701 1084.97
R18003 VDD.n701 VDD.n652 1084.97
R18004 VDD.n652 VDD.n644 1084.97
R18005 VDD.n702 VDD.n644 1084.97
R18006 VDD.n712 VDD.n711 1084.97
R18007 VDD.n711 VDD.n641 1084.97
R18008 VDD.n641 VDD.n631 1084.97
R18009 VDD.n712 VDD.n631 1084.97
R18010 VDD.n722 VDD.n721 1084.97
R18011 VDD.n721 VDD.n628 1084.97
R18012 VDD.n628 VDD.n619 1084.97
R18013 VDD.n722 VDD.n619 1084.97
R18014 VDD.n729 VDD.n616 1084.97
R18015 VDD.n729 VDD.n617 1084.97
R18016 VDD.n733 VDD.n617 1084.97
R18017 VDD.n733 VDD.n616 1084.97
R18018 VDD.n739 VDD.n738 1084.97
R18019 VDD.n738 VDD.n613 1084.97
R18020 VDD.n613 VDD.n603 1084.97
R18021 VDD.n739 VDD.n603 1084.97
R18022 VDD.n749 VDD.n748 1084.97
R18023 VDD.n748 VDD.n600 1084.97
R18024 VDD.n600 VDD.n593 1084.97
R18025 VDD.n749 VDD.n593 1084.97
R18026 VDD.n759 VDD.n758 1084.97
R18027 VDD.n758 VDD.n590 1084.97
R18028 VDD.n590 VDD.n582 1084.97
R18029 VDD.n759 VDD.n582 1084.97
R18030 VDD.n769 VDD.n768 1084.97
R18031 VDD.n768 VDD.n579 1084.97
R18032 VDD.n579 VDD.n569 1084.97
R18033 VDD.n769 VDD.n569 1084.97
R18034 VDD.n779 VDD.n778 1084.97
R18035 VDD.n778 VDD.n566 1084.97
R18036 VDD.n566 VDD.n559 1084.97
R18037 VDD.n779 VDD.n559 1084.97
R18038 VDD.n789 VDD.n788 1084.97
R18039 VDD.n788 VDD.n556 1084.97
R18040 VDD.n556 VDD.n548 1084.97
R18041 VDD.n789 VDD.n548 1084.97
R18042 VDD.n546 VDD.n545 1084.97
R18043 VDD.n796 VDD.n545 1084.97
R18044 VDD.n796 VDD.n543 1084.97
R18045 VDD.n419 VDD.n406 1084.97
R18046 VDD.n419 VDD.n407 1084.97
R18047 VDD.n426 VDD.n407 1084.97
R18048 VDD.n426 VDD.n406 1084.97
R18049 VDD.n429 VDD.n396 1084.97
R18050 VDD.n429 VDD.n397 1084.97
R18051 VDD.n436 VDD.n397 1084.97
R18052 VDD.n436 VDD.n396 1084.97
R18053 VDD.n439 VDD.n385 1084.97
R18054 VDD.n439 VDD.n386 1084.97
R18055 VDD.n446 VDD.n386 1084.97
R18056 VDD.n446 VDD.n385 1084.97
R18057 VDD.n449 VDD.n372 1084.97
R18058 VDD.n449 VDD.n373 1084.97
R18059 VDD.n456 VDD.n373 1084.97
R18060 VDD.n456 VDD.n372 1084.97
R18061 VDD.n459 VDD.n360 1084.97
R18062 VDD.n459 VDD.n361 1084.97
R18063 VDD.n466 VDD.n361 1084.97
R18064 VDD.n466 VDD.n360 1084.97
R18065 VDD.n476 VDD.n344 1084.97
R18066 VDD.n476 VDD.n345 1084.97
R18067 VDD.n483 VDD.n345 1084.97
R18068 VDD.n483 VDD.n344 1084.97
R18069 VDD.n486 VDD.n334 1084.97
R18070 VDD.n486 VDD.n335 1084.97
R18071 VDD.n493 VDD.n335 1084.97
R18072 VDD.n493 VDD.n334 1084.97
R18073 VDD.n496 VDD.n323 1084.97
R18074 VDD.n496 VDD.n324 1084.97
R18075 VDD.n503 VDD.n324 1084.97
R18076 VDD.n503 VDD.n323 1084.97
R18077 VDD.n506 VDD.n310 1084.97
R18078 VDD.n506 VDD.n311 1084.97
R18079 VDD.n513 VDD.n311 1084.97
R18080 VDD.n513 VDD.n310 1084.97
R18081 VDD.n516 VDD.n300 1084.97
R18082 VDD.n516 VDD.n301 1084.97
R18083 VDD.n523 VDD.n301 1084.97
R18084 VDD.n523 VDD.n300 1084.97
R18085 VDD.n526 VDD.n289 1084.97
R18086 VDD.n526 VDD.n290 1084.97
R18087 VDD.n533 VDD.n290 1084.97
R18088 VDD.n533 VDD.n289 1084.97
R18089 VDD.n422 VDD.n421 1084.97
R18090 VDD.n421 VDD.n415 1084.97
R18091 VDD.n415 VDD.n405 1084.97
R18092 VDD.n422 VDD.n405 1084.97
R18093 VDD.n432 VDD.n431 1084.97
R18094 VDD.n431 VDD.n402 1084.97
R18095 VDD.n402 VDD.n395 1084.97
R18096 VDD.n432 VDD.n395 1084.97
R18097 VDD.n442 VDD.n441 1084.97
R18098 VDD.n441 VDD.n392 1084.97
R18099 VDD.n392 VDD.n384 1084.97
R18100 VDD.n442 VDD.n384 1084.97
R18101 VDD.n452 VDD.n451 1084.97
R18102 VDD.n451 VDD.n381 1084.97
R18103 VDD.n381 VDD.n371 1084.97
R18104 VDD.n452 VDD.n371 1084.97
R18105 VDD.n462 VDD.n461 1084.97
R18106 VDD.n461 VDD.n368 1084.97
R18107 VDD.n368 VDD.n359 1084.97
R18108 VDD.n462 VDD.n359 1084.97
R18109 VDD.n469 VDD.n356 1084.97
R18110 VDD.n469 VDD.n357 1084.97
R18111 VDD.n473 VDD.n357 1084.97
R18112 VDD.n473 VDD.n356 1084.97
R18113 VDD.n479 VDD.n478 1084.97
R18114 VDD.n478 VDD.n353 1084.97
R18115 VDD.n353 VDD.n343 1084.97
R18116 VDD.n479 VDD.n343 1084.97
R18117 VDD.n489 VDD.n488 1084.97
R18118 VDD.n488 VDD.n340 1084.97
R18119 VDD.n340 VDD.n333 1084.97
R18120 VDD.n489 VDD.n333 1084.97
R18121 VDD.n499 VDD.n498 1084.97
R18122 VDD.n498 VDD.n330 1084.97
R18123 VDD.n330 VDD.n322 1084.97
R18124 VDD.n499 VDD.n322 1084.97
R18125 VDD.n509 VDD.n508 1084.97
R18126 VDD.n508 VDD.n319 1084.97
R18127 VDD.n319 VDD.n309 1084.97
R18128 VDD.n509 VDD.n309 1084.97
R18129 VDD.n519 VDD.n518 1084.97
R18130 VDD.n518 VDD.n306 1084.97
R18131 VDD.n306 VDD.n299 1084.97
R18132 VDD.n519 VDD.n299 1084.97
R18133 VDD.n529 VDD.n528 1084.97
R18134 VDD.n528 VDD.n296 1084.97
R18135 VDD.n296 VDD.n288 1084.97
R18136 VDD.n529 VDD.n288 1084.97
R18137 VDD.n286 VDD.n285 1084.97
R18138 VDD.n536 VDD.n285 1084.97
R18139 VDD.n536 VDD.n283 1084.97
R18140 VDD.n103 VDD.n98 1084.97
R18141 VDD.n107 VDD.n99 1084.97
R18142 VDD.n107 VDD.n98 1084.97
R18143 VDD.n110 VDD.n93 1084.97
R18144 VDD.n96 VDD.n95 1084.97
R18145 VDD.n110 VDD.n95 1084.97
R18146 VDD.n117 VDD.n85 1084.97
R18147 VDD.n121 VDD.n86 1084.97
R18148 VDD.n121 VDD.n85 1084.97
R18149 VDD.n124 VDD.n82 1084.97
R18150 VDD.n124 VDD.n83 1084.97
R18151 VDD.n128 VDD.n83 1084.97
R18152 VDD.n128 VDD.n82 1084.97
R18153 VDD.n131 VDD.n77 1084.97
R18154 VDD.n80 VDD.n79 1084.97
R18155 VDD.n131 VDD.n79 1084.97
R18156 VDD.n138 VDD.n73 1084.97
R18157 VDD.n142 VDD.n74 1084.97
R18158 VDD.n142 VDD.n73 1084.97
R18159 VDD.n145 VDD.n68 1084.97
R18160 VDD.n71 VDD.n70 1084.97
R18161 VDD.n145 VDD.n70 1084.97
R18162 VDD.n152 VDD.n60 1084.97
R18163 VDD.n156 VDD.n61 1084.97
R18164 VDD.n156 VDD.n60 1084.97
R18165 VDD.n159 VDD.n57 1084.97
R18166 VDD.n159 VDD.n58 1084.97
R18167 VDD.n163 VDD.n58 1084.97
R18168 VDD.n163 VDD.n57 1084.97
R18169 VDD.n166 VDD.n52 1084.97
R18170 VDD.n55 VDD.n54 1084.97
R18171 VDD.n166 VDD.n54 1084.97
R18172 VDD.n173 VDD.n48 1084.97
R18173 VDD.n177 VDD.n49 1084.97
R18174 VDD.n177 VDD.n48 1084.97
R18175 VDD.n180 VDD.n43 1084.97
R18176 VDD.n46 VDD.n45 1084.97
R18177 VDD.n180 VDD.n45 1084.97
R18178 VDD.n187 VDD.n35 1084.97
R18179 VDD.n191 VDD.n36 1084.97
R18180 VDD.n191 VDD.n35 1084.97
R18181 VDD.n194 VDD.n32 1084.97
R18182 VDD.n194 VDD.n33 1084.97
R18183 VDD.n198 VDD.n33 1084.97
R18184 VDD.n198 VDD.n32 1084.97
R18185 VDD.n201 VDD.n27 1084.97
R18186 VDD.n30 VDD.n29 1084.97
R18187 VDD.n201 VDD.n29 1084.97
R18188 VDD.n208 VDD.n23 1084.97
R18189 VDD.n212 VDD.n24 1084.97
R18190 VDD.n212 VDD.n23 1084.97
R18191 VDD.n215 VDD.n18 1084.97
R18192 VDD.n21 VDD.n20 1084.97
R18193 VDD.n215 VDD.n20 1084.97
R18194 VDD.n222 VDD.n10 1084.97
R18195 VDD.n226 VDD.n11 1084.97
R18196 VDD.n226 VDD.n10 1084.97
R18197 VDD.n229 VDD.n7 1084.97
R18198 VDD.n229 VDD.n8 1084.97
R18199 VDD.n233 VDD.n8 1084.97
R18200 VDD.n233 VDD.n7 1084.97
R18201 VDD.n236 VDD.n2 1084.97
R18202 VDD.n5 VDD.n4 1084.97
R18203 VDD.n236 VDD.n4 1084.97
R18204 VDD.n7335 VDD.n7322 1084.97
R18205 VDD.n7335 VDD.n7323 1084.97
R18206 VDD.n7342 VDD.n7323 1084.97
R18207 VDD.n7342 VDD.n7322 1084.97
R18208 VDD.n7345 VDD.n7312 1084.97
R18209 VDD.n7345 VDD.n7313 1084.97
R18210 VDD.n7352 VDD.n7313 1084.97
R18211 VDD.n7352 VDD.n7312 1084.97
R18212 VDD.n7355 VDD.n7301 1084.97
R18213 VDD.n7355 VDD.n7302 1084.97
R18214 VDD.n7362 VDD.n7302 1084.97
R18215 VDD.n7362 VDD.n7301 1084.97
R18216 VDD.n7365 VDD.n7288 1084.97
R18217 VDD.n7365 VDD.n7289 1084.97
R18218 VDD.n7372 VDD.n7289 1084.97
R18219 VDD.n7372 VDD.n7288 1084.97
R18220 VDD.n7375 VDD.n7276 1084.97
R18221 VDD.n7375 VDD.n7277 1084.97
R18222 VDD.n7382 VDD.n7277 1084.97
R18223 VDD.n7382 VDD.n7276 1084.97
R18224 VDD.n7392 VDD.n7260 1084.97
R18225 VDD.n7392 VDD.n7261 1084.97
R18226 VDD.n7399 VDD.n7261 1084.97
R18227 VDD.n7399 VDD.n7260 1084.97
R18228 VDD.n7402 VDD.n7250 1084.97
R18229 VDD.n7402 VDD.n7251 1084.97
R18230 VDD.n7409 VDD.n7251 1084.97
R18231 VDD.n7409 VDD.n7250 1084.97
R18232 VDD.n7412 VDD.n7239 1084.97
R18233 VDD.n7412 VDD.n7240 1084.97
R18234 VDD.n7419 VDD.n7240 1084.97
R18235 VDD.n7419 VDD.n7239 1084.97
R18236 VDD.n7422 VDD.n7226 1084.97
R18237 VDD.n7422 VDD.n7227 1084.97
R18238 VDD.n7429 VDD.n7227 1084.97
R18239 VDD.n7429 VDD.n7226 1084.97
R18240 VDD.n7432 VDD.n7216 1084.97
R18241 VDD.n7432 VDD.n7217 1084.97
R18242 VDD.n7439 VDD.n7217 1084.97
R18243 VDD.n7439 VDD.n7216 1084.97
R18244 VDD.n7442 VDD.n7205 1084.97
R18245 VDD.n7442 VDD.n7206 1084.97
R18246 VDD.n7449 VDD.n7206 1084.97
R18247 VDD.n7449 VDD.n7205 1084.97
R18248 VDD.n7338 VDD.n7337 1084.97
R18249 VDD.n7337 VDD.n7331 1084.97
R18250 VDD.n7331 VDD.n7321 1084.97
R18251 VDD.n7338 VDD.n7321 1084.97
R18252 VDD.n7348 VDD.n7347 1084.97
R18253 VDD.n7347 VDD.n7318 1084.97
R18254 VDD.n7318 VDD.n7311 1084.97
R18255 VDD.n7348 VDD.n7311 1084.97
R18256 VDD.n7358 VDD.n7357 1084.97
R18257 VDD.n7357 VDD.n7308 1084.97
R18258 VDD.n7308 VDD.n7300 1084.97
R18259 VDD.n7358 VDD.n7300 1084.97
R18260 VDD.n7368 VDD.n7367 1084.97
R18261 VDD.n7367 VDD.n7297 1084.97
R18262 VDD.n7297 VDD.n7287 1084.97
R18263 VDD.n7368 VDD.n7287 1084.97
R18264 VDD.n7378 VDD.n7377 1084.97
R18265 VDD.n7377 VDD.n7284 1084.97
R18266 VDD.n7284 VDD.n7275 1084.97
R18267 VDD.n7378 VDD.n7275 1084.97
R18268 VDD.n7385 VDD.n7272 1084.97
R18269 VDD.n7385 VDD.n7273 1084.97
R18270 VDD.n7389 VDD.n7273 1084.97
R18271 VDD.n7389 VDD.n7272 1084.97
R18272 VDD.n7395 VDD.n7394 1084.97
R18273 VDD.n7394 VDD.n7269 1084.97
R18274 VDD.n7269 VDD.n7259 1084.97
R18275 VDD.n7395 VDD.n7259 1084.97
R18276 VDD.n7405 VDD.n7404 1084.97
R18277 VDD.n7404 VDD.n7256 1084.97
R18278 VDD.n7256 VDD.n7249 1084.97
R18279 VDD.n7405 VDD.n7249 1084.97
R18280 VDD.n7415 VDD.n7414 1084.97
R18281 VDD.n7414 VDD.n7246 1084.97
R18282 VDD.n7246 VDD.n7238 1084.97
R18283 VDD.n7415 VDD.n7238 1084.97
R18284 VDD.n7425 VDD.n7424 1084.97
R18285 VDD.n7424 VDD.n7235 1084.97
R18286 VDD.n7235 VDD.n7225 1084.97
R18287 VDD.n7425 VDD.n7225 1084.97
R18288 VDD.n7435 VDD.n7434 1084.97
R18289 VDD.n7434 VDD.n7222 1084.97
R18290 VDD.n7222 VDD.n7215 1084.97
R18291 VDD.n7435 VDD.n7215 1084.97
R18292 VDD.n7445 VDD.n7444 1084.97
R18293 VDD.n7444 VDD.n7212 1084.97
R18294 VDD.n7212 VDD.n7204 1084.97
R18295 VDD.n7445 VDD.n7204 1084.97
R18296 VDD.n7202 VDD.n7201 1084.97
R18297 VDD.n7452 VDD.n7201 1084.97
R18298 VDD.n7452 VDD.n7199 1084.97
R18299 VDD.n7078 VDD.n1971 1084.97
R18300 VDD.n7078 VDD.n1972 1084.97
R18301 VDD.n7085 VDD.n1972 1084.97
R18302 VDD.n7085 VDD.n1971 1084.97
R18303 VDD.n7088 VDD.n1961 1084.97
R18304 VDD.n7088 VDD.n1962 1084.97
R18305 VDD.n7095 VDD.n1962 1084.97
R18306 VDD.n7095 VDD.n1961 1084.97
R18307 VDD.n7098 VDD.n1950 1084.97
R18308 VDD.n7098 VDD.n1951 1084.97
R18309 VDD.n7105 VDD.n1951 1084.97
R18310 VDD.n7105 VDD.n1950 1084.97
R18311 VDD.n7108 VDD.n1937 1084.97
R18312 VDD.n7108 VDD.n1938 1084.97
R18313 VDD.n7115 VDD.n1938 1084.97
R18314 VDD.n7115 VDD.n1937 1084.97
R18315 VDD.n7118 VDD.n1925 1084.97
R18316 VDD.n7118 VDD.n1926 1084.97
R18317 VDD.n7125 VDD.n1926 1084.97
R18318 VDD.n7125 VDD.n1925 1084.97
R18319 VDD.n7140 VDD.n7136 1084.97
R18320 VDD.n7136 VDD.n1905 1084.97
R18321 VDD.n7135 VDD.n1905 1084.97
R18322 VDD.n7140 VDD.n7135 1084.97
R18323 VDD.n7152 VDD.n1883 1084.97
R18324 VDD.n7152 VDD.n1884 1084.97
R18325 VDD.n7159 VDD.n1884 1084.97
R18326 VDD.n7159 VDD.n1883 1084.97
R18327 VDD.n7162 VDD.n1870 1084.97
R18328 VDD.n7162 VDD.n1871 1084.97
R18329 VDD.n7169 VDD.n1871 1084.97
R18330 VDD.n7169 VDD.n1870 1084.97
R18331 VDD.n7172 VDD.n1860 1084.97
R18332 VDD.n7172 VDD.n1861 1084.97
R18333 VDD.n7179 VDD.n1861 1084.97
R18334 VDD.n7179 VDD.n1860 1084.97
R18335 VDD.n7182 VDD.n1849 1084.97
R18336 VDD.n7182 VDD.n1850 1084.97
R18337 VDD.n7189 VDD.n1850 1084.97
R18338 VDD.n7189 VDD.n1849 1084.97
R18339 VDD.n7192 VDD.n1845 1084.97
R18340 VDD.n7192 VDD.n1843 1084.97
R18341 VDD.n1846 VDD.n1845 1084.97
R18342 VDD.n7081 VDD.n7080 1084.97
R18343 VDD.n7080 VDD.n7074 1084.97
R18344 VDD.n7074 VDD.n1970 1084.97
R18345 VDD.n7081 VDD.n1970 1084.97
R18346 VDD.n7091 VDD.n7090 1084.97
R18347 VDD.n7090 VDD.n1967 1084.97
R18348 VDD.n1967 VDD.n1960 1084.97
R18349 VDD.n7091 VDD.n1960 1084.97
R18350 VDD.n7101 VDD.n7100 1084.97
R18351 VDD.n7100 VDD.n1957 1084.97
R18352 VDD.n1957 VDD.n1949 1084.97
R18353 VDD.n7101 VDD.n1949 1084.97
R18354 VDD.n7111 VDD.n7110 1084.97
R18355 VDD.n7110 VDD.n1946 1084.97
R18356 VDD.n1946 VDD.n1936 1084.97
R18357 VDD.n7111 VDD.n1936 1084.97
R18358 VDD.n7121 VDD.n7120 1084.97
R18359 VDD.n7120 VDD.n1933 1084.97
R18360 VDD.n1933 VDD.n1924 1084.97
R18361 VDD.n7121 VDD.n1924 1084.97
R18362 VDD.n7128 VDD.n1921 1084.97
R18363 VDD.n7128 VDD.n1922 1084.97
R18364 VDD.n7132 VDD.n1922 1084.97
R18365 VDD.n7132 VDD.n1921 1084.97
R18366 VDD.n7141 VDD.n1908 1084.97
R18367 VDD.n1920 VDD.n1908 1084.97
R18368 VDD.n1920 VDD.n1907 1084.97
R18369 VDD.n7141 VDD.n1907 1084.97
R18370 VDD.n1900 VDD.n1894 1084.97
R18371 VDD.n1912 VDD.n1900 1084.97
R18372 VDD.n1912 VDD.n1909 1084.97
R18373 VDD.n1909 VDD.n1894 1084.97
R18374 VDD.n7155 VDD.n7154 1084.97
R18375 VDD.n7154 VDD.n1891 1084.97
R18376 VDD.n1891 VDD.n1882 1084.97
R18377 VDD.n7155 VDD.n1882 1084.97
R18378 VDD.n7165 VDD.n7164 1084.97
R18379 VDD.n7164 VDD.n1879 1084.97
R18380 VDD.n1879 VDD.n1869 1084.97
R18381 VDD.n7165 VDD.n1869 1084.97
R18382 VDD.n7175 VDD.n7174 1084.97
R18383 VDD.n7174 VDD.n1866 1084.97
R18384 VDD.n1866 VDD.n1859 1084.97
R18385 VDD.n7175 VDD.n1859 1084.97
R18386 VDD.n7185 VDD.n7184 1084.97
R18387 VDD.n7184 VDD.n1856 1084.97
R18388 VDD.n1856 VDD.n1848 1084.97
R18389 VDD.n7185 VDD.n1848 1084.97
R18390 VDD.n7149 VDD.n1895 1084.97
R18391 VDD.n1914 VDD.n1895 1084.97
R18392 VDD.n7149 VDD.n1896 1084.97
R18393 VDD.n1914 VDD.n1896 1084.97
R18394 VDD.n7056 VDD.n6847 1084.97
R18395 VDD.n7060 VDD.n6848 1084.97
R18396 VDD.n7060 VDD.n6847 1084.97
R18397 VDD.n7065 VDD.n6834 1084.97
R18398 VDD.n7064 VDD.n6834 1084.97
R18399 VDD.n7064 VDD.n6833 1084.97
R18400 VDD.n7065 VDD.n6833 1084.97
R18401 VDD.n6937 VDD.n6932 1084.97
R18402 VDD.n6941 VDD.n6933 1084.97
R18403 VDD.n6941 VDD.n6932 1084.97
R18404 VDD.n6944 VDD.n6927 1084.97
R18405 VDD.n6930 VDD.n6929 1084.97
R18406 VDD.n6944 VDD.n6929 1084.97
R18407 VDD.n6951 VDD.n6919 1084.97
R18408 VDD.n6955 VDD.n6920 1084.97
R18409 VDD.n6955 VDD.n6919 1084.97
R18410 VDD.n6958 VDD.n6916 1084.97
R18411 VDD.n6958 VDD.n6917 1084.97
R18412 VDD.n6962 VDD.n6917 1084.97
R18413 VDD.n6962 VDD.n6916 1084.97
R18414 VDD.n6965 VDD.n6911 1084.97
R18415 VDD.n6914 VDD.n6913 1084.97
R18416 VDD.n6965 VDD.n6913 1084.97
R18417 VDD.n6972 VDD.n6907 1084.97
R18418 VDD.n6976 VDD.n6908 1084.97
R18419 VDD.n6976 VDD.n6907 1084.97
R18420 VDD.n6979 VDD.n6902 1084.97
R18421 VDD.n6905 VDD.n6904 1084.97
R18422 VDD.n6979 VDD.n6904 1084.97
R18423 VDD.n6986 VDD.n6894 1084.97
R18424 VDD.n6990 VDD.n6895 1084.97
R18425 VDD.n6990 VDD.n6894 1084.97
R18426 VDD.n6993 VDD.n6891 1084.97
R18427 VDD.n6993 VDD.n6892 1084.97
R18428 VDD.n6997 VDD.n6892 1084.97
R18429 VDD.n6997 VDD.n6891 1084.97
R18430 VDD.n7000 VDD.n6886 1084.97
R18431 VDD.n6889 VDD.n6888 1084.97
R18432 VDD.n7000 VDD.n6888 1084.97
R18433 VDD.n7007 VDD.n6882 1084.97
R18434 VDD.n7011 VDD.n6883 1084.97
R18435 VDD.n7011 VDD.n6882 1084.97
R18436 VDD.n7014 VDD.n6877 1084.97
R18437 VDD.n6880 VDD.n6879 1084.97
R18438 VDD.n7014 VDD.n6879 1084.97
R18439 VDD.n7021 VDD.n6869 1084.97
R18440 VDD.n7025 VDD.n6870 1084.97
R18441 VDD.n7025 VDD.n6869 1084.97
R18442 VDD.n7028 VDD.n6866 1084.97
R18443 VDD.n7028 VDD.n6867 1084.97
R18444 VDD.n7032 VDD.n6867 1084.97
R18445 VDD.n7032 VDD.n6866 1084.97
R18446 VDD.n7035 VDD.n6861 1084.97
R18447 VDD.n6864 VDD.n6863 1084.97
R18448 VDD.n7035 VDD.n6863 1084.97
R18449 VDD.n7042 VDD.n6857 1084.97
R18450 VDD.n7046 VDD.n6858 1084.97
R18451 VDD.n7046 VDD.n6857 1084.97
R18452 VDD.n7049 VDD.n6852 1084.97
R18453 VDD.n6855 VDD.n6854 1084.97
R18454 VDD.n7049 VDD.n6854 1084.97
R18455 VDD.n6844 VDD.n6835 1084.97
R18456 VDD.n6840 VDD.n6836 1084.97
R18457 VDD.n6844 VDD.n6836 1084.97
R18458 VDD.n5963 VDD.n5959 1084.97
R18459 VDD.n5970 VDD.n5960 1084.97
R18460 VDD.n5970 VDD.n5959 1084.97
R18461 VDD.n5973 VDD.n5950 1084.97
R18462 VDD.n5973 VDD.n5951 1084.97
R18463 VDD.n5980 VDD.n5951 1084.97
R18464 VDD.n5980 VDD.n5950 1084.97
R18465 VDD.n5983 VDD.n5937 1084.97
R18466 VDD.n5983 VDD.n5938 1084.97
R18467 VDD.n5990 VDD.n5938 1084.97
R18468 VDD.n5990 VDD.n5937 1084.97
R18469 VDD.n5993 VDD.n5926 1084.97
R18470 VDD.n5993 VDD.n5927 1084.97
R18471 VDD.n6000 VDD.n5927 1084.97
R18472 VDD.n6000 VDD.n5926 1084.97
R18473 VDD.n6003 VDD.n5916 1084.97
R18474 VDD.n6003 VDD.n5917 1084.97
R18475 VDD.n6010 VDD.n5917 1084.97
R18476 VDD.n6010 VDD.n5916 1084.97
R18477 VDD.n6013 VDD.n5903 1084.97
R18478 VDD.n6013 VDD.n5904 1084.97
R18479 VDD.n6020 VDD.n5904 1084.97
R18480 VDD.n6020 VDD.n5903 1084.97
R18481 VDD.n6023 VDD.n5891 1084.97
R18482 VDD.n6023 VDD.n5892 1084.97
R18483 VDD.n6030 VDD.n5892 1084.97
R18484 VDD.n6030 VDD.n5891 1084.97
R18485 VDD.n6040 VDD.n5875 1084.97
R18486 VDD.n6040 VDD.n5876 1084.97
R18487 VDD.n6047 VDD.n5876 1084.97
R18488 VDD.n6047 VDD.n5875 1084.97
R18489 VDD.n6050 VDD.n5864 1084.97
R18490 VDD.n6050 VDD.n5865 1084.97
R18491 VDD.n6057 VDD.n5865 1084.97
R18492 VDD.n6057 VDD.n5864 1084.97
R18493 VDD.n6060 VDD.n5854 1084.97
R18494 VDD.n6060 VDD.n5855 1084.97
R18495 VDD.n6067 VDD.n5855 1084.97
R18496 VDD.n6067 VDD.n5854 1084.97
R18497 VDD.n6070 VDD.n5844 1084.97
R18498 VDD.n6070 VDD.n5845 1084.97
R18499 VDD.n6077 VDD.n5845 1084.97
R18500 VDD.n6077 VDD.n5844 1084.97
R18501 VDD.n5976 VDD.n5975 1084.97
R18502 VDD.n5975 VDD.n5956 1084.97
R18503 VDD.n5956 VDD.n5949 1084.97
R18504 VDD.n5976 VDD.n5949 1084.97
R18505 VDD.n5986 VDD.n5985 1084.97
R18506 VDD.n5985 VDD.n5946 1084.97
R18507 VDD.n5946 VDD.n5936 1084.97
R18508 VDD.n5986 VDD.n5936 1084.97
R18509 VDD.n5996 VDD.n5995 1084.97
R18510 VDD.n5995 VDD.n5933 1084.97
R18511 VDD.n5933 VDD.n5925 1084.97
R18512 VDD.n5996 VDD.n5925 1084.97
R18513 VDD.n6006 VDD.n6005 1084.97
R18514 VDD.n6005 VDD.n5922 1084.97
R18515 VDD.n5922 VDD.n5915 1084.97
R18516 VDD.n6006 VDD.n5915 1084.97
R18517 VDD.n6016 VDD.n6015 1084.97
R18518 VDD.n6015 VDD.n5912 1084.97
R18519 VDD.n5912 VDD.n5902 1084.97
R18520 VDD.n6016 VDD.n5902 1084.97
R18521 VDD.n6026 VDD.n6025 1084.97
R18522 VDD.n6025 VDD.n5899 1084.97
R18523 VDD.n5899 VDD.n5890 1084.97
R18524 VDD.n6026 VDD.n5890 1084.97
R18525 VDD.n6033 VDD.n5887 1084.97
R18526 VDD.n6033 VDD.n5888 1084.97
R18527 VDD.n6037 VDD.n5888 1084.97
R18528 VDD.n6037 VDD.n5887 1084.97
R18529 VDD.n6043 VDD.n6042 1084.97
R18530 VDD.n6042 VDD.n5884 1084.97
R18531 VDD.n5884 VDD.n5874 1084.97
R18532 VDD.n6043 VDD.n5874 1084.97
R18533 VDD.n6053 VDD.n6052 1084.97
R18534 VDD.n6052 VDD.n5871 1084.97
R18535 VDD.n5871 VDD.n5863 1084.97
R18536 VDD.n6053 VDD.n5863 1084.97
R18537 VDD.n6063 VDD.n6062 1084.97
R18538 VDD.n6062 VDD.n5860 1084.97
R18539 VDD.n5860 VDD.n5853 1084.97
R18540 VDD.n6063 VDD.n5853 1084.97
R18541 VDD.n6073 VDD.n6072 1084.97
R18542 VDD.n6072 VDD.n5850 1084.97
R18543 VDD.n5850 VDD.n5843 1084.97
R18544 VDD.n6073 VDD.n5843 1084.97
R18545 VDD.n6086 VDD.n5836 1084.97
R18546 VDD.n6086 VDD.n5837 1084.97
R18547 VDD.n5842 VDD.n5837 1084.97
R18548 VDD.n5842 VDD.n5836 1084.97
R18549 VDD.n6085 VDD.n6080 1084.97
R18550 VDD.n6085 VDD.n6081 1084.97
R18551 VDD.n6080 VDD.n5834 1084.97
R18552 VDD.n6081 VDD.n5834 1084.97
R18553 VDD.n5827 VDD.n5823 1084.97
R18554 VDD.n6093 VDD.n5824 1084.97
R18555 VDD.n6093 VDD.n5823 1084.97
R18556 VDD.n6096 VDD.n5814 1084.97
R18557 VDD.n6096 VDD.n5815 1084.97
R18558 VDD.n6103 VDD.n5815 1084.97
R18559 VDD.n6103 VDD.n5814 1084.97
R18560 VDD.n6106 VDD.n5801 1084.97
R18561 VDD.n6106 VDD.n5802 1084.97
R18562 VDD.n6113 VDD.n5802 1084.97
R18563 VDD.n6113 VDD.n5801 1084.97
R18564 VDD.n6116 VDD.n5790 1084.97
R18565 VDD.n6116 VDD.n5791 1084.97
R18566 VDD.n6123 VDD.n5791 1084.97
R18567 VDD.n6123 VDD.n5790 1084.97
R18568 VDD.n6126 VDD.n5780 1084.97
R18569 VDD.n6126 VDD.n5781 1084.97
R18570 VDD.n6133 VDD.n5781 1084.97
R18571 VDD.n6133 VDD.n5780 1084.97
R18572 VDD.n6136 VDD.n5767 1084.97
R18573 VDD.n6136 VDD.n5768 1084.97
R18574 VDD.n6143 VDD.n5768 1084.97
R18575 VDD.n6143 VDD.n5767 1084.97
R18576 VDD.n6146 VDD.n5755 1084.97
R18577 VDD.n6146 VDD.n5756 1084.97
R18578 VDD.n6153 VDD.n5756 1084.97
R18579 VDD.n6153 VDD.n5755 1084.97
R18580 VDD.n6163 VDD.n5739 1084.97
R18581 VDD.n6163 VDD.n5740 1084.97
R18582 VDD.n6170 VDD.n5740 1084.97
R18583 VDD.n6170 VDD.n5739 1084.97
R18584 VDD.n6173 VDD.n5728 1084.97
R18585 VDD.n6173 VDD.n5729 1084.97
R18586 VDD.n6180 VDD.n5729 1084.97
R18587 VDD.n6180 VDD.n5728 1084.97
R18588 VDD.n6183 VDD.n5718 1084.97
R18589 VDD.n6183 VDD.n5719 1084.97
R18590 VDD.n6190 VDD.n5719 1084.97
R18591 VDD.n6190 VDD.n5718 1084.97
R18592 VDD.n6193 VDD.n5708 1084.97
R18593 VDD.n6193 VDD.n5709 1084.97
R18594 VDD.n6200 VDD.n5709 1084.97
R18595 VDD.n6200 VDD.n5708 1084.97
R18596 VDD.n6099 VDD.n6098 1084.97
R18597 VDD.n6098 VDD.n5820 1084.97
R18598 VDD.n5820 VDD.n5813 1084.97
R18599 VDD.n6099 VDD.n5813 1084.97
R18600 VDD.n6109 VDD.n6108 1084.97
R18601 VDD.n6108 VDD.n5810 1084.97
R18602 VDD.n5810 VDD.n5800 1084.97
R18603 VDD.n6109 VDD.n5800 1084.97
R18604 VDD.n6119 VDD.n6118 1084.97
R18605 VDD.n6118 VDD.n5797 1084.97
R18606 VDD.n5797 VDD.n5789 1084.97
R18607 VDD.n6119 VDD.n5789 1084.97
R18608 VDD.n6129 VDD.n6128 1084.97
R18609 VDD.n6128 VDD.n5786 1084.97
R18610 VDD.n5786 VDD.n5779 1084.97
R18611 VDD.n6129 VDD.n5779 1084.97
R18612 VDD.n6139 VDD.n6138 1084.97
R18613 VDD.n6138 VDD.n5776 1084.97
R18614 VDD.n5776 VDD.n5766 1084.97
R18615 VDD.n6139 VDD.n5766 1084.97
R18616 VDD.n6149 VDD.n6148 1084.97
R18617 VDD.n6148 VDD.n5763 1084.97
R18618 VDD.n5763 VDD.n5754 1084.97
R18619 VDD.n6149 VDD.n5754 1084.97
R18620 VDD.n6156 VDD.n5751 1084.97
R18621 VDD.n6156 VDD.n5752 1084.97
R18622 VDD.n6160 VDD.n5752 1084.97
R18623 VDD.n6160 VDD.n5751 1084.97
R18624 VDD.n6166 VDD.n6165 1084.97
R18625 VDD.n6165 VDD.n5748 1084.97
R18626 VDD.n5748 VDD.n5738 1084.97
R18627 VDD.n6166 VDD.n5738 1084.97
R18628 VDD.n6176 VDD.n6175 1084.97
R18629 VDD.n6175 VDD.n5735 1084.97
R18630 VDD.n5735 VDD.n5727 1084.97
R18631 VDD.n6176 VDD.n5727 1084.97
R18632 VDD.n6186 VDD.n6185 1084.97
R18633 VDD.n6185 VDD.n5724 1084.97
R18634 VDD.n5724 VDD.n5717 1084.97
R18635 VDD.n6186 VDD.n5717 1084.97
R18636 VDD.n6196 VDD.n6195 1084.97
R18637 VDD.n6195 VDD.n5714 1084.97
R18638 VDD.n5714 VDD.n5707 1084.97
R18639 VDD.n6196 VDD.n5707 1084.97
R18640 VDD.n6209 VDD.n5700 1084.97
R18641 VDD.n6209 VDD.n5701 1084.97
R18642 VDD.n5706 VDD.n5701 1084.97
R18643 VDD.n5706 VDD.n5700 1084.97
R18644 VDD.n6208 VDD.n6203 1084.97
R18645 VDD.n6208 VDD.n6204 1084.97
R18646 VDD.n6203 VDD.n5698 1084.97
R18647 VDD.n6204 VDD.n5698 1084.97
R18648 VDD.n5691 VDD.n5687 1084.97
R18649 VDD.n6216 VDD.n5688 1084.97
R18650 VDD.n6216 VDD.n5687 1084.97
R18651 VDD.n6219 VDD.n5678 1084.97
R18652 VDD.n6219 VDD.n5679 1084.97
R18653 VDD.n6226 VDD.n5679 1084.97
R18654 VDD.n6226 VDD.n5678 1084.97
R18655 VDD.n6229 VDD.n5665 1084.97
R18656 VDD.n6229 VDD.n5666 1084.97
R18657 VDD.n6236 VDD.n5666 1084.97
R18658 VDD.n6236 VDD.n5665 1084.97
R18659 VDD.n6239 VDD.n5654 1084.97
R18660 VDD.n6239 VDD.n5655 1084.97
R18661 VDD.n6246 VDD.n5655 1084.97
R18662 VDD.n6246 VDD.n5654 1084.97
R18663 VDD.n6249 VDD.n5644 1084.97
R18664 VDD.n6249 VDD.n5645 1084.97
R18665 VDD.n6256 VDD.n5645 1084.97
R18666 VDD.n6256 VDD.n5644 1084.97
R18667 VDD.n6259 VDD.n5631 1084.97
R18668 VDD.n6259 VDD.n5632 1084.97
R18669 VDD.n6266 VDD.n5632 1084.97
R18670 VDD.n6266 VDD.n5631 1084.97
R18671 VDD.n6269 VDD.n5619 1084.97
R18672 VDD.n6269 VDD.n5620 1084.97
R18673 VDD.n6276 VDD.n5620 1084.97
R18674 VDD.n6276 VDD.n5619 1084.97
R18675 VDD.n6286 VDD.n5603 1084.97
R18676 VDD.n6286 VDD.n5604 1084.97
R18677 VDD.n6293 VDD.n5604 1084.97
R18678 VDD.n6293 VDD.n5603 1084.97
R18679 VDD.n6296 VDD.n5592 1084.97
R18680 VDD.n6296 VDD.n5593 1084.97
R18681 VDD.n6303 VDD.n5593 1084.97
R18682 VDD.n6303 VDD.n5592 1084.97
R18683 VDD.n6306 VDD.n5582 1084.97
R18684 VDD.n6306 VDD.n5583 1084.97
R18685 VDD.n6313 VDD.n5583 1084.97
R18686 VDD.n6313 VDD.n5582 1084.97
R18687 VDD.n6316 VDD.n5572 1084.97
R18688 VDD.n6316 VDD.n5573 1084.97
R18689 VDD.n6323 VDD.n5573 1084.97
R18690 VDD.n6323 VDD.n5572 1084.97
R18691 VDD.n6222 VDD.n6221 1084.97
R18692 VDD.n6221 VDD.n5684 1084.97
R18693 VDD.n5684 VDD.n5677 1084.97
R18694 VDD.n6222 VDD.n5677 1084.97
R18695 VDD.n6232 VDD.n6231 1084.97
R18696 VDD.n6231 VDD.n5674 1084.97
R18697 VDD.n5674 VDD.n5664 1084.97
R18698 VDD.n6232 VDD.n5664 1084.97
R18699 VDD.n6242 VDD.n6241 1084.97
R18700 VDD.n6241 VDD.n5661 1084.97
R18701 VDD.n5661 VDD.n5653 1084.97
R18702 VDD.n6242 VDD.n5653 1084.97
R18703 VDD.n6252 VDD.n6251 1084.97
R18704 VDD.n6251 VDD.n5650 1084.97
R18705 VDD.n5650 VDD.n5643 1084.97
R18706 VDD.n6252 VDD.n5643 1084.97
R18707 VDD.n6262 VDD.n6261 1084.97
R18708 VDD.n6261 VDD.n5640 1084.97
R18709 VDD.n5640 VDD.n5630 1084.97
R18710 VDD.n6262 VDD.n5630 1084.97
R18711 VDD.n6272 VDD.n6271 1084.97
R18712 VDD.n6271 VDD.n5627 1084.97
R18713 VDD.n5627 VDD.n5618 1084.97
R18714 VDD.n6272 VDD.n5618 1084.97
R18715 VDD.n6279 VDD.n5615 1084.97
R18716 VDD.n6279 VDD.n5616 1084.97
R18717 VDD.n6283 VDD.n5616 1084.97
R18718 VDD.n6283 VDD.n5615 1084.97
R18719 VDD.n6289 VDD.n6288 1084.97
R18720 VDD.n6288 VDD.n5612 1084.97
R18721 VDD.n5612 VDD.n5602 1084.97
R18722 VDD.n6289 VDD.n5602 1084.97
R18723 VDD.n6299 VDD.n6298 1084.97
R18724 VDD.n6298 VDD.n5599 1084.97
R18725 VDD.n5599 VDD.n5591 1084.97
R18726 VDD.n6299 VDD.n5591 1084.97
R18727 VDD.n6309 VDD.n6308 1084.97
R18728 VDD.n6308 VDD.n5588 1084.97
R18729 VDD.n5588 VDD.n5581 1084.97
R18730 VDD.n6309 VDD.n5581 1084.97
R18731 VDD.n6319 VDD.n6318 1084.97
R18732 VDD.n6318 VDD.n5578 1084.97
R18733 VDD.n5578 VDD.n5571 1084.97
R18734 VDD.n6319 VDD.n5571 1084.97
R18735 VDD.n6332 VDD.n5564 1084.97
R18736 VDD.n6332 VDD.n5565 1084.97
R18737 VDD.n5570 VDD.n5565 1084.97
R18738 VDD.n5570 VDD.n5564 1084.97
R18739 VDD.n6331 VDD.n6326 1084.97
R18740 VDD.n6331 VDD.n6327 1084.97
R18741 VDD.n6326 VDD.n5562 1084.97
R18742 VDD.n6327 VDD.n5562 1084.97
R18743 VDD.n5555 VDD.n5551 1084.97
R18744 VDD.n6339 VDD.n5552 1084.97
R18745 VDD.n6339 VDD.n5551 1084.97
R18746 VDD.n6342 VDD.n5542 1084.97
R18747 VDD.n6342 VDD.n5543 1084.97
R18748 VDD.n6349 VDD.n5543 1084.97
R18749 VDD.n6349 VDD.n5542 1084.97
R18750 VDD.n6352 VDD.n5529 1084.97
R18751 VDD.n6352 VDD.n5530 1084.97
R18752 VDD.n6359 VDD.n5530 1084.97
R18753 VDD.n6359 VDD.n5529 1084.97
R18754 VDD.n6362 VDD.n5518 1084.97
R18755 VDD.n6362 VDD.n5519 1084.97
R18756 VDD.n6369 VDD.n5519 1084.97
R18757 VDD.n6369 VDD.n5518 1084.97
R18758 VDD.n6372 VDD.n5508 1084.97
R18759 VDD.n6372 VDD.n5509 1084.97
R18760 VDD.n6379 VDD.n5509 1084.97
R18761 VDD.n6379 VDD.n5508 1084.97
R18762 VDD.n6382 VDD.n5495 1084.97
R18763 VDD.n6382 VDD.n5496 1084.97
R18764 VDD.n6389 VDD.n5496 1084.97
R18765 VDD.n6389 VDD.n5495 1084.97
R18766 VDD.n6392 VDD.n5483 1084.97
R18767 VDD.n6392 VDD.n5484 1084.97
R18768 VDD.n6399 VDD.n5484 1084.97
R18769 VDD.n6399 VDD.n5483 1084.97
R18770 VDD.n6409 VDD.n5467 1084.97
R18771 VDD.n6409 VDD.n5468 1084.97
R18772 VDD.n6416 VDD.n5468 1084.97
R18773 VDD.n6416 VDD.n5467 1084.97
R18774 VDD.n6419 VDD.n5456 1084.97
R18775 VDD.n6419 VDD.n5457 1084.97
R18776 VDD.n6426 VDD.n5457 1084.97
R18777 VDD.n6426 VDD.n5456 1084.97
R18778 VDD.n6429 VDD.n5446 1084.97
R18779 VDD.n6429 VDD.n5447 1084.97
R18780 VDD.n6436 VDD.n5447 1084.97
R18781 VDD.n6436 VDD.n5446 1084.97
R18782 VDD.n6439 VDD.n5436 1084.97
R18783 VDD.n6439 VDD.n5437 1084.97
R18784 VDD.n6446 VDD.n5437 1084.97
R18785 VDD.n6446 VDD.n5436 1084.97
R18786 VDD.n6345 VDD.n6344 1084.97
R18787 VDD.n6344 VDD.n5548 1084.97
R18788 VDD.n5548 VDD.n5541 1084.97
R18789 VDD.n6345 VDD.n5541 1084.97
R18790 VDD.n6355 VDD.n6354 1084.97
R18791 VDD.n6354 VDD.n5538 1084.97
R18792 VDD.n5538 VDD.n5528 1084.97
R18793 VDD.n6355 VDD.n5528 1084.97
R18794 VDD.n6365 VDD.n6364 1084.97
R18795 VDD.n6364 VDD.n5525 1084.97
R18796 VDD.n5525 VDD.n5517 1084.97
R18797 VDD.n6365 VDD.n5517 1084.97
R18798 VDD.n6375 VDD.n6374 1084.97
R18799 VDD.n6374 VDD.n5514 1084.97
R18800 VDD.n5514 VDD.n5507 1084.97
R18801 VDD.n6375 VDD.n5507 1084.97
R18802 VDD.n6385 VDD.n6384 1084.97
R18803 VDD.n6384 VDD.n5504 1084.97
R18804 VDD.n5504 VDD.n5494 1084.97
R18805 VDD.n6385 VDD.n5494 1084.97
R18806 VDD.n6395 VDD.n6394 1084.97
R18807 VDD.n6394 VDD.n5491 1084.97
R18808 VDD.n5491 VDD.n5482 1084.97
R18809 VDD.n6395 VDD.n5482 1084.97
R18810 VDD.n6402 VDD.n5479 1084.97
R18811 VDD.n6402 VDD.n5480 1084.97
R18812 VDD.n6406 VDD.n5480 1084.97
R18813 VDD.n6406 VDD.n5479 1084.97
R18814 VDD.n6412 VDD.n6411 1084.97
R18815 VDD.n6411 VDD.n5476 1084.97
R18816 VDD.n5476 VDD.n5466 1084.97
R18817 VDD.n6412 VDD.n5466 1084.97
R18818 VDD.n6422 VDD.n6421 1084.97
R18819 VDD.n6421 VDD.n5463 1084.97
R18820 VDD.n5463 VDD.n5455 1084.97
R18821 VDD.n6422 VDD.n5455 1084.97
R18822 VDD.n6432 VDD.n6431 1084.97
R18823 VDD.n6431 VDD.n5452 1084.97
R18824 VDD.n5452 VDD.n5445 1084.97
R18825 VDD.n6432 VDD.n5445 1084.97
R18826 VDD.n6442 VDD.n6441 1084.97
R18827 VDD.n6441 VDD.n5442 1084.97
R18828 VDD.n5442 VDD.n5435 1084.97
R18829 VDD.n6442 VDD.n5435 1084.97
R18830 VDD.n6455 VDD.n5428 1084.97
R18831 VDD.n6455 VDD.n5429 1084.97
R18832 VDD.n5434 VDD.n5429 1084.97
R18833 VDD.n5434 VDD.n5428 1084.97
R18834 VDD.n6454 VDD.n6449 1084.97
R18835 VDD.n6454 VDD.n6450 1084.97
R18836 VDD.n6449 VDD.n5426 1084.97
R18837 VDD.n6450 VDD.n5426 1084.97
R18838 VDD.n5419 VDD.n5415 1084.97
R18839 VDD.n6462 VDD.n5416 1084.97
R18840 VDD.n6462 VDD.n5415 1084.97
R18841 VDD.n6465 VDD.n5406 1084.97
R18842 VDD.n6465 VDD.n5407 1084.97
R18843 VDD.n6472 VDD.n5407 1084.97
R18844 VDD.n6472 VDD.n5406 1084.97
R18845 VDD.n6475 VDD.n5393 1084.97
R18846 VDD.n6475 VDD.n5394 1084.97
R18847 VDD.n6482 VDD.n5394 1084.97
R18848 VDD.n6482 VDD.n5393 1084.97
R18849 VDD.n6485 VDD.n5382 1084.97
R18850 VDD.n6485 VDD.n5383 1084.97
R18851 VDD.n6492 VDD.n5383 1084.97
R18852 VDD.n6492 VDD.n5382 1084.97
R18853 VDD.n6495 VDD.n5372 1084.97
R18854 VDD.n6495 VDD.n5373 1084.97
R18855 VDD.n6502 VDD.n5373 1084.97
R18856 VDD.n6502 VDD.n5372 1084.97
R18857 VDD.n6505 VDD.n5359 1084.97
R18858 VDD.n6505 VDD.n5360 1084.97
R18859 VDD.n6512 VDD.n5360 1084.97
R18860 VDD.n6512 VDD.n5359 1084.97
R18861 VDD.n6515 VDD.n5347 1084.97
R18862 VDD.n6515 VDD.n5348 1084.97
R18863 VDD.n6522 VDD.n5348 1084.97
R18864 VDD.n6522 VDD.n5347 1084.97
R18865 VDD.n6532 VDD.n5331 1084.97
R18866 VDD.n6532 VDD.n5332 1084.97
R18867 VDD.n6539 VDD.n5332 1084.97
R18868 VDD.n6539 VDD.n5331 1084.97
R18869 VDD.n6542 VDD.n5320 1084.97
R18870 VDD.n6542 VDD.n5321 1084.97
R18871 VDD.n6549 VDD.n5321 1084.97
R18872 VDD.n6549 VDD.n5320 1084.97
R18873 VDD.n6552 VDD.n5310 1084.97
R18874 VDD.n6552 VDD.n5311 1084.97
R18875 VDD.n6559 VDD.n5311 1084.97
R18876 VDD.n6559 VDD.n5310 1084.97
R18877 VDD.n6562 VDD.n5300 1084.97
R18878 VDD.n6562 VDD.n5301 1084.97
R18879 VDD.n6569 VDD.n5301 1084.97
R18880 VDD.n6569 VDD.n5300 1084.97
R18881 VDD.n6468 VDD.n6467 1084.97
R18882 VDD.n6467 VDD.n5412 1084.97
R18883 VDD.n5412 VDD.n5405 1084.97
R18884 VDD.n6468 VDD.n5405 1084.97
R18885 VDD.n6478 VDD.n6477 1084.97
R18886 VDD.n6477 VDD.n5402 1084.97
R18887 VDD.n5402 VDD.n5392 1084.97
R18888 VDD.n6478 VDD.n5392 1084.97
R18889 VDD.n6488 VDD.n6487 1084.97
R18890 VDD.n6487 VDD.n5389 1084.97
R18891 VDD.n5389 VDD.n5381 1084.97
R18892 VDD.n6488 VDD.n5381 1084.97
R18893 VDD.n6498 VDD.n6497 1084.97
R18894 VDD.n6497 VDD.n5378 1084.97
R18895 VDD.n5378 VDD.n5371 1084.97
R18896 VDD.n6498 VDD.n5371 1084.97
R18897 VDD.n6508 VDD.n6507 1084.97
R18898 VDD.n6507 VDD.n5368 1084.97
R18899 VDD.n5368 VDD.n5358 1084.97
R18900 VDD.n6508 VDD.n5358 1084.97
R18901 VDD.n6518 VDD.n6517 1084.97
R18902 VDD.n6517 VDD.n5355 1084.97
R18903 VDD.n5355 VDD.n5346 1084.97
R18904 VDD.n6518 VDD.n5346 1084.97
R18905 VDD.n6525 VDD.n5343 1084.97
R18906 VDD.n6525 VDD.n5344 1084.97
R18907 VDD.n6529 VDD.n5344 1084.97
R18908 VDD.n6529 VDD.n5343 1084.97
R18909 VDD.n6535 VDD.n6534 1084.97
R18910 VDD.n6534 VDD.n5340 1084.97
R18911 VDD.n5340 VDD.n5330 1084.97
R18912 VDD.n6535 VDD.n5330 1084.97
R18913 VDD.n6545 VDD.n6544 1084.97
R18914 VDD.n6544 VDD.n5327 1084.97
R18915 VDD.n5327 VDD.n5319 1084.97
R18916 VDD.n6545 VDD.n5319 1084.97
R18917 VDD.n6555 VDD.n6554 1084.97
R18918 VDD.n6554 VDD.n5316 1084.97
R18919 VDD.n5316 VDD.n5309 1084.97
R18920 VDD.n6555 VDD.n5309 1084.97
R18921 VDD.n6565 VDD.n6564 1084.97
R18922 VDD.n6564 VDD.n5306 1084.97
R18923 VDD.n5306 VDD.n5299 1084.97
R18924 VDD.n6565 VDD.n5299 1084.97
R18925 VDD.n6578 VDD.n5292 1084.97
R18926 VDD.n6578 VDD.n5293 1084.97
R18927 VDD.n5298 VDD.n5293 1084.97
R18928 VDD.n5298 VDD.n5292 1084.97
R18929 VDD.n6577 VDD.n6572 1084.97
R18930 VDD.n6577 VDD.n6573 1084.97
R18931 VDD.n6572 VDD.n5290 1084.97
R18932 VDD.n6573 VDD.n5290 1084.97
R18933 VDD.n5283 VDD.n5279 1084.97
R18934 VDD.n6585 VDD.n5280 1084.97
R18935 VDD.n6585 VDD.n5279 1084.97
R18936 VDD.n6588 VDD.n5270 1084.97
R18937 VDD.n6588 VDD.n5271 1084.97
R18938 VDD.n6595 VDD.n5271 1084.97
R18939 VDD.n6595 VDD.n5270 1084.97
R18940 VDD.n6598 VDD.n5257 1084.97
R18941 VDD.n6598 VDD.n5258 1084.97
R18942 VDD.n6605 VDD.n5258 1084.97
R18943 VDD.n6605 VDD.n5257 1084.97
R18944 VDD.n6608 VDD.n5246 1084.97
R18945 VDD.n6608 VDD.n5247 1084.97
R18946 VDD.n6615 VDD.n5247 1084.97
R18947 VDD.n6615 VDD.n5246 1084.97
R18948 VDD.n6618 VDD.n5236 1084.97
R18949 VDD.n6618 VDD.n5237 1084.97
R18950 VDD.n6625 VDD.n5237 1084.97
R18951 VDD.n6625 VDD.n5236 1084.97
R18952 VDD.n6628 VDD.n5223 1084.97
R18953 VDD.n6628 VDD.n5224 1084.97
R18954 VDD.n6635 VDD.n5224 1084.97
R18955 VDD.n6635 VDD.n5223 1084.97
R18956 VDD.n6638 VDD.n5211 1084.97
R18957 VDD.n6638 VDD.n5212 1084.97
R18958 VDD.n6645 VDD.n5212 1084.97
R18959 VDD.n6645 VDD.n5211 1084.97
R18960 VDD.n6655 VDD.n5195 1084.97
R18961 VDD.n6655 VDD.n5196 1084.97
R18962 VDD.n6662 VDD.n5196 1084.97
R18963 VDD.n6662 VDD.n5195 1084.97
R18964 VDD.n6665 VDD.n5184 1084.97
R18965 VDD.n6665 VDD.n5185 1084.97
R18966 VDD.n6672 VDD.n5185 1084.97
R18967 VDD.n6672 VDD.n5184 1084.97
R18968 VDD.n6675 VDD.n5174 1084.97
R18969 VDD.n6675 VDD.n5175 1084.97
R18970 VDD.n6682 VDD.n5175 1084.97
R18971 VDD.n6682 VDD.n5174 1084.97
R18972 VDD.n6685 VDD.n5164 1084.97
R18973 VDD.n6685 VDD.n5165 1084.97
R18974 VDD.n6692 VDD.n5165 1084.97
R18975 VDD.n6692 VDD.n5164 1084.97
R18976 VDD.n6591 VDD.n6590 1084.97
R18977 VDD.n6590 VDD.n5276 1084.97
R18978 VDD.n5276 VDD.n5269 1084.97
R18979 VDD.n6591 VDD.n5269 1084.97
R18980 VDD.n6601 VDD.n6600 1084.97
R18981 VDD.n6600 VDD.n5266 1084.97
R18982 VDD.n5266 VDD.n5256 1084.97
R18983 VDD.n6601 VDD.n5256 1084.97
R18984 VDD.n6611 VDD.n6610 1084.97
R18985 VDD.n6610 VDD.n5253 1084.97
R18986 VDD.n5253 VDD.n5245 1084.97
R18987 VDD.n6611 VDD.n5245 1084.97
R18988 VDD.n6621 VDD.n6620 1084.97
R18989 VDD.n6620 VDD.n5242 1084.97
R18990 VDD.n5242 VDD.n5235 1084.97
R18991 VDD.n6621 VDD.n5235 1084.97
R18992 VDD.n6631 VDD.n6630 1084.97
R18993 VDD.n6630 VDD.n5232 1084.97
R18994 VDD.n5232 VDD.n5222 1084.97
R18995 VDD.n6631 VDD.n5222 1084.97
R18996 VDD.n6641 VDD.n6640 1084.97
R18997 VDD.n6640 VDD.n5219 1084.97
R18998 VDD.n5219 VDD.n5210 1084.97
R18999 VDD.n6641 VDD.n5210 1084.97
R19000 VDD.n6648 VDD.n5207 1084.97
R19001 VDD.n6648 VDD.n5208 1084.97
R19002 VDD.n6652 VDD.n5208 1084.97
R19003 VDD.n6652 VDD.n5207 1084.97
R19004 VDD.n6658 VDD.n6657 1084.97
R19005 VDD.n6657 VDD.n5204 1084.97
R19006 VDD.n5204 VDD.n5194 1084.97
R19007 VDD.n6658 VDD.n5194 1084.97
R19008 VDD.n6668 VDD.n6667 1084.97
R19009 VDD.n6667 VDD.n5191 1084.97
R19010 VDD.n5191 VDD.n5183 1084.97
R19011 VDD.n6668 VDD.n5183 1084.97
R19012 VDD.n6678 VDD.n6677 1084.97
R19013 VDD.n6677 VDD.n5180 1084.97
R19014 VDD.n5180 VDD.n5173 1084.97
R19015 VDD.n6678 VDD.n5173 1084.97
R19016 VDD.n6688 VDD.n6687 1084.97
R19017 VDD.n6687 VDD.n5170 1084.97
R19018 VDD.n5170 VDD.n5163 1084.97
R19019 VDD.n6688 VDD.n5163 1084.97
R19020 VDD.n6701 VDD.n5156 1084.97
R19021 VDD.n6701 VDD.n5157 1084.97
R19022 VDD.n5162 VDD.n5157 1084.97
R19023 VDD.n5162 VDD.n5156 1084.97
R19024 VDD.n6700 VDD.n6695 1084.97
R19025 VDD.n6700 VDD.n6696 1084.97
R19026 VDD.n6695 VDD.n5154 1084.97
R19027 VDD.n6696 VDD.n5154 1084.97
R19028 VDD.n5147 VDD.n5143 1084.97
R19029 VDD.n6708 VDD.n5144 1084.97
R19030 VDD.n6708 VDD.n5143 1084.97
R19031 VDD.n6711 VDD.n5134 1084.97
R19032 VDD.n6711 VDD.n5135 1084.97
R19033 VDD.n6718 VDD.n5135 1084.97
R19034 VDD.n6718 VDD.n5134 1084.97
R19035 VDD.n6721 VDD.n5121 1084.97
R19036 VDD.n6721 VDD.n5122 1084.97
R19037 VDD.n6728 VDD.n5122 1084.97
R19038 VDD.n6728 VDD.n5121 1084.97
R19039 VDD.n6731 VDD.n5110 1084.97
R19040 VDD.n6731 VDD.n5111 1084.97
R19041 VDD.n6738 VDD.n5111 1084.97
R19042 VDD.n6738 VDD.n5110 1084.97
R19043 VDD.n6741 VDD.n5100 1084.97
R19044 VDD.n6741 VDD.n5101 1084.97
R19045 VDD.n6748 VDD.n5101 1084.97
R19046 VDD.n6748 VDD.n5100 1084.97
R19047 VDD.n6751 VDD.n5087 1084.97
R19048 VDD.n6751 VDD.n5088 1084.97
R19049 VDD.n6758 VDD.n5088 1084.97
R19050 VDD.n6758 VDD.n5087 1084.97
R19051 VDD.n6761 VDD.n5075 1084.97
R19052 VDD.n6761 VDD.n5076 1084.97
R19053 VDD.n6768 VDD.n5076 1084.97
R19054 VDD.n6768 VDD.n5075 1084.97
R19055 VDD.n6778 VDD.n5059 1084.97
R19056 VDD.n6778 VDD.n5060 1084.97
R19057 VDD.n6785 VDD.n5060 1084.97
R19058 VDD.n6785 VDD.n5059 1084.97
R19059 VDD.n6788 VDD.n5048 1084.97
R19060 VDD.n6788 VDD.n5049 1084.97
R19061 VDD.n6795 VDD.n5049 1084.97
R19062 VDD.n6795 VDD.n5048 1084.97
R19063 VDD.n6798 VDD.n5038 1084.97
R19064 VDD.n6798 VDD.n5039 1084.97
R19065 VDD.n6805 VDD.n5039 1084.97
R19066 VDD.n6805 VDD.n5038 1084.97
R19067 VDD.n6808 VDD.n5028 1084.97
R19068 VDD.n6808 VDD.n5029 1084.97
R19069 VDD.n6815 VDD.n5029 1084.97
R19070 VDD.n6815 VDD.n5028 1084.97
R19071 VDD.n6714 VDD.n6713 1084.97
R19072 VDD.n6713 VDD.n5140 1084.97
R19073 VDD.n5140 VDD.n5133 1084.97
R19074 VDD.n6714 VDD.n5133 1084.97
R19075 VDD.n6724 VDD.n6723 1084.97
R19076 VDD.n6723 VDD.n5130 1084.97
R19077 VDD.n5130 VDD.n5120 1084.97
R19078 VDD.n6724 VDD.n5120 1084.97
R19079 VDD.n6734 VDD.n6733 1084.97
R19080 VDD.n6733 VDD.n5117 1084.97
R19081 VDD.n5117 VDD.n5109 1084.97
R19082 VDD.n6734 VDD.n5109 1084.97
R19083 VDD.n6744 VDD.n6743 1084.97
R19084 VDD.n6743 VDD.n5106 1084.97
R19085 VDD.n5106 VDD.n5099 1084.97
R19086 VDD.n6744 VDD.n5099 1084.97
R19087 VDD.n6754 VDD.n6753 1084.97
R19088 VDD.n6753 VDD.n5096 1084.97
R19089 VDD.n5096 VDD.n5086 1084.97
R19090 VDD.n6754 VDD.n5086 1084.97
R19091 VDD.n6764 VDD.n6763 1084.97
R19092 VDD.n6763 VDD.n5083 1084.97
R19093 VDD.n5083 VDD.n5074 1084.97
R19094 VDD.n6764 VDD.n5074 1084.97
R19095 VDD.n6771 VDD.n5071 1084.97
R19096 VDD.n6771 VDD.n5072 1084.97
R19097 VDD.n6775 VDD.n5072 1084.97
R19098 VDD.n6775 VDD.n5071 1084.97
R19099 VDD.n6781 VDD.n6780 1084.97
R19100 VDD.n6780 VDD.n5068 1084.97
R19101 VDD.n5068 VDD.n5058 1084.97
R19102 VDD.n6781 VDD.n5058 1084.97
R19103 VDD.n6791 VDD.n6790 1084.97
R19104 VDD.n6790 VDD.n5055 1084.97
R19105 VDD.n5055 VDD.n5047 1084.97
R19106 VDD.n6791 VDD.n5047 1084.97
R19107 VDD.n6801 VDD.n6800 1084.97
R19108 VDD.n6800 VDD.n5044 1084.97
R19109 VDD.n5044 VDD.n5037 1084.97
R19110 VDD.n6801 VDD.n5037 1084.97
R19111 VDD.n6811 VDD.n6810 1084.97
R19112 VDD.n6810 VDD.n5034 1084.97
R19113 VDD.n5034 VDD.n5027 1084.97
R19114 VDD.n6811 VDD.n5027 1084.97
R19115 VDD.n6824 VDD.n5020 1084.97
R19116 VDD.n6824 VDD.n5021 1084.97
R19117 VDD.n5026 VDD.n5021 1084.97
R19118 VDD.n5026 VDD.n5020 1084.97
R19119 VDD.n6823 VDD.n6818 1084.97
R19120 VDD.n6823 VDD.n6819 1084.97
R19121 VDD.n6818 VDD.n5018 1084.97
R19122 VDD.n6819 VDD.n5018 1084.97
R19123 VDD.n5009 VDD.n4759 1084.97
R19124 VDD.n5006 VDD.n4757 1084.97
R19125 VDD.n5006 VDD.n4759 1084.97
R19126 VDD.n5004 VDD.n4761 1084.97
R19127 VDD.n5004 VDD.n4762 1084.97
R19128 VDD.n4997 VDD.n4762 1084.97
R19129 VDD.n4997 VDD.n4761 1084.97
R19130 VDD.n4994 VDD.n4772 1084.97
R19131 VDD.n4994 VDD.n4773 1084.97
R19132 VDD.n4987 VDD.n4773 1084.97
R19133 VDD.n4987 VDD.n4772 1084.97
R19134 VDD.n4984 VDD.n4782 1084.97
R19135 VDD.n4984 VDD.n4783 1084.97
R19136 VDD.n4977 VDD.n4783 1084.97
R19137 VDD.n4977 VDD.n4782 1084.97
R19138 VDD.n4974 VDD.n4795 1084.97
R19139 VDD.n4974 VDD.n4796 1084.97
R19140 VDD.n4967 VDD.n4796 1084.97
R19141 VDD.n4967 VDD.n4795 1084.97
R19142 VDD.n4964 VDD.n4806 1084.97
R19143 VDD.n4964 VDD.n4807 1084.97
R19144 VDD.n4957 VDD.n4807 1084.97
R19145 VDD.n4957 VDD.n4806 1084.97
R19146 VDD.n4954 VDD.n4816 1084.97
R19147 VDD.n4954 VDD.n4817 1084.97
R19148 VDD.n4947 VDD.n4817 1084.97
R19149 VDD.n4947 VDD.n4816 1084.97
R19150 VDD.n4937 VDD.n4832 1084.97
R19151 VDD.n4937 VDD.n4833 1084.97
R19152 VDD.n4930 VDD.n4833 1084.97
R19153 VDD.n4930 VDD.n4832 1084.97
R19154 VDD.n4927 VDD.n4844 1084.97
R19155 VDD.n4927 VDD.n4845 1084.97
R19156 VDD.n4920 VDD.n4845 1084.97
R19157 VDD.n4920 VDD.n4844 1084.97
R19158 VDD.n4917 VDD.n4857 1084.97
R19159 VDD.n4917 VDD.n4858 1084.97
R19160 VDD.n4910 VDD.n4858 1084.97
R19161 VDD.n4910 VDD.n4857 1084.97
R19162 VDD.n4907 VDD.n4868 1084.97
R19163 VDD.n4907 VDD.n4869 1084.97
R19164 VDD.n4900 VDD.n4869 1084.97
R19165 VDD.n4900 VDD.n4868 1084.97
R19166 VDD.n5000 VDD.n4760 1084.97
R19167 VDD.n4768 VDD.n4760 1084.97
R19168 VDD.n4999 VDD.n4768 1084.97
R19169 VDD.n5000 VDD.n4999 1084.97
R19170 VDD.n4990 VDD.n4771 1084.97
R19171 VDD.n4778 VDD.n4771 1084.97
R19172 VDD.n4989 VDD.n4778 1084.97
R19173 VDD.n4990 VDD.n4989 1084.97
R19174 VDD.n4980 VDD.n4781 1084.97
R19175 VDD.n4791 VDD.n4781 1084.97
R19176 VDD.n4979 VDD.n4791 1084.97
R19177 VDD.n4980 VDD.n4979 1084.97
R19178 VDD.n4970 VDD.n4794 1084.97
R19179 VDD.n4802 VDD.n4794 1084.97
R19180 VDD.n4969 VDD.n4802 1084.97
R19181 VDD.n4970 VDD.n4969 1084.97
R19182 VDD.n4960 VDD.n4805 1084.97
R19183 VDD.n4812 VDD.n4805 1084.97
R19184 VDD.n4959 VDD.n4812 1084.97
R19185 VDD.n4960 VDD.n4959 1084.97
R19186 VDD.n4950 VDD.n4815 1084.97
R19187 VDD.n4825 VDD.n4815 1084.97
R19188 VDD.n4949 VDD.n4825 1084.97
R19189 VDD.n4950 VDD.n4949 1084.97
R19190 VDD.n4944 VDD.n4828 1084.97
R19191 VDD.n4944 VDD.n4829 1084.97
R19192 VDD.n4940 VDD.n4829 1084.97
R19193 VDD.n4940 VDD.n4828 1084.97
R19194 VDD.n4933 VDD.n4831 1084.97
R19195 VDD.n4840 VDD.n4831 1084.97
R19196 VDD.n4932 VDD.n4840 1084.97
R19197 VDD.n4933 VDD.n4932 1084.97
R19198 VDD.n4923 VDD.n4843 1084.97
R19199 VDD.n4853 VDD.n4843 1084.97
R19200 VDD.n4922 VDD.n4853 1084.97
R19201 VDD.n4923 VDD.n4922 1084.97
R19202 VDD.n4913 VDD.n4856 1084.97
R19203 VDD.n4864 VDD.n4856 1084.97
R19204 VDD.n4912 VDD.n4864 1084.97
R19205 VDD.n4913 VDD.n4912 1084.97
R19206 VDD.n4903 VDD.n4867 1084.97
R19207 VDD.n4874 VDD.n4867 1084.97
R19208 VDD.n4902 VDD.n4874 1084.97
R19209 VDD.n4903 VDD.n4902 1084.97
R19210 VDD.n4890 VDD.n4889 1084.97
R19211 VDD.n4890 VDD.n4877 1084.97
R19212 VDD.n4883 VDD.n4877 1084.97
R19213 VDD.n4889 VDD.n4883 1084.97
R19214 VDD.n4887 VDD.n4878 1084.97
R19215 VDD.n4897 VDD.n4878 1084.97
R19216 VDD.n4887 VDD.n4879 1084.97
R19217 VDD.n4897 VDD.n4879 1084.97
R19218 VDD.n4637 VDD.n2107 1084.97
R19219 VDD.n4637 VDD.n2108 1084.97
R19220 VDD.n4644 VDD.n2108 1084.97
R19221 VDD.n4644 VDD.n2107 1084.97
R19222 VDD.n4647 VDD.n2097 1084.97
R19223 VDD.n4647 VDD.n2098 1084.97
R19224 VDD.n4654 VDD.n2098 1084.97
R19225 VDD.n4654 VDD.n2097 1084.97
R19226 VDD.n4657 VDD.n2086 1084.97
R19227 VDD.n4657 VDD.n2087 1084.97
R19228 VDD.n4664 VDD.n2087 1084.97
R19229 VDD.n4664 VDD.n2086 1084.97
R19230 VDD.n4667 VDD.n2073 1084.97
R19231 VDD.n4667 VDD.n2074 1084.97
R19232 VDD.n4674 VDD.n2074 1084.97
R19233 VDD.n4674 VDD.n2073 1084.97
R19234 VDD.n4677 VDD.n2061 1084.97
R19235 VDD.n4677 VDD.n2062 1084.97
R19236 VDD.n4684 VDD.n2062 1084.97
R19237 VDD.n4684 VDD.n2061 1084.97
R19238 VDD.n4699 VDD.n4695 1084.97
R19239 VDD.n4695 VDD.n2041 1084.97
R19240 VDD.n4694 VDD.n2041 1084.97
R19241 VDD.n4699 VDD.n4694 1084.97
R19242 VDD.n4711 VDD.n2019 1084.97
R19243 VDD.n4711 VDD.n2020 1084.97
R19244 VDD.n4718 VDD.n2020 1084.97
R19245 VDD.n4718 VDD.n2019 1084.97
R19246 VDD.n4721 VDD.n2006 1084.97
R19247 VDD.n4721 VDD.n2007 1084.97
R19248 VDD.n4728 VDD.n2007 1084.97
R19249 VDD.n4728 VDD.n2006 1084.97
R19250 VDD.n4731 VDD.n1996 1084.97
R19251 VDD.n4731 VDD.n1997 1084.97
R19252 VDD.n4738 VDD.n1997 1084.97
R19253 VDD.n4738 VDD.n1996 1084.97
R19254 VDD.n4741 VDD.n1985 1084.97
R19255 VDD.n4741 VDD.n1986 1084.97
R19256 VDD.n4748 VDD.n1986 1084.97
R19257 VDD.n4748 VDD.n1985 1084.97
R19258 VDD.n4751 VDD.n1981 1084.97
R19259 VDD.n4751 VDD.n1979 1084.97
R19260 VDD.n1982 VDD.n1981 1084.97
R19261 VDD.n4640 VDD.n4639 1084.97
R19262 VDD.n4639 VDD.n4633 1084.97
R19263 VDD.n4633 VDD.n2106 1084.97
R19264 VDD.n4640 VDD.n2106 1084.97
R19265 VDD.n4650 VDD.n4649 1084.97
R19266 VDD.n4649 VDD.n2103 1084.97
R19267 VDD.n2103 VDD.n2096 1084.97
R19268 VDD.n4650 VDD.n2096 1084.97
R19269 VDD.n4660 VDD.n4659 1084.97
R19270 VDD.n4659 VDD.n2093 1084.97
R19271 VDD.n2093 VDD.n2085 1084.97
R19272 VDD.n4660 VDD.n2085 1084.97
R19273 VDD.n4670 VDD.n4669 1084.97
R19274 VDD.n4669 VDD.n2082 1084.97
R19275 VDD.n2082 VDD.n2072 1084.97
R19276 VDD.n4670 VDD.n2072 1084.97
R19277 VDD.n4680 VDD.n4679 1084.97
R19278 VDD.n4679 VDD.n2069 1084.97
R19279 VDD.n2069 VDD.n2060 1084.97
R19280 VDD.n4680 VDD.n2060 1084.97
R19281 VDD.n4687 VDD.n2057 1084.97
R19282 VDD.n4687 VDD.n2058 1084.97
R19283 VDD.n4691 VDD.n2058 1084.97
R19284 VDD.n4691 VDD.n2057 1084.97
R19285 VDD.n4700 VDD.n2044 1084.97
R19286 VDD.n2056 VDD.n2044 1084.97
R19287 VDD.n2056 VDD.n2043 1084.97
R19288 VDD.n4700 VDD.n2043 1084.97
R19289 VDD.n2036 VDD.n2030 1084.97
R19290 VDD.n2048 VDD.n2036 1084.97
R19291 VDD.n2048 VDD.n2045 1084.97
R19292 VDD.n2045 VDD.n2030 1084.97
R19293 VDD.n4714 VDD.n4713 1084.97
R19294 VDD.n4713 VDD.n2027 1084.97
R19295 VDD.n2027 VDD.n2018 1084.97
R19296 VDD.n4714 VDD.n2018 1084.97
R19297 VDD.n4724 VDD.n4723 1084.97
R19298 VDD.n4723 VDD.n2015 1084.97
R19299 VDD.n2015 VDD.n2005 1084.97
R19300 VDD.n4724 VDD.n2005 1084.97
R19301 VDD.n4734 VDD.n4733 1084.97
R19302 VDD.n4733 VDD.n2002 1084.97
R19303 VDD.n2002 VDD.n1995 1084.97
R19304 VDD.n4734 VDD.n1995 1084.97
R19305 VDD.n4744 VDD.n4743 1084.97
R19306 VDD.n4743 VDD.n1992 1084.97
R19307 VDD.n1992 VDD.n1984 1084.97
R19308 VDD.n4744 VDD.n1984 1084.97
R19309 VDD.n4708 VDD.n2031 1084.97
R19310 VDD.n2050 VDD.n2031 1084.97
R19311 VDD.n4708 VDD.n2032 1084.97
R19312 VDD.n2050 VDD.n2032 1084.97
R19313 VDD.n4512 VDD.n2243 1084.97
R19314 VDD.n4512 VDD.n2244 1084.97
R19315 VDD.n4519 VDD.n2244 1084.97
R19316 VDD.n4519 VDD.n2243 1084.97
R19317 VDD.n4522 VDD.n2233 1084.97
R19318 VDD.n4522 VDD.n2234 1084.97
R19319 VDD.n4529 VDD.n2234 1084.97
R19320 VDD.n4529 VDD.n2233 1084.97
R19321 VDD.n4532 VDD.n2222 1084.97
R19322 VDD.n4532 VDD.n2223 1084.97
R19323 VDD.n4539 VDD.n2223 1084.97
R19324 VDD.n4539 VDD.n2222 1084.97
R19325 VDD.n4542 VDD.n2209 1084.97
R19326 VDD.n4542 VDD.n2210 1084.97
R19327 VDD.n4549 VDD.n2210 1084.97
R19328 VDD.n4549 VDD.n2209 1084.97
R19329 VDD.n4552 VDD.n2197 1084.97
R19330 VDD.n4552 VDD.n2198 1084.97
R19331 VDD.n4559 VDD.n2198 1084.97
R19332 VDD.n4559 VDD.n2197 1084.97
R19333 VDD.n4574 VDD.n4570 1084.97
R19334 VDD.n4570 VDD.n2177 1084.97
R19335 VDD.n4569 VDD.n2177 1084.97
R19336 VDD.n4574 VDD.n4569 1084.97
R19337 VDD.n4586 VDD.n2155 1084.97
R19338 VDD.n4586 VDD.n2156 1084.97
R19339 VDD.n4593 VDD.n2156 1084.97
R19340 VDD.n4593 VDD.n2155 1084.97
R19341 VDD.n4596 VDD.n2142 1084.97
R19342 VDD.n4596 VDD.n2143 1084.97
R19343 VDD.n4603 VDD.n2143 1084.97
R19344 VDD.n4603 VDD.n2142 1084.97
R19345 VDD.n4606 VDD.n2132 1084.97
R19346 VDD.n4606 VDD.n2133 1084.97
R19347 VDD.n4613 VDD.n2133 1084.97
R19348 VDD.n4613 VDD.n2132 1084.97
R19349 VDD.n4616 VDD.n2121 1084.97
R19350 VDD.n4616 VDD.n2122 1084.97
R19351 VDD.n4623 VDD.n2122 1084.97
R19352 VDD.n4623 VDD.n2121 1084.97
R19353 VDD.n4626 VDD.n2117 1084.97
R19354 VDD.n4626 VDD.n2115 1084.97
R19355 VDD.n2118 VDD.n2117 1084.97
R19356 VDD.n4515 VDD.n4514 1084.97
R19357 VDD.n4514 VDD.n4508 1084.97
R19358 VDD.n4508 VDD.n2242 1084.97
R19359 VDD.n4515 VDD.n2242 1084.97
R19360 VDD.n4525 VDD.n4524 1084.97
R19361 VDD.n4524 VDD.n2239 1084.97
R19362 VDD.n2239 VDD.n2232 1084.97
R19363 VDD.n4525 VDD.n2232 1084.97
R19364 VDD.n4535 VDD.n4534 1084.97
R19365 VDD.n4534 VDD.n2229 1084.97
R19366 VDD.n2229 VDD.n2221 1084.97
R19367 VDD.n4535 VDD.n2221 1084.97
R19368 VDD.n4545 VDD.n4544 1084.97
R19369 VDD.n4544 VDD.n2218 1084.97
R19370 VDD.n2218 VDD.n2208 1084.97
R19371 VDD.n4545 VDD.n2208 1084.97
R19372 VDD.n4555 VDD.n4554 1084.97
R19373 VDD.n4554 VDD.n2205 1084.97
R19374 VDD.n2205 VDD.n2196 1084.97
R19375 VDD.n4555 VDD.n2196 1084.97
R19376 VDD.n4562 VDD.n2193 1084.97
R19377 VDD.n4562 VDD.n2194 1084.97
R19378 VDD.n4566 VDD.n2194 1084.97
R19379 VDD.n4566 VDD.n2193 1084.97
R19380 VDD.n4575 VDD.n2180 1084.97
R19381 VDD.n2192 VDD.n2180 1084.97
R19382 VDD.n2192 VDD.n2179 1084.97
R19383 VDD.n4575 VDD.n2179 1084.97
R19384 VDD.n2172 VDD.n2166 1084.97
R19385 VDD.n2184 VDD.n2172 1084.97
R19386 VDD.n2184 VDD.n2181 1084.97
R19387 VDD.n2181 VDD.n2166 1084.97
R19388 VDD.n4589 VDD.n4588 1084.97
R19389 VDD.n4588 VDD.n2163 1084.97
R19390 VDD.n2163 VDD.n2154 1084.97
R19391 VDD.n4589 VDD.n2154 1084.97
R19392 VDD.n4599 VDD.n4598 1084.97
R19393 VDD.n4598 VDD.n2151 1084.97
R19394 VDD.n2151 VDD.n2141 1084.97
R19395 VDD.n4599 VDD.n2141 1084.97
R19396 VDD.n4609 VDD.n4608 1084.97
R19397 VDD.n4608 VDD.n2138 1084.97
R19398 VDD.n2138 VDD.n2131 1084.97
R19399 VDD.n4609 VDD.n2131 1084.97
R19400 VDD.n4619 VDD.n4618 1084.97
R19401 VDD.n4618 VDD.n2128 1084.97
R19402 VDD.n2128 VDD.n2120 1084.97
R19403 VDD.n4619 VDD.n2120 1084.97
R19404 VDD.n4583 VDD.n2167 1084.97
R19405 VDD.n2186 VDD.n2167 1084.97
R19406 VDD.n4583 VDD.n2168 1084.97
R19407 VDD.n2186 VDD.n2168 1084.97
R19408 VDD.n4387 VDD.n2379 1084.97
R19409 VDD.n4387 VDD.n2380 1084.97
R19410 VDD.n4394 VDD.n2380 1084.97
R19411 VDD.n4394 VDD.n2379 1084.97
R19412 VDD.n4397 VDD.n2369 1084.97
R19413 VDD.n4397 VDD.n2370 1084.97
R19414 VDD.n4404 VDD.n2370 1084.97
R19415 VDD.n4404 VDD.n2369 1084.97
R19416 VDD.n4407 VDD.n2358 1084.97
R19417 VDD.n4407 VDD.n2359 1084.97
R19418 VDD.n4414 VDD.n2359 1084.97
R19419 VDD.n4414 VDD.n2358 1084.97
R19420 VDD.n4417 VDD.n2345 1084.97
R19421 VDD.n4417 VDD.n2346 1084.97
R19422 VDD.n4424 VDD.n2346 1084.97
R19423 VDD.n4424 VDD.n2345 1084.97
R19424 VDD.n4427 VDD.n2333 1084.97
R19425 VDD.n4427 VDD.n2334 1084.97
R19426 VDD.n4434 VDD.n2334 1084.97
R19427 VDD.n4434 VDD.n2333 1084.97
R19428 VDD.n4449 VDD.n4445 1084.97
R19429 VDD.n4445 VDD.n2313 1084.97
R19430 VDD.n4444 VDD.n2313 1084.97
R19431 VDD.n4449 VDD.n4444 1084.97
R19432 VDD.n4461 VDD.n2291 1084.97
R19433 VDD.n4461 VDD.n2292 1084.97
R19434 VDD.n4468 VDD.n2292 1084.97
R19435 VDD.n4468 VDD.n2291 1084.97
R19436 VDD.n4471 VDD.n2278 1084.97
R19437 VDD.n4471 VDD.n2279 1084.97
R19438 VDD.n4478 VDD.n2279 1084.97
R19439 VDD.n4478 VDD.n2278 1084.97
R19440 VDD.n4481 VDD.n2268 1084.97
R19441 VDD.n4481 VDD.n2269 1084.97
R19442 VDD.n4488 VDD.n2269 1084.97
R19443 VDD.n4488 VDD.n2268 1084.97
R19444 VDD.n4491 VDD.n2257 1084.97
R19445 VDD.n4491 VDD.n2258 1084.97
R19446 VDD.n4498 VDD.n2258 1084.97
R19447 VDD.n4498 VDD.n2257 1084.97
R19448 VDD.n4501 VDD.n2253 1084.97
R19449 VDD.n4501 VDD.n2251 1084.97
R19450 VDD.n2254 VDD.n2253 1084.97
R19451 VDD.n4390 VDD.n4389 1084.97
R19452 VDD.n4389 VDD.n4383 1084.97
R19453 VDD.n4383 VDD.n2378 1084.97
R19454 VDD.n4390 VDD.n2378 1084.97
R19455 VDD.n4400 VDD.n4399 1084.97
R19456 VDD.n4399 VDD.n2375 1084.97
R19457 VDD.n2375 VDD.n2368 1084.97
R19458 VDD.n4400 VDD.n2368 1084.97
R19459 VDD.n4410 VDD.n4409 1084.97
R19460 VDD.n4409 VDD.n2365 1084.97
R19461 VDD.n2365 VDD.n2357 1084.97
R19462 VDD.n4410 VDD.n2357 1084.97
R19463 VDD.n4420 VDD.n4419 1084.97
R19464 VDD.n4419 VDD.n2354 1084.97
R19465 VDD.n2354 VDD.n2344 1084.97
R19466 VDD.n4420 VDD.n2344 1084.97
R19467 VDD.n4430 VDD.n4429 1084.97
R19468 VDD.n4429 VDD.n2341 1084.97
R19469 VDD.n2341 VDD.n2332 1084.97
R19470 VDD.n4430 VDD.n2332 1084.97
R19471 VDD.n4437 VDD.n2329 1084.97
R19472 VDD.n4437 VDD.n2330 1084.97
R19473 VDD.n4441 VDD.n2330 1084.97
R19474 VDD.n4441 VDD.n2329 1084.97
R19475 VDD.n4450 VDD.n2316 1084.97
R19476 VDD.n2328 VDD.n2316 1084.97
R19477 VDD.n2328 VDD.n2315 1084.97
R19478 VDD.n4450 VDD.n2315 1084.97
R19479 VDD.n2308 VDD.n2302 1084.97
R19480 VDD.n2320 VDD.n2308 1084.97
R19481 VDD.n2320 VDD.n2317 1084.97
R19482 VDD.n2317 VDD.n2302 1084.97
R19483 VDD.n4464 VDD.n4463 1084.97
R19484 VDD.n4463 VDD.n2299 1084.97
R19485 VDD.n2299 VDD.n2290 1084.97
R19486 VDD.n4464 VDD.n2290 1084.97
R19487 VDD.n4474 VDD.n4473 1084.97
R19488 VDD.n4473 VDD.n2287 1084.97
R19489 VDD.n2287 VDD.n2277 1084.97
R19490 VDD.n4474 VDD.n2277 1084.97
R19491 VDD.n4484 VDD.n4483 1084.97
R19492 VDD.n4483 VDD.n2274 1084.97
R19493 VDD.n2274 VDD.n2267 1084.97
R19494 VDD.n4484 VDD.n2267 1084.97
R19495 VDD.n4494 VDD.n4493 1084.97
R19496 VDD.n4493 VDD.n2264 1084.97
R19497 VDD.n2264 VDD.n2256 1084.97
R19498 VDD.n4494 VDD.n2256 1084.97
R19499 VDD.n4458 VDD.n2303 1084.97
R19500 VDD.n2322 VDD.n2303 1084.97
R19501 VDD.n4458 VDD.n2304 1084.97
R19502 VDD.n2322 VDD.n2304 1084.97
R19503 VDD.n4262 VDD.n2515 1084.97
R19504 VDD.n4262 VDD.n2516 1084.97
R19505 VDD.n4269 VDD.n2516 1084.97
R19506 VDD.n4269 VDD.n2515 1084.97
R19507 VDD.n4272 VDD.n2505 1084.97
R19508 VDD.n4272 VDD.n2506 1084.97
R19509 VDD.n4279 VDD.n2506 1084.97
R19510 VDD.n4279 VDD.n2505 1084.97
R19511 VDD.n4282 VDD.n2494 1084.97
R19512 VDD.n4282 VDD.n2495 1084.97
R19513 VDD.n4289 VDD.n2495 1084.97
R19514 VDD.n4289 VDD.n2494 1084.97
R19515 VDD.n4292 VDD.n2481 1084.97
R19516 VDD.n4292 VDD.n2482 1084.97
R19517 VDD.n4299 VDD.n2482 1084.97
R19518 VDD.n4299 VDD.n2481 1084.97
R19519 VDD.n4302 VDD.n2469 1084.97
R19520 VDD.n4302 VDD.n2470 1084.97
R19521 VDD.n4309 VDD.n2470 1084.97
R19522 VDD.n4309 VDD.n2469 1084.97
R19523 VDD.n4324 VDD.n4320 1084.97
R19524 VDD.n4320 VDD.n2449 1084.97
R19525 VDD.n4319 VDD.n2449 1084.97
R19526 VDD.n4324 VDD.n4319 1084.97
R19527 VDD.n4336 VDD.n2427 1084.97
R19528 VDD.n4336 VDD.n2428 1084.97
R19529 VDD.n4343 VDD.n2428 1084.97
R19530 VDD.n4343 VDD.n2427 1084.97
R19531 VDD.n4346 VDD.n2414 1084.97
R19532 VDD.n4346 VDD.n2415 1084.97
R19533 VDD.n4353 VDD.n2415 1084.97
R19534 VDD.n4353 VDD.n2414 1084.97
R19535 VDD.n4356 VDD.n2404 1084.97
R19536 VDD.n4356 VDD.n2405 1084.97
R19537 VDD.n4363 VDD.n2405 1084.97
R19538 VDD.n4363 VDD.n2404 1084.97
R19539 VDD.n4366 VDD.n2393 1084.97
R19540 VDD.n4366 VDD.n2394 1084.97
R19541 VDD.n4373 VDD.n2394 1084.97
R19542 VDD.n4373 VDD.n2393 1084.97
R19543 VDD.n4376 VDD.n2389 1084.97
R19544 VDD.n4376 VDD.n2387 1084.97
R19545 VDD.n2390 VDD.n2389 1084.97
R19546 VDD.n4265 VDD.n4264 1084.97
R19547 VDD.n4264 VDD.n4258 1084.97
R19548 VDD.n4258 VDD.n2514 1084.97
R19549 VDD.n4265 VDD.n2514 1084.97
R19550 VDD.n4275 VDD.n4274 1084.97
R19551 VDD.n4274 VDD.n2511 1084.97
R19552 VDD.n2511 VDD.n2504 1084.97
R19553 VDD.n4275 VDD.n2504 1084.97
R19554 VDD.n4285 VDD.n4284 1084.97
R19555 VDD.n4284 VDD.n2501 1084.97
R19556 VDD.n2501 VDD.n2493 1084.97
R19557 VDD.n4285 VDD.n2493 1084.97
R19558 VDD.n4295 VDD.n4294 1084.97
R19559 VDD.n4294 VDD.n2490 1084.97
R19560 VDD.n2490 VDD.n2480 1084.97
R19561 VDD.n4295 VDD.n2480 1084.97
R19562 VDD.n4305 VDD.n4304 1084.97
R19563 VDD.n4304 VDD.n2477 1084.97
R19564 VDD.n2477 VDD.n2468 1084.97
R19565 VDD.n4305 VDD.n2468 1084.97
R19566 VDD.n4312 VDD.n2465 1084.97
R19567 VDD.n4312 VDD.n2466 1084.97
R19568 VDD.n4316 VDD.n2466 1084.97
R19569 VDD.n4316 VDD.n2465 1084.97
R19570 VDD.n4325 VDD.n2452 1084.97
R19571 VDD.n2464 VDD.n2452 1084.97
R19572 VDD.n2464 VDD.n2451 1084.97
R19573 VDD.n4325 VDD.n2451 1084.97
R19574 VDD.n2444 VDD.n2438 1084.97
R19575 VDD.n2456 VDD.n2444 1084.97
R19576 VDD.n2456 VDD.n2453 1084.97
R19577 VDD.n2453 VDD.n2438 1084.97
R19578 VDD.n4339 VDD.n4338 1084.97
R19579 VDD.n4338 VDD.n2435 1084.97
R19580 VDD.n2435 VDD.n2426 1084.97
R19581 VDD.n4339 VDD.n2426 1084.97
R19582 VDD.n4349 VDD.n4348 1084.97
R19583 VDD.n4348 VDD.n2423 1084.97
R19584 VDD.n2423 VDD.n2413 1084.97
R19585 VDD.n4349 VDD.n2413 1084.97
R19586 VDD.n4359 VDD.n4358 1084.97
R19587 VDD.n4358 VDD.n2410 1084.97
R19588 VDD.n2410 VDD.n2403 1084.97
R19589 VDD.n4359 VDD.n2403 1084.97
R19590 VDD.n4369 VDD.n4368 1084.97
R19591 VDD.n4368 VDD.n2400 1084.97
R19592 VDD.n2400 VDD.n2392 1084.97
R19593 VDD.n4369 VDD.n2392 1084.97
R19594 VDD.n4333 VDD.n2439 1084.97
R19595 VDD.n2458 VDD.n2439 1084.97
R19596 VDD.n4333 VDD.n2440 1084.97
R19597 VDD.n2458 VDD.n2440 1084.97
R19598 VDD.n4137 VDD.n2651 1084.97
R19599 VDD.n4137 VDD.n2652 1084.97
R19600 VDD.n4144 VDD.n2652 1084.97
R19601 VDD.n4144 VDD.n2651 1084.97
R19602 VDD.n4147 VDD.n2641 1084.97
R19603 VDD.n4147 VDD.n2642 1084.97
R19604 VDD.n4154 VDD.n2642 1084.97
R19605 VDD.n4154 VDD.n2641 1084.97
R19606 VDD.n4157 VDD.n2630 1084.97
R19607 VDD.n4157 VDD.n2631 1084.97
R19608 VDD.n4164 VDD.n2631 1084.97
R19609 VDD.n4164 VDD.n2630 1084.97
R19610 VDD.n4167 VDD.n2617 1084.97
R19611 VDD.n4167 VDD.n2618 1084.97
R19612 VDD.n4174 VDD.n2618 1084.97
R19613 VDD.n4174 VDD.n2617 1084.97
R19614 VDD.n4177 VDD.n2605 1084.97
R19615 VDD.n4177 VDD.n2606 1084.97
R19616 VDD.n4184 VDD.n2606 1084.97
R19617 VDD.n4184 VDD.n2605 1084.97
R19618 VDD.n4199 VDD.n4195 1084.97
R19619 VDD.n4195 VDD.n2585 1084.97
R19620 VDD.n4194 VDD.n2585 1084.97
R19621 VDD.n4199 VDD.n4194 1084.97
R19622 VDD.n4211 VDD.n2563 1084.97
R19623 VDD.n4211 VDD.n2564 1084.97
R19624 VDD.n4218 VDD.n2564 1084.97
R19625 VDD.n4218 VDD.n2563 1084.97
R19626 VDD.n4221 VDD.n2550 1084.97
R19627 VDD.n4221 VDD.n2551 1084.97
R19628 VDD.n4228 VDD.n2551 1084.97
R19629 VDD.n4228 VDD.n2550 1084.97
R19630 VDD.n4231 VDD.n2540 1084.97
R19631 VDD.n4231 VDD.n2541 1084.97
R19632 VDD.n4238 VDD.n2541 1084.97
R19633 VDD.n4238 VDD.n2540 1084.97
R19634 VDD.n4241 VDD.n2529 1084.97
R19635 VDD.n4241 VDD.n2530 1084.97
R19636 VDD.n4248 VDD.n2530 1084.97
R19637 VDD.n4248 VDD.n2529 1084.97
R19638 VDD.n4251 VDD.n2525 1084.97
R19639 VDD.n4251 VDD.n2523 1084.97
R19640 VDD.n2526 VDD.n2525 1084.97
R19641 VDD.n4140 VDD.n4139 1084.97
R19642 VDD.n4139 VDD.n4133 1084.97
R19643 VDD.n4133 VDD.n2650 1084.97
R19644 VDD.n4140 VDD.n2650 1084.97
R19645 VDD.n4150 VDD.n4149 1084.97
R19646 VDD.n4149 VDD.n2647 1084.97
R19647 VDD.n2647 VDD.n2640 1084.97
R19648 VDD.n4150 VDD.n2640 1084.97
R19649 VDD.n4160 VDD.n4159 1084.97
R19650 VDD.n4159 VDD.n2637 1084.97
R19651 VDD.n2637 VDD.n2629 1084.97
R19652 VDD.n4160 VDD.n2629 1084.97
R19653 VDD.n4170 VDD.n4169 1084.97
R19654 VDD.n4169 VDD.n2626 1084.97
R19655 VDD.n2626 VDD.n2616 1084.97
R19656 VDD.n4170 VDD.n2616 1084.97
R19657 VDD.n4180 VDD.n4179 1084.97
R19658 VDD.n4179 VDD.n2613 1084.97
R19659 VDD.n2613 VDD.n2604 1084.97
R19660 VDD.n4180 VDD.n2604 1084.97
R19661 VDD.n4187 VDD.n2601 1084.97
R19662 VDD.n4187 VDD.n2602 1084.97
R19663 VDD.n4191 VDD.n2602 1084.97
R19664 VDD.n4191 VDD.n2601 1084.97
R19665 VDD.n4200 VDD.n2588 1084.97
R19666 VDD.n2600 VDD.n2588 1084.97
R19667 VDD.n2600 VDD.n2587 1084.97
R19668 VDD.n4200 VDD.n2587 1084.97
R19669 VDD.n2580 VDD.n2574 1084.97
R19670 VDD.n2592 VDD.n2580 1084.97
R19671 VDD.n2592 VDD.n2589 1084.97
R19672 VDD.n2589 VDD.n2574 1084.97
R19673 VDD.n4214 VDD.n4213 1084.97
R19674 VDD.n4213 VDD.n2571 1084.97
R19675 VDD.n2571 VDD.n2562 1084.97
R19676 VDD.n4214 VDD.n2562 1084.97
R19677 VDD.n4224 VDD.n4223 1084.97
R19678 VDD.n4223 VDD.n2559 1084.97
R19679 VDD.n2559 VDD.n2549 1084.97
R19680 VDD.n4224 VDD.n2549 1084.97
R19681 VDD.n4234 VDD.n4233 1084.97
R19682 VDD.n4233 VDD.n2546 1084.97
R19683 VDD.n2546 VDD.n2539 1084.97
R19684 VDD.n4234 VDD.n2539 1084.97
R19685 VDD.n4244 VDD.n4243 1084.97
R19686 VDD.n4243 VDD.n2536 1084.97
R19687 VDD.n2536 VDD.n2528 1084.97
R19688 VDD.n4244 VDD.n2528 1084.97
R19689 VDD.n4208 VDD.n2575 1084.97
R19690 VDD.n2594 VDD.n2575 1084.97
R19691 VDD.n4208 VDD.n2576 1084.97
R19692 VDD.n2594 VDD.n2576 1084.97
R19693 VDD.n4012 VDD.n2787 1084.97
R19694 VDD.n4012 VDD.n2788 1084.97
R19695 VDD.n4019 VDD.n2788 1084.97
R19696 VDD.n4019 VDD.n2787 1084.97
R19697 VDD.n4022 VDD.n2777 1084.97
R19698 VDD.n4022 VDD.n2778 1084.97
R19699 VDD.n4029 VDD.n2778 1084.97
R19700 VDD.n4029 VDD.n2777 1084.97
R19701 VDD.n4032 VDD.n2766 1084.97
R19702 VDD.n4032 VDD.n2767 1084.97
R19703 VDD.n4039 VDD.n2767 1084.97
R19704 VDD.n4039 VDD.n2766 1084.97
R19705 VDD.n4042 VDD.n2753 1084.97
R19706 VDD.n4042 VDD.n2754 1084.97
R19707 VDD.n4049 VDD.n2754 1084.97
R19708 VDD.n4049 VDD.n2753 1084.97
R19709 VDD.n4052 VDD.n2741 1084.97
R19710 VDD.n4052 VDD.n2742 1084.97
R19711 VDD.n4059 VDD.n2742 1084.97
R19712 VDD.n4059 VDD.n2741 1084.97
R19713 VDD.n4074 VDD.n4070 1084.97
R19714 VDD.n4070 VDD.n2721 1084.97
R19715 VDD.n4069 VDD.n2721 1084.97
R19716 VDD.n4074 VDD.n4069 1084.97
R19717 VDD.n4086 VDD.n2699 1084.97
R19718 VDD.n4086 VDD.n2700 1084.97
R19719 VDD.n4093 VDD.n2700 1084.97
R19720 VDD.n4093 VDD.n2699 1084.97
R19721 VDD.n4096 VDD.n2686 1084.97
R19722 VDD.n4096 VDD.n2687 1084.97
R19723 VDD.n4103 VDD.n2687 1084.97
R19724 VDD.n4103 VDD.n2686 1084.97
R19725 VDD.n4106 VDD.n2676 1084.97
R19726 VDD.n4106 VDD.n2677 1084.97
R19727 VDD.n4113 VDD.n2677 1084.97
R19728 VDD.n4113 VDD.n2676 1084.97
R19729 VDD.n4116 VDD.n2665 1084.97
R19730 VDD.n4116 VDD.n2666 1084.97
R19731 VDD.n4123 VDD.n2666 1084.97
R19732 VDD.n4123 VDD.n2665 1084.97
R19733 VDD.n4126 VDD.n2661 1084.97
R19734 VDD.n4126 VDD.n2659 1084.97
R19735 VDD.n2662 VDD.n2661 1084.97
R19736 VDD.n4015 VDD.n4014 1084.97
R19737 VDD.n4014 VDD.n4008 1084.97
R19738 VDD.n4008 VDD.n2786 1084.97
R19739 VDD.n4015 VDD.n2786 1084.97
R19740 VDD.n4025 VDD.n4024 1084.97
R19741 VDD.n4024 VDD.n2783 1084.97
R19742 VDD.n2783 VDD.n2776 1084.97
R19743 VDD.n4025 VDD.n2776 1084.97
R19744 VDD.n4035 VDD.n4034 1084.97
R19745 VDD.n4034 VDD.n2773 1084.97
R19746 VDD.n2773 VDD.n2765 1084.97
R19747 VDD.n4035 VDD.n2765 1084.97
R19748 VDD.n4045 VDD.n4044 1084.97
R19749 VDD.n4044 VDD.n2762 1084.97
R19750 VDD.n2762 VDD.n2752 1084.97
R19751 VDD.n4045 VDD.n2752 1084.97
R19752 VDD.n4055 VDD.n4054 1084.97
R19753 VDD.n4054 VDD.n2749 1084.97
R19754 VDD.n2749 VDD.n2740 1084.97
R19755 VDD.n4055 VDD.n2740 1084.97
R19756 VDD.n4062 VDD.n2737 1084.97
R19757 VDD.n4062 VDD.n2738 1084.97
R19758 VDD.n4066 VDD.n2738 1084.97
R19759 VDD.n4066 VDD.n2737 1084.97
R19760 VDD.n4075 VDD.n2724 1084.97
R19761 VDD.n2736 VDD.n2724 1084.97
R19762 VDD.n2736 VDD.n2723 1084.97
R19763 VDD.n4075 VDD.n2723 1084.97
R19764 VDD.n2716 VDD.n2710 1084.97
R19765 VDD.n2728 VDD.n2716 1084.97
R19766 VDD.n2728 VDD.n2725 1084.97
R19767 VDD.n2725 VDD.n2710 1084.97
R19768 VDD.n4089 VDD.n4088 1084.97
R19769 VDD.n4088 VDD.n2707 1084.97
R19770 VDD.n2707 VDD.n2698 1084.97
R19771 VDD.n4089 VDD.n2698 1084.97
R19772 VDD.n4099 VDD.n4098 1084.97
R19773 VDD.n4098 VDD.n2695 1084.97
R19774 VDD.n2695 VDD.n2685 1084.97
R19775 VDD.n4099 VDD.n2685 1084.97
R19776 VDD.n4109 VDD.n4108 1084.97
R19777 VDD.n4108 VDD.n2682 1084.97
R19778 VDD.n2682 VDD.n2675 1084.97
R19779 VDD.n4109 VDD.n2675 1084.97
R19780 VDD.n4119 VDD.n4118 1084.97
R19781 VDD.n4118 VDD.n2672 1084.97
R19782 VDD.n2672 VDD.n2664 1084.97
R19783 VDD.n4119 VDD.n2664 1084.97
R19784 VDD.n4083 VDD.n2711 1084.97
R19785 VDD.n2730 VDD.n2711 1084.97
R19786 VDD.n4083 VDD.n2712 1084.97
R19787 VDD.n2730 VDD.n2712 1084.97
R19788 VDD.n3887 VDD.n2923 1084.97
R19789 VDD.n3887 VDD.n2924 1084.97
R19790 VDD.n3894 VDD.n2924 1084.97
R19791 VDD.n3894 VDD.n2923 1084.97
R19792 VDD.n3897 VDD.n2913 1084.97
R19793 VDD.n3897 VDD.n2914 1084.97
R19794 VDD.n3904 VDD.n2914 1084.97
R19795 VDD.n3904 VDD.n2913 1084.97
R19796 VDD.n3907 VDD.n2902 1084.97
R19797 VDD.n3907 VDD.n2903 1084.97
R19798 VDD.n3914 VDD.n2903 1084.97
R19799 VDD.n3914 VDD.n2902 1084.97
R19800 VDD.n3917 VDD.n2889 1084.97
R19801 VDD.n3917 VDD.n2890 1084.97
R19802 VDD.n3924 VDD.n2890 1084.97
R19803 VDD.n3924 VDD.n2889 1084.97
R19804 VDD.n3927 VDD.n2877 1084.97
R19805 VDD.n3927 VDD.n2878 1084.97
R19806 VDD.n3934 VDD.n2878 1084.97
R19807 VDD.n3934 VDD.n2877 1084.97
R19808 VDD.n3949 VDD.n3945 1084.97
R19809 VDD.n3945 VDD.n2857 1084.97
R19810 VDD.n3944 VDD.n2857 1084.97
R19811 VDD.n3949 VDD.n3944 1084.97
R19812 VDD.n3961 VDD.n2835 1084.97
R19813 VDD.n3961 VDD.n2836 1084.97
R19814 VDD.n3968 VDD.n2836 1084.97
R19815 VDD.n3968 VDD.n2835 1084.97
R19816 VDD.n3971 VDD.n2822 1084.97
R19817 VDD.n3971 VDD.n2823 1084.97
R19818 VDD.n3978 VDD.n2823 1084.97
R19819 VDD.n3978 VDD.n2822 1084.97
R19820 VDD.n3981 VDD.n2812 1084.97
R19821 VDD.n3981 VDD.n2813 1084.97
R19822 VDD.n3988 VDD.n2813 1084.97
R19823 VDD.n3988 VDD.n2812 1084.97
R19824 VDD.n3991 VDD.n2801 1084.97
R19825 VDD.n3991 VDD.n2802 1084.97
R19826 VDD.n3998 VDD.n2802 1084.97
R19827 VDD.n3998 VDD.n2801 1084.97
R19828 VDD.n4001 VDD.n2797 1084.97
R19829 VDD.n4001 VDD.n2795 1084.97
R19830 VDD.n2798 VDD.n2797 1084.97
R19831 VDD.n3890 VDD.n3889 1084.97
R19832 VDD.n3889 VDD.n3883 1084.97
R19833 VDD.n3883 VDD.n2922 1084.97
R19834 VDD.n3890 VDD.n2922 1084.97
R19835 VDD.n3900 VDD.n3899 1084.97
R19836 VDD.n3899 VDD.n2919 1084.97
R19837 VDD.n2919 VDD.n2912 1084.97
R19838 VDD.n3900 VDD.n2912 1084.97
R19839 VDD.n3910 VDD.n3909 1084.97
R19840 VDD.n3909 VDD.n2909 1084.97
R19841 VDD.n2909 VDD.n2901 1084.97
R19842 VDD.n3910 VDD.n2901 1084.97
R19843 VDD.n3920 VDD.n3919 1084.97
R19844 VDD.n3919 VDD.n2898 1084.97
R19845 VDD.n2898 VDD.n2888 1084.97
R19846 VDD.n3920 VDD.n2888 1084.97
R19847 VDD.n3930 VDD.n3929 1084.97
R19848 VDD.n3929 VDD.n2885 1084.97
R19849 VDD.n2885 VDD.n2876 1084.97
R19850 VDD.n3930 VDD.n2876 1084.97
R19851 VDD.n3937 VDD.n2873 1084.97
R19852 VDD.n3937 VDD.n2874 1084.97
R19853 VDD.n3941 VDD.n2874 1084.97
R19854 VDD.n3941 VDD.n2873 1084.97
R19855 VDD.n3950 VDD.n2860 1084.97
R19856 VDD.n2872 VDD.n2860 1084.97
R19857 VDD.n2872 VDD.n2859 1084.97
R19858 VDD.n3950 VDD.n2859 1084.97
R19859 VDD.n2852 VDD.n2846 1084.97
R19860 VDD.n2864 VDD.n2852 1084.97
R19861 VDD.n2864 VDD.n2861 1084.97
R19862 VDD.n2861 VDD.n2846 1084.97
R19863 VDD.n3964 VDD.n3963 1084.97
R19864 VDD.n3963 VDD.n2843 1084.97
R19865 VDD.n2843 VDD.n2834 1084.97
R19866 VDD.n3964 VDD.n2834 1084.97
R19867 VDD.n3974 VDD.n3973 1084.97
R19868 VDD.n3973 VDD.n2831 1084.97
R19869 VDD.n2831 VDD.n2821 1084.97
R19870 VDD.n3974 VDD.n2821 1084.97
R19871 VDD.n3984 VDD.n3983 1084.97
R19872 VDD.n3983 VDD.n2818 1084.97
R19873 VDD.n2818 VDD.n2811 1084.97
R19874 VDD.n3984 VDD.n2811 1084.97
R19875 VDD.n3994 VDD.n3993 1084.97
R19876 VDD.n3993 VDD.n2808 1084.97
R19877 VDD.n2808 VDD.n2800 1084.97
R19878 VDD.n3994 VDD.n2800 1084.97
R19879 VDD.n3958 VDD.n2847 1084.97
R19880 VDD.n2866 VDD.n2847 1084.97
R19881 VDD.n3958 VDD.n2848 1084.97
R19882 VDD.n2866 VDD.n2848 1084.97
R19883 VDD.n3539 VDD.n3217 1084.97
R19884 VDD.n3539 VDD.n3218 1084.97
R19885 VDD.n3546 VDD.n3218 1084.97
R19886 VDD.n3546 VDD.n3217 1084.97
R19887 VDD.n3554 VDD.n3550 1084.97
R19888 VDD.n3550 VDD.n3207 1084.97
R19889 VDD.n3549 VDD.n3207 1084.97
R19890 VDD.n3554 VDD.n3549 1084.97
R19891 VDD.n3239 VDD.n3226 1084.97
R19892 VDD.n3239 VDD.n3238 1084.97
R19893 VDD.n3238 VDD.n3232 1084.97
R19894 VDD.n3232 VDD.n3226 1084.97
R19895 VDD.n3542 VDD.n3541 1084.97
R19896 VDD.n3541 VDD.n3223 1084.97
R19897 VDD.n3223 VDD.n3216 1084.97
R19898 VDD.n3542 VDD.n3216 1084.97
R19899 VDD.n3555 VDD.n3210 1084.97
R19900 VDD.n3215 VDD.n3210 1084.97
R19901 VDD.n3215 VDD.n3209 1084.97
R19902 VDD.n3555 VDD.n3209 1084.97
R19903 VDD.n3536 VDD.n3227 1084.97
R19904 VDD.n3236 VDD.n3227 1084.97
R19905 VDD.n3536 VDD.n3228 1084.97
R19906 VDD.n3236 VDD.n3228 1084.97
R19907 VDD.n3386 VDD.n3286 1084.97
R19908 VDD.n3383 VDD.n3284 1084.97
R19909 VDD.n3383 VDD.n3286 1084.97
R19910 VDD.n3381 VDD.n3287 1084.97
R19911 VDD.n3381 VDD.n3288 1084.97
R19912 VDD.n3369 VDD.n3288 1084.97
R19913 VDD.n3369 VDD.n3287 1084.97
R19914 VDD.n3367 VDD.n3366 1084.97
R19915 VDD.n3372 VDD.n3366 1084.97
R19916 VDD.n3372 VDD.n3364 1084.97
R19917 VDD.n3423 VDD.n3395 1084.97
R19918 VDD.n3420 VDD.n3393 1084.97
R19919 VDD.n3420 VDD.n3395 1084.97
R19920 VDD.n3418 VDD.n3396 1084.97
R19921 VDD.n3418 VDD.n3397 1084.97
R19922 VDD.n3407 VDD.n3397 1084.97
R19923 VDD.n3407 VDD.n3396 1084.97
R19924 VDD.n3405 VDD.n3404 1084.97
R19925 VDD.n3410 VDD.n3404 1084.97
R19926 VDD.n3410 VDD.n3402 1084.97
R19927 VDD.n3275 VDD.n3269 1084.97
R19928 VDD.n3272 VDD.n3267 1084.97
R19929 VDD.n3272 VDD.n3269 1084.97
R19930 VDD.n3270 VDD.n3262 1084.97
R19931 VDD.n3270 VDD.n3263 1084.97
R19932 VDD.n3447 VDD.n3263 1084.97
R19933 VDD.n3447 VDD.n3262 1084.97
R19934 VDD.n3260 VDD.n3259 1084.97
R19935 VDD.n3450 VDD.n3259 1084.97
R19936 VDD.n3450 VDD.n3257 1084.97
R19937 VDD.n3481 VDD.n3249 1084.97
R19938 VDD.n3478 VDD.n3247 1084.97
R19939 VDD.n3478 VDD.n3249 1084.97
R19940 VDD.n3476 VDD.n3250 1084.97
R19941 VDD.n3476 VDD.n3251 1084.97
R19942 VDD.n3464 VDD.n3251 1084.97
R19943 VDD.n3464 VDD.n3250 1084.97
R19944 VDD.n3462 VDD.n3461 1084.97
R19945 VDD.n3467 VDD.n3461 1084.97
R19946 VDD.n3467 VDD.n3459 1084.97
R19947 VDD.n3517 VDD.n3489 1084.97
R19948 VDD.n3514 VDD.n3487 1084.97
R19949 VDD.n3514 VDD.n3489 1084.97
R19950 VDD.n3512 VDD.n3490 1084.97
R19951 VDD.n3512 VDD.n3491 1084.97
R19952 VDD.n3501 VDD.n3491 1084.97
R19953 VDD.n3501 VDD.n3490 1084.97
R19954 VDD.n3499 VDD.n3498 1084.97
R19955 VDD.n3504 VDD.n3498 1084.97
R19956 VDD.n3504 VDD.n3496 1084.97
R19957 VDD.n3331 VDD.n3325 1084.97
R19958 VDD.n3328 VDD.n3323 1084.97
R19959 VDD.n3328 VDD.n3325 1084.97
R19960 VDD.n3326 VDD.n3318 1084.97
R19961 VDD.n3326 VDD.n3319 1084.97
R19962 VDD.n3352 VDD.n3319 1084.97
R19963 VDD.n3352 VDD.n3318 1084.97
R19964 VDD.n3316 VDD.n3315 1084.97
R19965 VDD.n3355 VDD.n3315 1084.97
R19966 VDD.n3355 VDD.n3313 1084.97
R19967 VDD.n3762 VDD.n3749 1084.97
R19968 VDD.n3762 VDD.n3750 1084.97
R19969 VDD.n3769 VDD.n3750 1084.97
R19970 VDD.n3769 VDD.n3749 1084.97
R19971 VDD.n3772 VDD.n3739 1084.97
R19972 VDD.n3772 VDD.n3740 1084.97
R19973 VDD.n3779 VDD.n3740 1084.97
R19974 VDD.n3779 VDD.n3739 1084.97
R19975 VDD.n3782 VDD.n3728 1084.97
R19976 VDD.n3782 VDD.n3729 1084.97
R19977 VDD.n3789 VDD.n3729 1084.97
R19978 VDD.n3789 VDD.n3728 1084.97
R19979 VDD.n3792 VDD.n3715 1084.97
R19980 VDD.n3792 VDD.n3716 1084.97
R19981 VDD.n3799 VDD.n3716 1084.97
R19982 VDD.n3799 VDD.n3715 1084.97
R19983 VDD.n3802 VDD.n3703 1084.97
R19984 VDD.n3802 VDD.n3704 1084.97
R19985 VDD.n3809 VDD.n3704 1084.97
R19986 VDD.n3809 VDD.n3703 1084.97
R19987 VDD.n3824 VDD.n3820 1084.97
R19988 VDD.n3820 VDD.n3683 1084.97
R19989 VDD.n3819 VDD.n3683 1084.97
R19990 VDD.n3824 VDD.n3819 1084.97
R19991 VDD.n3836 VDD.n2971 1084.97
R19992 VDD.n3836 VDD.n2972 1084.97
R19993 VDD.n3843 VDD.n2972 1084.97
R19994 VDD.n3843 VDD.n2971 1084.97
R19995 VDD.n3846 VDD.n2958 1084.97
R19996 VDD.n3846 VDD.n2959 1084.97
R19997 VDD.n3853 VDD.n2959 1084.97
R19998 VDD.n3853 VDD.n2958 1084.97
R19999 VDD.n3856 VDD.n2948 1084.97
R20000 VDD.n3856 VDD.n2949 1084.97
R20001 VDD.n3863 VDD.n2949 1084.97
R20002 VDD.n3863 VDD.n2948 1084.97
R20003 VDD.n3866 VDD.n2937 1084.97
R20004 VDD.n3866 VDD.n2938 1084.97
R20005 VDD.n3873 VDD.n2938 1084.97
R20006 VDD.n3873 VDD.n2937 1084.97
R20007 VDD.n3876 VDD.n2933 1084.97
R20008 VDD.n3876 VDD.n2931 1084.97
R20009 VDD.n2934 VDD.n2933 1084.97
R20010 VDD.n3765 VDD.n3764 1084.97
R20011 VDD.n3764 VDD.n3758 1084.97
R20012 VDD.n3758 VDD.n3748 1084.97
R20013 VDD.n3765 VDD.n3748 1084.97
R20014 VDD.n3775 VDD.n3774 1084.97
R20015 VDD.n3774 VDD.n3745 1084.97
R20016 VDD.n3745 VDD.n3738 1084.97
R20017 VDD.n3775 VDD.n3738 1084.97
R20018 VDD.n3785 VDD.n3784 1084.97
R20019 VDD.n3784 VDD.n3735 1084.97
R20020 VDD.n3735 VDD.n3727 1084.97
R20021 VDD.n3785 VDD.n3727 1084.97
R20022 VDD.n3795 VDD.n3794 1084.97
R20023 VDD.n3794 VDD.n3724 1084.97
R20024 VDD.n3724 VDD.n3714 1084.97
R20025 VDD.n3795 VDD.n3714 1084.97
R20026 VDD.n3805 VDD.n3804 1084.97
R20027 VDD.n3804 VDD.n3711 1084.97
R20028 VDD.n3711 VDD.n3702 1084.97
R20029 VDD.n3805 VDD.n3702 1084.97
R20030 VDD.n3812 VDD.n3699 1084.97
R20031 VDD.n3812 VDD.n3700 1084.97
R20032 VDD.n3816 VDD.n3700 1084.97
R20033 VDD.n3816 VDD.n3699 1084.97
R20034 VDD.n3825 VDD.n3686 1084.97
R20035 VDD.n3698 VDD.n3686 1084.97
R20036 VDD.n3698 VDD.n3685 1084.97
R20037 VDD.n3825 VDD.n3685 1084.97
R20038 VDD.n3678 VDD.n3672 1084.97
R20039 VDD.n3690 VDD.n3678 1084.97
R20040 VDD.n3690 VDD.n3687 1084.97
R20041 VDD.n3687 VDD.n3672 1084.97
R20042 VDD.n3839 VDD.n3838 1084.97
R20043 VDD.n3838 VDD.n3669 1084.97
R20044 VDD.n3669 VDD.n2970 1084.97
R20045 VDD.n3839 VDD.n2970 1084.97
R20046 VDD.n3849 VDD.n3848 1084.97
R20047 VDD.n3848 VDD.n2967 1084.97
R20048 VDD.n2967 VDD.n2957 1084.97
R20049 VDD.n3849 VDD.n2957 1084.97
R20050 VDD.n3859 VDD.n3858 1084.97
R20051 VDD.n3858 VDD.n2954 1084.97
R20052 VDD.n2954 VDD.n2947 1084.97
R20053 VDD.n3859 VDD.n2947 1084.97
R20054 VDD.n3869 VDD.n3868 1084.97
R20055 VDD.n3868 VDD.n2944 1084.97
R20056 VDD.n2944 VDD.n2936 1084.97
R20057 VDD.n3869 VDD.n2936 1084.97
R20058 VDD.n3833 VDD.n3673 1084.97
R20059 VDD.n3692 VDD.n3673 1084.97
R20060 VDD.n3833 VDD.n3674 1084.97
R20061 VDD.n3692 VDD.n3674 1084.97
R20062 VDD.n255 VDD.n248 516.932
R20063 VDD.n263 VDD.n248 516.932
R20064 VDD.n257 VDD.n252 516.932
R20065 VDD.n261 VDD.n252 516.932
R20066 VDD.n130 VDD.n129 295.125
R20067 VDD.n165 VDD.n164 295.125
R20068 VDD.n200 VDD.n199 295.125
R20069 VDD.n235 VDD.n234 295.125
R20070 VDD.n6964 VDD.n6963 295.125
R20071 VDD.n6999 VDD.n6998 295.125
R20072 VDD.n7034 VDD.n7033 295.125
R20073 VDD.n6846 VDD.n6845 295.125
R20074 VDD.n109 VDD.t379 253.119
R20075 VDD.n108 VDD.t197 253.119
R20076 VDD.n130 VDD.t859 253.119
R20077 VDD.n129 VDD.t1071 253.119
R20078 VDD.n123 VDD.t1071 253.119
R20079 VDD.n122 VDD.t250 253.119
R20080 VDD.n144 VDD.t993 253.119
R20081 VDD.n143 VDD.t827 253.119
R20082 VDD.n165 VDD.t326 253.119
R20083 VDD.n164 VDD.t1026 253.119
R20084 VDD.n158 VDD.t1026 253.119
R20085 VDD.n157 VDD.t7 253.119
R20086 VDD.n179 VDD.t568 253.119
R20087 VDD.n178 VDD.t153 253.119
R20088 VDD.n200 VDD.t637 253.119
R20089 VDD.n199 VDD.t1065 253.119
R20090 VDD.n193 VDD.t1065 253.119
R20091 VDD.n192 VDD.t821 253.119
R20092 VDD.n214 VDD.t910 253.119
R20093 VDD.n213 VDD.t201 253.119
R20094 VDD.n235 VDD.t834 253.119
R20095 VDD.n234 VDD.t1092 253.119
R20096 VDD.n228 VDD.t1092 253.119
R20097 VDD.n227 VDD.t539 253.119
R20098 VDD.n6943 VDD.t329 253.119
R20099 VDD.n6942 VDD.t694 253.119
R20100 VDD.n6964 VDD.t324 253.119
R20101 VDD.n6963 VDD.t339 253.119
R20102 VDD.n6957 VDD.t339 253.119
R20103 VDD.n6956 VDD.t1036 253.119
R20104 VDD.n6978 VDD.t357 253.119
R20105 VDD.n6977 VDD.t878 253.119
R20106 VDD.n6999 VDD.t576 253.119
R20107 VDD.n6998 VDD.t620 253.119
R20108 VDD.n6992 VDD.t620 253.119
R20109 VDD.n6991 VDD.t1012 253.119
R20110 VDD.n7013 VDD.t582 253.119
R20111 VDD.n7012 VDD.t905 253.119
R20112 VDD.n7034 VDD.t600 253.119
R20113 VDD.n7033 VDD.t958 253.119
R20114 VDD.n7027 VDD.t958 253.119
R20115 VDD.n7026 VDD.t1040 253.119
R20116 VDD.n7048 VDD.t367 253.119
R20117 VDD.n7047 VDD.t870 253.119
R20118 VDD.n6845 VDD.t589 253.119
R20119 VDD.t409 VDD.n6846 253.119
R20120 VDD.t409 VDD.n7062 253.119
R20121 VDD.n7061 VDD.t1008 253.119
R20122 VDD.n3371 VDD.t384 253.119
R20123 VDD.n3370 VDD.t386 253.119
R20124 VDD.n3382 VDD.t386 253.119
R20125 VDD.t307 VDD.n3384 253.119
R20126 VDD.n3409 VDD.t990 253.119
R20127 VDD.n3408 VDD.t992 253.119
R20128 VDD.n3419 VDD.t992 253.119
R20129 VDD.t618 VDD.n3421 253.119
R20130 VDD.n3449 VDD.t464 253.119
R20131 VDD.n3448 VDD.t225 253.119
R20132 VDD.n3271 VDD.t225 253.119
R20133 VDD.t381 VDD.n3273 253.119
R20134 VDD.n3466 VDD.t405 253.119
R20135 VDD.n3465 VDD.t407 253.119
R20136 VDD.n3477 VDD.t407 253.119
R20137 VDD.t867 VDD.n3479 253.119
R20138 VDD.n3503 VDD.t640 253.119
R20139 VDD.n3502 VDD.t642 253.119
R20140 VDD.n3513 VDD.t642 253.119
R20141 VDD.t966 VDD.n3515 253.119
R20142 VDD.n3354 VDD.t211 253.119
R20143 VDD.n3353 VDD.t213 253.119
R20144 VDD.n3327 VDD.t213 253.119
R20145 VDD.t533 VDD.n3329 253.119
R20146 VDD.n103 VDD.n102 214.357
R20147 VDD.n97 VDD.n96 214.357
R20148 VDD.n117 VDD.n116 214.357
R20149 VDD.n81 VDD.n80 214.357
R20150 VDD.n138 VDD.n137 214.357
R20151 VDD.n72 VDD.n71 214.357
R20152 VDD.n152 VDD.n151 214.357
R20153 VDD.n56 VDD.n55 214.357
R20154 VDD.n173 VDD.n172 214.357
R20155 VDD.n47 VDD.n46 214.357
R20156 VDD.n187 VDD.n186 214.357
R20157 VDD.n31 VDD.n30 214.357
R20158 VDD.n208 VDD.n207 214.357
R20159 VDD.n22 VDD.n21 214.357
R20160 VDD.n222 VDD.n221 214.357
R20161 VDD.n6 VDD.n5 214.357
R20162 VDD.n7056 VDD.n7055 214.357
R20163 VDD.n6937 VDD.n6936 214.357
R20164 VDD.n6931 VDD.n6930 214.357
R20165 VDD.n6951 VDD.n6950 214.357
R20166 VDD.n6915 VDD.n6914 214.357
R20167 VDD.n6972 VDD.n6971 214.357
R20168 VDD.n6906 VDD.n6905 214.357
R20169 VDD.n6986 VDD.n6985 214.357
R20170 VDD.n6890 VDD.n6889 214.357
R20171 VDD.n7007 VDD.n7006 214.357
R20172 VDD.n6881 VDD.n6880 214.357
R20173 VDD.n7021 VDD.n7020 214.357
R20174 VDD.n6865 VDD.n6864 214.357
R20175 VDD.n7042 VDD.n7041 214.357
R20176 VDD.n6856 VDD.n6855 214.357
R20177 VDD.n6840 VDD.n6839 214.357
R20178 VDD.n3386 VDD.n3385 214.357
R20179 VDD.n3368 VDD.n3367 214.357
R20180 VDD.n3423 VDD.n3422 214.357
R20181 VDD.n3406 VDD.n3405 214.357
R20182 VDD.n3275 VDD.n3274 214.357
R20183 VDD.n3261 VDD.n3260 214.357
R20184 VDD.n3481 VDD.n3480 214.357
R20185 VDD.n3463 VDD.n3462 214.357
R20186 VDD.n3517 VDD.n3516 214.357
R20187 VDD.n3500 VDD.n3499 214.357
R20188 VDD.n3331 VDD.n3330 214.357
R20189 VDD.n3317 VDD.n3316 214.357
R20190 VDD.n7599 VDD.n7598 212.329
R20191 VDD.n7598 VDD.n7591 212.329
R20192 VDD.n7600 VDD.n7590 212.329
R20193 VDD.n7607 VDD.n7590 212.329
R20194 VDD.n7586 VDD.n7585 212.329
R20195 VDD.n7585 VDD.n7581 212.329
R20196 VDD.n7610 VDD.n7580 212.329
R20197 VDD.n7617 VDD.n7580 212.329
R20198 VDD.n7576 VDD.n7575 212.329
R20199 VDD.n7575 VDD.n7570 212.329
R20200 VDD.n7620 VDD.n7569 212.329
R20201 VDD.n7627 VDD.n7569 212.329
R20202 VDD.n7565 VDD.n7564 212.329
R20203 VDD.n7564 VDD.n7557 212.329
R20204 VDD.n7630 VDD.n7556 212.329
R20205 VDD.n7637 VDD.n7556 212.329
R20206 VDD.n7552 VDD.n7551 212.329
R20207 VDD.n7551 VDD.n7545 212.329
R20208 VDD.n7640 VDD.n7544 212.329
R20209 VDD.n7647 VDD.n7544 212.329
R20210 VDD.n7653 VDD.n7652 212.329
R20211 VDD.n7654 VDD.n7653 212.329
R20212 VDD.n7537 VDD.n7536 212.329
R20213 VDD.n7536 VDD.n7529 212.329
R20214 VDD.n7657 VDD.n7528 212.329
R20215 VDD.n7664 VDD.n7528 212.329
R20216 VDD.n7524 VDD.n7523 212.329
R20217 VDD.n7523 VDD.n7519 212.329
R20218 VDD.n7667 VDD.n7518 212.329
R20219 VDD.n7674 VDD.n7518 212.329
R20220 VDD.n7514 VDD.n7513 212.329
R20221 VDD.n7513 VDD.n7508 212.329
R20222 VDD.n7677 VDD.n7507 212.329
R20223 VDD.n7684 VDD.n7507 212.329
R20224 VDD.n7503 VDD.n7502 212.329
R20225 VDD.n7502 VDD.n7495 212.329
R20226 VDD.n7687 VDD.n7494 212.329
R20227 VDD.n7694 VDD.n7494 212.329
R20228 VDD.n7490 VDD.n7489 212.329
R20229 VDD.n7489 VDD.n7486 212.329
R20230 VDD.n7697 VDD.n7485 212.329
R20231 VDD.n7704 VDD.n7485 212.329
R20232 VDD.n7480 VDD.n7479 212.329
R20233 VDD.n7480 VDD.n7478 212.329
R20234 VDD.n7712 VDD.n7711 212.329
R20235 VDD.n7712 VDD.n7710 212.329
R20236 VDD.n7474 VDD.n7469 212.329
R20237 VDD.n7472 VDD.n7469 212.329
R20238 VDD.n1717 VDD.n1716 212.329
R20239 VDD.n1716 VDD.n1709 212.329
R20240 VDD.n1718 VDD.n1708 212.329
R20241 VDD.n1725 VDD.n1708 212.329
R20242 VDD.n1704 VDD.n1703 212.329
R20243 VDD.n1703 VDD.n1699 212.329
R20244 VDD.n1728 VDD.n1698 212.329
R20245 VDD.n1735 VDD.n1698 212.329
R20246 VDD.n1694 VDD.n1693 212.329
R20247 VDD.n1693 VDD.n1688 212.329
R20248 VDD.n1738 VDD.n1687 212.329
R20249 VDD.n1745 VDD.n1687 212.329
R20250 VDD.n1683 VDD.n1682 212.329
R20251 VDD.n1682 VDD.n1675 212.329
R20252 VDD.n1748 VDD.n1674 212.329
R20253 VDD.n1755 VDD.n1674 212.329
R20254 VDD.n1670 VDD.n1669 212.329
R20255 VDD.n1669 VDD.n1663 212.329
R20256 VDD.n1758 VDD.n1662 212.329
R20257 VDD.n1765 VDD.n1662 212.329
R20258 VDD.n1771 VDD.n1770 212.329
R20259 VDD.n1772 VDD.n1771 212.329
R20260 VDD.n1655 VDD.n1654 212.329
R20261 VDD.n1654 VDD.n1647 212.329
R20262 VDD.n1775 VDD.n1646 212.329
R20263 VDD.n1782 VDD.n1646 212.329
R20264 VDD.n1642 VDD.n1641 212.329
R20265 VDD.n1641 VDD.n1637 212.329
R20266 VDD.n1785 VDD.n1636 212.329
R20267 VDD.n1792 VDD.n1636 212.329
R20268 VDD.n1632 VDD.n1631 212.329
R20269 VDD.n1631 VDD.n1626 212.329
R20270 VDD.n1795 VDD.n1625 212.329
R20271 VDD.n1802 VDD.n1625 212.329
R20272 VDD.n1621 VDD.n1620 212.329
R20273 VDD.n1620 VDD.n1613 212.329
R20274 VDD.n1805 VDD.n1612 212.329
R20275 VDD.n1812 VDD.n1612 212.329
R20276 VDD.n1608 VDD.n1607 212.329
R20277 VDD.n1607 VDD.n1603 212.329
R20278 VDD.n1815 VDD.n1602 212.329
R20279 VDD.n1822 VDD.n1602 212.329
R20280 VDD.n1598 VDD.n1597 212.329
R20281 VDD.n1597 VDD.n1592 212.329
R20282 VDD.n1825 VDD.n1591 212.329
R20283 VDD.n1832 VDD.n1591 212.329
R20284 VDD.n1837 VDD.n1584 212.329
R20285 VDD.n1584 VDD.n1582 212.329
R20286 VDD.n1457 VDD.n1456 212.329
R20287 VDD.n1456 VDD.n1449 212.329
R20288 VDD.n1458 VDD.n1448 212.329
R20289 VDD.n1465 VDD.n1448 212.329
R20290 VDD.n1444 VDD.n1443 212.329
R20291 VDD.n1443 VDD.n1439 212.329
R20292 VDD.n1468 VDD.n1438 212.329
R20293 VDD.n1475 VDD.n1438 212.329
R20294 VDD.n1434 VDD.n1433 212.329
R20295 VDD.n1433 VDD.n1428 212.329
R20296 VDD.n1478 VDD.n1427 212.329
R20297 VDD.n1485 VDD.n1427 212.329
R20298 VDD.n1423 VDD.n1422 212.329
R20299 VDD.n1422 VDD.n1415 212.329
R20300 VDD.n1488 VDD.n1414 212.329
R20301 VDD.n1495 VDD.n1414 212.329
R20302 VDD.n1410 VDD.n1409 212.329
R20303 VDD.n1409 VDD.n1403 212.329
R20304 VDD.n1498 VDD.n1402 212.329
R20305 VDD.n1505 VDD.n1402 212.329
R20306 VDD.n1511 VDD.n1510 212.329
R20307 VDD.n1512 VDD.n1511 212.329
R20308 VDD.n1395 VDD.n1394 212.329
R20309 VDD.n1394 VDD.n1387 212.329
R20310 VDD.n1515 VDD.n1386 212.329
R20311 VDD.n1522 VDD.n1386 212.329
R20312 VDD.n1382 VDD.n1381 212.329
R20313 VDD.n1381 VDD.n1377 212.329
R20314 VDD.n1525 VDD.n1376 212.329
R20315 VDD.n1532 VDD.n1376 212.329
R20316 VDD.n1372 VDD.n1371 212.329
R20317 VDD.n1371 VDD.n1366 212.329
R20318 VDD.n1535 VDD.n1365 212.329
R20319 VDD.n1542 VDD.n1365 212.329
R20320 VDD.n1361 VDD.n1360 212.329
R20321 VDD.n1360 VDD.n1353 212.329
R20322 VDD.n1545 VDD.n1352 212.329
R20323 VDD.n1552 VDD.n1352 212.329
R20324 VDD.n1348 VDD.n1347 212.329
R20325 VDD.n1347 VDD.n1343 212.329
R20326 VDD.n1555 VDD.n1342 212.329
R20327 VDD.n1562 VDD.n1342 212.329
R20328 VDD.n1338 VDD.n1337 212.329
R20329 VDD.n1337 VDD.n1332 212.329
R20330 VDD.n1565 VDD.n1331 212.329
R20331 VDD.n1572 VDD.n1331 212.329
R20332 VDD.n1577 VDD.n1324 212.329
R20333 VDD.n1324 VDD.n1322 212.329
R20334 VDD.n1197 VDD.n1196 212.329
R20335 VDD.n1196 VDD.n1189 212.329
R20336 VDD.n1198 VDD.n1188 212.329
R20337 VDD.n1205 VDD.n1188 212.329
R20338 VDD.n1184 VDD.n1183 212.329
R20339 VDD.n1183 VDD.n1179 212.329
R20340 VDD.n1208 VDD.n1178 212.329
R20341 VDD.n1215 VDD.n1178 212.329
R20342 VDD.n1174 VDD.n1173 212.329
R20343 VDD.n1173 VDD.n1168 212.329
R20344 VDD.n1218 VDD.n1167 212.329
R20345 VDD.n1225 VDD.n1167 212.329
R20346 VDD.n1163 VDD.n1162 212.329
R20347 VDD.n1162 VDD.n1155 212.329
R20348 VDD.n1228 VDD.n1154 212.329
R20349 VDD.n1235 VDD.n1154 212.329
R20350 VDD.n1150 VDD.n1149 212.329
R20351 VDD.n1149 VDD.n1143 212.329
R20352 VDD.n1238 VDD.n1142 212.329
R20353 VDD.n1245 VDD.n1142 212.329
R20354 VDD.n1251 VDD.n1250 212.329
R20355 VDD.n1252 VDD.n1251 212.329
R20356 VDD.n1135 VDD.n1134 212.329
R20357 VDD.n1134 VDD.n1127 212.329
R20358 VDD.n1255 VDD.n1126 212.329
R20359 VDD.n1262 VDD.n1126 212.329
R20360 VDD.n1122 VDD.n1121 212.329
R20361 VDD.n1121 VDD.n1117 212.329
R20362 VDD.n1265 VDD.n1116 212.329
R20363 VDD.n1272 VDD.n1116 212.329
R20364 VDD.n1112 VDD.n1111 212.329
R20365 VDD.n1111 VDD.n1106 212.329
R20366 VDD.n1275 VDD.n1105 212.329
R20367 VDD.n1282 VDD.n1105 212.329
R20368 VDD.n1101 VDD.n1100 212.329
R20369 VDD.n1100 VDD.n1093 212.329
R20370 VDD.n1285 VDD.n1092 212.329
R20371 VDD.n1292 VDD.n1092 212.329
R20372 VDD.n1088 VDD.n1087 212.329
R20373 VDD.n1087 VDD.n1083 212.329
R20374 VDD.n1295 VDD.n1082 212.329
R20375 VDD.n1302 VDD.n1082 212.329
R20376 VDD.n1078 VDD.n1077 212.329
R20377 VDD.n1077 VDD.n1072 212.329
R20378 VDD.n1305 VDD.n1071 212.329
R20379 VDD.n1312 VDD.n1071 212.329
R20380 VDD.n1317 VDD.n1064 212.329
R20381 VDD.n1064 VDD.n1062 212.329
R20382 VDD.n937 VDD.n936 212.329
R20383 VDD.n936 VDD.n929 212.329
R20384 VDD.n938 VDD.n928 212.329
R20385 VDD.n945 VDD.n928 212.329
R20386 VDD.n924 VDD.n923 212.329
R20387 VDD.n923 VDD.n919 212.329
R20388 VDD.n948 VDD.n918 212.329
R20389 VDD.n955 VDD.n918 212.329
R20390 VDD.n914 VDD.n913 212.329
R20391 VDD.n913 VDD.n908 212.329
R20392 VDD.n958 VDD.n907 212.329
R20393 VDD.n965 VDD.n907 212.329
R20394 VDD.n903 VDD.n902 212.329
R20395 VDD.n902 VDD.n895 212.329
R20396 VDD.n968 VDD.n894 212.329
R20397 VDD.n975 VDD.n894 212.329
R20398 VDD.n890 VDD.n889 212.329
R20399 VDD.n889 VDD.n883 212.329
R20400 VDD.n978 VDD.n882 212.329
R20401 VDD.n985 VDD.n882 212.329
R20402 VDD.n991 VDD.n990 212.329
R20403 VDD.n992 VDD.n991 212.329
R20404 VDD.n875 VDD.n874 212.329
R20405 VDD.n874 VDD.n867 212.329
R20406 VDD.n995 VDD.n866 212.329
R20407 VDD.n1002 VDD.n866 212.329
R20408 VDD.n862 VDD.n861 212.329
R20409 VDD.n861 VDD.n857 212.329
R20410 VDD.n1005 VDD.n856 212.329
R20411 VDD.n1012 VDD.n856 212.329
R20412 VDD.n852 VDD.n851 212.329
R20413 VDD.n851 VDD.n846 212.329
R20414 VDD.n1015 VDD.n845 212.329
R20415 VDD.n1022 VDD.n845 212.329
R20416 VDD.n841 VDD.n840 212.329
R20417 VDD.n840 VDD.n833 212.329
R20418 VDD.n1025 VDD.n832 212.329
R20419 VDD.n1032 VDD.n832 212.329
R20420 VDD.n828 VDD.n827 212.329
R20421 VDD.n827 VDD.n823 212.329
R20422 VDD.n1035 VDD.n822 212.329
R20423 VDD.n1042 VDD.n822 212.329
R20424 VDD.n818 VDD.n817 212.329
R20425 VDD.n817 VDD.n812 212.329
R20426 VDD.n1045 VDD.n811 212.329
R20427 VDD.n1052 VDD.n811 212.329
R20428 VDD.n1057 VDD.n804 212.329
R20429 VDD.n804 VDD.n802 212.329
R20430 VDD.n677 VDD.n676 212.329
R20431 VDD.n676 VDD.n669 212.329
R20432 VDD.n678 VDD.n668 212.329
R20433 VDD.n685 VDD.n668 212.329
R20434 VDD.n664 VDD.n663 212.329
R20435 VDD.n663 VDD.n659 212.329
R20436 VDD.n688 VDD.n658 212.329
R20437 VDD.n695 VDD.n658 212.329
R20438 VDD.n654 VDD.n653 212.329
R20439 VDD.n653 VDD.n648 212.329
R20440 VDD.n698 VDD.n647 212.329
R20441 VDD.n705 VDD.n647 212.329
R20442 VDD.n643 VDD.n642 212.329
R20443 VDD.n642 VDD.n635 212.329
R20444 VDD.n708 VDD.n634 212.329
R20445 VDD.n715 VDD.n634 212.329
R20446 VDD.n630 VDD.n629 212.329
R20447 VDD.n629 VDD.n623 212.329
R20448 VDD.n718 VDD.n622 212.329
R20449 VDD.n725 VDD.n622 212.329
R20450 VDD.n731 VDD.n730 212.329
R20451 VDD.n732 VDD.n731 212.329
R20452 VDD.n615 VDD.n614 212.329
R20453 VDD.n614 VDD.n607 212.329
R20454 VDD.n735 VDD.n606 212.329
R20455 VDD.n742 VDD.n606 212.329
R20456 VDD.n602 VDD.n601 212.329
R20457 VDD.n601 VDD.n597 212.329
R20458 VDD.n745 VDD.n596 212.329
R20459 VDD.n752 VDD.n596 212.329
R20460 VDD.n592 VDD.n591 212.329
R20461 VDD.n591 VDD.n586 212.329
R20462 VDD.n755 VDD.n585 212.329
R20463 VDD.n762 VDD.n585 212.329
R20464 VDD.n581 VDD.n580 212.329
R20465 VDD.n580 VDD.n573 212.329
R20466 VDD.n765 VDD.n572 212.329
R20467 VDD.n772 VDD.n572 212.329
R20468 VDD.n568 VDD.n567 212.329
R20469 VDD.n567 VDD.n563 212.329
R20470 VDD.n775 VDD.n562 212.329
R20471 VDD.n782 VDD.n562 212.329
R20472 VDD.n558 VDD.n557 212.329
R20473 VDD.n557 VDD.n552 212.329
R20474 VDD.n785 VDD.n551 212.329
R20475 VDD.n792 VDD.n551 212.329
R20476 VDD.n797 VDD.n544 212.329
R20477 VDD.n544 VDD.n542 212.329
R20478 VDD.n417 VDD.n416 212.329
R20479 VDD.n416 VDD.n409 212.329
R20480 VDD.n418 VDD.n408 212.329
R20481 VDD.n425 VDD.n408 212.329
R20482 VDD.n404 VDD.n403 212.329
R20483 VDD.n403 VDD.n399 212.329
R20484 VDD.n428 VDD.n398 212.329
R20485 VDD.n435 VDD.n398 212.329
R20486 VDD.n394 VDD.n393 212.329
R20487 VDD.n393 VDD.n388 212.329
R20488 VDD.n438 VDD.n387 212.329
R20489 VDD.n445 VDD.n387 212.329
R20490 VDD.n383 VDD.n382 212.329
R20491 VDD.n382 VDD.n375 212.329
R20492 VDD.n448 VDD.n374 212.329
R20493 VDD.n455 VDD.n374 212.329
R20494 VDD.n370 VDD.n369 212.329
R20495 VDD.n369 VDD.n363 212.329
R20496 VDD.n458 VDD.n362 212.329
R20497 VDD.n465 VDD.n362 212.329
R20498 VDD.n471 VDD.n470 212.329
R20499 VDD.n472 VDD.n471 212.329
R20500 VDD.n355 VDD.n354 212.329
R20501 VDD.n354 VDD.n347 212.329
R20502 VDD.n475 VDD.n346 212.329
R20503 VDD.n482 VDD.n346 212.329
R20504 VDD.n342 VDD.n341 212.329
R20505 VDD.n341 VDD.n337 212.329
R20506 VDD.n485 VDD.n336 212.329
R20507 VDD.n492 VDD.n336 212.329
R20508 VDD.n332 VDD.n331 212.329
R20509 VDD.n331 VDD.n326 212.329
R20510 VDD.n495 VDD.n325 212.329
R20511 VDD.n502 VDD.n325 212.329
R20512 VDD.n321 VDD.n320 212.329
R20513 VDD.n320 VDD.n313 212.329
R20514 VDD.n505 VDD.n312 212.329
R20515 VDD.n512 VDD.n312 212.329
R20516 VDD.n308 VDD.n307 212.329
R20517 VDD.n307 VDD.n303 212.329
R20518 VDD.n515 VDD.n302 212.329
R20519 VDD.n522 VDD.n302 212.329
R20520 VDD.n298 VDD.n297 212.329
R20521 VDD.n297 VDD.n292 212.329
R20522 VDD.n525 VDD.n291 212.329
R20523 VDD.n532 VDD.n291 212.329
R20524 VDD.n537 VDD.n284 212.329
R20525 VDD.n284 VDD.n282 212.329
R20526 VDD.n105 VDD.n104 212.329
R20527 VDD.n106 VDD.n105 212.329
R20528 VDD.n111 VDD.n94 212.329
R20529 VDD.n94 VDD.n92 212.329
R20530 VDD.n119 VDD.n118 212.329
R20531 VDD.n120 VDD.n119 212.329
R20532 VDD.n126 VDD.n125 212.329
R20533 VDD.n127 VDD.n126 212.329
R20534 VDD.n132 VDD.n78 212.329
R20535 VDD.n78 VDD.n76 212.329
R20536 VDD.n140 VDD.n139 212.329
R20537 VDD.n141 VDD.n140 212.329
R20538 VDD.n146 VDD.n69 212.329
R20539 VDD.n69 VDD.n67 212.329
R20540 VDD.n154 VDD.n153 212.329
R20541 VDD.n155 VDD.n154 212.329
R20542 VDD.n161 VDD.n160 212.329
R20543 VDD.n162 VDD.n161 212.329
R20544 VDD.n167 VDD.n53 212.329
R20545 VDD.n53 VDD.n51 212.329
R20546 VDD.n175 VDD.n174 212.329
R20547 VDD.n176 VDD.n175 212.329
R20548 VDD.n181 VDD.n44 212.329
R20549 VDD.n44 VDD.n42 212.329
R20550 VDD.n189 VDD.n188 212.329
R20551 VDD.n190 VDD.n189 212.329
R20552 VDD.n196 VDD.n195 212.329
R20553 VDD.n197 VDD.n196 212.329
R20554 VDD.n202 VDD.n28 212.329
R20555 VDD.n28 VDD.n26 212.329
R20556 VDD.n210 VDD.n209 212.329
R20557 VDD.n211 VDD.n210 212.329
R20558 VDD.n216 VDD.n19 212.329
R20559 VDD.n19 VDD.n17 212.329
R20560 VDD.n224 VDD.n223 212.329
R20561 VDD.n225 VDD.n224 212.329
R20562 VDD.n231 VDD.n230 212.329
R20563 VDD.n232 VDD.n231 212.329
R20564 VDD.n237 VDD.n3 212.329
R20565 VDD.n3 VDD.n1 212.329
R20566 VDD.n7333 VDD.n7332 212.329
R20567 VDD.n7332 VDD.n7325 212.329
R20568 VDD.n7334 VDD.n7324 212.329
R20569 VDD.n7341 VDD.n7324 212.329
R20570 VDD.n7320 VDD.n7319 212.329
R20571 VDD.n7319 VDD.n7315 212.329
R20572 VDD.n7344 VDD.n7314 212.329
R20573 VDD.n7351 VDD.n7314 212.329
R20574 VDD.n7310 VDD.n7309 212.329
R20575 VDD.n7309 VDD.n7304 212.329
R20576 VDD.n7354 VDD.n7303 212.329
R20577 VDD.n7361 VDD.n7303 212.329
R20578 VDD.n7299 VDD.n7298 212.329
R20579 VDD.n7298 VDD.n7291 212.329
R20580 VDD.n7364 VDD.n7290 212.329
R20581 VDD.n7371 VDD.n7290 212.329
R20582 VDD.n7286 VDD.n7285 212.329
R20583 VDD.n7285 VDD.n7279 212.329
R20584 VDD.n7374 VDD.n7278 212.329
R20585 VDD.n7381 VDD.n7278 212.329
R20586 VDD.n7387 VDD.n7386 212.329
R20587 VDD.n7388 VDD.n7387 212.329
R20588 VDD.n7271 VDD.n7270 212.329
R20589 VDD.n7270 VDD.n7263 212.329
R20590 VDD.n7391 VDD.n7262 212.329
R20591 VDD.n7398 VDD.n7262 212.329
R20592 VDD.n7258 VDD.n7257 212.329
R20593 VDD.n7257 VDD.n7253 212.329
R20594 VDD.n7401 VDD.n7252 212.329
R20595 VDD.n7408 VDD.n7252 212.329
R20596 VDD.n7248 VDD.n7247 212.329
R20597 VDD.n7247 VDD.n7242 212.329
R20598 VDD.n7411 VDD.n7241 212.329
R20599 VDD.n7418 VDD.n7241 212.329
R20600 VDD.n7237 VDD.n7236 212.329
R20601 VDD.n7236 VDD.n7229 212.329
R20602 VDD.n7421 VDD.n7228 212.329
R20603 VDD.n7428 VDD.n7228 212.329
R20604 VDD.n7224 VDD.n7223 212.329
R20605 VDD.n7223 VDD.n7219 212.329
R20606 VDD.n7431 VDD.n7218 212.329
R20607 VDD.n7438 VDD.n7218 212.329
R20608 VDD.n7214 VDD.n7213 212.329
R20609 VDD.n7213 VDD.n7208 212.329
R20610 VDD.n7441 VDD.n7207 212.329
R20611 VDD.n7448 VDD.n7207 212.329
R20612 VDD.n7453 VDD.n7200 212.329
R20613 VDD.n7200 VDD.n7198 212.329
R20614 VDD.n7193 VDD.n1844 212.329
R20615 VDD.n1844 VDD.n1842 212.329
R20616 VDD.n7076 VDD.n7075 212.329
R20617 VDD.n7075 VDD.n1974 212.329
R20618 VDD.n7077 VDD.n1973 212.329
R20619 VDD.n7084 VDD.n1973 212.329
R20620 VDD.n1969 VDD.n1968 212.329
R20621 VDD.n1968 VDD.n1964 212.329
R20622 VDD.n7087 VDD.n1963 212.329
R20623 VDD.n7094 VDD.n1963 212.329
R20624 VDD.n1959 VDD.n1958 212.329
R20625 VDD.n1958 VDD.n1953 212.329
R20626 VDD.n7097 VDD.n1952 212.329
R20627 VDD.n7104 VDD.n1952 212.329
R20628 VDD.n1948 VDD.n1947 212.329
R20629 VDD.n1947 VDD.n1940 212.329
R20630 VDD.n7107 VDD.n1939 212.329
R20631 VDD.n7114 VDD.n1939 212.329
R20632 VDD.n1935 VDD.n1934 212.329
R20633 VDD.n1934 VDD.n1928 212.329
R20634 VDD.n7117 VDD.n1927 212.329
R20635 VDD.n7124 VDD.n1927 212.329
R20636 VDD.n7130 VDD.n7129 212.329
R20637 VDD.n7131 VDD.n7130 212.329
R20638 VDD.n1919 VDD.n1918 212.329
R20639 VDD.n1919 VDD.n1917 212.329
R20640 VDD.n7139 VDD.n7138 212.329
R20641 VDD.n7139 VDD.n7137 212.329
R20642 VDD.n1911 VDD.n1910 212.329
R20643 VDD.n1910 VDD.n1898 212.329
R20644 VDD.n1893 VDD.n1892 212.329
R20645 VDD.n1892 VDD.n1886 212.329
R20646 VDD.n7151 VDD.n1885 212.329
R20647 VDD.n7158 VDD.n1885 212.329
R20648 VDD.n1881 VDD.n1880 212.329
R20649 VDD.n1880 VDD.n1873 212.329
R20650 VDD.n7161 VDD.n1872 212.329
R20651 VDD.n7168 VDD.n1872 212.329
R20652 VDD.n1868 VDD.n1867 212.329
R20653 VDD.n1867 VDD.n1863 212.329
R20654 VDD.n7171 VDD.n1862 212.329
R20655 VDD.n7178 VDD.n1862 212.329
R20656 VDD.n1858 VDD.n1857 212.329
R20657 VDD.n1857 VDD.n1852 212.329
R20658 VDD.n7181 VDD.n1851 212.329
R20659 VDD.n7188 VDD.n1851 212.329
R20660 VDD.n1913 VDD.n1897 212.329
R20661 VDD.n7148 VDD.n1897 212.329
R20662 VDD.n6939 VDD.n6938 212.329
R20663 VDD.n6940 VDD.n6939 212.329
R20664 VDD.n6945 VDD.n6928 212.329
R20665 VDD.n6928 VDD.n6926 212.329
R20666 VDD.n6953 VDD.n6952 212.329
R20667 VDD.n6954 VDD.n6953 212.329
R20668 VDD.n6960 VDD.n6959 212.329
R20669 VDD.n6961 VDD.n6960 212.329
R20670 VDD.n6966 VDD.n6912 212.329
R20671 VDD.n6912 VDD.n6910 212.329
R20672 VDD.n6974 VDD.n6973 212.329
R20673 VDD.n6975 VDD.n6974 212.329
R20674 VDD.n6980 VDD.n6903 212.329
R20675 VDD.n6903 VDD.n6901 212.329
R20676 VDD.n6988 VDD.n6987 212.329
R20677 VDD.n6989 VDD.n6988 212.329
R20678 VDD.n6995 VDD.n6994 212.329
R20679 VDD.n6996 VDD.n6995 212.329
R20680 VDD.n7001 VDD.n6887 212.329
R20681 VDD.n6887 VDD.n6885 212.329
R20682 VDD.n7009 VDD.n7008 212.329
R20683 VDD.n7010 VDD.n7009 212.329
R20684 VDD.n7015 VDD.n6878 212.329
R20685 VDD.n6878 VDD.n6876 212.329
R20686 VDD.n7023 VDD.n7022 212.329
R20687 VDD.n7024 VDD.n7023 212.329
R20688 VDD.n7030 VDD.n7029 212.329
R20689 VDD.n7031 VDD.n7030 212.329
R20690 VDD.n7036 VDD.n6862 212.329
R20691 VDD.n6862 VDD.n6860 212.329
R20692 VDD.n7044 VDD.n7043 212.329
R20693 VDD.n7045 VDD.n7044 212.329
R20694 VDD.n7050 VDD.n6853 212.329
R20695 VDD.n6853 VDD.n6851 212.329
R20696 VDD.n7058 VDD.n7057 212.329
R20697 VDD.n7059 VDD.n7058 212.329
R20698 VDD.n7063 VDD.n6832 212.329
R20699 VDD.n7063 VDD.n6831 212.329
R20700 VDD.n6843 VDD.n6842 212.329
R20701 VDD.n6842 VDD.n6841 212.329
R20702 VDD.n5964 VDD.n5961 212.329
R20703 VDD.n5969 VDD.n5961 212.329
R20704 VDD.n5958 VDD.n5957 212.329
R20705 VDD.n5957 VDD.n5953 212.329
R20706 VDD.n5972 VDD.n5952 212.329
R20707 VDD.n5979 VDD.n5952 212.329
R20708 VDD.n5948 VDD.n5947 212.329
R20709 VDD.n5947 VDD.n5940 212.329
R20710 VDD.n5982 VDD.n5939 212.329
R20711 VDD.n5989 VDD.n5939 212.329
R20712 VDD.n5935 VDD.n5934 212.329
R20713 VDD.n5934 VDD.n5929 212.329
R20714 VDD.n5992 VDD.n5928 212.329
R20715 VDD.n5999 VDD.n5928 212.329
R20716 VDD.n5924 VDD.n5923 212.329
R20717 VDD.n5923 VDD.n5919 212.329
R20718 VDD.n6002 VDD.n5918 212.329
R20719 VDD.n6009 VDD.n5918 212.329
R20720 VDD.n5914 VDD.n5913 212.329
R20721 VDD.n5913 VDD.n5906 212.329
R20722 VDD.n6012 VDD.n5905 212.329
R20723 VDD.n6019 VDD.n5905 212.329
R20724 VDD.n5901 VDD.n5900 212.329
R20725 VDD.n5900 VDD.n5894 212.329
R20726 VDD.n6022 VDD.n5893 212.329
R20727 VDD.n6029 VDD.n5893 212.329
R20728 VDD.n6035 VDD.n6034 212.329
R20729 VDD.n6036 VDD.n6035 212.329
R20730 VDD.n5886 VDD.n5885 212.329
R20731 VDD.n5885 VDD.n5878 212.329
R20732 VDD.n6039 VDD.n5877 212.329
R20733 VDD.n6046 VDD.n5877 212.329
R20734 VDD.n5873 VDD.n5872 212.329
R20735 VDD.n5872 VDD.n5867 212.329
R20736 VDD.n6049 VDD.n5866 212.329
R20737 VDD.n6056 VDD.n5866 212.329
R20738 VDD.n5862 VDD.n5861 212.329
R20739 VDD.n5861 VDD.n5857 212.329
R20740 VDD.n6059 VDD.n5856 212.329
R20741 VDD.n6066 VDD.n5856 212.329
R20742 VDD.n5852 VDD.n5851 212.329
R20743 VDD.n5851 VDD.n5847 212.329
R20744 VDD.n6069 VDD.n5846 212.329
R20745 VDD.n6076 VDD.n5846 212.329
R20746 VDD.n5841 VDD.n5840 212.329
R20747 VDD.n5841 VDD.n5839 212.329
R20748 VDD.n6084 VDD.n6083 212.329
R20749 VDD.n6084 VDD.n6082 212.329
R20750 VDD.n5828 VDD.n5825 212.329
R20751 VDD.n6092 VDD.n5825 212.329
R20752 VDD.n5822 VDD.n5821 212.329
R20753 VDD.n5821 VDD.n5817 212.329
R20754 VDD.n6095 VDD.n5816 212.329
R20755 VDD.n6102 VDD.n5816 212.329
R20756 VDD.n5812 VDD.n5811 212.329
R20757 VDD.n5811 VDD.n5804 212.329
R20758 VDD.n6105 VDD.n5803 212.329
R20759 VDD.n6112 VDD.n5803 212.329
R20760 VDD.n5799 VDD.n5798 212.329
R20761 VDD.n5798 VDD.n5793 212.329
R20762 VDD.n6115 VDD.n5792 212.329
R20763 VDD.n6122 VDD.n5792 212.329
R20764 VDD.n5788 VDD.n5787 212.329
R20765 VDD.n5787 VDD.n5783 212.329
R20766 VDD.n6125 VDD.n5782 212.329
R20767 VDD.n6132 VDD.n5782 212.329
R20768 VDD.n5778 VDD.n5777 212.329
R20769 VDD.n5777 VDD.n5770 212.329
R20770 VDD.n6135 VDD.n5769 212.329
R20771 VDD.n6142 VDD.n5769 212.329
R20772 VDD.n5765 VDD.n5764 212.329
R20773 VDD.n5764 VDD.n5758 212.329
R20774 VDD.n6145 VDD.n5757 212.329
R20775 VDD.n6152 VDD.n5757 212.329
R20776 VDD.n6158 VDD.n6157 212.329
R20777 VDD.n6159 VDD.n6158 212.329
R20778 VDD.n5750 VDD.n5749 212.329
R20779 VDD.n5749 VDD.n5742 212.329
R20780 VDD.n6162 VDD.n5741 212.329
R20781 VDD.n6169 VDD.n5741 212.329
R20782 VDD.n5737 VDD.n5736 212.329
R20783 VDD.n5736 VDD.n5731 212.329
R20784 VDD.n6172 VDD.n5730 212.329
R20785 VDD.n6179 VDD.n5730 212.329
R20786 VDD.n5726 VDD.n5725 212.329
R20787 VDD.n5725 VDD.n5721 212.329
R20788 VDD.n6182 VDD.n5720 212.329
R20789 VDD.n6189 VDD.n5720 212.329
R20790 VDD.n5716 VDD.n5715 212.329
R20791 VDD.n5715 VDD.n5711 212.329
R20792 VDD.n6192 VDD.n5710 212.329
R20793 VDD.n6199 VDD.n5710 212.329
R20794 VDD.n5705 VDD.n5704 212.329
R20795 VDD.n5705 VDD.n5703 212.329
R20796 VDD.n6207 VDD.n6206 212.329
R20797 VDD.n6207 VDD.n6205 212.329
R20798 VDD.n5692 VDD.n5689 212.329
R20799 VDD.n6215 VDD.n5689 212.329
R20800 VDD.n5686 VDD.n5685 212.329
R20801 VDD.n5685 VDD.n5681 212.329
R20802 VDD.n6218 VDD.n5680 212.329
R20803 VDD.n6225 VDD.n5680 212.329
R20804 VDD.n5676 VDD.n5675 212.329
R20805 VDD.n5675 VDD.n5668 212.329
R20806 VDD.n6228 VDD.n5667 212.329
R20807 VDD.n6235 VDD.n5667 212.329
R20808 VDD.n5663 VDD.n5662 212.329
R20809 VDD.n5662 VDD.n5657 212.329
R20810 VDD.n6238 VDD.n5656 212.329
R20811 VDD.n6245 VDD.n5656 212.329
R20812 VDD.n5652 VDD.n5651 212.329
R20813 VDD.n5651 VDD.n5647 212.329
R20814 VDD.n6248 VDD.n5646 212.329
R20815 VDD.n6255 VDD.n5646 212.329
R20816 VDD.n5642 VDD.n5641 212.329
R20817 VDD.n5641 VDD.n5634 212.329
R20818 VDD.n6258 VDD.n5633 212.329
R20819 VDD.n6265 VDD.n5633 212.329
R20820 VDD.n5629 VDD.n5628 212.329
R20821 VDD.n5628 VDD.n5622 212.329
R20822 VDD.n6268 VDD.n5621 212.329
R20823 VDD.n6275 VDD.n5621 212.329
R20824 VDD.n6281 VDD.n6280 212.329
R20825 VDD.n6282 VDD.n6281 212.329
R20826 VDD.n5614 VDD.n5613 212.329
R20827 VDD.n5613 VDD.n5606 212.329
R20828 VDD.n6285 VDD.n5605 212.329
R20829 VDD.n6292 VDD.n5605 212.329
R20830 VDD.n5601 VDD.n5600 212.329
R20831 VDD.n5600 VDD.n5595 212.329
R20832 VDD.n6295 VDD.n5594 212.329
R20833 VDD.n6302 VDD.n5594 212.329
R20834 VDD.n5590 VDD.n5589 212.329
R20835 VDD.n5589 VDD.n5585 212.329
R20836 VDD.n6305 VDD.n5584 212.329
R20837 VDD.n6312 VDD.n5584 212.329
R20838 VDD.n5580 VDD.n5579 212.329
R20839 VDD.n5579 VDD.n5575 212.329
R20840 VDD.n6315 VDD.n5574 212.329
R20841 VDD.n6322 VDD.n5574 212.329
R20842 VDD.n5569 VDD.n5568 212.329
R20843 VDD.n5569 VDD.n5567 212.329
R20844 VDD.n6330 VDD.n6329 212.329
R20845 VDD.n6330 VDD.n6328 212.329
R20846 VDD.n5556 VDD.n5553 212.329
R20847 VDD.n6338 VDD.n5553 212.329
R20848 VDD.n5550 VDD.n5549 212.329
R20849 VDD.n5549 VDD.n5545 212.329
R20850 VDD.n6341 VDD.n5544 212.329
R20851 VDD.n6348 VDD.n5544 212.329
R20852 VDD.n5540 VDD.n5539 212.329
R20853 VDD.n5539 VDD.n5532 212.329
R20854 VDD.n6351 VDD.n5531 212.329
R20855 VDD.n6358 VDD.n5531 212.329
R20856 VDD.n5527 VDD.n5526 212.329
R20857 VDD.n5526 VDD.n5521 212.329
R20858 VDD.n6361 VDD.n5520 212.329
R20859 VDD.n6368 VDD.n5520 212.329
R20860 VDD.n5516 VDD.n5515 212.329
R20861 VDD.n5515 VDD.n5511 212.329
R20862 VDD.n6371 VDD.n5510 212.329
R20863 VDD.n6378 VDD.n5510 212.329
R20864 VDD.n5506 VDD.n5505 212.329
R20865 VDD.n5505 VDD.n5498 212.329
R20866 VDD.n6381 VDD.n5497 212.329
R20867 VDD.n6388 VDD.n5497 212.329
R20868 VDD.n5493 VDD.n5492 212.329
R20869 VDD.n5492 VDD.n5486 212.329
R20870 VDD.n6391 VDD.n5485 212.329
R20871 VDD.n6398 VDD.n5485 212.329
R20872 VDD.n6404 VDD.n6403 212.329
R20873 VDD.n6405 VDD.n6404 212.329
R20874 VDD.n5478 VDD.n5477 212.329
R20875 VDD.n5477 VDD.n5470 212.329
R20876 VDD.n6408 VDD.n5469 212.329
R20877 VDD.n6415 VDD.n5469 212.329
R20878 VDD.n5465 VDD.n5464 212.329
R20879 VDD.n5464 VDD.n5459 212.329
R20880 VDD.n6418 VDD.n5458 212.329
R20881 VDD.n6425 VDD.n5458 212.329
R20882 VDD.n5454 VDD.n5453 212.329
R20883 VDD.n5453 VDD.n5449 212.329
R20884 VDD.n6428 VDD.n5448 212.329
R20885 VDD.n6435 VDD.n5448 212.329
R20886 VDD.n5444 VDD.n5443 212.329
R20887 VDD.n5443 VDD.n5439 212.329
R20888 VDD.n6438 VDD.n5438 212.329
R20889 VDD.n6445 VDD.n5438 212.329
R20890 VDD.n5433 VDD.n5432 212.329
R20891 VDD.n5433 VDD.n5431 212.329
R20892 VDD.n6453 VDD.n6452 212.329
R20893 VDD.n6453 VDD.n6451 212.329
R20894 VDD.n5420 VDD.n5417 212.329
R20895 VDD.n6461 VDD.n5417 212.329
R20896 VDD.n5414 VDD.n5413 212.329
R20897 VDD.n5413 VDD.n5409 212.329
R20898 VDD.n6464 VDD.n5408 212.329
R20899 VDD.n6471 VDD.n5408 212.329
R20900 VDD.n5404 VDD.n5403 212.329
R20901 VDD.n5403 VDD.n5396 212.329
R20902 VDD.n6474 VDD.n5395 212.329
R20903 VDD.n6481 VDD.n5395 212.329
R20904 VDD.n5391 VDD.n5390 212.329
R20905 VDD.n5390 VDD.n5385 212.329
R20906 VDD.n6484 VDD.n5384 212.329
R20907 VDD.n6491 VDD.n5384 212.329
R20908 VDD.n5380 VDD.n5379 212.329
R20909 VDD.n5379 VDD.n5375 212.329
R20910 VDD.n6494 VDD.n5374 212.329
R20911 VDD.n6501 VDD.n5374 212.329
R20912 VDD.n5370 VDD.n5369 212.329
R20913 VDD.n5369 VDD.n5362 212.329
R20914 VDD.n6504 VDD.n5361 212.329
R20915 VDD.n6511 VDD.n5361 212.329
R20916 VDD.n5357 VDD.n5356 212.329
R20917 VDD.n5356 VDD.n5350 212.329
R20918 VDD.n6514 VDD.n5349 212.329
R20919 VDD.n6521 VDD.n5349 212.329
R20920 VDD.n6527 VDD.n6526 212.329
R20921 VDD.n6528 VDD.n6527 212.329
R20922 VDD.n5342 VDD.n5341 212.329
R20923 VDD.n5341 VDD.n5334 212.329
R20924 VDD.n6531 VDD.n5333 212.329
R20925 VDD.n6538 VDD.n5333 212.329
R20926 VDD.n5329 VDD.n5328 212.329
R20927 VDD.n5328 VDD.n5323 212.329
R20928 VDD.n6541 VDD.n5322 212.329
R20929 VDD.n6548 VDD.n5322 212.329
R20930 VDD.n5318 VDD.n5317 212.329
R20931 VDD.n5317 VDD.n5313 212.329
R20932 VDD.n6551 VDD.n5312 212.329
R20933 VDD.n6558 VDD.n5312 212.329
R20934 VDD.n5308 VDD.n5307 212.329
R20935 VDD.n5307 VDD.n5303 212.329
R20936 VDD.n6561 VDD.n5302 212.329
R20937 VDD.n6568 VDD.n5302 212.329
R20938 VDD.n5297 VDD.n5296 212.329
R20939 VDD.n5297 VDD.n5295 212.329
R20940 VDD.n6576 VDD.n6575 212.329
R20941 VDD.n6576 VDD.n6574 212.329
R20942 VDD.n5284 VDD.n5281 212.329
R20943 VDD.n6584 VDD.n5281 212.329
R20944 VDD.n5278 VDD.n5277 212.329
R20945 VDD.n5277 VDD.n5273 212.329
R20946 VDD.n6587 VDD.n5272 212.329
R20947 VDD.n6594 VDD.n5272 212.329
R20948 VDD.n5268 VDD.n5267 212.329
R20949 VDD.n5267 VDD.n5260 212.329
R20950 VDD.n6597 VDD.n5259 212.329
R20951 VDD.n6604 VDD.n5259 212.329
R20952 VDD.n5255 VDD.n5254 212.329
R20953 VDD.n5254 VDD.n5249 212.329
R20954 VDD.n6607 VDD.n5248 212.329
R20955 VDD.n6614 VDD.n5248 212.329
R20956 VDD.n5244 VDD.n5243 212.329
R20957 VDD.n5243 VDD.n5239 212.329
R20958 VDD.n6617 VDD.n5238 212.329
R20959 VDD.n6624 VDD.n5238 212.329
R20960 VDD.n5234 VDD.n5233 212.329
R20961 VDD.n5233 VDD.n5226 212.329
R20962 VDD.n6627 VDD.n5225 212.329
R20963 VDD.n6634 VDD.n5225 212.329
R20964 VDD.n5221 VDD.n5220 212.329
R20965 VDD.n5220 VDD.n5214 212.329
R20966 VDD.n6637 VDD.n5213 212.329
R20967 VDD.n6644 VDD.n5213 212.329
R20968 VDD.n6650 VDD.n6649 212.329
R20969 VDD.n6651 VDD.n6650 212.329
R20970 VDD.n5206 VDD.n5205 212.329
R20971 VDD.n5205 VDD.n5198 212.329
R20972 VDD.n6654 VDD.n5197 212.329
R20973 VDD.n6661 VDD.n5197 212.329
R20974 VDD.n5193 VDD.n5192 212.329
R20975 VDD.n5192 VDD.n5187 212.329
R20976 VDD.n6664 VDD.n5186 212.329
R20977 VDD.n6671 VDD.n5186 212.329
R20978 VDD.n5182 VDD.n5181 212.329
R20979 VDD.n5181 VDD.n5177 212.329
R20980 VDD.n6674 VDD.n5176 212.329
R20981 VDD.n6681 VDD.n5176 212.329
R20982 VDD.n5172 VDD.n5171 212.329
R20983 VDD.n5171 VDD.n5167 212.329
R20984 VDD.n6684 VDD.n5166 212.329
R20985 VDD.n6691 VDD.n5166 212.329
R20986 VDD.n5161 VDD.n5160 212.329
R20987 VDD.n5161 VDD.n5159 212.329
R20988 VDD.n6699 VDD.n6698 212.329
R20989 VDD.n6699 VDD.n6697 212.329
R20990 VDD.n5148 VDD.n5145 212.329
R20991 VDD.n6707 VDD.n5145 212.329
R20992 VDD.n5142 VDD.n5141 212.329
R20993 VDD.n5141 VDD.n5137 212.329
R20994 VDD.n6710 VDD.n5136 212.329
R20995 VDD.n6717 VDD.n5136 212.329
R20996 VDD.n5132 VDD.n5131 212.329
R20997 VDD.n5131 VDD.n5124 212.329
R20998 VDD.n6720 VDD.n5123 212.329
R20999 VDD.n6727 VDD.n5123 212.329
R21000 VDD.n5119 VDD.n5118 212.329
R21001 VDD.n5118 VDD.n5113 212.329
R21002 VDD.n6730 VDD.n5112 212.329
R21003 VDD.n6737 VDD.n5112 212.329
R21004 VDD.n5108 VDD.n5107 212.329
R21005 VDD.n5107 VDD.n5103 212.329
R21006 VDD.n6740 VDD.n5102 212.329
R21007 VDD.n6747 VDD.n5102 212.329
R21008 VDD.n5098 VDD.n5097 212.329
R21009 VDD.n5097 VDD.n5090 212.329
R21010 VDD.n6750 VDD.n5089 212.329
R21011 VDD.n6757 VDD.n5089 212.329
R21012 VDD.n5085 VDD.n5084 212.329
R21013 VDD.n5084 VDD.n5078 212.329
R21014 VDD.n6760 VDD.n5077 212.329
R21015 VDD.n6767 VDD.n5077 212.329
R21016 VDD.n6773 VDD.n6772 212.329
R21017 VDD.n6774 VDD.n6773 212.329
R21018 VDD.n5070 VDD.n5069 212.329
R21019 VDD.n5069 VDD.n5062 212.329
R21020 VDD.n6777 VDD.n5061 212.329
R21021 VDD.n6784 VDD.n5061 212.329
R21022 VDD.n5057 VDD.n5056 212.329
R21023 VDD.n5056 VDD.n5051 212.329
R21024 VDD.n6787 VDD.n5050 212.329
R21025 VDD.n6794 VDD.n5050 212.329
R21026 VDD.n5046 VDD.n5045 212.329
R21027 VDD.n5045 VDD.n5041 212.329
R21028 VDD.n6797 VDD.n5040 212.329
R21029 VDD.n6804 VDD.n5040 212.329
R21030 VDD.n5036 VDD.n5035 212.329
R21031 VDD.n5035 VDD.n5031 212.329
R21032 VDD.n6807 VDD.n5030 212.329
R21033 VDD.n6814 VDD.n5030 212.329
R21034 VDD.n5025 VDD.n5024 212.329
R21035 VDD.n5025 VDD.n5023 212.329
R21036 VDD.n6822 VDD.n6821 212.329
R21037 VDD.n6822 VDD.n6820 212.329
R21038 VDD.n5010 VDD.n4758 212.329
R21039 VDD.n4758 VDD.n4756 212.329
R21040 VDD.n4769 VDD.n4764 212.329
R21041 VDD.n4770 VDD.n4769 212.329
R21042 VDD.n5003 VDD.n4763 212.329
R21043 VDD.n4996 VDD.n4763 212.329
R21044 VDD.n4779 VDD.n4775 212.329
R21045 VDD.n4780 VDD.n4779 212.329
R21046 VDD.n4993 VDD.n4774 212.329
R21047 VDD.n4986 VDD.n4774 212.329
R21048 VDD.n4792 VDD.n4785 212.329
R21049 VDD.n4793 VDD.n4792 212.329
R21050 VDD.n4983 VDD.n4784 212.329
R21051 VDD.n4976 VDD.n4784 212.329
R21052 VDD.n4803 VDD.n4798 212.329
R21053 VDD.n4804 VDD.n4803 212.329
R21054 VDD.n4973 VDD.n4797 212.329
R21055 VDD.n4966 VDD.n4797 212.329
R21056 VDD.n4813 VDD.n4809 212.329
R21057 VDD.n4814 VDD.n4813 212.329
R21058 VDD.n4963 VDD.n4808 212.329
R21059 VDD.n4956 VDD.n4808 212.329
R21060 VDD.n4826 VDD.n4819 212.329
R21061 VDD.n4827 VDD.n4826 212.329
R21062 VDD.n4953 VDD.n4818 212.329
R21063 VDD.n4946 VDD.n4818 212.329
R21064 VDD.n4943 VDD.n4942 212.329
R21065 VDD.n4942 VDD.n4941 212.329
R21066 VDD.n4841 VDD.n4835 212.329
R21067 VDD.n4842 VDD.n4841 212.329
R21068 VDD.n4936 VDD.n4834 212.329
R21069 VDD.n4929 VDD.n4834 212.329
R21070 VDD.n4854 VDD.n4847 212.329
R21071 VDD.n4855 VDD.n4854 212.329
R21072 VDD.n4926 VDD.n4846 212.329
R21073 VDD.n4919 VDD.n4846 212.329
R21074 VDD.n4865 VDD.n4860 212.329
R21075 VDD.n4866 VDD.n4865 212.329
R21076 VDD.n4916 VDD.n4859 212.329
R21077 VDD.n4909 VDD.n4859 212.329
R21078 VDD.n4875 VDD.n4871 212.329
R21079 VDD.n4876 VDD.n4875 212.329
R21080 VDD.n4906 VDD.n4870 212.329
R21081 VDD.n4899 VDD.n4870 212.329
R21082 VDD.n4884 VDD.n4881 212.329
R21083 VDD.n4885 VDD.n4884 212.329
R21084 VDD.n4896 VDD.n4880 212.329
R21085 VDD.n4886 VDD.n4880 212.329
R21086 VDD.n4752 VDD.n1980 212.329
R21087 VDD.n1980 VDD.n1978 212.329
R21088 VDD.n4635 VDD.n4634 212.329
R21089 VDD.n4634 VDD.n2110 212.329
R21090 VDD.n4636 VDD.n2109 212.329
R21091 VDD.n4643 VDD.n2109 212.329
R21092 VDD.n2105 VDD.n2104 212.329
R21093 VDD.n2104 VDD.n2100 212.329
R21094 VDD.n4646 VDD.n2099 212.329
R21095 VDD.n4653 VDD.n2099 212.329
R21096 VDD.n2095 VDD.n2094 212.329
R21097 VDD.n2094 VDD.n2089 212.329
R21098 VDD.n4656 VDD.n2088 212.329
R21099 VDD.n4663 VDD.n2088 212.329
R21100 VDD.n2084 VDD.n2083 212.329
R21101 VDD.n2083 VDD.n2076 212.329
R21102 VDD.n4666 VDD.n2075 212.329
R21103 VDD.n4673 VDD.n2075 212.329
R21104 VDD.n2071 VDD.n2070 212.329
R21105 VDD.n2070 VDD.n2064 212.329
R21106 VDD.n4676 VDD.n2063 212.329
R21107 VDD.n4683 VDD.n2063 212.329
R21108 VDD.n4689 VDD.n4688 212.329
R21109 VDD.n4690 VDD.n4689 212.329
R21110 VDD.n2055 VDD.n2054 212.329
R21111 VDD.n2055 VDD.n2053 212.329
R21112 VDD.n4698 VDD.n4697 212.329
R21113 VDD.n4698 VDD.n4696 212.329
R21114 VDD.n2047 VDD.n2046 212.329
R21115 VDD.n2046 VDD.n2034 212.329
R21116 VDD.n2029 VDD.n2028 212.329
R21117 VDD.n2028 VDD.n2022 212.329
R21118 VDD.n4710 VDD.n2021 212.329
R21119 VDD.n4717 VDD.n2021 212.329
R21120 VDD.n2017 VDD.n2016 212.329
R21121 VDD.n2016 VDD.n2009 212.329
R21122 VDD.n4720 VDD.n2008 212.329
R21123 VDD.n4727 VDD.n2008 212.329
R21124 VDD.n2004 VDD.n2003 212.329
R21125 VDD.n2003 VDD.n1999 212.329
R21126 VDD.n4730 VDD.n1998 212.329
R21127 VDD.n4737 VDD.n1998 212.329
R21128 VDD.n1994 VDD.n1993 212.329
R21129 VDD.n1993 VDD.n1988 212.329
R21130 VDD.n4740 VDD.n1987 212.329
R21131 VDD.n4747 VDD.n1987 212.329
R21132 VDD.n2049 VDD.n2033 212.329
R21133 VDD.n4707 VDD.n2033 212.329
R21134 VDD.n4627 VDD.n2116 212.329
R21135 VDD.n2116 VDD.n2114 212.329
R21136 VDD.n4510 VDD.n4509 212.329
R21137 VDD.n4509 VDD.n2246 212.329
R21138 VDD.n4511 VDD.n2245 212.329
R21139 VDD.n4518 VDD.n2245 212.329
R21140 VDD.n2241 VDD.n2240 212.329
R21141 VDD.n2240 VDD.n2236 212.329
R21142 VDD.n4521 VDD.n2235 212.329
R21143 VDD.n4528 VDD.n2235 212.329
R21144 VDD.n2231 VDD.n2230 212.329
R21145 VDD.n2230 VDD.n2225 212.329
R21146 VDD.n4531 VDD.n2224 212.329
R21147 VDD.n4538 VDD.n2224 212.329
R21148 VDD.n2220 VDD.n2219 212.329
R21149 VDD.n2219 VDD.n2212 212.329
R21150 VDD.n4541 VDD.n2211 212.329
R21151 VDD.n4548 VDD.n2211 212.329
R21152 VDD.n2207 VDD.n2206 212.329
R21153 VDD.n2206 VDD.n2200 212.329
R21154 VDD.n4551 VDD.n2199 212.329
R21155 VDD.n4558 VDD.n2199 212.329
R21156 VDD.n4564 VDD.n4563 212.329
R21157 VDD.n4565 VDD.n4564 212.329
R21158 VDD.n2191 VDD.n2190 212.329
R21159 VDD.n2191 VDD.n2189 212.329
R21160 VDD.n4573 VDD.n4572 212.329
R21161 VDD.n4573 VDD.n4571 212.329
R21162 VDD.n2183 VDD.n2182 212.329
R21163 VDD.n2182 VDD.n2170 212.329
R21164 VDD.n2165 VDD.n2164 212.329
R21165 VDD.n2164 VDD.n2158 212.329
R21166 VDD.n4585 VDD.n2157 212.329
R21167 VDD.n4592 VDD.n2157 212.329
R21168 VDD.n2153 VDD.n2152 212.329
R21169 VDD.n2152 VDD.n2145 212.329
R21170 VDD.n4595 VDD.n2144 212.329
R21171 VDD.n4602 VDD.n2144 212.329
R21172 VDD.n2140 VDD.n2139 212.329
R21173 VDD.n2139 VDD.n2135 212.329
R21174 VDD.n4605 VDD.n2134 212.329
R21175 VDD.n4612 VDD.n2134 212.329
R21176 VDD.n2130 VDD.n2129 212.329
R21177 VDD.n2129 VDD.n2124 212.329
R21178 VDD.n4615 VDD.n2123 212.329
R21179 VDD.n4622 VDD.n2123 212.329
R21180 VDD.n2185 VDD.n2169 212.329
R21181 VDD.n4582 VDD.n2169 212.329
R21182 VDD.n4502 VDD.n2252 212.329
R21183 VDD.n2252 VDD.n2250 212.329
R21184 VDD.n4385 VDD.n4384 212.329
R21185 VDD.n4384 VDD.n2382 212.329
R21186 VDD.n4386 VDD.n2381 212.329
R21187 VDD.n4393 VDD.n2381 212.329
R21188 VDD.n2377 VDD.n2376 212.329
R21189 VDD.n2376 VDD.n2372 212.329
R21190 VDD.n4396 VDD.n2371 212.329
R21191 VDD.n4403 VDD.n2371 212.329
R21192 VDD.n2367 VDD.n2366 212.329
R21193 VDD.n2366 VDD.n2361 212.329
R21194 VDD.n4406 VDD.n2360 212.329
R21195 VDD.n4413 VDD.n2360 212.329
R21196 VDD.n2356 VDD.n2355 212.329
R21197 VDD.n2355 VDD.n2348 212.329
R21198 VDD.n4416 VDD.n2347 212.329
R21199 VDD.n4423 VDD.n2347 212.329
R21200 VDD.n2343 VDD.n2342 212.329
R21201 VDD.n2342 VDD.n2336 212.329
R21202 VDD.n4426 VDD.n2335 212.329
R21203 VDD.n4433 VDD.n2335 212.329
R21204 VDD.n4439 VDD.n4438 212.329
R21205 VDD.n4440 VDD.n4439 212.329
R21206 VDD.n2327 VDD.n2326 212.329
R21207 VDD.n2327 VDD.n2325 212.329
R21208 VDD.n4448 VDD.n4447 212.329
R21209 VDD.n4448 VDD.n4446 212.329
R21210 VDD.n2319 VDD.n2318 212.329
R21211 VDD.n2318 VDD.n2306 212.329
R21212 VDD.n2301 VDD.n2300 212.329
R21213 VDD.n2300 VDD.n2294 212.329
R21214 VDD.n4460 VDD.n2293 212.329
R21215 VDD.n4467 VDD.n2293 212.329
R21216 VDD.n2289 VDD.n2288 212.329
R21217 VDD.n2288 VDD.n2281 212.329
R21218 VDD.n4470 VDD.n2280 212.329
R21219 VDD.n4477 VDD.n2280 212.329
R21220 VDD.n2276 VDD.n2275 212.329
R21221 VDD.n2275 VDD.n2271 212.329
R21222 VDD.n4480 VDD.n2270 212.329
R21223 VDD.n4487 VDD.n2270 212.329
R21224 VDD.n2266 VDD.n2265 212.329
R21225 VDD.n2265 VDD.n2260 212.329
R21226 VDD.n4490 VDD.n2259 212.329
R21227 VDD.n4497 VDD.n2259 212.329
R21228 VDD.n2321 VDD.n2305 212.329
R21229 VDD.n4457 VDD.n2305 212.329
R21230 VDD.n4377 VDD.n2388 212.329
R21231 VDD.n2388 VDD.n2386 212.329
R21232 VDD.n4260 VDD.n4259 212.329
R21233 VDD.n4259 VDD.n2518 212.329
R21234 VDD.n4261 VDD.n2517 212.329
R21235 VDD.n4268 VDD.n2517 212.329
R21236 VDD.n2513 VDD.n2512 212.329
R21237 VDD.n2512 VDD.n2508 212.329
R21238 VDD.n4271 VDD.n2507 212.329
R21239 VDD.n4278 VDD.n2507 212.329
R21240 VDD.n2503 VDD.n2502 212.329
R21241 VDD.n2502 VDD.n2497 212.329
R21242 VDD.n4281 VDD.n2496 212.329
R21243 VDD.n4288 VDD.n2496 212.329
R21244 VDD.n2492 VDD.n2491 212.329
R21245 VDD.n2491 VDD.n2484 212.329
R21246 VDD.n4291 VDD.n2483 212.329
R21247 VDD.n4298 VDD.n2483 212.329
R21248 VDD.n2479 VDD.n2478 212.329
R21249 VDD.n2478 VDD.n2472 212.329
R21250 VDD.n4301 VDD.n2471 212.329
R21251 VDD.n4308 VDD.n2471 212.329
R21252 VDD.n4314 VDD.n4313 212.329
R21253 VDD.n4315 VDD.n4314 212.329
R21254 VDD.n2463 VDD.n2462 212.329
R21255 VDD.n2463 VDD.n2461 212.329
R21256 VDD.n4323 VDD.n4322 212.329
R21257 VDD.n4323 VDD.n4321 212.329
R21258 VDD.n2455 VDD.n2454 212.329
R21259 VDD.n2454 VDD.n2442 212.329
R21260 VDD.n2437 VDD.n2436 212.329
R21261 VDD.n2436 VDD.n2430 212.329
R21262 VDD.n4335 VDD.n2429 212.329
R21263 VDD.n4342 VDD.n2429 212.329
R21264 VDD.n2425 VDD.n2424 212.329
R21265 VDD.n2424 VDD.n2417 212.329
R21266 VDD.n4345 VDD.n2416 212.329
R21267 VDD.n4352 VDD.n2416 212.329
R21268 VDD.n2412 VDD.n2411 212.329
R21269 VDD.n2411 VDD.n2407 212.329
R21270 VDD.n4355 VDD.n2406 212.329
R21271 VDD.n4362 VDD.n2406 212.329
R21272 VDD.n2402 VDD.n2401 212.329
R21273 VDD.n2401 VDD.n2396 212.329
R21274 VDD.n4365 VDD.n2395 212.329
R21275 VDD.n4372 VDD.n2395 212.329
R21276 VDD.n2457 VDD.n2441 212.329
R21277 VDD.n4332 VDD.n2441 212.329
R21278 VDD.n4252 VDD.n2524 212.329
R21279 VDD.n2524 VDD.n2522 212.329
R21280 VDD.n4135 VDD.n4134 212.329
R21281 VDD.n4134 VDD.n2654 212.329
R21282 VDD.n4136 VDD.n2653 212.329
R21283 VDD.n4143 VDD.n2653 212.329
R21284 VDD.n2649 VDD.n2648 212.329
R21285 VDD.n2648 VDD.n2644 212.329
R21286 VDD.n4146 VDD.n2643 212.329
R21287 VDD.n4153 VDD.n2643 212.329
R21288 VDD.n2639 VDD.n2638 212.329
R21289 VDD.n2638 VDD.n2633 212.329
R21290 VDD.n4156 VDD.n2632 212.329
R21291 VDD.n4163 VDD.n2632 212.329
R21292 VDD.n2628 VDD.n2627 212.329
R21293 VDD.n2627 VDD.n2620 212.329
R21294 VDD.n4166 VDD.n2619 212.329
R21295 VDD.n4173 VDD.n2619 212.329
R21296 VDD.n2615 VDD.n2614 212.329
R21297 VDD.n2614 VDD.n2608 212.329
R21298 VDD.n4176 VDD.n2607 212.329
R21299 VDD.n4183 VDD.n2607 212.329
R21300 VDD.n4189 VDD.n4188 212.329
R21301 VDD.n4190 VDD.n4189 212.329
R21302 VDD.n2599 VDD.n2598 212.329
R21303 VDD.n2599 VDD.n2597 212.329
R21304 VDD.n4198 VDD.n4197 212.329
R21305 VDD.n4198 VDD.n4196 212.329
R21306 VDD.n2591 VDD.n2590 212.329
R21307 VDD.n2590 VDD.n2578 212.329
R21308 VDD.n2573 VDD.n2572 212.329
R21309 VDD.n2572 VDD.n2566 212.329
R21310 VDD.n4210 VDD.n2565 212.329
R21311 VDD.n4217 VDD.n2565 212.329
R21312 VDD.n2561 VDD.n2560 212.329
R21313 VDD.n2560 VDD.n2553 212.329
R21314 VDD.n4220 VDD.n2552 212.329
R21315 VDD.n4227 VDD.n2552 212.329
R21316 VDD.n2548 VDD.n2547 212.329
R21317 VDD.n2547 VDD.n2543 212.329
R21318 VDD.n4230 VDD.n2542 212.329
R21319 VDD.n4237 VDD.n2542 212.329
R21320 VDD.n2538 VDD.n2537 212.329
R21321 VDD.n2537 VDD.n2532 212.329
R21322 VDD.n4240 VDD.n2531 212.329
R21323 VDD.n4247 VDD.n2531 212.329
R21324 VDD.n2593 VDD.n2577 212.329
R21325 VDD.n4207 VDD.n2577 212.329
R21326 VDD.n4127 VDD.n2660 212.329
R21327 VDD.n2660 VDD.n2658 212.329
R21328 VDD.n4010 VDD.n4009 212.329
R21329 VDD.n4009 VDD.n2790 212.329
R21330 VDD.n4011 VDD.n2789 212.329
R21331 VDD.n4018 VDD.n2789 212.329
R21332 VDD.n2785 VDD.n2784 212.329
R21333 VDD.n2784 VDD.n2780 212.329
R21334 VDD.n4021 VDD.n2779 212.329
R21335 VDD.n4028 VDD.n2779 212.329
R21336 VDD.n2775 VDD.n2774 212.329
R21337 VDD.n2774 VDD.n2769 212.329
R21338 VDD.n4031 VDD.n2768 212.329
R21339 VDD.n4038 VDD.n2768 212.329
R21340 VDD.n2764 VDD.n2763 212.329
R21341 VDD.n2763 VDD.n2756 212.329
R21342 VDD.n4041 VDD.n2755 212.329
R21343 VDD.n4048 VDD.n2755 212.329
R21344 VDD.n2751 VDD.n2750 212.329
R21345 VDD.n2750 VDD.n2744 212.329
R21346 VDD.n4051 VDD.n2743 212.329
R21347 VDD.n4058 VDD.n2743 212.329
R21348 VDD.n4064 VDD.n4063 212.329
R21349 VDD.n4065 VDD.n4064 212.329
R21350 VDD.n2735 VDD.n2734 212.329
R21351 VDD.n2735 VDD.n2733 212.329
R21352 VDD.n4073 VDD.n4072 212.329
R21353 VDD.n4073 VDD.n4071 212.329
R21354 VDD.n2727 VDD.n2726 212.329
R21355 VDD.n2726 VDD.n2714 212.329
R21356 VDD.n2709 VDD.n2708 212.329
R21357 VDD.n2708 VDD.n2702 212.329
R21358 VDD.n4085 VDD.n2701 212.329
R21359 VDD.n4092 VDD.n2701 212.329
R21360 VDD.n2697 VDD.n2696 212.329
R21361 VDD.n2696 VDD.n2689 212.329
R21362 VDD.n4095 VDD.n2688 212.329
R21363 VDD.n4102 VDD.n2688 212.329
R21364 VDD.n2684 VDD.n2683 212.329
R21365 VDD.n2683 VDD.n2679 212.329
R21366 VDD.n4105 VDD.n2678 212.329
R21367 VDD.n4112 VDD.n2678 212.329
R21368 VDD.n2674 VDD.n2673 212.329
R21369 VDD.n2673 VDD.n2668 212.329
R21370 VDD.n4115 VDD.n2667 212.329
R21371 VDD.n4122 VDD.n2667 212.329
R21372 VDD.n2729 VDD.n2713 212.329
R21373 VDD.n4082 VDD.n2713 212.329
R21374 VDD.n4002 VDD.n2796 212.329
R21375 VDD.n2796 VDD.n2794 212.329
R21376 VDD.n3885 VDD.n3884 212.329
R21377 VDD.n3884 VDD.n2926 212.329
R21378 VDD.n3886 VDD.n2925 212.329
R21379 VDD.n3893 VDD.n2925 212.329
R21380 VDD.n2921 VDD.n2920 212.329
R21381 VDD.n2920 VDD.n2916 212.329
R21382 VDD.n3896 VDD.n2915 212.329
R21383 VDD.n3903 VDD.n2915 212.329
R21384 VDD.n2911 VDD.n2910 212.329
R21385 VDD.n2910 VDD.n2905 212.329
R21386 VDD.n3906 VDD.n2904 212.329
R21387 VDD.n3913 VDD.n2904 212.329
R21388 VDD.n2900 VDD.n2899 212.329
R21389 VDD.n2899 VDD.n2892 212.329
R21390 VDD.n3916 VDD.n2891 212.329
R21391 VDD.n3923 VDD.n2891 212.329
R21392 VDD.n2887 VDD.n2886 212.329
R21393 VDD.n2886 VDD.n2880 212.329
R21394 VDD.n3926 VDD.n2879 212.329
R21395 VDD.n3933 VDD.n2879 212.329
R21396 VDD.n3939 VDD.n3938 212.329
R21397 VDD.n3940 VDD.n3939 212.329
R21398 VDD.n2871 VDD.n2870 212.329
R21399 VDD.n2871 VDD.n2869 212.329
R21400 VDD.n3948 VDD.n3947 212.329
R21401 VDD.n3948 VDD.n3946 212.329
R21402 VDD.n2863 VDD.n2862 212.329
R21403 VDD.n2862 VDD.n2850 212.329
R21404 VDD.n2845 VDD.n2844 212.329
R21405 VDD.n2844 VDD.n2838 212.329
R21406 VDD.n3960 VDD.n2837 212.329
R21407 VDD.n3967 VDD.n2837 212.329
R21408 VDD.n2833 VDD.n2832 212.329
R21409 VDD.n2832 VDD.n2825 212.329
R21410 VDD.n3970 VDD.n2824 212.329
R21411 VDD.n3977 VDD.n2824 212.329
R21412 VDD.n2820 VDD.n2819 212.329
R21413 VDD.n2819 VDD.n2815 212.329
R21414 VDD.n3980 VDD.n2814 212.329
R21415 VDD.n3987 VDD.n2814 212.329
R21416 VDD.n2810 VDD.n2809 212.329
R21417 VDD.n2809 VDD.n2804 212.329
R21418 VDD.n3990 VDD.n2803 212.329
R21419 VDD.n3997 VDD.n2803 212.329
R21420 VDD.n2865 VDD.n2849 212.329
R21421 VDD.n3957 VDD.n2849 212.329
R21422 VDD.n3234 VDD.n3233 212.329
R21423 VDD.n3233 VDD.n3230 212.329
R21424 VDD.n3225 VDD.n3224 212.329
R21425 VDD.n3224 VDD.n3220 212.329
R21426 VDD.n3538 VDD.n3219 212.329
R21427 VDD.n3545 VDD.n3219 212.329
R21428 VDD.n3214 VDD.n3213 212.329
R21429 VDD.n3214 VDD.n3212 212.329
R21430 VDD.n3553 VDD.n3552 212.329
R21431 VDD.n3553 VDD.n3551 212.329
R21432 VDD.n3235 VDD.n3229 212.329
R21433 VDD.n3535 VDD.n3229 212.329
R21434 VDD.n3387 VDD.n3285 212.329
R21435 VDD.n3285 VDD.n3283 212.329
R21436 VDD.n3380 VDD.n3289 212.329
R21437 VDD.n3290 VDD.n3289 212.329
R21438 VDD.n3373 VDD.n3365 212.329
R21439 VDD.n3365 VDD.n3363 212.329
R21440 VDD.n3424 VDD.n3394 212.329
R21441 VDD.n3394 VDD.n3392 212.329
R21442 VDD.n3417 VDD.n3398 212.329
R21443 VDD.n3399 VDD.n3398 212.329
R21444 VDD.n3411 VDD.n3403 212.329
R21445 VDD.n3403 VDD.n3401 212.329
R21446 VDD.n3276 VDD.n3268 212.329
R21447 VDD.n3268 VDD.n3266 212.329
R21448 VDD.n3265 VDD.n3264 212.329
R21449 VDD.n3446 VDD.n3264 212.329
R21450 VDD.n3451 VDD.n3258 212.329
R21451 VDD.n3258 VDD.n3256 212.329
R21452 VDD.n3482 VDD.n3248 212.329
R21453 VDD.n3248 VDD.n3246 212.329
R21454 VDD.n3475 VDD.n3252 212.329
R21455 VDD.n3253 VDD.n3252 212.329
R21456 VDD.n3468 VDD.n3460 212.329
R21457 VDD.n3460 VDD.n3458 212.329
R21458 VDD.n3518 VDD.n3488 212.329
R21459 VDD.n3488 VDD.n3486 212.329
R21460 VDD.n3511 VDD.n3492 212.329
R21461 VDD.n3493 VDD.n3492 212.329
R21462 VDD.n3505 VDD.n3497 212.329
R21463 VDD.n3497 VDD.n3495 212.329
R21464 VDD.n3332 VDD.n3324 212.329
R21465 VDD.n3324 VDD.n3322 212.329
R21466 VDD.n3321 VDD.n3320 212.329
R21467 VDD.n3351 VDD.n3320 212.329
R21468 VDD.n3356 VDD.n3314 212.329
R21469 VDD.n3314 VDD.n3312 212.329
R21470 VDD.n3877 VDD.n2932 212.329
R21471 VDD.n2932 VDD.n2930 212.329
R21472 VDD.n3760 VDD.n3759 212.329
R21473 VDD.n3759 VDD.n3752 212.329
R21474 VDD.n3761 VDD.n3751 212.329
R21475 VDD.n3768 VDD.n3751 212.329
R21476 VDD.n3747 VDD.n3746 212.329
R21477 VDD.n3746 VDD.n3742 212.329
R21478 VDD.n3771 VDD.n3741 212.329
R21479 VDD.n3778 VDD.n3741 212.329
R21480 VDD.n3737 VDD.n3736 212.329
R21481 VDD.n3736 VDD.n3731 212.329
R21482 VDD.n3781 VDD.n3730 212.329
R21483 VDD.n3788 VDD.n3730 212.329
R21484 VDD.n3726 VDD.n3725 212.329
R21485 VDD.n3725 VDD.n3718 212.329
R21486 VDD.n3791 VDD.n3717 212.329
R21487 VDD.n3798 VDD.n3717 212.329
R21488 VDD.n3713 VDD.n3712 212.329
R21489 VDD.n3712 VDD.n3706 212.329
R21490 VDD.n3801 VDD.n3705 212.329
R21491 VDD.n3808 VDD.n3705 212.329
R21492 VDD.n3814 VDD.n3813 212.329
R21493 VDD.n3815 VDD.n3814 212.329
R21494 VDD.n3697 VDD.n3696 212.329
R21495 VDD.n3697 VDD.n3695 212.329
R21496 VDD.n3823 VDD.n3822 212.329
R21497 VDD.n3823 VDD.n3821 212.329
R21498 VDD.n3689 VDD.n3688 212.329
R21499 VDD.n3688 VDD.n3676 212.329
R21500 VDD.n3671 VDD.n3670 212.329
R21501 VDD.n3670 VDD.n2974 212.329
R21502 VDD.n3835 VDD.n2973 212.329
R21503 VDD.n3842 VDD.n2973 212.329
R21504 VDD.n2969 VDD.n2968 212.329
R21505 VDD.n2968 VDD.n2961 212.329
R21506 VDD.n3845 VDD.n2960 212.329
R21507 VDD.n3852 VDD.n2960 212.329
R21508 VDD.n2956 VDD.n2955 212.329
R21509 VDD.n2955 VDD.n2951 212.329
R21510 VDD.n3855 VDD.n2950 212.329
R21511 VDD.n3862 VDD.n2950 212.329
R21512 VDD.n2946 VDD.n2945 212.329
R21513 VDD.n2945 VDD.n2940 212.329
R21514 VDD.n3865 VDD.n2939 212.329
R21515 VDD.n3872 VDD.n2939 212.329
R21516 VDD.n3691 VDD.n3675 212.329
R21517 VDD.n3832 VDD.n3675 212.329
R21518 VDD.n3337 VDD.t534 176.65
R21519 VDD.n3342 VDD.t308 176.65
R21520 VDD.n3279 VDD.t619 176.65
R21521 VDD.n3432 VDD.t382 176.65
R21522 VDD.n3437 VDD.t868 176.65
R21523 VDD.n3242 VDD.t967 176.65
R21524 VDD.n3526 VDD.t557 176.65
R21525 VDD.n3529 VDD.t283 176.65
R21526 VDD.n1840 VDD.t940 169.018
R21527 VDD.n1593 VDD.t290 169.018
R21528 VDD.n1593 VDD.t389 169.018
R21529 VDD.n1627 VDD.t654 169.018
R21530 VDD.n1627 VDD.t581 169.018
R21531 VDD.n1689 VDD.t483 169.018
R21532 VDD.n1689 VDD.t294 169.018
R21533 VDD.n1664 VDD.t134 169.018
R21534 VDD.n1580 VDD.t853 169.018
R21535 VDD.n1333 VDD.t883 169.018
R21536 VDD.n1333 VDD.t433 169.018
R21537 VDD.n1367 VDD.t987 169.018
R21538 VDD.n1367 VDD.t882 169.018
R21539 VDD.n1429 VDD.t437 169.018
R21540 VDD.n1429 VDD.t535 169.018
R21541 VDD.n1404 VDD.t419 169.018
R21542 VDD.n1320 VDD.t977 169.018
R21543 VDD.n1073 VDD.t948 169.018
R21544 VDD.n1073 VDD.t72 169.018
R21545 VDD.n1107 VDD.t130 169.018
R21546 VDD.n1107 VDD.t945 169.018
R21547 VDD.n1169 VDD.t68 169.018
R21548 VDD.n1169 VDD.t196 169.018
R21549 VDD.n1144 VDD.t143 169.018
R21550 VDD.n1060 VDD.t942 169.018
R21551 VDD.n813 VDD.t573 169.018
R21552 VDD.n813 VDD.t393 169.018
R21553 VDD.n847 VDD.t435 169.018
R21554 VDD.n847 VDD.t826 169.018
R21555 VDD.n909 VDD.t983 169.018
R21556 VDD.n909 VDD.t575 169.018
R21557 VDD.n884 VDD.t179 169.018
R21558 VDD.n800 VDD.t849 169.018
R21559 VDD.n553 VDD.t709 169.018
R21560 VDD.n553 VDD.t649 169.018
R21561 VDD.n587 VDD.t485 169.018
R21562 VDD.n587 VDD.t708 169.018
R21563 VDD.n649 VDD.t653 169.018
R21564 VDD.n649 VDD.t710 169.018
R21565 VDD.n624 VDD.t517 169.018
R21566 VDD.n540 VDD.t979 169.018
R21567 VDD.n293 VDD.t934 169.018
R21568 VDD.n293 VDD.t984 169.018
R21569 VDD.n327 VDD.t395 169.018
R21570 VDD.n327 VDD.t932 169.018
R21571 VDD.n389 VDD.t467 169.018
R21572 VDD.n389 VDD.t936 169.018
R21573 VDD.n364 VDD.t415 169.018
R21574 VDD.n75 VDD.t860 169.018
R21575 VDD.n50 VDD.t327 169.018
R21576 VDD.n25 VDD.t638 169.018
R21577 VDD.n0 VDD.t835 169.018
R21578 VDD.n7456 VDD.t851 169.018
R21579 VDD.n7209 VDD.t1104 169.018
R21580 VDD.n7209 VDD.t651 169.018
R21581 VDD.n7243 VDD.t986 169.018
R21582 VDD.n7243 VDD.t1101 169.018
R21583 VDD.n7305 VDD.t431 169.018
R21584 VDD.n7305 VDD.t332 169.018
R21585 VDD.n7280 VDD.t272 169.018
R21586 VDD.n6909 VDD.t325 169.018
R21587 VDD.n6884 VDD.t577 169.018
R21588 VDD.n6859 VDD.t601 169.018
R21589 VDD.n6837 VDD.t590 169.018
R21590 VDD.n5052 VDD.t757 169.018
R21591 VDD.n5052 VDD.t24 169.018
R21592 VDD.n5114 VDD.t727 169.018
R21593 VDD.n5114 VDD.t100 169.018
R21594 VDD.n5149 VDD.t48 169.018
R21595 VDD.n5149 VDD.t805 169.018
R21596 VDD.n6704 VDD.t567 169.018
R21597 VDD.n5188 VDD.t809 169.018
R21598 VDD.n5188 VDD.t74 169.018
R21599 VDD.n5250 VDD.t733 169.018
R21600 VDD.n5250 VDD.t112 169.018
R21601 VDD.n5285 VDD.t56 169.018
R21602 VDD.n5285 VDD.t811 169.018
R21603 VDD.n6581 VDD.t156 169.018
R21604 VDD.n5324 VDD.t715 169.018
R21605 VDD.n5324 VDD.t84 169.018
R21606 VDD.n5386 VDD.t797 169.018
R21607 VDD.n5386 VDD.t66 169.018
R21608 VDD.n5421 VDD.t70 169.018
R21609 VDD.n5421 VDD.t725 169.018
R21610 VDD.n6458 VDD.t838 169.018
R21611 VDD.n5460 VDD.t787 169.018
R21612 VDD.n5460 VDD.t50 169.018
R21613 VDD.n5522 VDD.t815 169.018
R21614 VDD.n5522 VDD.t82 169.018
R21615 VDD.n5557 VDD.t34 169.018
R21616 VDD.n5557 VDD.t789 169.018
R21617 VDD.n6335 VDD.t830 169.018
R21618 VDD.n5596 VDD.t731 169.018
R21619 VDD.n5596 VDD.t104 169.018
R21620 VDD.n5658 VDD.t773 169.018
R21621 VDD.n5658 VDD.t44 169.018
R21622 VDD.n5693 VDD.t54 169.018
R21623 VDD.n5693 VDD.t807 169.018
R21624 VDD.n6212 VDD.t210 169.018
R21625 VDD.n5732 VDD.t759 169.018
R21626 VDD.n5732 VDD.t26 169.018
R21627 VDD.n5794 VDD.t793 169.018
R21628 VDD.n5794 VDD.t62 169.018
R21629 VDD.n5829 VDD.t108 169.018
R21630 VDD.n5829 VDD.t761 169.018
R21631 VDD.n6089 VDD.t947 169.018
R21632 VDD.n5868 VDD.t122 169.018
R21633 VDD.n5868 VDD.t779 169.018
R21634 VDD.n5930 VDD.t126 169.018
R21635 VDD.n5930 VDD.t781 169.018
R21636 VDD.n5965 VDD.t719 169.018
R21637 VDD.n5965 VDD.t86 169.018
R21638 VDD.n5966 VDD.t346 169.018
R21639 VDD.n5896 VDD.t1025 169.018
R21640 VDD.n5760 VDD.t1080 169.018
R21641 VDD.n5624 VDD.t1055 169.018
R21642 VDD.n5488 VDD.t1090 169.018
R21643 VDD.n5352 VDD.t1085 169.018
R21644 VDD.n5216 VDD.t1059 169.018
R21645 VDD.n5080 VDD.t1077 169.018
R21646 VDD.n4862 VDD.t729 169.018
R21647 VDD.n4862 VDD.t102 169.018
R21648 VDD.n4800 VDD.t813 169.018
R21649 VDD.n4800 VDD.t78 169.018
R21650 VDD.n4766 VDD.t88 169.018
R21651 VDD.n4766 VDD.t745 169.018
R21652 VDD.n5013 VDD.t204 169.018
R21653 VDD.n4837 VDD.t1053 169.018
R21654 VDD.n3732 VDD.t771 169.018
R21655 VDD.n3732 VDD.t36 169.018
R21656 VDD.n3707 VDD.t1095 169.018
R21657 VDD.n2906 VDD.t775 169.018
R21658 VDD.n2906 VDD.t38 169.018
R21659 VDD.n3880 VDD.t697 169.018
R21660 VDD.n2941 VDD.t120 169.018
R21661 VDD.n2941 VDD.t765 169.018
R21662 VDD.n2975 VDD.t717 169.018
R21663 VDD.n2975 VDD.t76 169.018
R21664 VDD.n2881 VDD.t1035 169.018
R21665 VDD.n2770 VDD.t751 169.018
R21666 VDD.n2770 VDD.t116 169.018
R21667 VDD.n4005 VDD.t1103 169.018
R21668 VDD.n2805 VDD.t94 169.018
R21669 VDD.n2805 VDD.t739 169.018
R21670 VDD.n2839 VDD.t763 169.018
R21671 VDD.n2839 VDD.t28 169.018
R21672 VDD.n2745 VDD.t1007 169.018
R21673 VDD.n2634 VDD.t799 169.018
R21674 VDD.n2634 VDD.t60 169.018
R21675 VDD.n4130 VDD.t877 169.018
R21676 VDD.n2669 VDD.t46 169.018
R21677 VDD.n2669 VDD.t791 169.018
R21678 VDD.n2703 VDD.t735 169.018
R21679 VDD.n2703 VDD.t106 169.018
R21680 VDD.n2609 VDD.t1063 169.018
R21681 VDD.n2498 VDD.t783 169.018
R21682 VDD.n2498 VDD.t42 169.018
R21683 VDD.n4255 VDD.t572 169.018
R21684 VDD.n2533 VDD.t128 169.018
R21685 VDD.n2533 VDD.t769 169.018
R21686 VDD.n2567 VDD.t721 169.018
R21687 VDD.n2567 VDD.t80 169.018
R21688 VDD.n2473 VDD.t1039 169.018
R21689 VDD.n2362 VDD.t755 169.018
R21690 VDD.n2362 VDD.t124 169.018
R21691 VDD.n4380 VDD.t904 169.018
R21692 VDD.n2397 VDD.t96 169.018
R21693 VDD.n2397 VDD.t743 169.018
R21694 VDD.n2431 VDD.t767 169.018
R21695 VDD.n2431 VDD.t32 169.018
R21696 VDD.n2337 VDD.t1011 169.018
R21697 VDD.n2226 VDD.t803 169.018
R21698 VDD.n2226 VDD.t64 169.018
R21699 VDD.n4505 VDD.t292 169.018
R21700 VDD.n2261 VDD.t98 169.018
R21701 VDD.n2261 VDD.t749 169.018
R21702 VDD.n2295 VDD.t741 169.018
R21703 VDD.n2295 VDD.t110 169.018
R21704 VDD.n2201 VDD.t1083 169.018
R21705 VDD.n2090 VDD.t795 169.018
R21706 VDD.n2090 VDD.t58 169.018
R21707 VDD.n4630 VDD.t921 169.018
R21708 VDD.n2125 VDD.t90 169.018
R21709 VDD.n2125 VDD.t737 169.018
R21710 VDD.n2159 VDD.t777 169.018
R21711 VDD.n2159 VDD.t40 169.018
R21712 VDD.n2065 VDD.t1069 169.018
R21713 VDD.n4755 VDD.t3 169.018
R21714 VDD.n1989 VDD.t52 169.018
R21715 VDD.n1989 VDD.t801 169.018
R21716 VDD.n2023 VDD.t753 169.018
R21717 VDD.n2023 VDD.t118 169.018
R21718 VDD.n1954 VDD.t747 169.018
R21719 VDD.n1954 VDD.t114 169.018
R21720 VDD.n1929 VDD.t1075 169.018
R21721 VDD.n7196 VDD.t914 169.018
R21722 VDD.n1853 VDD.t30 169.018
R21723 VDD.n1853 VDD.t785 169.018
R21724 VDD.n1887 VDD.t723 169.018
R21725 VDD.n1887 VDD.t92 169.018
R21726 VDD.n7459 VDD.t944 169.018
R21727 VDD.n7717 VDD.t521 169.018
R21728 VDD.n7717 VDD.t397 169.018
R21729 VDD.n7509 VDD.t471 169.018
R21730 VDD.n7509 VDD.t520 169.018
R21731 VDD.n7571 VDD.t195 169.018
R21732 VDD.n7571 VDD.t359 169.018
R21733 VDD.n7546 VDD.t149 169.018
R21734 VDD.n3376 VDD.t385 169.012
R21735 VDD.n3414 VDD.t991 169.012
R21736 VDD.n3255 VDD.t465 169.012
R21737 VDD.n3471 VDD.t406 169.012
R21738 VDD.n3508 VDD.t641 169.012
R21739 VDD.n3311 VDD.t212 169.012
R21740 VDD.n3205 VDD.t673 169.012
R21741 VDD.n3205 VDD.t161 169.012
R21742 VDD.n1615 VDD.t135 168.635
R21743 VDD.n1615 VDD.t917 168.635
R21744 VDD.n1614 VDD.t844 168.635
R21745 VDD.n1614 VDD.t132 168.635
R21746 VDD.n1649 VDD.t372 168.635
R21747 VDD.n1649 VDD.t594 168.635
R21748 VDD.n1648 VDD.t681 168.635
R21749 VDD.n1648 VDD.t400 168.635
R21750 VDD.n1677 VDD.t672 168.635
R21751 VDD.n1677 VDD.t401 168.635
R21752 VDD.n1676 VDD.t370 168.635
R21753 VDD.n1676 VDD.t671 168.635
R21754 VDD.n1711 VDD.t6 168.635
R21755 VDD.n1711 VDD.t963 168.635
R21756 VDD.n1710 VDD.t588 168.635
R21757 VDD.n1710 VDD.t425 168.635
R21758 VDD.n1355 VDD.t420 168.635
R21759 VDD.n1355 VDD.t265 168.635
R21760 VDD.n1354 VDD.t631 168.635
R21761 VDD.n1354 VDD.t417 168.635
R21762 VDD.n1389 VDD.t688 168.635
R21763 VDD.n1389 VDD.t691 168.635
R21764 VDD.n1388 VDD.t524 168.635
R21765 VDD.n1388 VDD.t864 168.635
R21766 VDD.n1417 VDD.t505 168.635
R21767 VDD.n1417 VDD.t361 168.635
R21768 VDD.n1416 VDD.t680 168.635
R21769 VDD.n1416 VDD.t506 168.635
R21770 VDD.n1451 VDD.t404 168.635
R21771 VDD.n1451 VDD.t888 168.635
R21772 VDD.n1450 VDD.t996 168.635
R21773 VDD.n1450 VDD.t901 168.635
R21774 VDD.n1095 VDD.t458 168.635
R21775 VDD.n1095 VDD.t227 168.635
R21776 VDD.n1094 VDD.t545 168.635
R21777 VDD.n1094 VDD.t141 168.635
R21778 VDD.n1129 VDD.t239 168.635
R21779 VDD.n1129 VDD.t191 168.635
R21780 VDD.n1128 VDD.t682 168.635
R21781 VDD.n1128 VDD.t284 168.635
R21782 VDD.n1157 VDD.t443 168.635
R21783 VDD.n1157 VDD.t231 168.635
R21784 VDD.n1156 VDD.t503 168.635
R21785 VDD.n1156 VDD.t444 168.635
R21786 VDD.n1191 VDD.t973 168.635
R21787 VDD.n1191 VDD.t14 168.635
R21788 VDD.n1190 VDD.t362 168.635
R21789 VDD.n1190 VDD.t189 168.635
R21790 VDD.n835 VDD.t613 168.635
R21791 VDD.n835 VDD.t586 168.635
R21792 VDD.n834 VDD.t845 168.635
R21793 VDD.n834 VDD.t614 168.635
R21794 VDD.n869 VDD.t962 168.635
R21795 VDD.n869 VDD.t558 168.635
R21796 VDD.n868 VDD.t169 168.635
R21797 VDD.n868 VDD.t139 168.635
R21798 VDD.n897 VDD.t677 168.635
R21799 VDD.n897 VDD.t137 168.635
R21800 VDD.n896 VDD.t961 168.635
R21801 VDD.n896 VDD.t676 168.635
R21802 VDD.n931 VDD.t989 168.635
R21803 VDD.n931 VDD.t328 168.635
R21804 VDD.n930 VDD.t314 168.635
R21805 VDD.n930 VDD.t886 168.635
R21806 VDD.n575 VDD.t518 168.635
R21807 VDD.n575 VDD.t317 168.635
R21808 VDD.n574 VDD.t980 168.635
R21809 VDD.n574 VDD.t515 168.635
R21810 VDD.n609 VDD.t288 168.635
R21811 VDD.n609 VDD.t636 168.635
R21812 VDD.n608 VDD.t982 168.635
R21813 VDD.n608 VDD.t177 168.635
R21814 VDD.n637 VDD.t267 168.635
R21815 VDD.n637 VDD.t217 168.635
R21816 VDD.n636 VDD.t287 168.635
R21817 VDD.n636 VDD.t268 168.635
R21818 VDD.n671 VDD.t896 168.635
R21819 VDD.n671 VDD.t350 168.635
R21820 VDD.n670 VDD.t253 168.635
R21821 VDD.n670 VDD.t241 168.635
R21822 VDD.n315 VDD.t412 168.635
R21823 VDD.n315 VDD.t336 168.635
R21824 VDD.n314 VDD.t546 168.635
R21825 VDD.n314 VDD.t413 168.635
R21826 VDD.n349 VDD.t383 168.635
R21827 VDD.n349 VDD.t597 168.635
R21828 VDD.n348 VDD.t606 168.635
R21829 VDD.n348 VDD.t175 168.635
R21830 VDD.n377 VDD.t629 168.635
R21831 VDD.n377 VDD.t479 168.635
R21832 VDD.n376 VDD.t674 168.635
R21833 VDD.n376 VDD.t630 168.635
R21834 VDD.n411 VDD.t215 168.635
R21835 VDD.n411 VDD.t964 168.635
R21836 VDD.n410 VDD.t193 168.635
R21837 VDD.n410 VDD.t218 168.635
R21838 VDD.n90 VDD.t198 168.635
R21839 VDD.n90 VDD.t380 168.635
R21840 VDD.n87 VDD.t251 168.635
R21841 VDD.n87 VDD.t1072 168.635
R21842 VDD.n65 VDD.t828 168.635
R21843 VDD.n65 VDD.t994 168.635
R21844 VDD.n62 VDD.t8 168.635
R21845 VDD.n62 VDD.t1027 168.635
R21846 VDD.n40 VDD.t154 168.635
R21847 VDD.n40 VDD.t569 168.635
R21848 VDD.n37 VDD.t822 168.635
R21849 VDD.n37 VDD.t1066 168.635
R21850 VDD.n15 VDD.t202 168.635
R21851 VDD.n15 VDD.t911 168.635
R21852 VDD.n12 VDD.t540 168.635
R21853 VDD.n12 VDD.t1093 168.635
R21854 VDD.n7231 VDD.t273 168.635
R21855 VDD.n7231 VDD.t605 168.635
R21856 VDD.n7230 VDD.t981 168.635
R21857 VDD.n7230 VDD.t270 168.635
R21858 VDD.n7265 VDD.t923 168.635
R21859 VDD.n7265 VDD.t310 168.635
R21860 VDD.n7264 VDD.t669 168.635
R21861 VDD.n7264 VDD.t874 168.635
R21862 VDD.n7293 VDD.t259 168.635
R21863 VDD.n7293 VDD.t376 168.635
R21864 VDD.n7292 VDD.t922 168.635
R21865 VDD.n7292 VDD.t260 168.635
R21866 VDD.n7327 VDD.t499 168.635
R21867 VDD.n7327 VDD.t489 168.635
R21868 VDD.n7326 VDD.t473 168.635
R21869 VDD.n7326 VDD.t928 168.635
R21870 VDD.n6924 VDD.t695 168.635
R21871 VDD.n6924 VDD.t330 168.635
R21872 VDD.n6921 VDD.t1037 168.635
R21873 VDD.n6921 VDD.t340 168.635
R21874 VDD.n6899 VDD.t879 168.635
R21875 VDD.n6899 VDD.t358 168.635
R21876 VDD.n6896 VDD.t1013 168.635
R21877 VDD.n6896 VDD.t621 168.635
R21878 VDD.n6874 VDD.t906 168.635
R21879 VDD.n6874 VDD.t583 168.635
R21880 VDD.n6871 VDD.t1041 168.635
R21881 VDD.n6871 VDD.t959 168.635
R21882 VDD.n6849 VDD.t871 168.635
R21883 VDD.n6849 VDD.t368 168.635
R21884 VDD.n6829 VDD.t1009 168.635
R21885 VDD.n6829 VDD.t410 168.635
R21886 VDD.n5015 VDD.t145 168.635
R21887 VDD.n5015 VDD.t938 168.635
R21888 VDD.n5014 VDD.t960 168.635
R21889 VDD.n5014 VDD.t865 168.635
R21890 VDD.n5064 VDD.t10 168.635
R21891 VDD.n5064 VDD.t508 168.635
R21892 VDD.n5063 VDD.t509 168.635
R21893 VDD.n5063 VDD.t668 168.635
R21894 VDD.n5092 VDD.t824 168.635
R21895 VDD.n5092 VDD.t667 168.635
R21896 VDD.n5091 VDD.t12 168.635
R21897 VDD.n5091 VDD.t562 168.635
R21898 VDD.n5126 VDD.t599 168.635
R21899 VDD.n5126 VDD.t1031 168.635
R21900 VDD.n5125 VDD.t1097 168.635
R21901 VDD.n5125 VDD.t861 168.635
R21902 VDD.n5151 VDD.t459 168.635
R21903 VDD.n5151 VDD.t863 168.635
R21904 VDD.n5150 VDD.t869 168.635
R21905 VDD.n5150 VDD.t286 168.635
R21906 VDD.n5200 VDD.t666 168.635
R21907 VDD.n5200 VDD.t342 168.635
R21908 VDD.n5199 VDD.t711 168.635
R21909 VDD.n5199 VDD.t832 168.635
R21910 VDD.n5228 VDD.t522 168.635
R21911 VDD.n5228 VDD.t644 168.635
R21912 VDD.n5227 VDD.t664 168.635
R21913 VDD.n5227 VDD.t487 168.635
R21914 VDD.n5262 VDD.t1107 168.635
R21915 VDD.n5262 VDD.t1078 168.635
R21916 VDD.n5261 VDD.t1033 168.635
R21917 VDD.n5261 VDD.t399 168.635
R21918 VDD.n5287 VDD.t448 168.635
R21919 VDD.n5287 VDD.t152 168.635
R21920 VDD.n5286 VDD.t488 168.635
R21921 VDD.n5286 VDD.t610 168.635
R21922 VDD.n5336 VDD.t16 168.635
R21923 VDD.n5336 VDD.t364 168.635
R21924 VDD.n5335 VDD.t833 168.635
R21925 VDD.n5335 VDD.t679 168.635
R21926 VDD.n5364 VDD.t935 168.635
R21927 VDD.n5364 VDD.t678 168.635
R21928 VDD.n5363 VDD.t22 168.635
R21929 VDD.n5363 VDD.t616 168.635
R21930 VDD.n5398 VDD.t858 168.635
R21931 VDD.n5398 VDD.t1096 168.635
R21932 VDD.n5397 VDD.t1061 168.635
R21933 VDD.n5397 VDD.t173 168.635
R21934 VDD.n5423 VDD.t200 168.635
R21935 VDD.n5423 VDD.t995 168.635
R21936 VDD.n5422 VDD.t659 168.635
R21937 VDD.n5422 VDD.t541 168.635
R21938 VDD.n5472 VDD.t171 168.635
R21939 VDD.n5472 VDD.t972 168.635
R21940 VDD.n5471 VDD.t429 168.635
R21941 VDD.n5471 VDD.t279 168.635
R21942 VDD.n5500 VDD.t366 168.635
R21943 VDD.n5500 VDD.t281 168.635
R21944 VDD.n5499 VDD.t841 168.635
R21945 VDD.n5499 VDD.t965 168.635
R21946 VDD.n5534 VDD.t255 168.635
R21947 VDD.n5534 VDD.t1047 168.635
R21948 VDD.n5533 VDD.t1003 168.635
R21949 VDD.n5533 VDD.t825 168.635
R21950 VDD.n5559 VDD.t278 168.635
R21951 VDD.n5559 VDD.t831 168.635
R21952 VDD.n5558 VDD.t312 168.635
R21953 VDD.n5558 VDD.t185 168.635
R21954 VDD.n5608 VDD.t302 168.635
R21955 VDD.n5608 VDD.t857 168.635
R21956 VDD.n5607 VDD.t856 168.635
R21957 VDD.n5607 VDD.t449 168.635
R21958 VDD.n5636 VDD.t924 168.635
R21959 VDD.n5636 VDD.t450 168.635
R21960 VDD.n5635 VDD.t304 168.635
R21961 VDD.n5635 VDD.t549 168.635
R21962 VDD.n5670 VDD.t624 168.635
R21963 VDD.n5670 VDD.t1070 168.635
R21964 VDD.n5669 VDD.t1029 168.635
R21965 VDD.n5669 VDD.t378 168.635
R21966 VDD.n5695 VDD.t352 168.635
R21967 VDD.n5695 VDD.t208 168.635
R21968 VDD.n5694 VDD.t997 168.635
R21969 VDD.n5694 VDD.t570 168.635
R21970 VDD.n5744 VDD.t500 168.635
R21971 VDD.n5744 VDD.t530 168.635
R21972 VDD.n5743 VDD.t531 168.635
R21973 VDD.n5743 VDD.t491 168.635
R21974 VDD.n5772 VDD.t300 168.635
R21975 VDD.n5772 VDD.t816 168.635
R21976 VDD.n5771 VDD.t502 168.635
R21977 VDD.n5771 VDD.t333 168.635
R21978 VDD.n5806 VDD.t611 168.635
R21979 VDD.n5806 VDD.t1088 168.635
R21980 VDD.n5805 VDD.t1057 168.635
R21981 VDD.n5805 VDD.t469 168.635
R21982 VDD.n5831 VDD.t889 168.635
R21983 VDD.n5831 VDD.t391 168.635
R21984 VDD.n5830 VDD.t918 168.635
R21985 VDD.n5830 VDD.t707 168.635
R21986 VDD.n5880 VDD.t951 168.635
R21987 VDD.n5880 VDD.t298 168.635
R21988 VDD.n5879 VDD.t387 168.635
R21989 VDD.n5879 VDD.t275 168.635
R21990 VDD.n5908 VDD.t899 168.635
R21991 VDD.n5908 VDD.t277 168.635
R21992 VDD.n5907 VDD.t952 168.635
R21993 VDD.n5907 VDD.t220 168.635
R21994 VDD.n5942 VDD.t563 168.635
R21995 VDD.n5942 VDD.t1044 168.635
R21996 VDD.n5941 VDD.t1001 168.635
R21997 VDD.n5941 VDD.t344 168.635
R21998 VDD.n4892 VDD.t349 168.635
R21999 VDD.n4892 VDD.t912 168.635
R22000 VDD.n4891 VDD.t493 168.635
R22001 VDD.n4891 VDD.t249 168.635
R22002 VDD.n4850 VDD.t421 168.635
R22003 VDD.n4850 VDD.t657 168.635
R22004 VDD.n4849 VDD.t656 168.635
R22005 VDD.n4849 VDD.t243 168.635
R22006 VDD.n4822 VDD.t820 168.635
R22007 VDD.n4822 VDD.t245 168.635
R22008 VDD.n4821 VDD.t422 168.635
R22009 VDD.n4821 VDD.t446 168.635
R22010 VDD.n4788 VDD.t408 168.635
R22011 VDD.n4788 VDD.t1005 168.635
R22012 VDD.n4787 VDD.t1081 168.635
R22013 VDD.n4787 VDD.t206 168.635
R22014 VDD.n3681 VDD.t163 168.635
R22015 VDD.n3681 VDD.t165 168.635
R22016 VDD.n3680 VDD.t584 168.635
R22017 VDD.n3680 VDD.t683 168.635
R22018 VDD.n3720 VDD.t551 168.635
R22019 VDD.n3720 VDD.t684 168.635
R22020 VDD.n3719 VDD.t247 168.635
R22021 VDD.n3719 VDD.t552 168.635
R22022 VDD.n3754 VDD.t348 168.635
R22023 VDD.n3754 VDD.t634 168.635
R22024 VDD.n3753 VDD.t909 168.635
R22025 VDD.n3753 VDD.t537 168.635
R22026 VDD.n2855 VDD.t542 168.635
R22027 VDD.n2855 VDD.t1106 168.635
R22028 VDD.n2854 VDD.t374 168.635
R22029 VDD.n2854 VDD.t511 168.635
R22030 VDD.n2894 VDD.t167 168.635
R22031 VDD.n2894 VDD.t930 168.635
R22032 VDD.n2893 VDD.t544 168.635
R22033 VDD.n2893 VDD.t334 168.635
R22034 VDD.n2928 VDD.t698 168.635
R22035 VDD.n2928 VDD.t840 168.635
R22036 VDD.n2927 VDD.t705 168.635
R22037 VDD.n2927 VDD.t690 168.635
R22038 VDD.n2963 VDD.t1064 168.635
R22039 VDD.n2963 VDD.t975 168.635
R22040 VDD.n2962 VDD.t693 168.635
R22041 VDD.n2962 VDD.t1015 168.635
R22042 VDD.n2719 VDD.t526 168.635
R22043 VDD.n2719 VDD.t926 168.635
R22044 VDD.n2718 VDD.t953 168.635
R22045 VDD.n2718 VDD.t559 168.635
R22046 VDD.n2758 VDD.t839 168.635
R22047 VDD.n2758 VDD.t560 168.635
R22048 VDD.n2757 VDD.t528 168.635
R22049 VDD.n2757 VDD.t296 168.635
R22050 VDD.n2792 VDD.t183 168.635
R22051 VDD.n2792 VDD.t842 168.635
R22052 VDD.n2791 VDD.t1 168.635
R22053 VDD.n2791 VDD.t627 168.635
R22054 VDD.n2827 VDD.t1046 168.635
R22055 VDD.n2827 VDD.t547 168.635
R22056 VDD.n2826 VDD.t181 168.635
R22057 VDD.n2826 VDD.t1099 168.635
R22058 VDD.n2583 VDD.t439 168.635
R22059 VDD.n2583 VDD.t477 168.635
R22060 VDD.n2582 VDD.t854 168.635
R22061 VDD.n2582 VDD.t622 168.635
R22062 VDD.n2622 VDD.t818 168.635
R22063 VDD.n2622 VDD.t623 168.635
R22064 VDD.n2621 VDD.t441 168.635
R22065 VDD.n2621 VDD.t819 168.635
R22066 VDD.n2656 VDD.t321 168.635
R22067 VDD.n2656 VDD.t475 168.635
R22068 VDD.n2655 VDD.t482 168.635
R22069 VDD.n2655 VDD.t457 168.635
R22070 VDD.n2691 VDD.t1019 168.635
R22071 VDD.n2691 VDD.t632 168.635
R22072 VDD.n2690 VDD.t319 168.635
R22073 VDD.n2690 VDD.t1087 168.635
R22074 VDD.n2447 VDD.t237 168.635
R22075 VDD.n2447 VDD.t427 168.635
R22076 VDD.n2446 VDD.t894 168.635
R22077 VDD.n2446 VDD.t497 168.635
R22078 VDD.n2486 VDD.t496 168.635
R22079 VDD.n2486 VDD.t645 168.635
R22080 VDD.n2485 VDD.t235 168.635
R22081 VDD.n2485 VDD.t263 168.635
R22082 VDD.n2520 VDD.t356 168.635
R22083 VDD.n2520 VDD.t323 168.635
R22084 VDD.n2519 VDD.t494 168.635
R22085 VDD.n2519 VDD.t519 168.635
R22086 VDD.n2555 VDD.t1073 168.635
R22087 VDD.n2555 VDD.t595 168.635
R22088 VDD.n2554 VDD.t354 168.635
R22089 VDD.n2554 VDD.t1023 168.635
R22090 VDD.n2311 VDD.t955 168.635
R22091 VDD.n2311 VDD.t452 168.635
R22092 VDD.n2310 VDD.t875 168.635
R22093 VDD.n2310 VDD.t968 168.635
R22094 VDD.n2350 VDD.t956 168.635
R22095 VDD.n2350 VDD.t998 168.635
R22096 VDD.n2349 VDD.t661 168.635
R22097 VDD.n2349 VDD.t338 168.635
R22098 VDD.n2384 VDD.t908 168.635
R22099 VDD.n2384 VDD.t823 168.635
R22100 VDD.n2383 VDD.t626 168.635
R22101 VDD.n2383 VDD.t454 168.635
R22102 VDD.n2419 VDD.t1049 168.635
R22103 VDD.n2419 VDD.t592 168.635
R22104 VDD.n2418 VDD.t907 168.635
R22105 VDD.n2418 VDD.t1100 168.635
R22106 VDD.n2175 VDD.t222 168.635
R22107 VDD.n2175 VDD.t513 168.635
R22108 VDD.n2174 VDD.t957 168.635
R22109 VDD.n2174 VDD.t1105 168.635
R22110 VDD.n2214 VDD.t836 168.635
R22111 VDD.n2214 VDD.t430 168.635
R22112 VDD.n2213 VDD.t224 168.635
R22113 VDD.n2213 VDD.t686 168.635
R22114 VDD.n2248 VDD.t579 168.635
R22115 VDD.n2248 VDD.t461 168.635
R22116 VDD.n2247 VDD.t538 168.635
R22117 VDD.n2247 VDD.t617 168.635
R22118 VDD.n2283 VDD.t1091 168.635
R22119 VDD.n2283 VDD.t565 168.635
R22120 VDD.n2282 VDD.t931 168.635
R22121 VDD.n2282 VDD.t1051 168.635
R22122 VDD.n2039 VDD.t388 168.635
R22123 VDD.n2039 VDD.t919 168.635
R22124 VDD.n2038 VDD.t257 168.635
R22125 VDD.n2038 VDD.t18 168.635
R22126 VDD.n2078 VDD.t608 168.635
R22127 VDD.n2078 VDD.t20 168.635
R22128 VDD.n2077 VDD.t639 168.635
R22129 VDD.n2077 VDD.t609 168.635
R22130 VDD.n2112 VDD.t872 168.635
R22131 VDD.n2112 VDD.t999 168.635
R22132 VDD.n2111 VDD.t233 168.635
R22133 VDD.n2111 VDD.t603 168.635
R22134 VDD.n2147 VDD.t1043 168.635
R22135 VDD.n2147 VDD.t187 168.635
R22136 VDD.n2146 VDD.t884 168.635
R22137 VDD.n2146 VDD.t1098 168.635
R22138 VDD.n2011 VDD.t1017 168.635
R22139 VDD.n2011 VDD.t647 168.635
R22140 VDD.n2010 VDD.t880 168.635
R22141 VDD.n2010 VDD.t1086 168.635
R22142 VDD.n1903 VDD.t424 168.635
R22143 VDD.n1903 VDD.t261 168.635
R22144 VDD.n1902 VDD.t229 168.635
R22145 VDD.n1902 VDD.t929 168.635
R22146 VDD.n1942 VDD.t971 168.635
R22147 VDD.n1942 VDD.t495 168.635
R22148 VDD.n1941 VDD.t306 168.635
R22149 VDD.n1941 VDD.t970 168.635
R22150 VDD.n1976 VDD.t536 168.635
R22151 VDD.n1976 VDD.t898 168.635
R22152 VDD.n1975 VDD.t927 168.635
R22153 VDD.n1975 VDD.t481 168.635
R22154 VDD.n1875 VDD.t1067 168.635
R22155 VDD.n1875 VDD.t456 168.635
R22156 VDD.n1874 VDD.t902 168.635
R22157 VDD.n1874 VDD.t1021 168.635
R22158 VDD.n7497 VDD.t150 168.635
R22159 VDD.n7497 VDD.t866 168.635
R22160 VDD.n7496 VDD.t847 168.635
R22161 VDD.n7496 VDD.t147 168.635
R22162 VDD.n7531 VDD.t950 168.635
R22163 VDD.n7531 VDD.t713 168.635
R22164 VDD.n7530 VDD.t900 168.635
R22165 VDD.n7530 VDD.t554 168.635
R22166 VDD.n7559 VDD.t892 168.635
R22167 VDD.n7559 VDD.t556 168.635
R22168 VDD.n7558 VDD.t949 168.635
R22169 VDD.n7558 VDD.t891 168.635
R22170 VDD.n7593 VDD.t158 168.635
R22171 VDD.n7593 VDD.t893 168.635
R22172 VDD.n7592 VDD.t663 168.635
R22173 VDD.n7592 VDD.t915 168.635
R22174 VDD.n7652 VDD.n7540 166.238
R22175 VDD.n7654 VDD.n7540 166.238
R22176 VDD.n7474 VDD.n7473 166.238
R22177 VDD.n7473 VDD.n7472 166.238
R22178 VDD.n1770 VDD.n1658 166.238
R22179 VDD.n1772 VDD.n1658 166.238
R22180 VDD.n1838 VDD.n1837 166.238
R22181 VDD.n1838 VDD.n1582 166.238
R22182 VDD.n1510 VDD.n1398 166.238
R22183 VDD.n1512 VDD.n1398 166.238
R22184 VDD.n1578 VDD.n1577 166.238
R22185 VDD.n1578 VDD.n1322 166.238
R22186 VDD.n1250 VDD.n1138 166.238
R22187 VDD.n1252 VDD.n1138 166.238
R22188 VDD.n1318 VDD.n1317 166.238
R22189 VDD.n1318 VDD.n1062 166.238
R22190 VDD.n990 VDD.n878 166.238
R22191 VDD.n992 VDD.n878 166.238
R22192 VDD.n1058 VDD.n1057 166.238
R22193 VDD.n1058 VDD.n802 166.238
R22194 VDD.n730 VDD.n618 166.238
R22195 VDD.n732 VDD.n618 166.238
R22196 VDD.n798 VDD.n797 166.238
R22197 VDD.n798 VDD.n542 166.238
R22198 VDD.n470 VDD.n358 166.238
R22199 VDD.n472 VDD.n358 166.238
R22200 VDD.n538 VDD.n537 166.238
R22201 VDD.n538 VDD.n282 166.238
R22202 VDD.n104 VDD.n101 166.238
R22203 VDD.n106 VDD.n101 166.238
R22204 VDD.n112 VDD.n111 166.238
R22205 VDD.n112 VDD.n92 166.238
R22206 VDD.n118 VDD.n115 166.238
R22207 VDD.n120 VDD.n115 166.238
R22208 VDD.n125 VDD.n84 166.238
R22209 VDD.n127 VDD.n84 166.238
R22210 VDD.n133 VDD.n132 166.238
R22211 VDD.n133 VDD.n76 166.238
R22212 VDD.n139 VDD.n136 166.238
R22213 VDD.n141 VDD.n136 166.238
R22214 VDD.n147 VDD.n146 166.238
R22215 VDD.n147 VDD.n67 166.238
R22216 VDD.n153 VDD.n150 166.238
R22217 VDD.n155 VDD.n150 166.238
R22218 VDD.n160 VDD.n59 166.238
R22219 VDD.n162 VDD.n59 166.238
R22220 VDD.n168 VDD.n167 166.238
R22221 VDD.n168 VDD.n51 166.238
R22222 VDD.n174 VDD.n171 166.238
R22223 VDD.n176 VDD.n171 166.238
R22224 VDD.n182 VDD.n181 166.238
R22225 VDD.n182 VDD.n42 166.238
R22226 VDD.n188 VDD.n185 166.238
R22227 VDD.n190 VDD.n185 166.238
R22228 VDD.n195 VDD.n34 166.238
R22229 VDD.n197 VDD.n34 166.238
R22230 VDD.n203 VDD.n202 166.238
R22231 VDD.n203 VDD.n26 166.238
R22232 VDD.n209 VDD.n206 166.238
R22233 VDD.n211 VDD.n206 166.238
R22234 VDD.n217 VDD.n216 166.238
R22235 VDD.n217 VDD.n17 166.238
R22236 VDD.n223 VDD.n220 166.238
R22237 VDD.n225 VDD.n220 166.238
R22238 VDD.n230 VDD.n9 166.238
R22239 VDD.n232 VDD.n9 166.238
R22240 VDD.n238 VDD.n237 166.238
R22241 VDD.n238 VDD.n1 166.238
R22242 VDD.n7386 VDD.n7274 166.238
R22243 VDD.n7388 VDD.n7274 166.238
R22244 VDD.n7454 VDD.n7453 166.238
R22245 VDD.n7454 VDD.n7198 166.238
R22246 VDD.n7194 VDD.n7193 166.238
R22247 VDD.n7194 VDD.n1842 166.238
R22248 VDD.n7129 VDD.n1923 166.238
R22249 VDD.n7131 VDD.n1923 166.238
R22250 VDD.n6938 VDD.n6935 166.238
R22251 VDD.n6940 VDD.n6935 166.238
R22252 VDD.n6946 VDD.n6945 166.238
R22253 VDD.n6946 VDD.n6926 166.238
R22254 VDD.n6952 VDD.n6949 166.238
R22255 VDD.n6954 VDD.n6949 166.238
R22256 VDD.n6959 VDD.n6918 166.238
R22257 VDD.n6961 VDD.n6918 166.238
R22258 VDD.n6967 VDD.n6966 166.238
R22259 VDD.n6967 VDD.n6910 166.238
R22260 VDD.n6973 VDD.n6970 166.238
R22261 VDD.n6975 VDD.n6970 166.238
R22262 VDD.n6981 VDD.n6980 166.238
R22263 VDD.n6981 VDD.n6901 166.238
R22264 VDD.n6987 VDD.n6984 166.238
R22265 VDD.n6989 VDD.n6984 166.238
R22266 VDD.n6994 VDD.n6893 166.238
R22267 VDD.n6996 VDD.n6893 166.238
R22268 VDD.n7002 VDD.n7001 166.238
R22269 VDD.n7002 VDD.n6885 166.238
R22270 VDD.n7008 VDD.n7005 166.238
R22271 VDD.n7010 VDD.n7005 166.238
R22272 VDD.n7016 VDD.n7015 166.238
R22273 VDD.n7016 VDD.n6876 166.238
R22274 VDD.n7022 VDD.n7019 166.238
R22275 VDD.n7024 VDD.n7019 166.238
R22276 VDD.n7029 VDD.n6868 166.238
R22277 VDD.n7031 VDD.n6868 166.238
R22278 VDD.n7037 VDD.n7036 166.238
R22279 VDD.n7037 VDD.n6860 166.238
R22280 VDD.n7043 VDD.n7040 166.238
R22281 VDD.n7045 VDD.n7040 166.238
R22282 VDD.n7051 VDD.n7050 166.238
R22283 VDD.n7051 VDD.n6851 166.238
R22284 VDD.n7057 VDD.n7054 166.238
R22285 VDD.n7059 VDD.n7054 166.238
R22286 VDD.n7066 VDD.n6832 166.238
R22287 VDD.n7066 VDD.n6831 166.238
R22288 VDD.n6843 VDD.n6838 166.238
R22289 VDD.n6841 VDD.n6838 166.238
R22290 VDD.n5968 VDD.n5964 166.238
R22291 VDD.n5969 VDD.n5968 166.238
R22292 VDD.n6034 VDD.n5889 166.238
R22293 VDD.n6036 VDD.n5889 166.238
R22294 VDD.n6091 VDD.n5828 166.238
R22295 VDD.n6092 VDD.n6091 166.238
R22296 VDD.n6157 VDD.n5753 166.238
R22297 VDD.n6159 VDD.n5753 166.238
R22298 VDD.n6214 VDD.n5692 166.238
R22299 VDD.n6215 VDD.n6214 166.238
R22300 VDD.n6280 VDD.n5617 166.238
R22301 VDD.n6282 VDD.n5617 166.238
R22302 VDD.n6337 VDD.n5556 166.238
R22303 VDD.n6338 VDD.n6337 166.238
R22304 VDD.n6403 VDD.n5481 166.238
R22305 VDD.n6405 VDD.n5481 166.238
R22306 VDD.n6460 VDD.n5420 166.238
R22307 VDD.n6461 VDD.n6460 166.238
R22308 VDD.n6526 VDD.n5345 166.238
R22309 VDD.n6528 VDD.n5345 166.238
R22310 VDD.n6583 VDD.n5284 166.238
R22311 VDD.n6584 VDD.n6583 166.238
R22312 VDD.n6649 VDD.n5209 166.238
R22313 VDD.n6651 VDD.n5209 166.238
R22314 VDD.n6706 VDD.n5148 166.238
R22315 VDD.n6707 VDD.n6706 166.238
R22316 VDD.n6772 VDD.n5073 166.238
R22317 VDD.n6774 VDD.n5073 166.238
R22318 VDD.n5011 VDD.n5010 166.238
R22319 VDD.n5011 VDD.n4756 166.238
R22320 VDD.n4943 VDD.n4830 166.238
R22321 VDD.n4941 VDD.n4830 166.238
R22322 VDD.n4753 VDD.n4752 166.238
R22323 VDD.n4753 VDD.n1978 166.238
R22324 VDD.n4688 VDD.n2059 166.238
R22325 VDD.n4690 VDD.n2059 166.238
R22326 VDD.n4628 VDD.n4627 166.238
R22327 VDD.n4628 VDD.n2114 166.238
R22328 VDD.n4563 VDD.n2195 166.238
R22329 VDD.n4565 VDD.n2195 166.238
R22330 VDD.n4503 VDD.n4502 166.238
R22331 VDD.n4503 VDD.n2250 166.238
R22332 VDD.n4438 VDD.n2331 166.238
R22333 VDD.n4440 VDD.n2331 166.238
R22334 VDD.n4378 VDD.n4377 166.238
R22335 VDD.n4378 VDD.n2386 166.238
R22336 VDD.n4313 VDD.n2467 166.238
R22337 VDD.n4315 VDD.n2467 166.238
R22338 VDD.n4253 VDD.n4252 166.238
R22339 VDD.n4253 VDD.n2522 166.238
R22340 VDD.n4188 VDD.n2603 166.238
R22341 VDD.n4190 VDD.n2603 166.238
R22342 VDD.n4128 VDD.n4127 166.238
R22343 VDD.n4128 VDD.n2658 166.238
R22344 VDD.n4063 VDD.n2739 166.238
R22345 VDD.n4065 VDD.n2739 166.238
R22346 VDD.n4003 VDD.n4002 166.238
R22347 VDD.n4003 VDD.n2794 166.238
R22348 VDD.n3938 VDD.n2875 166.238
R22349 VDD.n3940 VDD.n2875 166.238
R22350 VDD.n3388 VDD.n3387 166.238
R22351 VDD.n3388 VDD.n3283 166.238
R22352 VDD.n3380 VDD.n3379 166.238
R22353 VDD.n3379 VDD.n3290 166.238
R22354 VDD.n3374 VDD.n3373 166.238
R22355 VDD.n3374 VDD.n3363 166.238
R22356 VDD.n3425 VDD.n3424 166.238
R22357 VDD.n3425 VDD.n3392 166.238
R22358 VDD.n3417 VDD.n3416 166.238
R22359 VDD.n3416 VDD.n3399 166.238
R22360 VDD.n3412 VDD.n3411 166.238
R22361 VDD.n3412 VDD.n3401 166.238
R22362 VDD.n3277 VDD.n3276 166.238
R22363 VDD.n3277 VDD.n3266 166.238
R22364 VDD.n3445 VDD.n3265 166.238
R22365 VDD.n3446 VDD.n3445 166.238
R22366 VDD.n3452 VDD.n3451 166.238
R22367 VDD.n3452 VDD.n3256 166.238
R22368 VDD.n3483 VDD.n3482 166.238
R22369 VDD.n3483 VDD.n3246 166.238
R22370 VDD.n3475 VDD.n3474 166.238
R22371 VDD.n3474 VDD.n3253 166.238
R22372 VDD.n3469 VDD.n3468 166.238
R22373 VDD.n3469 VDD.n3458 166.238
R22374 VDD.n3519 VDD.n3518 166.238
R22375 VDD.n3519 VDD.n3486 166.238
R22376 VDD.n3511 VDD.n3510 166.238
R22377 VDD.n3510 VDD.n3493 166.238
R22378 VDD.n3506 VDD.n3505 166.238
R22379 VDD.n3506 VDD.n3495 166.238
R22380 VDD.n3333 VDD.n3332 166.238
R22381 VDD.n3333 VDD.n3322 166.238
R22382 VDD.n3350 VDD.n3321 166.238
R22383 VDD.n3351 VDD.n3350 166.238
R22384 VDD.n3357 VDD.n3356 166.238
R22385 VDD.n3357 VDD.n3312 166.238
R22386 VDD.n3878 VDD.n3877 166.238
R22387 VDD.n3878 VDD.n2930 166.238
R22388 VDD.n3813 VDD.n3701 166.238
R22389 VDD.n3815 VDD.n3701 166.238
R22390 VDD.n3085 VDD.t804 158.988
R22391 VDD.n3101 VDD.t800 158.988
R22392 VDD.n3149 VDD.t810 158.988
R22393 VDD.n3165 VDD.t736 158.988
R22394 VDD.n3046 VDD.t724 158.988
R22395 VDD.n3189 VDD.t748 158.988
R22396 VDD.n3300 VDD.t788 158.988
R22397 VDD.n3566 VDD.t742 158.988
R22398 VDD.n3007 VDD.t806 158.988
R22399 VDD.n3023 VDD.t768 158.988
R22400 VDD.n3594 VDD.t760 158.988
R22401 VDD.n3610 VDD.t790 158.988
R22402 VDD.n3633 VDD.t738 158.988
R22403 VDD.n3065 VDD.t744 158.988
R22404 VDD.n3120 VDD.t784 158.988
R22405 VDD.n3654 VDD.t764 158.988
R22406 VDD VDD.t718 158.581
R22407 VDD.n3113 VDD.t752 158.379
R22408 VDD.n3177 VDD.t776 158.379
R22409 VDD.n3201 VDD.t740 158.379
R22410 VDD.n3578 VDD.t766 158.379
R22411 VDD.n3035 VDD.t720 158.379
R22412 VDD.n3622 VDD.t734 158.379
R22413 VDD.n3645 VDD.t762 158.379
R22414 VDD.n3132 VDD.t722 158.379
R22415 VDD.n3666 VDD.t716 158.379
R22416 VDD.n109 VDD.n108 155.102
R22417 VDD.n123 VDD.n122 155.102
R22418 VDD.n144 VDD.n143 155.102
R22419 VDD.n158 VDD.n157 155.102
R22420 VDD.n179 VDD.n178 155.102
R22421 VDD.n193 VDD.n192 155.102
R22422 VDD.n214 VDD.n213 155.102
R22423 VDD.n228 VDD.n227 155.102
R22424 VDD.n6943 VDD.n6942 155.102
R22425 VDD.n6957 VDD.n6956 155.102
R22426 VDD.n6978 VDD.n6977 155.102
R22427 VDD.n6992 VDD.n6991 155.102
R22428 VDD.n7013 VDD.n7012 155.102
R22429 VDD.n7027 VDD.n7026 155.102
R22430 VDD.n7048 VDD.n7047 155.102
R22431 VDD.n7062 VDD.n7061 155.102
R22432 VDD.n3371 VDD.n3370 155.102
R22433 VDD.n3384 VDD.n3382 155.102
R22434 VDD.n3409 VDD.n3408 155.102
R22435 VDD.n3421 VDD.n3419 155.102
R22436 VDD.n3449 VDD.n3448 155.102
R22437 VDD.n3273 VDD.n3271 155.102
R22438 VDD.n3466 VDD.n3465 155.102
R22439 VDD.n3479 VDD.n3477 155.102
R22440 VDD.n3503 VDD.n3502 155.102
R22441 VDD.n3515 VDD.n3513 155.102
R22442 VDD.n3354 VDD.n3353 155.102
R22443 VDD.n3329 VDD.n3327 155.102
R22444 VDD.n7599 VDD.n7596 153.601
R22445 VDD.n7606 VDD.n7591 153.601
R22446 VDD.n7600 VDD.n7596 153.601
R22447 VDD.n7607 VDD.n7606 153.601
R22448 VDD.n7586 VDD.n7583 153.601
R22449 VDD.n7616 VDD.n7581 153.601
R22450 VDD.n7610 VDD.n7583 153.601
R22451 VDD.n7617 VDD.n7616 153.601
R22452 VDD.n7576 VDD.n7573 153.601
R22453 VDD.n7626 VDD.n7570 153.601
R22454 VDD.n7620 VDD.n7573 153.601
R22455 VDD.n7627 VDD.n7626 153.601
R22456 VDD.n7565 VDD.n7562 153.601
R22457 VDD.n7636 VDD.n7557 153.601
R22458 VDD.n7630 VDD.n7562 153.601
R22459 VDD.n7637 VDD.n7636 153.601
R22460 VDD.n7552 VDD.n7549 153.601
R22461 VDD.n7646 VDD.n7545 153.601
R22462 VDD.n7640 VDD.n7549 153.601
R22463 VDD.n7647 VDD.n7646 153.601
R22464 VDD.n7537 VDD.n7534 153.601
R22465 VDD.n7663 VDD.n7529 153.601
R22466 VDD.n7657 VDD.n7534 153.601
R22467 VDD.n7664 VDD.n7663 153.601
R22468 VDD.n7524 VDD.n7521 153.601
R22469 VDD.n7673 VDD.n7519 153.601
R22470 VDD.n7667 VDD.n7521 153.601
R22471 VDD.n7674 VDD.n7673 153.601
R22472 VDD.n7514 VDD.n7511 153.601
R22473 VDD.n7683 VDD.n7508 153.601
R22474 VDD.n7677 VDD.n7511 153.601
R22475 VDD.n7684 VDD.n7683 153.601
R22476 VDD.n7503 VDD.n7500 153.601
R22477 VDD.n7693 VDD.n7495 153.601
R22478 VDD.n7687 VDD.n7500 153.601
R22479 VDD.n7694 VDD.n7693 153.601
R22480 VDD.n7490 VDD.n7487 153.601
R22481 VDD.n7703 VDD.n7486 153.601
R22482 VDD.n7697 VDD.n7487 153.601
R22483 VDD.n7704 VDD.n7703 153.601
R22484 VDD.n7479 VDD.n7464 153.601
R22485 VDD.n7478 VDD.n7462 153.601
R22486 VDD.n7711 VDD.n7464 153.601
R22487 VDD.n7710 VDD.n7462 153.601
R22488 VDD.n1717 VDD.n1714 153.601
R22489 VDD.n1724 VDD.n1709 153.601
R22490 VDD.n1718 VDD.n1714 153.601
R22491 VDD.n1725 VDD.n1724 153.601
R22492 VDD.n1704 VDD.n1701 153.601
R22493 VDD.n1734 VDD.n1699 153.601
R22494 VDD.n1728 VDD.n1701 153.601
R22495 VDD.n1735 VDD.n1734 153.601
R22496 VDD.n1694 VDD.n1691 153.601
R22497 VDD.n1744 VDD.n1688 153.601
R22498 VDD.n1738 VDD.n1691 153.601
R22499 VDD.n1745 VDD.n1744 153.601
R22500 VDD.n1683 VDD.n1680 153.601
R22501 VDD.n1754 VDD.n1675 153.601
R22502 VDD.n1748 VDD.n1680 153.601
R22503 VDD.n1755 VDD.n1754 153.601
R22504 VDD.n1670 VDD.n1667 153.601
R22505 VDD.n1764 VDD.n1663 153.601
R22506 VDD.n1758 VDD.n1667 153.601
R22507 VDD.n1765 VDD.n1764 153.601
R22508 VDD.n1655 VDD.n1652 153.601
R22509 VDD.n1781 VDD.n1647 153.601
R22510 VDD.n1775 VDD.n1652 153.601
R22511 VDD.n1782 VDD.n1781 153.601
R22512 VDD.n1642 VDD.n1639 153.601
R22513 VDD.n1791 VDD.n1637 153.601
R22514 VDD.n1785 VDD.n1639 153.601
R22515 VDD.n1792 VDD.n1791 153.601
R22516 VDD.n1632 VDD.n1629 153.601
R22517 VDD.n1801 VDD.n1626 153.601
R22518 VDD.n1795 VDD.n1629 153.601
R22519 VDD.n1802 VDD.n1801 153.601
R22520 VDD.n1621 VDD.n1618 153.601
R22521 VDD.n1811 VDD.n1613 153.601
R22522 VDD.n1805 VDD.n1618 153.601
R22523 VDD.n1812 VDD.n1811 153.601
R22524 VDD.n1608 VDD.n1605 153.601
R22525 VDD.n1821 VDD.n1603 153.601
R22526 VDD.n1815 VDD.n1605 153.601
R22527 VDD.n1822 VDD.n1821 153.601
R22528 VDD.n1598 VDD.n1595 153.601
R22529 VDD.n1831 VDD.n1592 153.601
R22530 VDD.n1825 VDD.n1595 153.601
R22531 VDD.n1832 VDD.n1831 153.601
R22532 VDD.n1457 VDD.n1454 153.601
R22533 VDD.n1464 VDD.n1449 153.601
R22534 VDD.n1458 VDD.n1454 153.601
R22535 VDD.n1465 VDD.n1464 153.601
R22536 VDD.n1444 VDD.n1441 153.601
R22537 VDD.n1474 VDD.n1439 153.601
R22538 VDD.n1468 VDD.n1441 153.601
R22539 VDD.n1475 VDD.n1474 153.601
R22540 VDD.n1434 VDD.n1431 153.601
R22541 VDD.n1484 VDD.n1428 153.601
R22542 VDD.n1478 VDD.n1431 153.601
R22543 VDD.n1485 VDD.n1484 153.601
R22544 VDD.n1423 VDD.n1420 153.601
R22545 VDD.n1494 VDD.n1415 153.601
R22546 VDD.n1488 VDD.n1420 153.601
R22547 VDD.n1495 VDD.n1494 153.601
R22548 VDD.n1410 VDD.n1407 153.601
R22549 VDD.n1504 VDD.n1403 153.601
R22550 VDD.n1498 VDD.n1407 153.601
R22551 VDD.n1505 VDD.n1504 153.601
R22552 VDD.n1395 VDD.n1392 153.601
R22553 VDD.n1521 VDD.n1387 153.601
R22554 VDD.n1515 VDD.n1392 153.601
R22555 VDD.n1522 VDD.n1521 153.601
R22556 VDD.n1382 VDD.n1379 153.601
R22557 VDD.n1531 VDD.n1377 153.601
R22558 VDD.n1525 VDD.n1379 153.601
R22559 VDD.n1532 VDD.n1531 153.601
R22560 VDD.n1372 VDD.n1369 153.601
R22561 VDD.n1541 VDD.n1366 153.601
R22562 VDD.n1535 VDD.n1369 153.601
R22563 VDD.n1542 VDD.n1541 153.601
R22564 VDD.n1361 VDD.n1358 153.601
R22565 VDD.n1551 VDD.n1353 153.601
R22566 VDD.n1545 VDD.n1358 153.601
R22567 VDD.n1552 VDD.n1551 153.601
R22568 VDD.n1348 VDD.n1345 153.601
R22569 VDD.n1561 VDD.n1343 153.601
R22570 VDD.n1555 VDD.n1345 153.601
R22571 VDD.n1562 VDD.n1561 153.601
R22572 VDD.n1338 VDD.n1335 153.601
R22573 VDD.n1571 VDD.n1332 153.601
R22574 VDD.n1565 VDD.n1335 153.601
R22575 VDD.n1572 VDD.n1571 153.601
R22576 VDD.n1197 VDD.n1194 153.601
R22577 VDD.n1204 VDD.n1189 153.601
R22578 VDD.n1198 VDD.n1194 153.601
R22579 VDD.n1205 VDD.n1204 153.601
R22580 VDD.n1184 VDD.n1181 153.601
R22581 VDD.n1214 VDD.n1179 153.601
R22582 VDD.n1208 VDD.n1181 153.601
R22583 VDD.n1215 VDD.n1214 153.601
R22584 VDD.n1174 VDD.n1171 153.601
R22585 VDD.n1224 VDD.n1168 153.601
R22586 VDD.n1218 VDD.n1171 153.601
R22587 VDD.n1225 VDD.n1224 153.601
R22588 VDD.n1163 VDD.n1160 153.601
R22589 VDD.n1234 VDD.n1155 153.601
R22590 VDD.n1228 VDD.n1160 153.601
R22591 VDD.n1235 VDD.n1234 153.601
R22592 VDD.n1150 VDD.n1147 153.601
R22593 VDD.n1244 VDD.n1143 153.601
R22594 VDD.n1238 VDD.n1147 153.601
R22595 VDD.n1245 VDD.n1244 153.601
R22596 VDD.n1135 VDD.n1132 153.601
R22597 VDD.n1261 VDD.n1127 153.601
R22598 VDD.n1255 VDD.n1132 153.601
R22599 VDD.n1262 VDD.n1261 153.601
R22600 VDD.n1122 VDD.n1119 153.601
R22601 VDD.n1271 VDD.n1117 153.601
R22602 VDD.n1265 VDD.n1119 153.601
R22603 VDD.n1272 VDD.n1271 153.601
R22604 VDD.n1112 VDD.n1109 153.601
R22605 VDD.n1281 VDD.n1106 153.601
R22606 VDD.n1275 VDD.n1109 153.601
R22607 VDD.n1282 VDD.n1281 153.601
R22608 VDD.n1101 VDD.n1098 153.601
R22609 VDD.n1291 VDD.n1093 153.601
R22610 VDD.n1285 VDD.n1098 153.601
R22611 VDD.n1292 VDD.n1291 153.601
R22612 VDD.n1088 VDD.n1085 153.601
R22613 VDD.n1301 VDD.n1083 153.601
R22614 VDD.n1295 VDD.n1085 153.601
R22615 VDD.n1302 VDD.n1301 153.601
R22616 VDD.n1078 VDD.n1075 153.601
R22617 VDD.n1311 VDD.n1072 153.601
R22618 VDD.n1305 VDD.n1075 153.601
R22619 VDD.n1312 VDD.n1311 153.601
R22620 VDD.n937 VDD.n934 153.601
R22621 VDD.n944 VDD.n929 153.601
R22622 VDD.n938 VDD.n934 153.601
R22623 VDD.n945 VDD.n944 153.601
R22624 VDD.n924 VDD.n921 153.601
R22625 VDD.n954 VDD.n919 153.601
R22626 VDD.n948 VDD.n921 153.601
R22627 VDD.n955 VDD.n954 153.601
R22628 VDD.n914 VDD.n911 153.601
R22629 VDD.n964 VDD.n908 153.601
R22630 VDD.n958 VDD.n911 153.601
R22631 VDD.n965 VDD.n964 153.601
R22632 VDD.n903 VDD.n900 153.601
R22633 VDD.n974 VDD.n895 153.601
R22634 VDD.n968 VDD.n900 153.601
R22635 VDD.n975 VDD.n974 153.601
R22636 VDD.n890 VDD.n887 153.601
R22637 VDD.n984 VDD.n883 153.601
R22638 VDD.n978 VDD.n887 153.601
R22639 VDD.n985 VDD.n984 153.601
R22640 VDD.n875 VDD.n872 153.601
R22641 VDD.n1001 VDD.n867 153.601
R22642 VDD.n995 VDD.n872 153.601
R22643 VDD.n1002 VDD.n1001 153.601
R22644 VDD.n862 VDD.n859 153.601
R22645 VDD.n1011 VDD.n857 153.601
R22646 VDD.n1005 VDD.n859 153.601
R22647 VDD.n1012 VDD.n1011 153.601
R22648 VDD.n852 VDD.n849 153.601
R22649 VDD.n1021 VDD.n846 153.601
R22650 VDD.n1015 VDD.n849 153.601
R22651 VDD.n1022 VDD.n1021 153.601
R22652 VDD.n841 VDD.n838 153.601
R22653 VDD.n1031 VDD.n833 153.601
R22654 VDD.n1025 VDD.n838 153.601
R22655 VDD.n1032 VDD.n1031 153.601
R22656 VDD.n828 VDD.n825 153.601
R22657 VDD.n1041 VDD.n823 153.601
R22658 VDD.n1035 VDD.n825 153.601
R22659 VDD.n1042 VDD.n1041 153.601
R22660 VDD.n818 VDD.n815 153.601
R22661 VDD.n1051 VDD.n812 153.601
R22662 VDD.n1045 VDD.n815 153.601
R22663 VDD.n1052 VDD.n1051 153.601
R22664 VDD.n677 VDD.n674 153.601
R22665 VDD.n684 VDD.n669 153.601
R22666 VDD.n678 VDD.n674 153.601
R22667 VDD.n685 VDD.n684 153.601
R22668 VDD.n664 VDD.n661 153.601
R22669 VDD.n694 VDD.n659 153.601
R22670 VDD.n688 VDD.n661 153.601
R22671 VDD.n695 VDD.n694 153.601
R22672 VDD.n654 VDD.n651 153.601
R22673 VDD.n704 VDD.n648 153.601
R22674 VDD.n698 VDD.n651 153.601
R22675 VDD.n705 VDD.n704 153.601
R22676 VDD.n643 VDD.n640 153.601
R22677 VDD.n714 VDD.n635 153.601
R22678 VDD.n708 VDD.n640 153.601
R22679 VDD.n715 VDD.n714 153.601
R22680 VDD.n630 VDD.n627 153.601
R22681 VDD.n724 VDD.n623 153.601
R22682 VDD.n718 VDD.n627 153.601
R22683 VDD.n725 VDD.n724 153.601
R22684 VDD.n615 VDD.n612 153.601
R22685 VDD.n741 VDD.n607 153.601
R22686 VDD.n735 VDD.n612 153.601
R22687 VDD.n742 VDD.n741 153.601
R22688 VDD.n602 VDD.n599 153.601
R22689 VDD.n751 VDD.n597 153.601
R22690 VDD.n745 VDD.n599 153.601
R22691 VDD.n752 VDD.n751 153.601
R22692 VDD.n592 VDD.n589 153.601
R22693 VDD.n761 VDD.n586 153.601
R22694 VDD.n755 VDD.n589 153.601
R22695 VDD.n762 VDD.n761 153.601
R22696 VDD.n581 VDD.n578 153.601
R22697 VDD.n771 VDD.n573 153.601
R22698 VDD.n765 VDD.n578 153.601
R22699 VDD.n772 VDD.n771 153.601
R22700 VDD.n568 VDD.n565 153.601
R22701 VDD.n781 VDD.n563 153.601
R22702 VDD.n775 VDD.n565 153.601
R22703 VDD.n782 VDD.n781 153.601
R22704 VDD.n558 VDD.n555 153.601
R22705 VDD.n791 VDD.n552 153.601
R22706 VDD.n785 VDD.n555 153.601
R22707 VDD.n792 VDD.n791 153.601
R22708 VDD.n417 VDD.n414 153.601
R22709 VDD.n424 VDD.n409 153.601
R22710 VDD.n418 VDD.n414 153.601
R22711 VDD.n425 VDD.n424 153.601
R22712 VDD.n404 VDD.n401 153.601
R22713 VDD.n434 VDD.n399 153.601
R22714 VDD.n428 VDD.n401 153.601
R22715 VDD.n435 VDD.n434 153.601
R22716 VDD.n394 VDD.n391 153.601
R22717 VDD.n444 VDD.n388 153.601
R22718 VDD.n438 VDD.n391 153.601
R22719 VDD.n445 VDD.n444 153.601
R22720 VDD.n383 VDD.n380 153.601
R22721 VDD.n454 VDD.n375 153.601
R22722 VDD.n448 VDD.n380 153.601
R22723 VDD.n455 VDD.n454 153.601
R22724 VDD.n370 VDD.n367 153.601
R22725 VDD.n464 VDD.n363 153.601
R22726 VDD.n458 VDD.n367 153.601
R22727 VDD.n465 VDD.n464 153.601
R22728 VDD.n355 VDD.n352 153.601
R22729 VDD.n481 VDD.n347 153.601
R22730 VDD.n475 VDD.n352 153.601
R22731 VDD.n482 VDD.n481 153.601
R22732 VDD.n342 VDD.n339 153.601
R22733 VDD.n491 VDD.n337 153.601
R22734 VDD.n485 VDD.n339 153.601
R22735 VDD.n492 VDD.n491 153.601
R22736 VDD.n332 VDD.n329 153.601
R22737 VDD.n501 VDD.n326 153.601
R22738 VDD.n495 VDD.n329 153.601
R22739 VDD.n502 VDD.n501 153.601
R22740 VDD.n321 VDD.n318 153.601
R22741 VDD.n511 VDD.n313 153.601
R22742 VDD.n505 VDD.n318 153.601
R22743 VDD.n512 VDD.n511 153.601
R22744 VDD.n308 VDD.n305 153.601
R22745 VDD.n521 VDD.n303 153.601
R22746 VDD.n515 VDD.n305 153.601
R22747 VDD.n522 VDD.n521 153.601
R22748 VDD.n298 VDD.n295 153.601
R22749 VDD.n531 VDD.n292 153.601
R22750 VDD.n525 VDD.n295 153.601
R22751 VDD.n532 VDD.n531 153.601
R22752 VDD.n7333 VDD.n7330 153.601
R22753 VDD.n7340 VDD.n7325 153.601
R22754 VDD.n7334 VDD.n7330 153.601
R22755 VDD.n7341 VDD.n7340 153.601
R22756 VDD.n7320 VDD.n7317 153.601
R22757 VDD.n7350 VDD.n7315 153.601
R22758 VDD.n7344 VDD.n7317 153.601
R22759 VDD.n7351 VDD.n7350 153.601
R22760 VDD.n7310 VDD.n7307 153.601
R22761 VDD.n7360 VDD.n7304 153.601
R22762 VDD.n7354 VDD.n7307 153.601
R22763 VDD.n7361 VDD.n7360 153.601
R22764 VDD.n7299 VDD.n7296 153.601
R22765 VDD.n7370 VDD.n7291 153.601
R22766 VDD.n7364 VDD.n7296 153.601
R22767 VDD.n7371 VDD.n7370 153.601
R22768 VDD.n7286 VDD.n7283 153.601
R22769 VDD.n7380 VDD.n7279 153.601
R22770 VDD.n7374 VDD.n7283 153.601
R22771 VDD.n7381 VDD.n7380 153.601
R22772 VDD.n7271 VDD.n7268 153.601
R22773 VDD.n7397 VDD.n7263 153.601
R22774 VDD.n7391 VDD.n7268 153.601
R22775 VDD.n7398 VDD.n7397 153.601
R22776 VDD.n7258 VDD.n7255 153.601
R22777 VDD.n7407 VDD.n7253 153.601
R22778 VDD.n7401 VDD.n7255 153.601
R22779 VDD.n7408 VDD.n7407 153.601
R22780 VDD.n7248 VDD.n7245 153.601
R22781 VDD.n7417 VDD.n7242 153.601
R22782 VDD.n7411 VDD.n7245 153.601
R22783 VDD.n7418 VDD.n7417 153.601
R22784 VDD.n7237 VDD.n7234 153.601
R22785 VDD.n7427 VDD.n7229 153.601
R22786 VDD.n7421 VDD.n7234 153.601
R22787 VDD.n7428 VDD.n7427 153.601
R22788 VDD.n7224 VDD.n7221 153.601
R22789 VDD.n7437 VDD.n7219 153.601
R22790 VDD.n7431 VDD.n7221 153.601
R22791 VDD.n7438 VDD.n7437 153.601
R22792 VDD.n7214 VDD.n7211 153.601
R22793 VDD.n7447 VDD.n7208 153.601
R22794 VDD.n7441 VDD.n7211 153.601
R22795 VDD.n7448 VDD.n7447 153.601
R22796 VDD.n7076 VDD.n7073 153.601
R22797 VDD.n7083 VDD.n1974 153.601
R22798 VDD.n7077 VDD.n7073 153.601
R22799 VDD.n7084 VDD.n7083 153.601
R22800 VDD.n1969 VDD.n1966 153.601
R22801 VDD.n7093 VDD.n1964 153.601
R22802 VDD.n7087 VDD.n1966 153.601
R22803 VDD.n7094 VDD.n7093 153.601
R22804 VDD.n1959 VDD.n1956 153.601
R22805 VDD.n7103 VDD.n1953 153.601
R22806 VDD.n7097 VDD.n1956 153.601
R22807 VDD.n7104 VDD.n7103 153.601
R22808 VDD.n1948 VDD.n1945 153.601
R22809 VDD.n7113 VDD.n1940 153.601
R22810 VDD.n7107 VDD.n1945 153.601
R22811 VDD.n7114 VDD.n7113 153.601
R22812 VDD.n1935 VDD.n1932 153.601
R22813 VDD.n7123 VDD.n1928 153.601
R22814 VDD.n7117 VDD.n1932 153.601
R22815 VDD.n7124 VDD.n7123 153.601
R22816 VDD.n1918 VDD.n1906 153.601
R22817 VDD.n1917 VDD.n1904 153.601
R22818 VDD.n7138 VDD.n1906 153.601
R22819 VDD.n7137 VDD.n1904 153.601
R22820 VDD.n1911 VDD.n1899 153.601
R22821 VDD.n7147 VDD.n1898 153.601
R22822 VDD.n1893 VDD.n1890 153.601
R22823 VDD.n7157 VDD.n1886 153.601
R22824 VDD.n7151 VDD.n1890 153.601
R22825 VDD.n7158 VDD.n7157 153.601
R22826 VDD.n1881 VDD.n1878 153.601
R22827 VDD.n7167 VDD.n1873 153.601
R22828 VDD.n7161 VDD.n1878 153.601
R22829 VDD.n7168 VDD.n7167 153.601
R22830 VDD.n1868 VDD.n1865 153.601
R22831 VDD.n7177 VDD.n1863 153.601
R22832 VDD.n7171 VDD.n1865 153.601
R22833 VDD.n7178 VDD.n7177 153.601
R22834 VDD.n1858 VDD.n1855 153.601
R22835 VDD.n7187 VDD.n1852 153.601
R22836 VDD.n7181 VDD.n1855 153.601
R22837 VDD.n7188 VDD.n7187 153.601
R22838 VDD.n1913 VDD.n1899 153.601
R22839 VDD.n7148 VDD.n7147 153.601
R22840 VDD.n5958 VDD.n5955 153.601
R22841 VDD.n5978 VDD.n5953 153.601
R22842 VDD.n5972 VDD.n5955 153.601
R22843 VDD.n5979 VDD.n5978 153.601
R22844 VDD.n5948 VDD.n5945 153.601
R22845 VDD.n5988 VDD.n5940 153.601
R22846 VDD.n5982 VDD.n5945 153.601
R22847 VDD.n5989 VDD.n5988 153.601
R22848 VDD.n5935 VDD.n5932 153.601
R22849 VDD.n5998 VDD.n5929 153.601
R22850 VDD.n5992 VDD.n5932 153.601
R22851 VDD.n5999 VDD.n5998 153.601
R22852 VDD.n5924 VDD.n5921 153.601
R22853 VDD.n6008 VDD.n5919 153.601
R22854 VDD.n6002 VDD.n5921 153.601
R22855 VDD.n6009 VDD.n6008 153.601
R22856 VDD.n5914 VDD.n5911 153.601
R22857 VDD.n6018 VDD.n5906 153.601
R22858 VDD.n6012 VDD.n5911 153.601
R22859 VDD.n6019 VDD.n6018 153.601
R22860 VDD.n5901 VDD.n5898 153.601
R22861 VDD.n6028 VDD.n5894 153.601
R22862 VDD.n6022 VDD.n5898 153.601
R22863 VDD.n6029 VDD.n6028 153.601
R22864 VDD.n5886 VDD.n5883 153.601
R22865 VDD.n6045 VDD.n5878 153.601
R22866 VDD.n6039 VDD.n5883 153.601
R22867 VDD.n6046 VDD.n6045 153.601
R22868 VDD.n5873 VDD.n5870 153.601
R22869 VDD.n6055 VDD.n5867 153.601
R22870 VDD.n6049 VDD.n5870 153.601
R22871 VDD.n6056 VDD.n6055 153.601
R22872 VDD.n5862 VDD.n5859 153.601
R22873 VDD.n6065 VDD.n5857 153.601
R22874 VDD.n6059 VDD.n5859 153.601
R22875 VDD.n6066 VDD.n6065 153.601
R22876 VDD.n5852 VDD.n5849 153.601
R22877 VDD.n6075 VDD.n5847 153.601
R22878 VDD.n6069 VDD.n5849 153.601
R22879 VDD.n6076 VDD.n6075 153.601
R22880 VDD.n5840 VDD.n5835 153.601
R22881 VDD.n5839 VDD.n5833 153.601
R22882 VDD.n6083 VDD.n5835 153.601
R22883 VDD.n6082 VDD.n5833 153.601
R22884 VDD.n5822 VDD.n5819 153.601
R22885 VDD.n6101 VDD.n5817 153.601
R22886 VDD.n6095 VDD.n5819 153.601
R22887 VDD.n6102 VDD.n6101 153.601
R22888 VDD.n5812 VDD.n5809 153.601
R22889 VDD.n6111 VDD.n5804 153.601
R22890 VDD.n6105 VDD.n5809 153.601
R22891 VDD.n6112 VDD.n6111 153.601
R22892 VDD.n5799 VDD.n5796 153.601
R22893 VDD.n6121 VDD.n5793 153.601
R22894 VDD.n6115 VDD.n5796 153.601
R22895 VDD.n6122 VDD.n6121 153.601
R22896 VDD.n5788 VDD.n5785 153.601
R22897 VDD.n6131 VDD.n5783 153.601
R22898 VDD.n6125 VDD.n5785 153.601
R22899 VDD.n6132 VDD.n6131 153.601
R22900 VDD.n5778 VDD.n5775 153.601
R22901 VDD.n6141 VDD.n5770 153.601
R22902 VDD.n6135 VDD.n5775 153.601
R22903 VDD.n6142 VDD.n6141 153.601
R22904 VDD.n5765 VDD.n5762 153.601
R22905 VDD.n6151 VDD.n5758 153.601
R22906 VDD.n6145 VDD.n5762 153.601
R22907 VDD.n6152 VDD.n6151 153.601
R22908 VDD.n5750 VDD.n5747 153.601
R22909 VDD.n6168 VDD.n5742 153.601
R22910 VDD.n6162 VDD.n5747 153.601
R22911 VDD.n6169 VDD.n6168 153.601
R22912 VDD.n5737 VDD.n5734 153.601
R22913 VDD.n6178 VDD.n5731 153.601
R22914 VDD.n6172 VDD.n5734 153.601
R22915 VDD.n6179 VDD.n6178 153.601
R22916 VDD.n5726 VDD.n5723 153.601
R22917 VDD.n6188 VDD.n5721 153.601
R22918 VDD.n6182 VDD.n5723 153.601
R22919 VDD.n6189 VDD.n6188 153.601
R22920 VDD.n5716 VDD.n5713 153.601
R22921 VDD.n6198 VDD.n5711 153.601
R22922 VDD.n6192 VDD.n5713 153.601
R22923 VDD.n6199 VDD.n6198 153.601
R22924 VDD.n5704 VDD.n5699 153.601
R22925 VDD.n5703 VDD.n5697 153.601
R22926 VDD.n6206 VDD.n5699 153.601
R22927 VDD.n6205 VDD.n5697 153.601
R22928 VDD.n5686 VDD.n5683 153.601
R22929 VDD.n6224 VDD.n5681 153.601
R22930 VDD.n6218 VDD.n5683 153.601
R22931 VDD.n6225 VDD.n6224 153.601
R22932 VDD.n5676 VDD.n5673 153.601
R22933 VDD.n6234 VDD.n5668 153.601
R22934 VDD.n6228 VDD.n5673 153.601
R22935 VDD.n6235 VDD.n6234 153.601
R22936 VDD.n5663 VDD.n5660 153.601
R22937 VDD.n6244 VDD.n5657 153.601
R22938 VDD.n6238 VDD.n5660 153.601
R22939 VDD.n6245 VDD.n6244 153.601
R22940 VDD.n5652 VDD.n5649 153.601
R22941 VDD.n6254 VDD.n5647 153.601
R22942 VDD.n6248 VDD.n5649 153.601
R22943 VDD.n6255 VDD.n6254 153.601
R22944 VDD.n5642 VDD.n5639 153.601
R22945 VDD.n6264 VDD.n5634 153.601
R22946 VDD.n6258 VDD.n5639 153.601
R22947 VDD.n6265 VDD.n6264 153.601
R22948 VDD.n5629 VDD.n5626 153.601
R22949 VDD.n6274 VDD.n5622 153.601
R22950 VDD.n6268 VDD.n5626 153.601
R22951 VDD.n6275 VDD.n6274 153.601
R22952 VDD.n5614 VDD.n5611 153.601
R22953 VDD.n6291 VDD.n5606 153.601
R22954 VDD.n6285 VDD.n5611 153.601
R22955 VDD.n6292 VDD.n6291 153.601
R22956 VDD.n5601 VDD.n5598 153.601
R22957 VDD.n6301 VDD.n5595 153.601
R22958 VDD.n6295 VDD.n5598 153.601
R22959 VDD.n6302 VDD.n6301 153.601
R22960 VDD.n5590 VDD.n5587 153.601
R22961 VDD.n6311 VDD.n5585 153.601
R22962 VDD.n6305 VDD.n5587 153.601
R22963 VDD.n6312 VDD.n6311 153.601
R22964 VDD.n5580 VDD.n5577 153.601
R22965 VDD.n6321 VDD.n5575 153.601
R22966 VDD.n6315 VDD.n5577 153.601
R22967 VDD.n6322 VDD.n6321 153.601
R22968 VDD.n5568 VDD.n5563 153.601
R22969 VDD.n5567 VDD.n5561 153.601
R22970 VDD.n6329 VDD.n5563 153.601
R22971 VDD.n6328 VDD.n5561 153.601
R22972 VDD.n5550 VDD.n5547 153.601
R22973 VDD.n6347 VDD.n5545 153.601
R22974 VDD.n6341 VDD.n5547 153.601
R22975 VDD.n6348 VDD.n6347 153.601
R22976 VDD.n5540 VDD.n5537 153.601
R22977 VDD.n6357 VDD.n5532 153.601
R22978 VDD.n6351 VDD.n5537 153.601
R22979 VDD.n6358 VDD.n6357 153.601
R22980 VDD.n5527 VDD.n5524 153.601
R22981 VDD.n6367 VDD.n5521 153.601
R22982 VDD.n6361 VDD.n5524 153.601
R22983 VDD.n6368 VDD.n6367 153.601
R22984 VDD.n5516 VDD.n5513 153.601
R22985 VDD.n6377 VDD.n5511 153.601
R22986 VDD.n6371 VDD.n5513 153.601
R22987 VDD.n6378 VDD.n6377 153.601
R22988 VDD.n5506 VDD.n5503 153.601
R22989 VDD.n6387 VDD.n5498 153.601
R22990 VDD.n6381 VDD.n5503 153.601
R22991 VDD.n6388 VDD.n6387 153.601
R22992 VDD.n5493 VDD.n5490 153.601
R22993 VDD.n6397 VDD.n5486 153.601
R22994 VDD.n6391 VDD.n5490 153.601
R22995 VDD.n6398 VDD.n6397 153.601
R22996 VDD.n5478 VDD.n5475 153.601
R22997 VDD.n6414 VDD.n5470 153.601
R22998 VDD.n6408 VDD.n5475 153.601
R22999 VDD.n6415 VDD.n6414 153.601
R23000 VDD.n5465 VDD.n5462 153.601
R23001 VDD.n6424 VDD.n5459 153.601
R23002 VDD.n6418 VDD.n5462 153.601
R23003 VDD.n6425 VDD.n6424 153.601
R23004 VDD.n5454 VDD.n5451 153.601
R23005 VDD.n6434 VDD.n5449 153.601
R23006 VDD.n6428 VDD.n5451 153.601
R23007 VDD.n6435 VDD.n6434 153.601
R23008 VDD.n5444 VDD.n5441 153.601
R23009 VDD.n6444 VDD.n5439 153.601
R23010 VDD.n6438 VDD.n5441 153.601
R23011 VDD.n6445 VDD.n6444 153.601
R23012 VDD.n5432 VDD.n5427 153.601
R23013 VDD.n5431 VDD.n5425 153.601
R23014 VDD.n6452 VDD.n5427 153.601
R23015 VDD.n6451 VDD.n5425 153.601
R23016 VDD.n5414 VDD.n5411 153.601
R23017 VDD.n6470 VDD.n5409 153.601
R23018 VDD.n6464 VDD.n5411 153.601
R23019 VDD.n6471 VDD.n6470 153.601
R23020 VDD.n5404 VDD.n5401 153.601
R23021 VDD.n6480 VDD.n5396 153.601
R23022 VDD.n6474 VDD.n5401 153.601
R23023 VDD.n6481 VDD.n6480 153.601
R23024 VDD.n5391 VDD.n5388 153.601
R23025 VDD.n6490 VDD.n5385 153.601
R23026 VDD.n6484 VDD.n5388 153.601
R23027 VDD.n6491 VDD.n6490 153.601
R23028 VDD.n5380 VDD.n5377 153.601
R23029 VDD.n6500 VDD.n5375 153.601
R23030 VDD.n6494 VDD.n5377 153.601
R23031 VDD.n6501 VDD.n6500 153.601
R23032 VDD.n5370 VDD.n5367 153.601
R23033 VDD.n6510 VDD.n5362 153.601
R23034 VDD.n6504 VDD.n5367 153.601
R23035 VDD.n6511 VDD.n6510 153.601
R23036 VDD.n5357 VDD.n5354 153.601
R23037 VDD.n6520 VDD.n5350 153.601
R23038 VDD.n6514 VDD.n5354 153.601
R23039 VDD.n6521 VDD.n6520 153.601
R23040 VDD.n5342 VDD.n5339 153.601
R23041 VDD.n6537 VDD.n5334 153.601
R23042 VDD.n6531 VDD.n5339 153.601
R23043 VDD.n6538 VDD.n6537 153.601
R23044 VDD.n5329 VDD.n5326 153.601
R23045 VDD.n6547 VDD.n5323 153.601
R23046 VDD.n6541 VDD.n5326 153.601
R23047 VDD.n6548 VDD.n6547 153.601
R23048 VDD.n5318 VDD.n5315 153.601
R23049 VDD.n6557 VDD.n5313 153.601
R23050 VDD.n6551 VDD.n5315 153.601
R23051 VDD.n6558 VDD.n6557 153.601
R23052 VDD.n5308 VDD.n5305 153.601
R23053 VDD.n6567 VDD.n5303 153.601
R23054 VDD.n6561 VDD.n5305 153.601
R23055 VDD.n6568 VDD.n6567 153.601
R23056 VDD.n5296 VDD.n5291 153.601
R23057 VDD.n5295 VDD.n5289 153.601
R23058 VDD.n6575 VDD.n5291 153.601
R23059 VDD.n6574 VDD.n5289 153.601
R23060 VDD.n5278 VDD.n5275 153.601
R23061 VDD.n6593 VDD.n5273 153.601
R23062 VDD.n6587 VDD.n5275 153.601
R23063 VDD.n6594 VDD.n6593 153.601
R23064 VDD.n5268 VDD.n5265 153.601
R23065 VDD.n6603 VDD.n5260 153.601
R23066 VDD.n6597 VDD.n5265 153.601
R23067 VDD.n6604 VDD.n6603 153.601
R23068 VDD.n5255 VDD.n5252 153.601
R23069 VDD.n6613 VDD.n5249 153.601
R23070 VDD.n6607 VDD.n5252 153.601
R23071 VDD.n6614 VDD.n6613 153.601
R23072 VDD.n5244 VDD.n5241 153.601
R23073 VDD.n6623 VDD.n5239 153.601
R23074 VDD.n6617 VDD.n5241 153.601
R23075 VDD.n6624 VDD.n6623 153.601
R23076 VDD.n5234 VDD.n5231 153.601
R23077 VDD.n6633 VDD.n5226 153.601
R23078 VDD.n6627 VDD.n5231 153.601
R23079 VDD.n6634 VDD.n6633 153.601
R23080 VDD.n5221 VDD.n5218 153.601
R23081 VDD.n6643 VDD.n5214 153.601
R23082 VDD.n6637 VDD.n5218 153.601
R23083 VDD.n6644 VDD.n6643 153.601
R23084 VDD.n5206 VDD.n5203 153.601
R23085 VDD.n6660 VDD.n5198 153.601
R23086 VDD.n6654 VDD.n5203 153.601
R23087 VDD.n6661 VDD.n6660 153.601
R23088 VDD.n5193 VDD.n5190 153.601
R23089 VDD.n6670 VDD.n5187 153.601
R23090 VDD.n6664 VDD.n5190 153.601
R23091 VDD.n6671 VDD.n6670 153.601
R23092 VDD.n5182 VDD.n5179 153.601
R23093 VDD.n6680 VDD.n5177 153.601
R23094 VDD.n6674 VDD.n5179 153.601
R23095 VDD.n6681 VDD.n6680 153.601
R23096 VDD.n5172 VDD.n5169 153.601
R23097 VDD.n6690 VDD.n5167 153.601
R23098 VDD.n6684 VDD.n5169 153.601
R23099 VDD.n6691 VDD.n6690 153.601
R23100 VDD.n5160 VDD.n5155 153.601
R23101 VDD.n5159 VDD.n5153 153.601
R23102 VDD.n6698 VDD.n5155 153.601
R23103 VDD.n6697 VDD.n5153 153.601
R23104 VDD.n5142 VDD.n5139 153.601
R23105 VDD.n6716 VDD.n5137 153.601
R23106 VDD.n6710 VDD.n5139 153.601
R23107 VDD.n6717 VDD.n6716 153.601
R23108 VDD.n5132 VDD.n5129 153.601
R23109 VDD.n6726 VDD.n5124 153.601
R23110 VDD.n6720 VDD.n5129 153.601
R23111 VDD.n6727 VDD.n6726 153.601
R23112 VDD.n5119 VDD.n5116 153.601
R23113 VDD.n6736 VDD.n5113 153.601
R23114 VDD.n6730 VDD.n5116 153.601
R23115 VDD.n6737 VDD.n6736 153.601
R23116 VDD.n5108 VDD.n5105 153.601
R23117 VDD.n6746 VDD.n5103 153.601
R23118 VDD.n6740 VDD.n5105 153.601
R23119 VDD.n6747 VDD.n6746 153.601
R23120 VDD.n5098 VDD.n5095 153.601
R23121 VDD.n6756 VDD.n5090 153.601
R23122 VDD.n6750 VDD.n5095 153.601
R23123 VDD.n6757 VDD.n6756 153.601
R23124 VDD.n5085 VDD.n5082 153.601
R23125 VDD.n6766 VDD.n5078 153.601
R23126 VDD.n6760 VDD.n5082 153.601
R23127 VDD.n6767 VDD.n6766 153.601
R23128 VDD.n5070 VDD.n5067 153.601
R23129 VDD.n6783 VDD.n5062 153.601
R23130 VDD.n6777 VDD.n5067 153.601
R23131 VDD.n6784 VDD.n6783 153.601
R23132 VDD.n5057 VDD.n5054 153.601
R23133 VDD.n6793 VDD.n5051 153.601
R23134 VDD.n6787 VDD.n5054 153.601
R23135 VDD.n6794 VDD.n6793 153.601
R23136 VDD.n5046 VDD.n5043 153.601
R23137 VDD.n6803 VDD.n5041 153.601
R23138 VDD.n6797 VDD.n5043 153.601
R23139 VDD.n6804 VDD.n6803 153.601
R23140 VDD.n5036 VDD.n5033 153.601
R23141 VDD.n6813 VDD.n5031 153.601
R23142 VDD.n6807 VDD.n5033 153.601
R23143 VDD.n6814 VDD.n6813 153.601
R23144 VDD.n5024 VDD.n5019 153.601
R23145 VDD.n5023 VDD.n5017 153.601
R23146 VDD.n6821 VDD.n5019 153.601
R23147 VDD.n6820 VDD.n5017 153.601
R23148 VDD.n5002 VDD.n4764 153.601
R23149 VDD.n4770 VDD.n4765 153.601
R23150 VDD.n5003 VDD.n5002 153.601
R23151 VDD.n4996 VDD.n4765 153.601
R23152 VDD.n4992 VDD.n4775 153.601
R23153 VDD.n4780 VDD.n4776 153.601
R23154 VDD.n4993 VDD.n4992 153.601
R23155 VDD.n4986 VDD.n4776 153.601
R23156 VDD.n4982 VDD.n4785 153.601
R23157 VDD.n4793 VDD.n4786 153.601
R23158 VDD.n4983 VDD.n4982 153.601
R23159 VDD.n4976 VDD.n4786 153.601
R23160 VDD.n4972 VDD.n4798 153.601
R23161 VDD.n4804 VDD.n4799 153.601
R23162 VDD.n4973 VDD.n4972 153.601
R23163 VDD.n4966 VDD.n4799 153.601
R23164 VDD.n4962 VDD.n4809 153.601
R23165 VDD.n4814 VDD.n4810 153.601
R23166 VDD.n4963 VDD.n4962 153.601
R23167 VDD.n4956 VDD.n4810 153.601
R23168 VDD.n4952 VDD.n4819 153.601
R23169 VDD.n4827 VDD.n4820 153.601
R23170 VDD.n4953 VDD.n4952 153.601
R23171 VDD.n4946 VDD.n4820 153.601
R23172 VDD.n4935 VDD.n4835 153.601
R23173 VDD.n4842 VDD.n4836 153.601
R23174 VDD.n4936 VDD.n4935 153.601
R23175 VDD.n4929 VDD.n4836 153.601
R23176 VDD.n4925 VDD.n4847 153.601
R23177 VDD.n4855 VDD.n4848 153.601
R23178 VDD.n4926 VDD.n4925 153.601
R23179 VDD.n4919 VDD.n4848 153.601
R23180 VDD.n4915 VDD.n4860 153.601
R23181 VDD.n4866 VDD.n4861 153.601
R23182 VDD.n4916 VDD.n4915 153.601
R23183 VDD.n4909 VDD.n4861 153.601
R23184 VDD.n4905 VDD.n4871 153.601
R23185 VDD.n4876 VDD.n4872 153.601
R23186 VDD.n4906 VDD.n4905 153.601
R23187 VDD.n4899 VDD.n4872 153.601
R23188 VDD.n4895 VDD.n4881 153.601
R23189 VDD.n4885 VDD.n4882 153.601
R23190 VDD.n4896 VDD.n4895 153.601
R23191 VDD.n4886 VDD.n4882 153.601
R23192 VDD.n4635 VDD.n4632 153.601
R23193 VDD.n4642 VDD.n2110 153.601
R23194 VDD.n4636 VDD.n4632 153.601
R23195 VDD.n4643 VDD.n4642 153.601
R23196 VDD.n2105 VDD.n2102 153.601
R23197 VDD.n4652 VDD.n2100 153.601
R23198 VDD.n4646 VDD.n2102 153.601
R23199 VDD.n4653 VDD.n4652 153.601
R23200 VDD.n2095 VDD.n2092 153.601
R23201 VDD.n4662 VDD.n2089 153.601
R23202 VDD.n4656 VDD.n2092 153.601
R23203 VDD.n4663 VDD.n4662 153.601
R23204 VDD.n2084 VDD.n2081 153.601
R23205 VDD.n4672 VDD.n2076 153.601
R23206 VDD.n4666 VDD.n2081 153.601
R23207 VDD.n4673 VDD.n4672 153.601
R23208 VDD.n2071 VDD.n2068 153.601
R23209 VDD.n4682 VDD.n2064 153.601
R23210 VDD.n4676 VDD.n2068 153.601
R23211 VDD.n4683 VDD.n4682 153.601
R23212 VDD.n2054 VDD.n2042 153.601
R23213 VDD.n2053 VDD.n2040 153.601
R23214 VDD.n4697 VDD.n2042 153.601
R23215 VDD.n4696 VDD.n2040 153.601
R23216 VDD.n2047 VDD.n2035 153.601
R23217 VDD.n4706 VDD.n2034 153.601
R23218 VDD.n2029 VDD.n2026 153.601
R23219 VDD.n4716 VDD.n2022 153.601
R23220 VDD.n4710 VDD.n2026 153.601
R23221 VDD.n4717 VDD.n4716 153.601
R23222 VDD.n2017 VDD.n2014 153.601
R23223 VDD.n4726 VDD.n2009 153.601
R23224 VDD.n4720 VDD.n2014 153.601
R23225 VDD.n4727 VDD.n4726 153.601
R23226 VDD.n2004 VDD.n2001 153.601
R23227 VDD.n4736 VDD.n1999 153.601
R23228 VDD.n4730 VDD.n2001 153.601
R23229 VDD.n4737 VDD.n4736 153.601
R23230 VDD.n1994 VDD.n1991 153.601
R23231 VDD.n4746 VDD.n1988 153.601
R23232 VDD.n4740 VDD.n1991 153.601
R23233 VDD.n4747 VDD.n4746 153.601
R23234 VDD.n2049 VDD.n2035 153.601
R23235 VDD.n4707 VDD.n4706 153.601
R23236 VDD.n4510 VDD.n4507 153.601
R23237 VDD.n4517 VDD.n2246 153.601
R23238 VDD.n4511 VDD.n4507 153.601
R23239 VDD.n4518 VDD.n4517 153.601
R23240 VDD.n2241 VDD.n2238 153.601
R23241 VDD.n4527 VDD.n2236 153.601
R23242 VDD.n4521 VDD.n2238 153.601
R23243 VDD.n4528 VDD.n4527 153.601
R23244 VDD.n2231 VDD.n2228 153.601
R23245 VDD.n4537 VDD.n2225 153.601
R23246 VDD.n4531 VDD.n2228 153.601
R23247 VDD.n4538 VDD.n4537 153.601
R23248 VDD.n2220 VDD.n2217 153.601
R23249 VDD.n4547 VDD.n2212 153.601
R23250 VDD.n4541 VDD.n2217 153.601
R23251 VDD.n4548 VDD.n4547 153.601
R23252 VDD.n2207 VDD.n2204 153.601
R23253 VDD.n4557 VDD.n2200 153.601
R23254 VDD.n4551 VDD.n2204 153.601
R23255 VDD.n4558 VDD.n4557 153.601
R23256 VDD.n2190 VDD.n2178 153.601
R23257 VDD.n2189 VDD.n2176 153.601
R23258 VDD.n4572 VDD.n2178 153.601
R23259 VDD.n4571 VDD.n2176 153.601
R23260 VDD.n2183 VDD.n2171 153.601
R23261 VDD.n4581 VDD.n2170 153.601
R23262 VDD.n2165 VDD.n2162 153.601
R23263 VDD.n4591 VDD.n2158 153.601
R23264 VDD.n4585 VDD.n2162 153.601
R23265 VDD.n4592 VDD.n4591 153.601
R23266 VDD.n2153 VDD.n2150 153.601
R23267 VDD.n4601 VDD.n2145 153.601
R23268 VDD.n4595 VDD.n2150 153.601
R23269 VDD.n4602 VDD.n4601 153.601
R23270 VDD.n2140 VDD.n2137 153.601
R23271 VDD.n4611 VDD.n2135 153.601
R23272 VDD.n4605 VDD.n2137 153.601
R23273 VDD.n4612 VDD.n4611 153.601
R23274 VDD.n2130 VDD.n2127 153.601
R23275 VDD.n4621 VDD.n2124 153.601
R23276 VDD.n4615 VDD.n2127 153.601
R23277 VDD.n4622 VDD.n4621 153.601
R23278 VDD.n2185 VDD.n2171 153.601
R23279 VDD.n4582 VDD.n4581 153.601
R23280 VDD.n4385 VDD.n4382 153.601
R23281 VDD.n4392 VDD.n2382 153.601
R23282 VDD.n4386 VDD.n4382 153.601
R23283 VDD.n4393 VDD.n4392 153.601
R23284 VDD.n2377 VDD.n2374 153.601
R23285 VDD.n4402 VDD.n2372 153.601
R23286 VDD.n4396 VDD.n2374 153.601
R23287 VDD.n4403 VDD.n4402 153.601
R23288 VDD.n2367 VDD.n2364 153.601
R23289 VDD.n4412 VDD.n2361 153.601
R23290 VDD.n4406 VDD.n2364 153.601
R23291 VDD.n4413 VDD.n4412 153.601
R23292 VDD.n2356 VDD.n2353 153.601
R23293 VDD.n4422 VDD.n2348 153.601
R23294 VDD.n4416 VDD.n2353 153.601
R23295 VDD.n4423 VDD.n4422 153.601
R23296 VDD.n2343 VDD.n2340 153.601
R23297 VDD.n4432 VDD.n2336 153.601
R23298 VDD.n4426 VDD.n2340 153.601
R23299 VDD.n4433 VDD.n4432 153.601
R23300 VDD.n2326 VDD.n2314 153.601
R23301 VDD.n2325 VDD.n2312 153.601
R23302 VDD.n4447 VDD.n2314 153.601
R23303 VDD.n4446 VDD.n2312 153.601
R23304 VDD.n2319 VDD.n2307 153.601
R23305 VDD.n4456 VDD.n2306 153.601
R23306 VDD.n2301 VDD.n2298 153.601
R23307 VDD.n4466 VDD.n2294 153.601
R23308 VDD.n4460 VDD.n2298 153.601
R23309 VDD.n4467 VDD.n4466 153.601
R23310 VDD.n2289 VDD.n2286 153.601
R23311 VDD.n4476 VDD.n2281 153.601
R23312 VDD.n4470 VDD.n2286 153.601
R23313 VDD.n4477 VDD.n4476 153.601
R23314 VDD.n2276 VDD.n2273 153.601
R23315 VDD.n4486 VDD.n2271 153.601
R23316 VDD.n4480 VDD.n2273 153.601
R23317 VDD.n4487 VDD.n4486 153.601
R23318 VDD.n2266 VDD.n2263 153.601
R23319 VDD.n4496 VDD.n2260 153.601
R23320 VDD.n4490 VDD.n2263 153.601
R23321 VDD.n4497 VDD.n4496 153.601
R23322 VDD.n2321 VDD.n2307 153.601
R23323 VDD.n4457 VDD.n4456 153.601
R23324 VDD.n4260 VDD.n4257 153.601
R23325 VDD.n4267 VDD.n2518 153.601
R23326 VDD.n4261 VDD.n4257 153.601
R23327 VDD.n4268 VDD.n4267 153.601
R23328 VDD.n2513 VDD.n2510 153.601
R23329 VDD.n4277 VDD.n2508 153.601
R23330 VDD.n4271 VDD.n2510 153.601
R23331 VDD.n4278 VDD.n4277 153.601
R23332 VDD.n2503 VDD.n2500 153.601
R23333 VDD.n4287 VDD.n2497 153.601
R23334 VDD.n4281 VDD.n2500 153.601
R23335 VDD.n4288 VDD.n4287 153.601
R23336 VDD.n2492 VDD.n2489 153.601
R23337 VDD.n4297 VDD.n2484 153.601
R23338 VDD.n4291 VDD.n2489 153.601
R23339 VDD.n4298 VDD.n4297 153.601
R23340 VDD.n2479 VDD.n2476 153.601
R23341 VDD.n4307 VDD.n2472 153.601
R23342 VDD.n4301 VDD.n2476 153.601
R23343 VDD.n4308 VDD.n4307 153.601
R23344 VDD.n2462 VDD.n2450 153.601
R23345 VDD.n2461 VDD.n2448 153.601
R23346 VDD.n4322 VDD.n2450 153.601
R23347 VDD.n4321 VDD.n2448 153.601
R23348 VDD.n2455 VDD.n2443 153.601
R23349 VDD.n4331 VDD.n2442 153.601
R23350 VDD.n2437 VDD.n2434 153.601
R23351 VDD.n4341 VDD.n2430 153.601
R23352 VDD.n4335 VDD.n2434 153.601
R23353 VDD.n4342 VDD.n4341 153.601
R23354 VDD.n2425 VDD.n2422 153.601
R23355 VDD.n4351 VDD.n2417 153.601
R23356 VDD.n4345 VDD.n2422 153.601
R23357 VDD.n4352 VDD.n4351 153.601
R23358 VDD.n2412 VDD.n2409 153.601
R23359 VDD.n4361 VDD.n2407 153.601
R23360 VDD.n4355 VDD.n2409 153.601
R23361 VDD.n4362 VDD.n4361 153.601
R23362 VDD.n2402 VDD.n2399 153.601
R23363 VDD.n4371 VDD.n2396 153.601
R23364 VDD.n4365 VDD.n2399 153.601
R23365 VDD.n4372 VDD.n4371 153.601
R23366 VDD.n2457 VDD.n2443 153.601
R23367 VDD.n4332 VDD.n4331 153.601
R23368 VDD.n4135 VDD.n4132 153.601
R23369 VDD.n4142 VDD.n2654 153.601
R23370 VDD.n4136 VDD.n4132 153.601
R23371 VDD.n4143 VDD.n4142 153.601
R23372 VDD.n2649 VDD.n2646 153.601
R23373 VDD.n4152 VDD.n2644 153.601
R23374 VDD.n4146 VDD.n2646 153.601
R23375 VDD.n4153 VDD.n4152 153.601
R23376 VDD.n2639 VDD.n2636 153.601
R23377 VDD.n4162 VDD.n2633 153.601
R23378 VDD.n4156 VDD.n2636 153.601
R23379 VDD.n4163 VDD.n4162 153.601
R23380 VDD.n2628 VDD.n2625 153.601
R23381 VDD.n4172 VDD.n2620 153.601
R23382 VDD.n4166 VDD.n2625 153.601
R23383 VDD.n4173 VDD.n4172 153.601
R23384 VDD.n2615 VDD.n2612 153.601
R23385 VDD.n4182 VDD.n2608 153.601
R23386 VDD.n4176 VDD.n2612 153.601
R23387 VDD.n4183 VDD.n4182 153.601
R23388 VDD.n2598 VDD.n2586 153.601
R23389 VDD.n2597 VDD.n2584 153.601
R23390 VDD.n4197 VDD.n2586 153.601
R23391 VDD.n4196 VDD.n2584 153.601
R23392 VDD.n2591 VDD.n2579 153.601
R23393 VDD.n4206 VDD.n2578 153.601
R23394 VDD.n2573 VDD.n2570 153.601
R23395 VDD.n4216 VDD.n2566 153.601
R23396 VDD.n4210 VDD.n2570 153.601
R23397 VDD.n4217 VDD.n4216 153.601
R23398 VDD.n2561 VDD.n2558 153.601
R23399 VDD.n4226 VDD.n2553 153.601
R23400 VDD.n4220 VDD.n2558 153.601
R23401 VDD.n4227 VDD.n4226 153.601
R23402 VDD.n2548 VDD.n2545 153.601
R23403 VDD.n4236 VDD.n2543 153.601
R23404 VDD.n4230 VDD.n2545 153.601
R23405 VDD.n4237 VDD.n4236 153.601
R23406 VDD.n2538 VDD.n2535 153.601
R23407 VDD.n4246 VDD.n2532 153.601
R23408 VDD.n4240 VDD.n2535 153.601
R23409 VDD.n4247 VDD.n4246 153.601
R23410 VDD.n2593 VDD.n2579 153.601
R23411 VDD.n4207 VDD.n4206 153.601
R23412 VDD.n4010 VDD.n4007 153.601
R23413 VDD.n4017 VDD.n2790 153.601
R23414 VDD.n4011 VDD.n4007 153.601
R23415 VDD.n4018 VDD.n4017 153.601
R23416 VDD.n2785 VDD.n2782 153.601
R23417 VDD.n4027 VDD.n2780 153.601
R23418 VDD.n4021 VDD.n2782 153.601
R23419 VDD.n4028 VDD.n4027 153.601
R23420 VDD.n2775 VDD.n2772 153.601
R23421 VDD.n4037 VDD.n2769 153.601
R23422 VDD.n4031 VDD.n2772 153.601
R23423 VDD.n4038 VDD.n4037 153.601
R23424 VDD.n2764 VDD.n2761 153.601
R23425 VDD.n4047 VDD.n2756 153.601
R23426 VDD.n4041 VDD.n2761 153.601
R23427 VDD.n4048 VDD.n4047 153.601
R23428 VDD.n2751 VDD.n2748 153.601
R23429 VDD.n4057 VDD.n2744 153.601
R23430 VDD.n4051 VDD.n2748 153.601
R23431 VDD.n4058 VDD.n4057 153.601
R23432 VDD.n2734 VDD.n2722 153.601
R23433 VDD.n2733 VDD.n2720 153.601
R23434 VDD.n4072 VDD.n2722 153.601
R23435 VDD.n4071 VDD.n2720 153.601
R23436 VDD.n2727 VDD.n2715 153.601
R23437 VDD.n4081 VDD.n2714 153.601
R23438 VDD.n2709 VDD.n2706 153.601
R23439 VDD.n4091 VDD.n2702 153.601
R23440 VDD.n4085 VDD.n2706 153.601
R23441 VDD.n4092 VDD.n4091 153.601
R23442 VDD.n2697 VDD.n2694 153.601
R23443 VDD.n4101 VDD.n2689 153.601
R23444 VDD.n4095 VDD.n2694 153.601
R23445 VDD.n4102 VDD.n4101 153.601
R23446 VDD.n2684 VDD.n2681 153.601
R23447 VDD.n4111 VDD.n2679 153.601
R23448 VDD.n4105 VDD.n2681 153.601
R23449 VDD.n4112 VDD.n4111 153.601
R23450 VDD.n2674 VDD.n2671 153.601
R23451 VDD.n4121 VDD.n2668 153.601
R23452 VDD.n4115 VDD.n2671 153.601
R23453 VDD.n4122 VDD.n4121 153.601
R23454 VDD.n2729 VDD.n2715 153.601
R23455 VDD.n4082 VDD.n4081 153.601
R23456 VDD.n3885 VDD.n3882 153.601
R23457 VDD.n3892 VDD.n2926 153.601
R23458 VDD.n3886 VDD.n3882 153.601
R23459 VDD.n3893 VDD.n3892 153.601
R23460 VDD.n2921 VDD.n2918 153.601
R23461 VDD.n3902 VDD.n2916 153.601
R23462 VDD.n3896 VDD.n2918 153.601
R23463 VDD.n3903 VDD.n3902 153.601
R23464 VDD.n2911 VDD.n2908 153.601
R23465 VDD.n3912 VDD.n2905 153.601
R23466 VDD.n3906 VDD.n2908 153.601
R23467 VDD.n3913 VDD.n3912 153.601
R23468 VDD.n2900 VDD.n2897 153.601
R23469 VDD.n3922 VDD.n2892 153.601
R23470 VDD.n3916 VDD.n2897 153.601
R23471 VDD.n3923 VDD.n3922 153.601
R23472 VDD.n2887 VDD.n2884 153.601
R23473 VDD.n3932 VDD.n2880 153.601
R23474 VDD.n3926 VDD.n2884 153.601
R23475 VDD.n3933 VDD.n3932 153.601
R23476 VDD.n2870 VDD.n2858 153.601
R23477 VDD.n2869 VDD.n2856 153.601
R23478 VDD.n3947 VDD.n2858 153.601
R23479 VDD.n3946 VDD.n2856 153.601
R23480 VDD.n2863 VDD.n2851 153.601
R23481 VDD.n3956 VDD.n2850 153.601
R23482 VDD.n2845 VDD.n2842 153.601
R23483 VDD.n3966 VDD.n2838 153.601
R23484 VDD.n3960 VDD.n2842 153.601
R23485 VDD.n3967 VDD.n3966 153.601
R23486 VDD.n2833 VDD.n2830 153.601
R23487 VDD.n3976 VDD.n2825 153.601
R23488 VDD.n3970 VDD.n2830 153.601
R23489 VDD.n3977 VDD.n3976 153.601
R23490 VDD.n2820 VDD.n2817 153.601
R23491 VDD.n3986 VDD.n2815 153.601
R23492 VDD.n3980 VDD.n2817 153.601
R23493 VDD.n3987 VDD.n3986 153.601
R23494 VDD.n2810 VDD.n2807 153.601
R23495 VDD.n3996 VDD.n2804 153.601
R23496 VDD.n3990 VDD.n2807 153.601
R23497 VDD.n3997 VDD.n3996 153.601
R23498 VDD.n2865 VDD.n2851 153.601
R23499 VDD.n3957 VDD.n3956 153.601
R23500 VDD.n3234 VDD.n3231 153.601
R23501 VDD.n3534 VDD.n3230 153.601
R23502 VDD.n3225 VDD.n3222 153.601
R23503 VDD.n3544 VDD.n3220 153.601
R23504 VDD.n3538 VDD.n3222 153.601
R23505 VDD.n3545 VDD.n3544 153.601
R23506 VDD.n3213 VDD.n3208 153.601
R23507 VDD.n3212 VDD.n3206 153.601
R23508 VDD.n3552 VDD.n3208 153.601
R23509 VDD.n3551 VDD.n3206 153.601
R23510 VDD.n3235 VDD.n3231 153.601
R23511 VDD.n3535 VDD.n3534 153.601
R23512 VDD.n3760 VDD.n3757 153.601
R23513 VDD.n3767 VDD.n3752 153.601
R23514 VDD.n3761 VDD.n3757 153.601
R23515 VDD.n3768 VDD.n3767 153.601
R23516 VDD.n3747 VDD.n3744 153.601
R23517 VDD.n3777 VDD.n3742 153.601
R23518 VDD.n3771 VDD.n3744 153.601
R23519 VDD.n3778 VDD.n3777 153.601
R23520 VDD.n3737 VDD.n3734 153.601
R23521 VDD.n3787 VDD.n3731 153.601
R23522 VDD.n3781 VDD.n3734 153.601
R23523 VDD.n3788 VDD.n3787 153.601
R23524 VDD.n3726 VDD.n3723 153.601
R23525 VDD.n3797 VDD.n3718 153.601
R23526 VDD.n3791 VDD.n3723 153.601
R23527 VDD.n3798 VDD.n3797 153.601
R23528 VDD.n3713 VDD.n3710 153.601
R23529 VDD.n3807 VDD.n3706 153.601
R23530 VDD.n3801 VDD.n3710 153.601
R23531 VDD.n3808 VDD.n3807 153.601
R23532 VDD.n3696 VDD.n3684 153.601
R23533 VDD.n3695 VDD.n3682 153.601
R23534 VDD.n3822 VDD.n3684 153.601
R23535 VDD.n3821 VDD.n3682 153.601
R23536 VDD.n3689 VDD.n3677 153.601
R23537 VDD.n3831 VDD.n3676 153.601
R23538 VDD.n3671 VDD.n3668 153.601
R23539 VDD.n3841 VDD.n2974 153.601
R23540 VDD.n3835 VDD.n3668 153.601
R23541 VDD.n3842 VDD.n3841 153.601
R23542 VDD.n2969 VDD.n2966 153.601
R23543 VDD.n3851 VDD.n2961 153.601
R23544 VDD.n3845 VDD.n2966 153.601
R23545 VDD.n3852 VDD.n3851 153.601
R23546 VDD.n2956 VDD.n2953 153.601
R23547 VDD.n3861 VDD.n2951 153.601
R23548 VDD.n3855 VDD.n2953 153.601
R23549 VDD.n3862 VDD.n3861 153.601
R23550 VDD.n2946 VDD.n2943 153.601
R23551 VDD.n3871 VDD.n2940 153.601
R23552 VDD.n3865 VDD.n2943 153.601
R23553 VDD.n3872 VDD.n3871 153.601
R23554 VDD.n3691 VDD.n3677 153.601
R23555 VDD.n3832 VDD.n3831 153.601
R23556 VDD.n3087 VDD.t726 150.293
R23557 VDD.n3076 VDD.t756 150.293
R23558 VDD.n3103 VDD.t794 150.293
R23559 VDD.t752 VDD.n3112 150.293
R23560 VDD.n3151 VDD.t732 150.293
R23561 VDD.n3140 VDD.t808 150.293
R23562 VDD.n3167 VDD.t802 150.293
R23563 VDD.t776 VDD.n3176 150.293
R23564 VDD.n3048 VDD.t796 150.293
R23565 VDD.n3037 VDD.t714 150.293
R23566 VDD.n3191 VDD.t754 150.293
R23567 VDD.t740 VDD.n3200 150.293
R23568 VDD.n3302 VDD.t814 150.293
R23569 VDD.n3291 VDD.t786 150.293
R23570 VDD.n3568 VDD.t782 150.293
R23571 VDD.t766 VDD.n3577 150.293
R23572 VDD.n3009 VDD.t772 150.293
R23573 VDD.n2998 VDD.t730 150.293
R23574 VDD.n3025 VDD.t798 150.293
R23575 VDD.t720 VDD.n3034 150.293
R23576 VDD.n3596 VDD.t792 150.293
R23577 VDD.n3585 VDD.t758 150.293
R23578 VDD.n3612 VDD.t750 150.293
R23579 VDD.t734 VDD.n3621 150.293
R23580 VDD.t718 VDD.n2986 150.293
R23581 VDD.n3635 VDD.t774 150.293
R23582 VDD.t762 VDD.n3644 150.293
R23583 VDD.n3067 VDD.t812 150.293
R23584 VDD.n3056 VDD.t728 150.293
R23585 VDD.n3122 VDD.t746 150.293
R23586 VDD.t722 VDD.n3131 150.293
R23587 VDD.n3656 VDD.t770 150.293
R23588 VDD.t716 VDD.n3665 150.293
R23589 VDD.t804 VDD.n3084 150.273
R23590 VDD.t800 VDD.n3100 150.273
R23591 VDD.t810 VDD.n3148 150.273
R23592 VDD.t736 VDD.n3164 150.273
R23593 VDD.t724 VDD.n3045 150.273
R23594 VDD.t748 VDD.n3188 150.273
R23595 VDD.t788 VDD.n3299 150.273
R23596 VDD.t742 VDD.n3565 150.273
R23597 VDD.t806 VDD.n3006 150.273
R23598 VDD.t768 VDD.n3022 150.273
R23599 VDD.t760 VDD.n3593 150.273
R23600 VDD.t790 VDD.n3609 150.273
R23601 VDD.n2991 VDD.t780 150.273
R23602 VDD.n2980 VDD.t778 150.273
R23603 VDD.t738 VDD.n3632 150.273
R23604 VDD.t744 VDD.n3064 150.273
R23605 VDD.t784 VDD.n3119 150.273
R23606 VDD.t764 VDD.n3653 150.273
R23607 VDD.n7477 VDD.n7476 143.812
R23608 VDD.n7689 VDD.n7686 143.812
R23609 VDD.n7659 VDD.n7656 143.812
R23610 VDD.n7650 VDD.n7649 143.812
R23611 VDD.n7632 VDD.n7629 143.812
R23612 VDD.n1835 VDD.n1834 143.812
R23613 VDD.n1807 VDD.n1804 143.812
R23614 VDD.n1777 VDD.n1774 143.812
R23615 VDD.n1768 VDD.n1767 143.812
R23616 VDD.n1750 VDD.n1747 143.812
R23617 VDD.n1575 VDD.n1574 143.812
R23618 VDD.n1547 VDD.n1544 143.812
R23619 VDD.n1517 VDD.n1514 143.812
R23620 VDD.n1508 VDD.n1507 143.812
R23621 VDD.n1490 VDD.n1487 143.812
R23622 VDD.n1315 VDD.n1314 143.812
R23623 VDD.n1287 VDD.n1284 143.812
R23624 VDD.n1257 VDD.n1254 143.812
R23625 VDD.n1248 VDD.n1247 143.812
R23626 VDD.n1230 VDD.n1227 143.812
R23627 VDD.n1055 VDD.n1054 143.812
R23628 VDD.n1027 VDD.n1024 143.812
R23629 VDD.n997 VDD.n994 143.812
R23630 VDD.n988 VDD.n987 143.812
R23631 VDD.n970 VDD.n967 143.812
R23632 VDD.n795 VDD.n794 143.812
R23633 VDD.n767 VDD.n764 143.812
R23634 VDD.n737 VDD.n734 143.812
R23635 VDD.n728 VDD.n727 143.812
R23636 VDD.n710 VDD.n707 143.812
R23637 VDD.n535 VDD.n534 143.812
R23638 VDD.n507 VDD.n504 143.812
R23639 VDD.n477 VDD.n474 143.812
R23640 VDD.n468 VDD.n467 143.812
R23641 VDD.n450 VDD.n447 143.812
R23642 VDD.n7451 VDD.n7450 143.812
R23643 VDD.n7423 VDD.n7420 143.812
R23644 VDD.n7393 VDD.n7390 143.812
R23645 VDD.n7384 VDD.n7383 143.812
R23646 VDD.n7366 VDD.n7363 143.812
R23647 VDD.n7191 VDD.n7190 143.812
R23648 VDD.n7163 VDD.n7160 143.812
R23649 VDD.n7134 VDD.n7133 143.812
R23650 VDD.n7127 VDD.n7126 143.812
R23651 VDD.n7109 VDD.n7106 143.812
R23652 VDD.n6061 VDD.n6058 143.812
R23653 VDD.n6041 VDD.n6038 143.812
R23654 VDD.n6032 VDD.n6031 143.812
R23655 VDD.n6004 VDD.n6001 143.812
R23656 VDD.n5974 VDD.n5971 143.812
R23657 VDD.n6184 VDD.n6181 143.812
R23658 VDD.n6164 VDD.n6161 143.812
R23659 VDD.n6155 VDD.n6154 143.812
R23660 VDD.n6127 VDD.n6124 143.812
R23661 VDD.n6097 VDD.n6094 143.812
R23662 VDD.n6307 VDD.n6304 143.812
R23663 VDD.n6287 VDD.n6284 143.812
R23664 VDD.n6278 VDD.n6277 143.812
R23665 VDD.n6250 VDD.n6247 143.812
R23666 VDD.n6220 VDD.n6217 143.812
R23667 VDD.n6430 VDD.n6427 143.812
R23668 VDD.n6410 VDD.n6407 143.812
R23669 VDD.n6401 VDD.n6400 143.812
R23670 VDD.n6373 VDD.n6370 143.812
R23671 VDD.n6343 VDD.n6340 143.812
R23672 VDD.n6553 VDD.n6550 143.812
R23673 VDD.n6533 VDD.n6530 143.812
R23674 VDD.n6524 VDD.n6523 143.812
R23675 VDD.n6496 VDD.n6493 143.812
R23676 VDD.n6466 VDD.n6463 143.812
R23677 VDD.n6676 VDD.n6673 143.812
R23678 VDD.n6656 VDD.n6653 143.812
R23679 VDD.n6647 VDD.n6646 143.812
R23680 VDD.n6619 VDD.n6616 143.812
R23681 VDD.n6589 VDD.n6586 143.812
R23682 VDD.n6799 VDD.n6796 143.812
R23683 VDD.n6779 VDD.n6776 143.812
R23684 VDD.n6770 VDD.n6769 143.812
R23685 VDD.n6742 VDD.n6739 143.812
R23686 VDD.n6712 VDD.n6709 143.812
R23687 VDD.n4921 VDD.n4918 143.812
R23688 VDD.n4939 VDD.n4938 143.812
R23689 VDD.n4948 VDD.n4945 143.812
R23690 VDD.n4978 VDD.n4975 143.812
R23691 VDD.n5007 VDD.n5005 143.812
R23692 VDD.n4750 VDD.n4749 143.812
R23693 VDD.n4722 VDD.n4719 143.812
R23694 VDD.n4693 VDD.n4692 143.812
R23695 VDD.n4686 VDD.n4685 143.812
R23696 VDD.n4668 VDD.n4665 143.812
R23697 VDD.n4625 VDD.n4624 143.812
R23698 VDD.n4597 VDD.n4594 143.812
R23699 VDD.n4568 VDD.n4567 143.812
R23700 VDD.n4561 VDD.n4560 143.812
R23701 VDD.n4543 VDD.n4540 143.812
R23702 VDD.n4500 VDD.n4499 143.812
R23703 VDD.n4472 VDD.n4469 143.812
R23704 VDD.n4443 VDD.n4442 143.812
R23705 VDD.n4436 VDD.n4435 143.812
R23706 VDD.n4418 VDD.n4415 143.812
R23707 VDD.n4375 VDD.n4374 143.812
R23708 VDD.n4347 VDD.n4344 143.812
R23709 VDD.n4318 VDD.n4317 143.812
R23710 VDD.n4311 VDD.n4310 143.812
R23711 VDD.n4293 VDD.n4290 143.812
R23712 VDD.n4250 VDD.n4249 143.812
R23713 VDD.n4222 VDD.n4219 143.812
R23714 VDD.n4193 VDD.n4192 143.812
R23715 VDD.n4186 VDD.n4185 143.812
R23716 VDD.n4168 VDD.n4165 143.812
R23717 VDD.n4125 VDD.n4124 143.812
R23718 VDD.n4097 VDD.n4094 143.812
R23719 VDD.n4068 VDD.n4067 143.812
R23720 VDD.n4061 VDD.n4060 143.812
R23721 VDD.n4043 VDD.n4040 143.812
R23722 VDD.n4000 VDD.n3999 143.812
R23723 VDD.n3972 VDD.n3969 143.812
R23724 VDD.n3943 VDD.n3942 143.812
R23725 VDD.n3936 VDD.n3935 143.812
R23726 VDD.n3918 VDD.n3915 143.812
R23727 VDD.n3875 VDD.n3874 143.812
R23728 VDD.n3847 VDD.n3844 143.812
R23729 VDD.n3818 VDD.n3817 143.812
R23730 VDD.n3811 VDD.n3810 143.812
R23731 VDD.n3793 VDD.n3790 143.812
R23732 VDD.n7471 VDD.n7470 125.284
R23733 VDD.n1587 VDD.n1586 125.284
R23734 VDD.n1327 VDD.n1326 125.284
R23735 VDD.n1067 VDD.n1066 125.284
R23736 VDD.n807 VDD.n806 125.284
R23737 VDD.n547 VDD.n546 125.284
R23738 VDD.n287 VDD.n286 125.284
R23739 VDD.n7203 VDD.n7202 125.284
R23740 VDD.n1847 VDD.n1846 125.284
R23741 VDD.n5963 VDD.n5962 125.284
R23742 VDD.n5827 VDD.n5826 125.284
R23743 VDD.n5691 VDD.n5690 125.284
R23744 VDD.n5555 VDD.n5554 125.284
R23745 VDD.n5419 VDD.n5418 125.284
R23746 VDD.n5283 VDD.n5282 125.284
R23747 VDD.n5147 VDD.n5146 125.284
R23748 VDD.n5009 VDD.n5008 125.284
R23749 VDD.n1983 VDD.n1982 125.284
R23750 VDD.n2119 VDD.n2118 125.284
R23751 VDD.n2255 VDD.n2254 125.284
R23752 VDD.n2391 VDD.n2390 125.284
R23753 VDD.n2527 VDD.n2526 125.284
R23754 VDD.n2663 VDD.n2662 125.284
R23755 VDD.n2799 VDD.n2798 125.284
R23756 VDD.n2935 VDD.n2934 125.284
R23757 VDD.n7476 VDD.t943 123.344
R23758 VDD.t396 VDD.n7477 123.344
R23759 VDD.t396 VDD.n7707 123.344
R23760 VDD.n7706 VDD.t846 123.344
R23761 VDD.n7699 VDD.t846 123.344
R23762 VDD.n7696 VDD.t146 123.344
R23763 VDD.n7689 VDD.t146 123.344
R23764 VDD.n7686 VDD.t470 123.344
R23765 VDD.n7679 VDD.t470 123.344
R23766 VDD.n7676 VDD.t712 123.344
R23767 VDD.n7669 VDD.t712 123.344
R23768 VDD.n7666 VDD.t553 123.344
R23769 VDD.n7659 VDD.t553 123.344
R23770 VDD.n7656 VDD.t148 123.344
R23771 VDD.n7650 VDD.t148 123.344
R23772 VDD.n7649 VDD.t555 123.344
R23773 VDD.n7642 VDD.t555 123.344
R23774 VDD.n7639 VDD.t890 123.344
R23775 VDD.n7632 VDD.t890 123.344
R23776 VDD.n7629 VDD.t194 123.344
R23777 VDD.n7622 VDD.t194 123.344
R23778 VDD.n7619 VDD.t662 123.344
R23779 VDD.n7612 VDD.t662 123.344
R23780 VDD.n7609 VDD.t157 123.344
R23781 VDD.n7602 VDD.t157 123.344
R23782 VDD.n1835 VDD.t939 123.344
R23783 VDD.n1834 VDD.t289 123.344
R23784 VDD.n1827 VDD.t289 123.344
R23785 VDD.n1824 VDD.t843 123.344
R23786 VDD.n1817 VDD.t843 123.344
R23787 VDD.n1814 VDD.t131 123.344
R23788 VDD.n1807 VDD.t131 123.344
R23789 VDD.n1804 VDD.t580 123.344
R23790 VDD.n1797 VDD.t580 123.344
R23791 VDD.n1794 VDD.t593 123.344
R23792 VDD.n1787 VDD.t593 123.344
R23793 VDD.n1784 VDD.t371 123.344
R23794 VDD.n1777 VDD.t371 123.344
R23795 VDD.n1774 VDD.t133 123.344
R23796 VDD.n1768 VDD.t133 123.344
R23797 VDD.n1767 VDD.t369 123.344
R23798 VDD.n1760 VDD.t369 123.344
R23799 VDD.n1757 VDD.t670 123.344
R23800 VDD.n1750 VDD.t670 123.344
R23801 VDD.n1747 VDD.t293 123.344
R23802 VDD.n1740 VDD.t293 123.344
R23803 VDD.n1737 VDD.t587 123.344
R23804 VDD.n1730 VDD.t587 123.344
R23805 VDD.n1727 VDD.t5 123.344
R23806 VDD.n1720 VDD.t5 123.344
R23807 VDD.n1575 VDD.t852 123.344
R23808 VDD.n1574 VDD.t432 123.344
R23809 VDD.n1567 VDD.t432 123.344
R23810 VDD.n1564 VDD.t264 123.344
R23811 VDD.n1557 VDD.t264 123.344
R23812 VDD.n1554 VDD.t416 123.344
R23813 VDD.n1547 VDD.t416 123.344
R23814 VDD.n1544 VDD.t881 123.344
R23815 VDD.n1537 VDD.t881 123.344
R23816 VDD.n1534 VDD.t523 123.344
R23817 VDD.n1527 VDD.t523 123.344
R23818 VDD.n1524 VDD.t687 123.344
R23819 VDD.n1517 VDD.t687 123.344
R23820 VDD.n1514 VDD.t418 123.344
R23821 VDD.n1508 VDD.t418 123.344
R23822 VDD.n1507 VDD.t360 123.344
R23823 VDD.n1500 VDD.t360 123.344
R23824 VDD.n1497 VDD.t504 123.344
R23825 VDD.n1490 VDD.t504 123.344
R23826 VDD.n1487 VDD.t436 123.344
R23827 VDD.n1480 VDD.t436 123.344
R23828 VDD.n1477 VDD.t887 123.344
R23829 VDD.n1470 VDD.t887 123.344
R23830 VDD.n1467 VDD.t403 123.344
R23831 VDD.n1460 VDD.t403 123.344
R23832 VDD.n1315 VDD.t976 123.344
R23833 VDD.n1314 VDD.t71 123.344
R23834 VDD.n1307 VDD.t71 123.344
R23835 VDD.n1304 VDD.t226 123.344
R23836 VDD.n1297 VDD.t226 123.344
R23837 VDD.n1294 VDD.t140 123.344
R23838 VDD.n1287 VDD.t140 123.344
R23839 VDD.n1284 VDD.t129 123.344
R23840 VDD.n1277 VDD.t129 123.344
R23841 VDD.n1274 VDD.t190 123.344
R23842 VDD.n1267 VDD.t190 123.344
R23843 VDD.n1264 VDD.t238 123.344
R23844 VDD.n1257 VDD.t238 123.344
R23845 VDD.n1254 VDD.t142 123.344
R23846 VDD.n1248 VDD.t142 123.344
R23847 VDD.n1247 VDD.t230 123.344
R23848 VDD.n1240 VDD.t230 123.344
R23849 VDD.n1237 VDD.t442 123.344
R23850 VDD.n1230 VDD.t442 123.344
R23851 VDD.n1227 VDD.t67 123.344
R23852 VDD.n1220 VDD.t67 123.344
R23853 VDD.n1217 VDD.t13 123.344
R23854 VDD.n1210 VDD.t13 123.344
R23855 VDD.n1207 VDD.t188 123.344
R23856 VDD.n1200 VDD.t188 123.344
R23857 VDD.n1055 VDD.t941 123.344
R23858 VDD.n1054 VDD.t392 123.344
R23859 VDD.n1047 VDD.t392 123.344
R23860 VDD.n1044 VDD.t585 123.344
R23861 VDD.n1037 VDD.t585 123.344
R23862 VDD.n1034 VDD.t612 123.344
R23863 VDD.n1027 VDD.t612 123.344
R23864 VDD.n1024 VDD.t434 123.344
R23865 VDD.n1017 VDD.t434 123.344
R23866 VDD.n1014 VDD.t168 123.344
R23867 VDD.n1007 VDD.t168 123.344
R23868 VDD.n1004 VDD.t138 123.344
R23869 VDD.n997 VDD.t138 123.344
R23870 VDD.n994 VDD.t178 123.344
R23871 VDD.n988 VDD.t178 123.344
R23872 VDD.n987 VDD.t136 123.344
R23873 VDD.n980 VDD.t136 123.344
R23874 VDD.n977 VDD.t675 123.344
R23875 VDD.n970 VDD.t675 123.344
R23876 VDD.n967 VDD.t574 123.344
R23877 VDD.n960 VDD.t574 123.344
R23878 VDD.n957 VDD.t313 123.344
R23879 VDD.n950 VDD.t313 123.344
R23880 VDD.n947 VDD.t885 123.344
R23881 VDD.n940 VDD.t885 123.344
R23882 VDD.n795 VDD.t848 123.344
R23883 VDD.n794 VDD.t648 123.344
R23884 VDD.n787 VDD.t648 123.344
R23885 VDD.n784 VDD.t316 123.344
R23886 VDD.n777 VDD.t316 123.344
R23887 VDD.n774 VDD.t514 123.344
R23888 VDD.n767 VDD.t514 123.344
R23889 VDD.n764 VDD.t484 123.344
R23890 VDD.n757 VDD.t484 123.344
R23891 VDD.n754 VDD.t635 123.344
R23892 VDD.n747 VDD.t635 123.344
R23893 VDD.n744 VDD.t176 123.344
R23894 VDD.n737 VDD.t176 123.344
R23895 VDD.n734 VDD.t516 123.344
R23896 VDD.n728 VDD.t516 123.344
R23897 VDD.n727 VDD.t216 123.344
R23898 VDD.n720 VDD.t216 123.344
R23899 VDD.n717 VDD.t266 123.344
R23900 VDD.n710 VDD.t266 123.344
R23901 VDD.n707 VDD.t652 123.344
R23902 VDD.n700 VDD.t652 123.344
R23903 VDD.n697 VDD.t252 123.344
R23904 VDD.n690 VDD.t252 123.344
R23905 VDD.n687 VDD.t240 123.344
R23906 VDD.n680 VDD.t240 123.344
R23907 VDD.n535 VDD.t978 123.344
R23908 VDD.n534 VDD.t933 123.344
R23909 VDD.n527 VDD.t933 123.344
R23910 VDD.n524 VDD.t335 123.344
R23911 VDD.n517 VDD.t335 123.344
R23912 VDD.n514 VDD.t411 123.344
R23913 VDD.n507 VDD.t411 123.344
R23914 VDD.n504 VDD.t394 123.344
R23915 VDD.n497 VDD.t394 123.344
R23916 VDD.n494 VDD.t596 123.344
R23917 VDD.n487 VDD.t596 123.344
R23918 VDD.n484 VDD.t174 123.344
R23919 VDD.n477 VDD.t174 123.344
R23920 VDD.n474 VDD.t414 123.344
R23921 VDD.n468 VDD.t414 123.344
R23922 VDD.n467 VDD.t478 123.344
R23923 VDD.n460 VDD.t478 123.344
R23924 VDD.n457 VDD.t628 123.344
R23925 VDD.n450 VDD.t628 123.344
R23926 VDD.n447 VDD.t466 123.344
R23927 VDD.n440 VDD.t466 123.344
R23928 VDD.n437 VDD.t192 123.344
R23929 VDD.n430 VDD.t192 123.344
R23930 VDD.n427 VDD.t214 123.344
R23931 VDD.n420 VDD.t214 123.344
R23932 VDD.n7451 VDD.t850 123.344
R23933 VDD.n7450 VDD.t650 123.344
R23934 VDD.n7443 VDD.t650 123.344
R23935 VDD.n7440 VDD.t604 123.344
R23936 VDD.n7433 VDD.t604 123.344
R23937 VDD.n7430 VDD.t269 123.344
R23938 VDD.n7423 VDD.t269 123.344
R23939 VDD.n7420 VDD.t985 123.344
R23940 VDD.n7413 VDD.t985 123.344
R23941 VDD.n7410 VDD.t309 123.344
R23942 VDD.n7403 VDD.t309 123.344
R23943 VDD.n7400 VDD.t873 123.344
R23944 VDD.n7393 VDD.t873 123.344
R23945 VDD.n7390 VDD.t271 123.344
R23946 VDD.n7384 VDD.t271 123.344
R23947 VDD.n7383 VDD.t375 123.344
R23948 VDD.n7376 VDD.t375 123.344
R23949 VDD.n7373 VDD.t258 123.344
R23950 VDD.n7366 VDD.t258 123.344
R23951 VDD.n7363 VDD.t331 123.344
R23952 VDD.n7356 VDD.t331 123.344
R23953 VDD.n7353 VDD.t472 123.344
R23954 VDD.n7346 VDD.t472 123.344
R23955 VDD.n7343 VDD.t498 123.344
R23956 VDD.n7336 VDD.t498 123.344
R23957 VDD.n7191 VDD.t913 123.344
R23958 VDD.n7190 VDD.t29 123.344
R23959 VDD.n7183 VDD.t29 123.344
R23960 VDD.n7180 VDD.t455 123.344
R23961 VDD.n7173 VDD.t455 123.344
R23962 VDD.n7170 VDD.t1020 123.344
R23963 VDD.n7163 VDD.t1020 123.344
R23964 VDD.n7160 VDD.t91 123.344
R23965 VDD.n7153 VDD.t91 123.344
R23966 VDD.n7150 VDD.t228 123.344
R23967 VDD.n1915 VDD.t228 123.344
R23968 VDD.t423 VDD.n1916 123.344
R23969 VDD.t423 VDD.n7134 123.344
R23970 VDD.n7133 VDD.t1074 123.344
R23971 VDD.n7127 VDD.t1074 123.344
R23972 VDD.n7126 VDD.t305 123.344
R23973 VDD.n7119 VDD.t305 123.344
R23974 VDD.n7116 VDD.t969 123.344
R23975 VDD.n7109 VDD.t969 123.344
R23976 VDD.n7106 VDD.t113 123.344
R23977 VDD.n7099 VDD.t113 123.344
R23978 VDD.n7096 VDD.t897 123.344
R23979 VDD.n7089 VDD.t897 123.344
R23980 VDD.n7086 VDD.t480 123.344
R23981 VDD.n7079 VDD.t480 123.344
R23982 VDD.t390 VDD.n5838 123.344
R23983 VDD.t390 VDD.n6079 123.344
R23984 VDD.n6078 VDD.t706 123.344
R23985 VDD.n6071 VDD.t706 123.344
R23986 VDD.n6068 VDD.t121 123.344
R23987 VDD.n6061 VDD.t121 123.344
R23988 VDD.n6058 VDD.t297 123.344
R23989 VDD.n6051 VDD.t297 123.344
R23990 VDD.n6048 VDD.t274 123.344
R23991 VDD.n6041 VDD.t274 123.344
R23992 VDD.n6038 VDD.t1024 123.344
R23993 VDD.n6032 VDD.t1024 123.344
R23994 VDD.n6031 VDD.t276 123.344
R23995 VDD.n6024 VDD.t276 123.344
R23996 VDD.n6021 VDD.t219 123.344
R23997 VDD.n6014 VDD.t219 123.344
R23998 VDD.n6011 VDD.t125 123.344
R23999 VDD.n6004 VDD.t125 123.344
R24000 VDD.n6001 VDD.t1000 123.344
R24001 VDD.n5994 VDD.t1000 123.344
R24002 VDD.n5991 VDD.t343 123.344
R24003 VDD.n5984 VDD.t343 123.344
R24004 VDD.n5981 VDD.t85 123.344
R24005 VDD.n5974 VDD.t85 123.344
R24006 VDD.n5971 VDD.t345 123.344
R24007 VDD.t207 VDD.n5702 123.344
R24008 VDD.t207 VDD.n6202 123.344
R24009 VDD.n6201 VDD.t351 123.344
R24010 VDD.n6194 VDD.t351 123.344
R24011 VDD.n6191 VDD.t25 123.344
R24012 VDD.n6184 VDD.t25 123.344
R24013 VDD.n6181 VDD.t529 123.344
R24014 VDD.n6174 VDD.t529 123.344
R24015 VDD.n6171 VDD.t490 123.344
R24016 VDD.n6164 VDD.t490 123.344
R24017 VDD.n6161 VDD.t1079 123.344
R24018 VDD.n6155 VDD.t1079 123.344
R24019 VDD.n6154 VDD.t501 123.344
R24020 VDD.n6147 VDD.t501 123.344
R24021 VDD.n6144 VDD.t299 123.344
R24022 VDD.n6137 VDD.t299 123.344
R24023 VDD.n6134 VDD.t61 123.344
R24024 VDD.n6127 VDD.t61 123.344
R24025 VDD.n6124 VDD.t1056 123.344
R24026 VDD.n6117 VDD.t1056 123.344
R24027 VDD.n6114 VDD.t468 123.344
R24028 VDD.n6107 VDD.t468 123.344
R24029 VDD.n6104 VDD.t107 123.344
R24030 VDD.n6097 VDD.t107 123.344
R24031 VDD.n6094 VDD.t946 123.344
R24032 VDD.t311 VDD.n5566 123.344
R24033 VDD.t311 VDD.n6325 123.344
R24034 VDD.n6324 VDD.t184 123.344
R24035 VDD.n6317 VDD.t184 123.344
R24036 VDD.n6314 VDD.t103 123.344
R24037 VDD.n6307 VDD.t103 123.344
R24038 VDD.n6304 VDD.t855 123.344
R24039 VDD.n6297 VDD.t855 123.344
R24040 VDD.n6294 VDD.t301 123.344
R24041 VDD.n6287 VDD.t301 123.344
R24042 VDD.n6284 VDD.t1054 123.344
R24043 VDD.n6278 VDD.t1054 123.344
R24044 VDD.n6277 VDD.t303 123.344
R24045 VDD.n6270 VDD.t303 123.344
R24046 VDD.n6267 VDD.t548 123.344
R24047 VDD.n6260 VDD.t548 123.344
R24048 VDD.n6257 VDD.t43 123.344
R24049 VDD.n6250 VDD.t43 123.344
R24050 VDD.n6247 VDD.t1028 123.344
R24051 VDD.n6240 VDD.t1028 123.344
R24052 VDD.n6237 VDD.t377 123.344
R24053 VDD.n6230 VDD.t377 123.344
R24054 VDD.n6227 VDD.t53 123.344
R24055 VDD.n6220 VDD.t53 123.344
R24056 VDD.n6217 VDD.t209 123.344
R24057 VDD.t658 VDD.n5430 123.344
R24058 VDD.t658 VDD.n6448 123.344
R24059 VDD.n6447 VDD.t199 123.344
R24060 VDD.n6440 VDD.t199 123.344
R24061 VDD.n6437 VDD.t49 123.344
R24062 VDD.n6430 VDD.t49 123.344
R24063 VDD.n6427 VDD.t428 123.344
R24064 VDD.n6420 VDD.t428 123.344
R24065 VDD.n6417 VDD.t170 123.344
R24066 VDD.n6410 VDD.t170 123.344
R24067 VDD.n6407 VDD.t1089 123.344
R24068 VDD.n6401 VDD.t1089 123.344
R24069 VDD.n6400 VDD.t280 123.344
R24070 VDD.n6393 VDD.t280 123.344
R24071 VDD.n6390 VDD.t365 123.344
R24072 VDD.n6383 VDD.t365 123.344
R24073 VDD.n6380 VDD.t81 123.344
R24074 VDD.n6373 VDD.t81 123.344
R24075 VDD.n6370 VDD.t1002 123.344
R24076 VDD.n6363 VDD.t1002 123.344
R24077 VDD.n6360 VDD.t254 123.344
R24078 VDD.n6353 VDD.t254 123.344
R24079 VDD.n6350 VDD.t33 123.344
R24080 VDD.n6343 VDD.t33 123.344
R24081 VDD.n6340 VDD.t829 123.344
R24082 VDD.t151 VDD.n5294 123.344
R24083 VDD.t151 VDD.n6571 123.344
R24084 VDD.n6570 VDD.t447 123.344
R24085 VDD.n6563 VDD.t447 123.344
R24086 VDD.n6560 VDD.t83 123.344
R24087 VDD.n6553 VDD.t83 123.344
R24088 VDD.n6550 VDD.t363 123.344
R24089 VDD.n6543 VDD.t363 123.344
R24090 VDD.n6540 VDD.t15 123.344
R24091 VDD.n6533 VDD.t15 123.344
R24092 VDD.n6530 VDD.t1084 123.344
R24093 VDD.n6524 VDD.t1084 123.344
R24094 VDD.n6523 VDD.t21 123.344
R24095 VDD.n6516 VDD.t21 123.344
R24096 VDD.n6513 VDD.t615 123.344
R24097 VDD.n6506 VDD.t615 123.344
R24098 VDD.n6503 VDD.t65 123.344
R24099 VDD.n6496 VDD.t65 123.344
R24100 VDD.n6493 VDD.t1060 123.344
R24101 VDD.n6486 VDD.t1060 123.344
R24102 VDD.n6483 VDD.t172 123.344
R24103 VDD.n6476 VDD.t172 123.344
R24104 VDD.n6473 VDD.t69 123.344
R24105 VDD.n6466 VDD.t69 123.344
R24106 VDD.n6463 VDD.t837 123.344
R24107 VDD.t862 VDD.n5158 123.344
R24108 VDD.t862 VDD.n6694 123.344
R24109 VDD.n6693 VDD.t285 123.344
R24110 VDD.n6686 VDD.t285 123.344
R24111 VDD.n6683 VDD.t73 123.344
R24112 VDD.n6676 VDD.t73 123.344
R24113 VDD.n6673 VDD.t341 123.344
R24114 VDD.n6666 VDD.t341 123.344
R24115 VDD.n6663 VDD.t665 123.344
R24116 VDD.n6656 VDD.t665 123.344
R24117 VDD.n6653 VDD.t1058 123.344
R24118 VDD.n6647 VDD.t1058 123.344
R24119 VDD.n6646 VDD.t643 123.344
R24120 VDD.n6639 VDD.t643 123.344
R24121 VDD.n6636 VDD.t486 123.344
R24122 VDD.n6629 VDD.t486 123.344
R24123 VDD.n6626 VDD.t111 123.344
R24124 VDD.n6619 VDD.t111 123.344
R24125 VDD.n6616 VDD.t1032 123.344
R24126 VDD.n6609 VDD.t1032 123.344
R24127 VDD.n6606 VDD.t398 123.344
R24128 VDD.n6599 VDD.t398 123.344
R24129 VDD.n6596 VDD.t55 123.344
R24130 VDD.n6589 VDD.t55 123.344
R24131 VDD.n6586 VDD.t155 123.344
R24132 VDD.t937 VDD.n5022 123.344
R24133 VDD.t937 VDD.n6817 123.344
R24134 VDD.n6816 VDD.t144 123.344
R24135 VDD.n6809 VDD.t144 123.344
R24136 VDD.n6806 VDD.t23 123.344
R24137 VDD.n6799 VDD.t23 123.344
R24138 VDD.n6796 VDD.t507 123.344
R24139 VDD.n6789 VDD.t507 123.344
R24140 VDD.n6786 VDD.t9 123.344
R24141 VDD.n6779 VDD.t9 123.344
R24142 VDD.n6776 VDD.t1076 123.344
R24143 VDD.n6770 VDD.t1076 123.344
R24144 VDD.n6769 VDD.t11 123.344
R24145 VDD.n6762 VDD.t11 123.344
R24146 VDD.n6759 VDD.t561 123.344
R24147 VDD.n6752 VDD.t561 123.344
R24148 VDD.n6749 VDD.t99 123.344
R24149 VDD.n6742 VDD.t99 123.344
R24150 VDD.n6739 VDD.t1030 123.344
R24151 VDD.n6732 VDD.t1030 123.344
R24152 VDD.n6729 VDD.t598 123.344
R24153 VDD.n6722 VDD.t598 123.344
R24154 VDD.n6719 VDD.t47 123.344
R24155 VDD.n6712 VDD.t47 123.344
R24156 VDD.n6709 VDD.t566 123.344
R24157 VDD.n4888 VDD.t492 123.344
R24158 VDD.n4898 VDD.t492 123.344
R24159 VDD.n4901 VDD.t248 123.344
R24160 VDD.n4908 VDD.t248 123.344
R24161 VDD.n4911 VDD.t101 123.344
R24162 VDD.n4918 VDD.t101 123.344
R24163 VDD.n4921 VDD.t655 123.344
R24164 VDD.n4928 VDD.t655 123.344
R24165 VDD.n4931 VDD.t242 123.344
R24166 VDD.n4938 VDD.t242 123.344
R24167 VDD.n4939 VDD.t1052 123.344
R24168 VDD.n4945 VDD.t1052 123.344
R24169 VDD.n4948 VDD.t244 123.344
R24170 VDD.n4955 VDD.t244 123.344
R24171 VDD.n4958 VDD.t445 123.344
R24172 VDD.n4965 VDD.t445 123.344
R24173 VDD.n4968 VDD.t77 123.344
R24174 VDD.n4975 VDD.t77 123.344
R24175 VDD.n4978 VDD.t1004 123.344
R24176 VDD.n4985 VDD.t1004 123.344
R24177 VDD.n4988 VDD.t205 123.344
R24178 VDD.n4995 VDD.t205 123.344
R24179 VDD.n4998 VDD.t87 123.344
R24180 VDD.n5005 VDD.t87 123.344
R24181 VDD.t203 VDD.n5007 123.344
R24182 VDD.n4750 VDD.t2 123.344
R24183 VDD.n4749 VDD.t51 123.344
R24184 VDD.n4742 VDD.t51 123.344
R24185 VDD.n4739 VDD.t646 123.344
R24186 VDD.n4732 VDD.t646 123.344
R24187 VDD.n4729 VDD.t1016 123.344
R24188 VDD.n4722 VDD.t1016 123.344
R24189 VDD.n4719 VDD.t117 123.344
R24190 VDD.n4712 VDD.t117 123.344
R24191 VDD.n4709 VDD.t256 123.344
R24192 VDD.n2051 VDD.t256 123.344
R24193 VDD.t17 VDD.n2052 123.344
R24194 VDD.t17 VDD.n4693 123.344
R24195 VDD.n4692 VDD.t1068 123.344
R24196 VDD.n4686 VDD.t1068 123.344
R24197 VDD.n4685 VDD.t19 123.344
R24198 VDD.n4678 VDD.t19 123.344
R24199 VDD.n4675 VDD.t607 123.344
R24200 VDD.n4668 VDD.t607 123.344
R24201 VDD.n4665 VDD.t57 123.344
R24202 VDD.n4658 VDD.t57 123.344
R24203 VDD.n4655 VDD.t232 123.344
R24204 VDD.n4648 VDD.t232 123.344
R24205 VDD.n4645 VDD.t602 123.344
R24206 VDD.n4638 VDD.t602 123.344
R24207 VDD.n4625 VDD.t920 123.344
R24208 VDD.n4624 VDD.t89 123.344
R24209 VDD.n4617 VDD.t89 123.344
R24210 VDD.n4614 VDD.t186 123.344
R24211 VDD.n4607 VDD.t186 123.344
R24212 VDD.n4604 VDD.t1042 123.344
R24213 VDD.n4597 VDD.t1042 123.344
R24214 VDD.n4594 VDD.t39 123.344
R24215 VDD.n4587 VDD.t39 123.344
R24216 VDD.n4584 VDD.t512 123.344
R24217 VDD.n2187 VDD.t512 123.344
R24218 VDD.t221 VDD.n2188 123.344
R24219 VDD.t221 VDD.n4568 123.344
R24220 VDD.n4567 VDD.t1082 123.344
R24221 VDD.n4561 VDD.t1082 123.344
R24222 VDD.n4560 VDD.t223 123.344
R24223 VDD.n4553 VDD.t223 123.344
R24224 VDD.n4550 VDD.t685 123.344
R24225 VDD.n4543 VDD.t685 123.344
R24226 VDD.n4540 VDD.t63 123.344
R24227 VDD.n4533 VDD.t63 123.344
R24228 VDD.n4530 VDD.t460 123.344
R24229 VDD.n4523 VDD.t460 123.344
R24230 VDD.n4520 VDD.t578 123.344
R24231 VDD.n4513 VDD.t578 123.344
R24232 VDD.n4500 VDD.t291 123.344
R24233 VDD.n4499 VDD.t97 123.344
R24234 VDD.n4492 VDD.t97 123.344
R24235 VDD.n4489 VDD.t564 123.344
R24236 VDD.n4482 VDD.t564 123.344
R24237 VDD.n4479 VDD.t1050 123.344
R24238 VDD.n4472 VDD.t1050 123.344
R24239 VDD.n4469 VDD.t109 123.344
R24240 VDD.n4462 VDD.t109 123.344
R24241 VDD.n4459 VDD.t451 123.344
R24242 VDD.n2323 VDD.t451 123.344
R24243 VDD.t954 VDD.n2324 123.344
R24244 VDD.t954 VDD.n4443 123.344
R24245 VDD.n4442 VDD.t1010 123.344
R24246 VDD.n4436 VDD.t1010 123.344
R24247 VDD.n4435 VDD.t660 123.344
R24248 VDD.n4428 VDD.t660 123.344
R24249 VDD.n4425 VDD.t337 123.344
R24250 VDD.n4418 VDD.t337 123.344
R24251 VDD.n4415 VDD.t123 123.344
R24252 VDD.n4408 VDD.t123 123.344
R24253 VDD.n4405 VDD.t625 123.344
R24254 VDD.n4398 VDD.t625 123.344
R24255 VDD.n4395 VDD.t453 123.344
R24256 VDD.n4388 VDD.t453 123.344
R24257 VDD.n4375 VDD.t903 123.344
R24258 VDD.n4374 VDD.t95 123.344
R24259 VDD.n4367 VDD.t95 123.344
R24260 VDD.n4364 VDD.t591 123.344
R24261 VDD.n4357 VDD.t591 123.344
R24262 VDD.n4354 VDD.t1048 123.344
R24263 VDD.n4347 VDD.t1048 123.344
R24264 VDD.n4344 VDD.t31 123.344
R24265 VDD.n4337 VDD.t31 123.344
R24266 VDD.n4334 VDD.t426 123.344
R24267 VDD.n2459 VDD.t426 123.344
R24268 VDD.t236 VDD.n2460 123.344
R24269 VDD.t236 VDD.n4318 123.344
R24270 VDD.n4317 VDD.t1038 123.344
R24271 VDD.n4311 VDD.t1038 123.344
R24272 VDD.n4310 VDD.t234 123.344
R24273 VDD.n4303 VDD.t234 123.344
R24274 VDD.n4300 VDD.t262 123.344
R24275 VDD.n4293 VDD.t262 123.344
R24276 VDD.n4290 VDD.t41 123.344
R24277 VDD.n4283 VDD.t41 123.344
R24278 VDD.n4280 VDD.t322 123.344
R24279 VDD.n4273 VDD.t322 123.344
R24280 VDD.n4270 VDD.t355 123.344
R24281 VDD.n4263 VDD.t355 123.344
R24282 VDD.n4250 VDD.t571 123.344
R24283 VDD.n4249 VDD.t127 123.344
R24284 VDD.n4242 VDD.t127 123.344
R24285 VDD.n4239 VDD.t353 123.344
R24286 VDD.n4232 VDD.t353 123.344
R24287 VDD.n4229 VDD.t1022 123.344
R24288 VDD.n4222 VDD.t1022 123.344
R24289 VDD.n4219 VDD.t79 123.344
R24290 VDD.n4212 VDD.t79 123.344
R24291 VDD.n4209 VDD.t476 123.344
R24292 VDD.n2595 VDD.t476 123.344
R24293 VDD.t438 VDD.n2596 123.344
R24294 VDD.t438 VDD.n4193 123.344
R24295 VDD.n4192 VDD.t1062 123.344
R24296 VDD.n4186 VDD.t1062 123.344
R24297 VDD.n4185 VDD.t440 123.344
R24298 VDD.n4178 VDD.t440 123.344
R24299 VDD.n4175 VDD.t817 123.344
R24300 VDD.n4168 VDD.t817 123.344
R24301 VDD.n4165 VDD.t59 123.344
R24302 VDD.n4158 VDD.t59 123.344
R24303 VDD.n4155 VDD.t474 123.344
R24304 VDD.n4148 VDD.t474 123.344
R24305 VDD.n4145 VDD.t320 123.344
R24306 VDD.n4138 VDD.t320 123.344
R24307 VDD.n4125 VDD.t876 123.344
R24308 VDD.n4124 VDD.t45 123.344
R24309 VDD.n4117 VDD.t45 123.344
R24310 VDD.n4114 VDD.t318 123.344
R24311 VDD.n4107 VDD.t318 123.344
R24312 VDD.n4104 VDD.t1018 123.344
R24313 VDD.n4097 VDD.t1018 123.344
R24314 VDD.n4094 VDD.t105 123.344
R24315 VDD.n4087 VDD.t105 123.344
R24316 VDD.n4084 VDD.t925 123.344
R24317 VDD.n2731 VDD.t925 123.344
R24318 VDD.t525 VDD.n2732 123.344
R24319 VDD.t525 VDD.n4068 123.344
R24320 VDD.n4067 VDD.t1006 123.344
R24321 VDD.n4061 VDD.t1006 123.344
R24322 VDD.n4060 VDD.t527 123.344
R24323 VDD.n4053 VDD.t527 123.344
R24324 VDD.n4050 VDD.t295 123.344
R24325 VDD.n4043 VDD.t295 123.344
R24326 VDD.n4040 VDD.t115 123.344
R24327 VDD.n4033 VDD.t115 123.344
R24328 VDD.n4030 VDD.t0 123.344
R24329 VDD.n4023 VDD.t0 123.344
R24330 VDD.n4020 VDD.t182 123.344
R24331 VDD.n4013 VDD.t182 123.344
R24332 VDD.n4000 VDD.t1102 123.344
R24333 VDD.n3999 VDD.t93 123.344
R24334 VDD.n3992 VDD.t93 123.344
R24335 VDD.n3989 VDD.t180 123.344
R24336 VDD.n3982 VDD.t180 123.344
R24337 VDD.n3979 VDD.t1045 123.344
R24338 VDD.n3972 VDD.t1045 123.344
R24339 VDD.n3969 VDD.t27 123.344
R24340 VDD.n3962 VDD.t27 123.344
R24341 VDD.n3959 VDD.t373 123.344
R24342 VDD.n2867 VDD.t373 123.344
R24343 VDD.t510 VDD.n2868 123.344
R24344 VDD.t510 VDD.n3943 123.344
R24345 VDD.n3942 VDD.t1034 123.344
R24346 VDD.n3936 VDD.t1034 123.344
R24347 VDD.n3935 VDD.t543 123.344
R24348 VDD.n3928 VDD.t543 123.344
R24349 VDD.n3925 VDD.t166 123.344
R24350 VDD.n3918 VDD.t166 123.344
R24351 VDD.n3915 VDD.t37 123.344
R24352 VDD.n3908 VDD.t37 123.344
R24353 VDD.n3905 VDD.t704 123.344
R24354 VDD.n3898 VDD.t704 123.344
R24355 VDD.n3895 VDD.t689 123.344
R24356 VDD.n3888 VDD.t689 123.344
R24357 VDD.t160 VDD.n3211 123.344
R24358 VDD.t160 VDD.n3548 123.344
R24359 VDD.n3547 VDD.t315 123.344
R24360 VDD.n3540 VDD.t315 123.344
R24361 VDD.n3537 VDD.t282 123.344
R24362 VDD.n3237 VDD.t282 123.344
R24363 VDD.n3875 VDD.t696 123.344
R24364 VDD.n3874 VDD.t119 123.344
R24365 VDD.n3867 VDD.t119 123.344
R24366 VDD.n3864 VDD.t692 123.344
R24367 VDD.n3857 VDD.t692 123.344
R24368 VDD.n3854 VDD.t1014 123.344
R24369 VDD.n3847 VDD.t1014 123.344
R24370 VDD.n3844 VDD.t75 123.344
R24371 VDD.n3837 VDD.t75 123.344
R24372 VDD.n3834 VDD.t164 123.344
R24373 VDD.n3693 VDD.t164 123.344
R24374 VDD.t162 VDD.n3694 123.344
R24375 VDD.t162 VDD.n3818 123.344
R24376 VDD.n3817 VDD.t1094 123.344
R24377 VDD.n3811 VDD.t1094 123.344
R24378 VDD.n3810 VDD.t246 123.344
R24379 VDD.n3803 VDD.t246 123.344
R24380 VDD.n3800 VDD.t550 123.344
R24381 VDD.n3793 VDD.t550 123.344
R24382 VDD.n3790 VDD.t35 123.344
R24383 VDD.n3783 VDD.t35 123.344
R24384 VDD.n3780 VDD.t633 123.344
R24385 VDD.n3773 VDD.t633 123.344
R24386 VDD.n3770 VDD.t347 123.344
R24387 VDD.n3763 VDD.t347 123.344
R24388 VDD.n259 VDD.n258 99.0123
R24389 VDD.n260 VDD.n259 99.0123
R24390 VDD.n7707 VDD.n7706 75.5806
R24391 VDD.n7699 VDD.n7696 75.5806
R24392 VDD.n7679 VDD.n7676 75.5806
R24393 VDD.n7669 VDD.n7666 75.5806
R24394 VDD.n7642 VDD.n7639 75.5806
R24395 VDD.n7622 VDD.n7619 75.5806
R24396 VDD.n7612 VDD.n7609 75.5806
R24397 VDD.n1827 VDD.n1824 75.5806
R24398 VDD.n1817 VDD.n1814 75.5806
R24399 VDD.n1797 VDD.n1794 75.5806
R24400 VDD.n1787 VDD.n1784 75.5806
R24401 VDD.n1760 VDD.n1757 75.5806
R24402 VDD.n1740 VDD.n1737 75.5806
R24403 VDD.n1730 VDD.n1727 75.5806
R24404 VDD.n1567 VDD.n1564 75.5806
R24405 VDD.n1557 VDD.n1554 75.5806
R24406 VDD.n1537 VDD.n1534 75.5806
R24407 VDD.n1527 VDD.n1524 75.5806
R24408 VDD.n1500 VDD.n1497 75.5806
R24409 VDD.n1480 VDD.n1477 75.5806
R24410 VDD.n1470 VDD.n1467 75.5806
R24411 VDD.n1307 VDD.n1304 75.5806
R24412 VDD.n1297 VDD.n1294 75.5806
R24413 VDD.n1277 VDD.n1274 75.5806
R24414 VDD.n1267 VDD.n1264 75.5806
R24415 VDD.n1240 VDD.n1237 75.5806
R24416 VDD.n1220 VDD.n1217 75.5806
R24417 VDD.n1210 VDD.n1207 75.5806
R24418 VDD.n1047 VDD.n1044 75.5806
R24419 VDD.n1037 VDD.n1034 75.5806
R24420 VDD.n1017 VDD.n1014 75.5806
R24421 VDD.n1007 VDD.n1004 75.5806
R24422 VDD.n980 VDD.n977 75.5806
R24423 VDD.n960 VDD.n957 75.5806
R24424 VDD.n950 VDD.n947 75.5806
R24425 VDD.n787 VDD.n784 75.5806
R24426 VDD.n777 VDD.n774 75.5806
R24427 VDD.n757 VDD.n754 75.5806
R24428 VDD.n747 VDD.n744 75.5806
R24429 VDD.n720 VDD.n717 75.5806
R24430 VDD.n700 VDD.n697 75.5806
R24431 VDD.n690 VDD.n687 75.5806
R24432 VDD.n527 VDD.n524 75.5806
R24433 VDD.n517 VDD.n514 75.5806
R24434 VDD.n497 VDD.n494 75.5806
R24435 VDD.n487 VDD.n484 75.5806
R24436 VDD.n460 VDD.n457 75.5806
R24437 VDD.n440 VDD.n437 75.5806
R24438 VDD.n430 VDD.n427 75.5806
R24439 VDD.n7443 VDD.n7440 75.5806
R24440 VDD.n7433 VDD.n7430 75.5806
R24441 VDD.n7413 VDD.n7410 75.5806
R24442 VDD.n7403 VDD.n7400 75.5806
R24443 VDD.n7376 VDD.n7373 75.5806
R24444 VDD.n7356 VDD.n7353 75.5806
R24445 VDD.n7346 VDD.n7343 75.5806
R24446 VDD.n7183 VDD.n7180 75.5806
R24447 VDD.n7173 VDD.n7170 75.5806
R24448 VDD.n7153 VDD.n7150 75.5806
R24449 VDD.n1916 VDD.n1915 75.5806
R24450 VDD.n7119 VDD.n7116 75.5806
R24451 VDD.n7099 VDD.n7096 75.5806
R24452 VDD.n7089 VDD.n7086 75.5806
R24453 VDD.n6079 VDD.n6078 75.5806
R24454 VDD.n6071 VDD.n6068 75.5806
R24455 VDD.n6051 VDD.n6048 75.5806
R24456 VDD.n6024 VDD.n6021 75.5806
R24457 VDD.n6014 VDD.n6011 75.5806
R24458 VDD.n5994 VDD.n5991 75.5806
R24459 VDD.n5984 VDD.n5981 75.5806
R24460 VDD.n6202 VDD.n6201 75.5806
R24461 VDD.n6194 VDD.n6191 75.5806
R24462 VDD.n6174 VDD.n6171 75.5806
R24463 VDD.n6147 VDD.n6144 75.5806
R24464 VDD.n6137 VDD.n6134 75.5806
R24465 VDD.n6117 VDD.n6114 75.5806
R24466 VDD.n6107 VDD.n6104 75.5806
R24467 VDD.n6325 VDD.n6324 75.5806
R24468 VDD.n6317 VDD.n6314 75.5806
R24469 VDD.n6297 VDD.n6294 75.5806
R24470 VDD.n6270 VDD.n6267 75.5806
R24471 VDD.n6260 VDD.n6257 75.5806
R24472 VDD.n6240 VDD.n6237 75.5806
R24473 VDD.n6230 VDD.n6227 75.5806
R24474 VDD.n6448 VDD.n6447 75.5806
R24475 VDD.n6440 VDD.n6437 75.5806
R24476 VDD.n6420 VDD.n6417 75.5806
R24477 VDD.n6393 VDD.n6390 75.5806
R24478 VDD.n6383 VDD.n6380 75.5806
R24479 VDD.n6363 VDD.n6360 75.5806
R24480 VDD.n6353 VDD.n6350 75.5806
R24481 VDD.n6571 VDD.n6570 75.5806
R24482 VDD.n6563 VDD.n6560 75.5806
R24483 VDD.n6543 VDD.n6540 75.5806
R24484 VDD.n6516 VDD.n6513 75.5806
R24485 VDD.n6506 VDD.n6503 75.5806
R24486 VDD.n6486 VDD.n6483 75.5806
R24487 VDD.n6476 VDD.n6473 75.5806
R24488 VDD.n6694 VDD.n6693 75.5806
R24489 VDD.n6686 VDD.n6683 75.5806
R24490 VDD.n6666 VDD.n6663 75.5806
R24491 VDD.n6639 VDD.n6636 75.5806
R24492 VDD.n6629 VDD.n6626 75.5806
R24493 VDD.n6609 VDD.n6606 75.5806
R24494 VDD.n6599 VDD.n6596 75.5806
R24495 VDD.n6817 VDD.n6816 75.5806
R24496 VDD.n6809 VDD.n6806 75.5806
R24497 VDD.n6789 VDD.n6786 75.5806
R24498 VDD.n6762 VDD.n6759 75.5806
R24499 VDD.n6752 VDD.n6749 75.5806
R24500 VDD.n6732 VDD.n6729 75.5806
R24501 VDD.n6722 VDD.n6719 75.5806
R24502 VDD.n4901 VDD.n4898 75.5806
R24503 VDD.n4911 VDD.n4908 75.5806
R24504 VDD.n4931 VDD.n4928 75.5806
R24505 VDD.n4958 VDD.n4955 75.5806
R24506 VDD.n4968 VDD.n4965 75.5806
R24507 VDD.n4988 VDD.n4985 75.5806
R24508 VDD.n4998 VDD.n4995 75.5806
R24509 VDD.n4742 VDD.n4739 75.5806
R24510 VDD.n4732 VDD.n4729 75.5806
R24511 VDD.n4712 VDD.n4709 75.5806
R24512 VDD.n2052 VDD.n2051 75.5806
R24513 VDD.n4678 VDD.n4675 75.5806
R24514 VDD.n4658 VDD.n4655 75.5806
R24515 VDD.n4648 VDD.n4645 75.5806
R24516 VDD.n4617 VDD.n4614 75.5806
R24517 VDD.n4607 VDD.n4604 75.5806
R24518 VDD.n4587 VDD.n4584 75.5806
R24519 VDD.n2188 VDD.n2187 75.5806
R24520 VDD.n4553 VDD.n4550 75.5806
R24521 VDD.n4533 VDD.n4530 75.5806
R24522 VDD.n4523 VDD.n4520 75.5806
R24523 VDD.n4492 VDD.n4489 75.5806
R24524 VDD.n4482 VDD.n4479 75.5806
R24525 VDD.n4462 VDD.n4459 75.5806
R24526 VDD.n2324 VDD.n2323 75.5806
R24527 VDD.n4428 VDD.n4425 75.5806
R24528 VDD.n4408 VDD.n4405 75.5806
R24529 VDD.n4398 VDD.n4395 75.5806
R24530 VDD.n4367 VDD.n4364 75.5806
R24531 VDD.n4357 VDD.n4354 75.5806
R24532 VDD.n4337 VDD.n4334 75.5806
R24533 VDD.n2460 VDD.n2459 75.5806
R24534 VDD.n4303 VDD.n4300 75.5806
R24535 VDD.n4283 VDD.n4280 75.5806
R24536 VDD.n4273 VDD.n4270 75.5806
R24537 VDD.n4242 VDD.n4239 75.5806
R24538 VDD.n4232 VDD.n4229 75.5806
R24539 VDD.n4212 VDD.n4209 75.5806
R24540 VDD.n2596 VDD.n2595 75.5806
R24541 VDD.n4178 VDD.n4175 75.5806
R24542 VDD.n4158 VDD.n4155 75.5806
R24543 VDD.n4148 VDD.n4145 75.5806
R24544 VDD.n4117 VDD.n4114 75.5806
R24545 VDD.n4107 VDD.n4104 75.5806
R24546 VDD.n4087 VDD.n4084 75.5806
R24547 VDD.n2732 VDD.n2731 75.5806
R24548 VDD.n4053 VDD.n4050 75.5806
R24549 VDD.n4033 VDD.n4030 75.5806
R24550 VDD.n4023 VDD.n4020 75.5806
R24551 VDD.n3992 VDD.n3989 75.5806
R24552 VDD.n3982 VDD.n3979 75.5806
R24553 VDD.n3962 VDD.n3959 75.5806
R24554 VDD.n2868 VDD.n2867 75.5806
R24555 VDD.n3928 VDD.n3925 75.5806
R24556 VDD.n3908 VDD.n3905 75.5806
R24557 VDD.n3898 VDD.n3895 75.5806
R24558 VDD.n3548 VDD.n3547 75.5806
R24559 VDD.n3540 VDD.n3537 75.5806
R24560 VDD.n3867 VDD.n3864 75.5806
R24561 VDD.n3857 VDD.n3854 75.5806
R24562 VDD.n3837 VDD.n3834 75.5806
R24563 VDD.n3694 VDD.n3693 75.5806
R24564 VDD.n3803 VDD.n3800 75.5806
R24565 VDD.n3783 VDD.n3780 75.5806
R24566 VDD.n3773 VDD.n3770 75.5806
R24567 VDD.n3082 VDD.t1124 73.6406
R24568 VDD.n3098 VDD.t1110 73.6406
R24569 VDD.n3146 VDD.t1154 73.6406
R24570 VDD.n3162 VDD.t1151 73.6406
R24571 VDD.n3043 VDD.t1143 73.6406
R24572 VDD.n3186 VDD.t1133 73.6406
R24573 VDD.n3297 VDD.t1114 73.6406
R24574 VDD.n3563 VDD.t1147 73.6406
R24575 VDD.n3004 VDD.t1157 73.6406
R24576 VDD.n3020 VDD.t1119 73.6406
R24577 VDD.n3591 VDD.t1144 73.6406
R24578 VDD.n3607 VDD.t1109 73.6406
R24579 VDD.n2989 VDD.t1120 73.6406
R24580 VDD.n2978 VDD.t1140 73.6406
R24581 VDD.n3630 VDD.t1150 73.6406
R24582 VDD.n3062 VDD.t1136 73.6406
R24583 VDD.n3117 VDD.t1121 73.6406
R24584 VDD.n3651 VDD.t1123 73.6406
R24585 VDD.n3089 VDD.t1128 73.6304
R24586 VDD.n3078 VDD.t1113 73.6304
R24587 VDD.n3105 VDD.t1141 73.6304
R24588 VDD.n3095 VDD.t1132 73.6304
R24589 VDD.n3153 VDD.t1122 73.6304
R24590 VDD.n3142 VDD.t1156 73.6304
R24591 VDD.n3169 VDD.t1138 73.6304
R24592 VDD.n3159 VDD.t1155 73.6304
R24593 VDD.n3050 VDD.t1111 73.6304
R24594 VDD.n3039 VDD.t1135 73.6304
R24595 VDD.n3193 VDD.t1129 73.6304
R24596 VDD.n3183 VDD.t1130 73.6304
R24597 VDD.n3304 VDD.t1137 73.6304
R24598 VDD.n3293 VDD.t1152 73.6304
R24599 VDD.n3570 VDD.t1146 73.6304
R24600 VDD.n3560 VDD.t1115 73.6304
R24601 VDD.n3011 VDD.t1125 73.6304
R24602 VDD.n3000 VDD.t1126 73.6304
R24603 VDD.n3027 VDD.t1139 73.6304
R24604 VDD.n3017 VDD.t1158 73.6304
R24605 VDD.n3598 VDD.t1145 73.6304
R24606 VDD.n3587 VDD.t1112 73.6304
R24607 VDD.n3614 VDD.t1108 73.6304
R24608 VDD.n3604 VDD.t1131 73.6304
R24609 VDD.n2984 VDD.t1134 73.6304
R24610 VDD.n3637 VDD.t1148 73.6304
R24611 VDD.n3627 VDD.t1117 73.6304
R24612 VDD.n3069 VDD.t1153 73.6304
R24613 VDD.n3058 VDD.t1127 73.6304
R24614 VDD.n3124 VDD.t1116 73.6304
R24615 VDD.n3114 VDD.t1149 73.6304
R24616 VDD.n3658 VDD.t1118 73.6304
R24617 VDD.n3648 VDD.t1142 73.6304
R24618 VDD.n3334 VDD 71.7309
R24619 VDD.n3335 VDD.t916 69.9039
R24620 VDD VDD.t532 69.9004
R24621 VDD.n3345 VDD.t895 69.8804
R24622 VDD.n3340 VDD.t988 69.8804
R24623 VDD.n3429 VDD.t974 69.8804
R24624 VDD.n3440 VDD.t402 69.8804
R24625 VDD.n3435 VDD.t4 69.8804
R24626 VDD.n3523 VDD.t159 69.8804
R24627 VDD.n3282 VDD 63.2179
R24628 VDD.n3390 VDD 53.5114
R24629 VDD.n3391 VDD 43.8048
R24630 VDD.n7457 VDD.n7197 42.18
R24631 VDD.n7715 VDD.n7714 37.0005
R24632 VDD.n7714 VDD.t396 37.0005
R24633 VDD.n7481 VDD.n7480 37.0005
R24634 VDD.t396 VDD.n7481 37.0005
R24635 VDD.n7702 VDD.n7701 37.0005
R24636 VDD.n7701 VDD.t846 37.0005
R24637 VDD.n7489 VDD.n7488 37.0005
R24638 VDD.n7488 VDD.t846 37.0005
R24639 VDD.n7692 VDD.n7691 37.0005
R24640 VDD.n7691 VDD.t146 37.0005
R24641 VDD.n7502 VDD.n7501 37.0005
R24642 VDD.n7501 VDD.t146 37.0005
R24643 VDD.n7682 VDD.n7681 37.0005
R24644 VDD.n7681 VDD.t470 37.0005
R24645 VDD.n7513 VDD.n7512 37.0005
R24646 VDD.n7512 VDD.t470 37.0005
R24647 VDD.n7672 VDD.n7671 37.0005
R24648 VDD.n7671 VDD.t712 37.0005
R24649 VDD.n7523 VDD.n7522 37.0005
R24650 VDD.n7522 VDD.t712 37.0005
R24651 VDD.n7662 VDD.n7661 37.0005
R24652 VDD.n7661 VDD.t553 37.0005
R24653 VDD.n7536 VDD.n7535 37.0005
R24654 VDD.n7535 VDD.t553 37.0005
R24655 VDD.n7540 VDD.n7538 37.0005
R24656 VDD.n7538 VDD.t148 37.0005
R24657 VDD.n7653 VDD.n7539 37.0005
R24658 VDD.n7539 VDD.t148 37.0005
R24659 VDD.n7645 VDD.n7644 37.0005
R24660 VDD.n7644 VDD.t555 37.0005
R24661 VDD.n7551 VDD.n7550 37.0005
R24662 VDD.n7550 VDD.t555 37.0005
R24663 VDD.n7635 VDD.n7634 37.0005
R24664 VDD.n7634 VDD.t890 37.0005
R24665 VDD.n7564 VDD.n7563 37.0005
R24666 VDD.n7563 VDD.t890 37.0005
R24667 VDD.n7625 VDD.n7624 37.0005
R24668 VDD.n7624 VDD.t194 37.0005
R24669 VDD.n7575 VDD.n7574 37.0005
R24670 VDD.n7574 VDD.t194 37.0005
R24671 VDD.n7615 VDD.n7614 37.0005
R24672 VDD.n7614 VDD.t662 37.0005
R24673 VDD.n7585 VDD.n7584 37.0005
R24674 VDD.n7584 VDD.t662 37.0005
R24675 VDD.n7605 VDD.n7604 37.0005
R24676 VDD.n7604 VDD.t157 37.0005
R24677 VDD.n7598 VDD.n7597 37.0005
R24678 VDD.n7597 VDD.t157 37.0005
R24679 VDD.n7713 VDD.n7712 37.0005
R24680 VDD.t396 VDD.n7713 37.0005
R24681 VDD.n7715 VDD.n7463 37.0005
R24682 VDD.t396 VDD.n7463 37.0005
R24683 VDD.n7485 VDD.n7483 37.0005
R24684 VDD.n7483 VDD.t846 37.0005
R24685 VDD.n7702 VDD.n7484 37.0005
R24686 VDD.n7484 VDD.t846 37.0005
R24687 VDD.n7494 VDD.n7492 37.0005
R24688 VDD.n7492 VDD.t146 37.0005
R24689 VDD.n7692 VDD.n7493 37.0005
R24690 VDD.n7493 VDD.t146 37.0005
R24691 VDD.n7507 VDD.n7505 37.0005
R24692 VDD.n7505 VDD.t470 37.0005
R24693 VDD.n7682 VDD.n7506 37.0005
R24694 VDD.n7506 VDD.t470 37.0005
R24695 VDD.n7518 VDD.n7516 37.0005
R24696 VDD.n7516 VDD.t712 37.0005
R24697 VDD.n7672 VDD.n7517 37.0005
R24698 VDD.n7517 VDD.t712 37.0005
R24699 VDD.n7528 VDD.n7526 37.0005
R24700 VDD.n7526 VDD.t553 37.0005
R24701 VDD.n7662 VDD.n7527 37.0005
R24702 VDD.n7527 VDD.t553 37.0005
R24703 VDD.n7544 VDD.n7542 37.0005
R24704 VDD.n7542 VDD.t555 37.0005
R24705 VDD.n7645 VDD.n7543 37.0005
R24706 VDD.n7543 VDD.t555 37.0005
R24707 VDD.n7556 VDD.n7554 37.0005
R24708 VDD.n7554 VDD.t890 37.0005
R24709 VDD.n7635 VDD.n7555 37.0005
R24710 VDD.n7555 VDD.t890 37.0005
R24711 VDD.n7569 VDD.n7567 37.0005
R24712 VDD.n7567 VDD.t194 37.0005
R24713 VDD.n7625 VDD.n7568 37.0005
R24714 VDD.n7568 VDD.t194 37.0005
R24715 VDD.n7580 VDD.n7578 37.0005
R24716 VDD.n7578 VDD.t662 37.0005
R24717 VDD.n7615 VDD.n7579 37.0005
R24718 VDD.n7579 VDD.t662 37.0005
R24719 VDD.n7590 VDD.n7588 37.0005
R24720 VDD.n7588 VDD.t157 37.0005
R24721 VDD.n7605 VDD.n7589 37.0005
R24722 VDD.n7589 VDD.t157 37.0005
R24723 VDD.n7469 VDD.n7467 37.0005
R24724 VDD.n7467 VDD.t943 37.0005
R24725 VDD.n7473 VDD.n7468 37.0005
R24726 VDD.n1830 VDD.n1829 37.0005
R24727 VDD.n1829 VDD.t289 37.0005
R24728 VDD.n1597 VDD.n1596 37.0005
R24729 VDD.n1596 VDD.t289 37.0005
R24730 VDD.n1820 VDD.n1819 37.0005
R24731 VDD.n1819 VDD.t843 37.0005
R24732 VDD.n1607 VDD.n1606 37.0005
R24733 VDD.n1606 VDD.t843 37.0005
R24734 VDD.n1810 VDD.n1809 37.0005
R24735 VDD.n1809 VDD.t131 37.0005
R24736 VDD.n1620 VDD.n1619 37.0005
R24737 VDD.n1619 VDD.t131 37.0005
R24738 VDD.n1800 VDD.n1799 37.0005
R24739 VDD.n1799 VDD.t580 37.0005
R24740 VDD.n1631 VDD.n1630 37.0005
R24741 VDD.n1630 VDD.t580 37.0005
R24742 VDD.n1790 VDD.n1789 37.0005
R24743 VDD.n1789 VDD.t593 37.0005
R24744 VDD.n1641 VDD.n1640 37.0005
R24745 VDD.n1640 VDD.t593 37.0005
R24746 VDD.n1780 VDD.n1779 37.0005
R24747 VDD.n1779 VDD.t371 37.0005
R24748 VDD.n1654 VDD.n1653 37.0005
R24749 VDD.n1653 VDD.t371 37.0005
R24750 VDD.n1658 VDD.n1656 37.0005
R24751 VDD.n1656 VDD.t133 37.0005
R24752 VDD.n1771 VDD.n1657 37.0005
R24753 VDD.n1657 VDD.t133 37.0005
R24754 VDD.n1763 VDD.n1762 37.0005
R24755 VDD.n1762 VDD.t369 37.0005
R24756 VDD.n1669 VDD.n1668 37.0005
R24757 VDD.n1668 VDD.t369 37.0005
R24758 VDD.n1753 VDD.n1752 37.0005
R24759 VDD.n1752 VDD.t670 37.0005
R24760 VDD.n1682 VDD.n1681 37.0005
R24761 VDD.n1681 VDD.t670 37.0005
R24762 VDD.n1743 VDD.n1742 37.0005
R24763 VDD.n1742 VDD.t293 37.0005
R24764 VDD.n1693 VDD.n1692 37.0005
R24765 VDD.n1692 VDD.t293 37.0005
R24766 VDD.n1733 VDD.n1732 37.0005
R24767 VDD.n1732 VDD.t587 37.0005
R24768 VDD.n1703 VDD.n1702 37.0005
R24769 VDD.n1702 VDD.t587 37.0005
R24770 VDD.n1723 VDD.n1722 37.0005
R24771 VDD.n1722 VDD.t5 37.0005
R24772 VDD.n1716 VDD.n1715 37.0005
R24773 VDD.n1715 VDD.t5 37.0005
R24774 VDD.n1591 VDD.n1589 37.0005
R24775 VDD.n1589 VDD.t289 37.0005
R24776 VDD.n1830 VDD.n1590 37.0005
R24777 VDD.n1590 VDD.t289 37.0005
R24778 VDD.n1602 VDD.n1600 37.0005
R24779 VDD.n1600 VDD.t843 37.0005
R24780 VDD.n1820 VDD.n1601 37.0005
R24781 VDD.n1601 VDD.t843 37.0005
R24782 VDD.n1612 VDD.n1610 37.0005
R24783 VDD.n1610 VDD.t131 37.0005
R24784 VDD.n1810 VDD.n1611 37.0005
R24785 VDD.n1611 VDD.t131 37.0005
R24786 VDD.n1625 VDD.n1623 37.0005
R24787 VDD.n1623 VDD.t580 37.0005
R24788 VDD.n1800 VDD.n1624 37.0005
R24789 VDD.n1624 VDD.t580 37.0005
R24790 VDD.n1636 VDD.n1634 37.0005
R24791 VDD.n1634 VDD.t593 37.0005
R24792 VDD.n1790 VDD.n1635 37.0005
R24793 VDD.n1635 VDD.t593 37.0005
R24794 VDD.n1646 VDD.n1644 37.0005
R24795 VDD.n1644 VDD.t371 37.0005
R24796 VDD.n1780 VDD.n1645 37.0005
R24797 VDD.n1645 VDD.t371 37.0005
R24798 VDD.n1662 VDD.n1660 37.0005
R24799 VDD.n1660 VDD.t369 37.0005
R24800 VDD.n1763 VDD.n1661 37.0005
R24801 VDD.n1661 VDD.t369 37.0005
R24802 VDD.n1674 VDD.n1672 37.0005
R24803 VDD.n1672 VDD.t670 37.0005
R24804 VDD.n1753 VDD.n1673 37.0005
R24805 VDD.n1673 VDD.t670 37.0005
R24806 VDD.n1687 VDD.n1685 37.0005
R24807 VDD.n1685 VDD.t293 37.0005
R24808 VDD.n1743 VDD.n1686 37.0005
R24809 VDD.n1686 VDD.t293 37.0005
R24810 VDD.n1698 VDD.n1696 37.0005
R24811 VDD.n1696 VDD.t587 37.0005
R24812 VDD.n1733 VDD.n1697 37.0005
R24813 VDD.n1697 VDD.t587 37.0005
R24814 VDD.n1708 VDD.n1706 37.0005
R24815 VDD.n1706 VDD.t5 37.0005
R24816 VDD.n1723 VDD.n1707 37.0005
R24817 VDD.n1707 VDD.t5 37.0005
R24818 VDD.n1585 VDD.n1584 37.0005
R24819 VDD.t939 VDD.n1585 37.0005
R24820 VDD.n1838 VDD.n1583 37.0005
R24821 VDD.n1570 VDD.n1569 37.0005
R24822 VDD.n1569 VDD.t432 37.0005
R24823 VDD.n1337 VDD.n1336 37.0005
R24824 VDD.n1336 VDD.t432 37.0005
R24825 VDD.n1560 VDD.n1559 37.0005
R24826 VDD.n1559 VDD.t264 37.0005
R24827 VDD.n1347 VDD.n1346 37.0005
R24828 VDD.n1346 VDD.t264 37.0005
R24829 VDD.n1550 VDD.n1549 37.0005
R24830 VDD.n1549 VDD.t416 37.0005
R24831 VDD.n1360 VDD.n1359 37.0005
R24832 VDD.n1359 VDD.t416 37.0005
R24833 VDD.n1540 VDD.n1539 37.0005
R24834 VDD.n1539 VDD.t881 37.0005
R24835 VDD.n1371 VDD.n1370 37.0005
R24836 VDD.n1370 VDD.t881 37.0005
R24837 VDD.n1530 VDD.n1529 37.0005
R24838 VDD.n1529 VDD.t523 37.0005
R24839 VDD.n1381 VDD.n1380 37.0005
R24840 VDD.n1380 VDD.t523 37.0005
R24841 VDD.n1520 VDD.n1519 37.0005
R24842 VDD.n1519 VDD.t687 37.0005
R24843 VDD.n1394 VDD.n1393 37.0005
R24844 VDD.n1393 VDD.t687 37.0005
R24845 VDD.n1398 VDD.n1396 37.0005
R24846 VDD.n1396 VDD.t418 37.0005
R24847 VDD.n1511 VDD.n1397 37.0005
R24848 VDD.n1397 VDD.t418 37.0005
R24849 VDD.n1503 VDD.n1502 37.0005
R24850 VDD.n1502 VDD.t360 37.0005
R24851 VDD.n1409 VDD.n1408 37.0005
R24852 VDD.n1408 VDD.t360 37.0005
R24853 VDD.n1493 VDD.n1492 37.0005
R24854 VDD.n1492 VDD.t504 37.0005
R24855 VDD.n1422 VDD.n1421 37.0005
R24856 VDD.n1421 VDD.t504 37.0005
R24857 VDD.n1483 VDD.n1482 37.0005
R24858 VDD.n1482 VDD.t436 37.0005
R24859 VDD.n1433 VDD.n1432 37.0005
R24860 VDD.n1432 VDD.t436 37.0005
R24861 VDD.n1473 VDD.n1472 37.0005
R24862 VDD.n1472 VDD.t887 37.0005
R24863 VDD.n1443 VDD.n1442 37.0005
R24864 VDD.n1442 VDD.t887 37.0005
R24865 VDD.n1463 VDD.n1462 37.0005
R24866 VDD.n1462 VDD.t403 37.0005
R24867 VDD.n1456 VDD.n1455 37.0005
R24868 VDD.n1455 VDD.t403 37.0005
R24869 VDD.n1331 VDD.n1329 37.0005
R24870 VDD.n1329 VDD.t432 37.0005
R24871 VDD.n1570 VDD.n1330 37.0005
R24872 VDD.n1330 VDD.t432 37.0005
R24873 VDD.n1342 VDD.n1340 37.0005
R24874 VDD.n1340 VDD.t264 37.0005
R24875 VDD.n1560 VDD.n1341 37.0005
R24876 VDD.n1341 VDD.t264 37.0005
R24877 VDD.n1352 VDD.n1350 37.0005
R24878 VDD.n1350 VDD.t416 37.0005
R24879 VDD.n1550 VDD.n1351 37.0005
R24880 VDD.n1351 VDD.t416 37.0005
R24881 VDD.n1365 VDD.n1363 37.0005
R24882 VDD.n1363 VDD.t881 37.0005
R24883 VDD.n1540 VDD.n1364 37.0005
R24884 VDD.n1364 VDD.t881 37.0005
R24885 VDD.n1376 VDD.n1374 37.0005
R24886 VDD.n1374 VDD.t523 37.0005
R24887 VDD.n1530 VDD.n1375 37.0005
R24888 VDD.n1375 VDD.t523 37.0005
R24889 VDD.n1386 VDD.n1384 37.0005
R24890 VDD.n1384 VDD.t687 37.0005
R24891 VDD.n1520 VDD.n1385 37.0005
R24892 VDD.n1385 VDD.t687 37.0005
R24893 VDD.n1402 VDD.n1400 37.0005
R24894 VDD.n1400 VDD.t360 37.0005
R24895 VDD.n1503 VDD.n1401 37.0005
R24896 VDD.n1401 VDD.t360 37.0005
R24897 VDD.n1414 VDD.n1412 37.0005
R24898 VDD.n1412 VDD.t504 37.0005
R24899 VDD.n1493 VDD.n1413 37.0005
R24900 VDD.n1413 VDD.t504 37.0005
R24901 VDD.n1427 VDD.n1425 37.0005
R24902 VDD.n1425 VDD.t436 37.0005
R24903 VDD.n1483 VDD.n1426 37.0005
R24904 VDD.n1426 VDD.t436 37.0005
R24905 VDD.n1438 VDD.n1436 37.0005
R24906 VDD.n1436 VDD.t887 37.0005
R24907 VDD.n1473 VDD.n1437 37.0005
R24908 VDD.n1437 VDD.t887 37.0005
R24909 VDD.n1448 VDD.n1446 37.0005
R24910 VDD.n1446 VDD.t403 37.0005
R24911 VDD.n1463 VDD.n1447 37.0005
R24912 VDD.n1447 VDD.t403 37.0005
R24913 VDD.n1325 VDD.n1324 37.0005
R24914 VDD.t852 VDD.n1325 37.0005
R24915 VDD.n1578 VDD.n1323 37.0005
R24916 VDD.n1310 VDD.n1309 37.0005
R24917 VDD.n1309 VDD.t71 37.0005
R24918 VDD.n1077 VDD.n1076 37.0005
R24919 VDD.n1076 VDD.t71 37.0005
R24920 VDD.n1300 VDD.n1299 37.0005
R24921 VDD.n1299 VDD.t226 37.0005
R24922 VDD.n1087 VDD.n1086 37.0005
R24923 VDD.n1086 VDD.t226 37.0005
R24924 VDD.n1290 VDD.n1289 37.0005
R24925 VDD.n1289 VDD.t140 37.0005
R24926 VDD.n1100 VDD.n1099 37.0005
R24927 VDD.n1099 VDD.t140 37.0005
R24928 VDD.n1280 VDD.n1279 37.0005
R24929 VDD.n1279 VDD.t129 37.0005
R24930 VDD.n1111 VDD.n1110 37.0005
R24931 VDD.n1110 VDD.t129 37.0005
R24932 VDD.n1270 VDD.n1269 37.0005
R24933 VDD.n1269 VDD.t190 37.0005
R24934 VDD.n1121 VDD.n1120 37.0005
R24935 VDD.n1120 VDD.t190 37.0005
R24936 VDD.n1260 VDD.n1259 37.0005
R24937 VDD.n1259 VDD.t238 37.0005
R24938 VDD.n1134 VDD.n1133 37.0005
R24939 VDD.n1133 VDD.t238 37.0005
R24940 VDD.n1138 VDD.n1136 37.0005
R24941 VDD.n1136 VDD.t142 37.0005
R24942 VDD.n1251 VDD.n1137 37.0005
R24943 VDD.n1137 VDD.t142 37.0005
R24944 VDD.n1243 VDD.n1242 37.0005
R24945 VDD.n1242 VDD.t230 37.0005
R24946 VDD.n1149 VDD.n1148 37.0005
R24947 VDD.n1148 VDD.t230 37.0005
R24948 VDD.n1233 VDD.n1232 37.0005
R24949 VDD.n1232 VDD.t442 37.0005
R24950 VDD.n1162 VDD.n1161 37.0005
R24951 VDD.n1161 VDD.t442 37.0005
R24952 VDD.n1223 VDD.n1222 37.0005
R24953 VDD.n1222 VDD.t67 37.0005
R24954 VDD.n1173 VDD.n1172 37.0005
R24955 VDD.n1172 VDD.t67 37.0005
R24956 VDD.n1213 VDD.n1212 37.0005
R24957 VDD.n1212 VDD.t13 37.0005
R24958 VDD.n1183 VDD.n1182 37.0005
R24959 VDD.n1182 VDD.t13 37.0005
R24960 VDD.n1203 VDD.n1202 37.0005
R24961 VDD.n1202 VDD.t188 37.0005
R24962 VDD.n1196 VDD.n1195 37.0005
R24963 VDD.n1195 VDD.t188 37.0005
R24964 VDD.n1071 VDD.n1069 37.0005
R24965 VDD.n1069 VDD.t71 37.0005
R24966 VDD.n1310 VDD.n1070 37.0005
R24967 VDD.n1070 VDD.t71 37.0005
R24968 VDD.n1082 VDD.n1080 37.0005
R24969 VDD.n1080 VDD.t226 37.0005
R24970 VDD.n1300 VDD.n1081 37.0005
R24971 VDD.n1081 VDD.t226 37.0005
R24972 VDD.n1092 VDD.n1090 37.0005
R24973 VDD.n1090 VDD.t140 37.0005
R24974 VDD.n1290 VDD.n1091 37.0005
R24975 VDD.n1091 VDD.t140 37.0005
R24976 VDD.n1105 VDD.n1103 37.0005
R24977 VDD.n1103 VDD.t129 37.0005
R24978 VDD.n1280 VDD.n1104 37.0005
R24979 VDD.n1104 VDD.t129 37.0005
R24980 VDD.n1116 VDD.n1114 37.0005
R24981 VDD.n1114 VDD.t190 37.0005
R24982 VDD.n1270 VDD.n1115 37.0005
R24983 VDD.n1115 VDD.t190 37.0005
R24984 VDD.n1126 VDD.n1124 37.0005
R24985 VDD.n1124 VDD.t238 37.0005
R24986 VDD.n1260 VDD.n1125 37.0005
R24987 VDD.n1125 VDD.t238 37.0005
R24988 VDD.n1142 VDD.n1140 37.0005
R24989 VDD.n1140 VDD.t230 37.0005
R24990 VDD.n1243 VDD.n1141 37.0005
R24991 VDD.n1141 VDD.t230 37.0005
R24992 VDD.n1154 VDD.n1152 37.0005
R24993 VDD.n1152 VDD.t442 37.0005
R24994 VDD.n1233 VDD.n1153 37.0005
R24995 VDD.n1153 VDD.t442 37.0005
R24996 VDD.n1167 VDD.n1165 37.0005
R24997 VDD.n1165 VDD.t67 37.0005
R24998 VDD.n1223 VDD.n1166 37.0005
R24999 VDD.n1166 VDD.t67 37.0005
R25000 VDD.n1178 VDD.n1176 37.0005
R25001 VDD.n1176 VDD.t13 37.0005
R25002 VDD.n1213 VDD.n1177 37.0005
R25003 VDD.n1177 VDD.t13 37.0005
R25004 VDD.n1188 VDD.n1186 37.0005
R25005 VDD.n1186 VDD.t188 37.0005
R25006 VDD.n1203 VDD.n1187 37.0005
R25007 VDD.n1187 VDD.t188 37.0005
R25008 VDD.n1065 VDD.n1064 37.0005
R25009 VDD.t976 VDD.n1065 37.0005
R25010 VDD.n1318 VDD.n1063 37.0005
R25011 VDD.n1050 VDD.n1049 37.0005
R25012 VDD.n1049 VDD.t392 37.0005
R25013 VDD.n817 VDD.n816 37.0005
R25014 VDD.n816 VDD.t392 37.0005
R25015 VDD.n1040 VDD.n1039 37.0005
R25016 VDD.n1039 VDD.t585 37.0005
R25017 VDD.n827 VDD.n826 37.0005
R25018 VDD.n826 VDD.t585 37.0005
R25019 VDD.n1030 VDD.n1029 37.0005
R25020 VDD.n1029 VDD.t612 37.0005
R25021 VDD.n840 VDD.n839 37.0005
R25022 VDD.n839 VDD.t612 37.0005
R25023 VDD.n1020 VDD.n1019 37.0005
R25024 VDD.n1019 VDD.t434 37.0005
R25025 VDD.n851 VDD.n850 37.0005
R25026 VDD.n850 VDD.t434 37.0005
R25027 VDD.n1010 VDD.n1009 37.0005
R25028 VDD.n1009 VDD.t168 37.0005
R25029 VDD.n861 VDD.n860 37.0005
R25030 VDD.n860 VDD.t168 37.0005
R25031 VDD.n1000 VDD.n999 37.0005
R25032 VDD.n999 VDD.t138 37.0005
R25033 VDD.n874 VDD.n873 37.0005
R25034 VDD.n873 VDD.t138 37.0005
R25035 VDD.n878 VDD.n876 37.0005
R25036 VDD.n876 VDD.t178 37.0005
R25037 VDD.n991 VDD.n877 37.0005
R25038 VDD.n877 VDD.t178 37.0005
R25039 VDD.n983 VDD.n982 37.0005
R25040 VDD.n982 VDD.t136 37.0005
R25041 VDD.n889 VDD.n888 37.0005
R25042 VDD.n888 VDD.t136 37.0005
R25043 VDD.n973 VDD.n972 37.0005
R25044 VDD.n972 VDD.t675 37.0005
R25045 VDD.n902 VDD.n901 37.0005
R25046 VDD.n901 VDD.t675 37.0005
R25047 VDD.n963 VDD.n962 37.0005
R25048 VDD.n962 VDD.t574 37.0005
R25049 VDD.n913 VDD.n912 37.0005
R25050 VDD.n912 VDD.t574 37.0005
R25051 VDD.n953 VDD.n952 37.0005
R25052 VDD.n952 VDD.t313 37.0005
R25053 VDD.n923 VDD.n922 37.0005
R25054 VDD.n922 VDD.t313 37.0005
R25055 VDD.n943 VDD.n942 37.0005
R25056 VDD.n942 VDD.t885 37.0005
R25057 VDD.n936 VDD.n935 37.0005
R25058 VDD.n935 VDD.t885 37.0005
R25059 VDD.n811 VDD.n809 37.0005
R25060 VDD.n809 VDD.t392 37.0005
R25061 VDD.n1050 VDD.n810 37.0005
R25062 VDD.n810 VDD.t392 37.0005
R25063 VDD.n822 VDD.n820 37.0005
R25064 VDD.n820 VDD.t585 37.0005
R25065 VDD.n1040 VDD.n821 37.0005
R25066 VDD.n821 VDD.t585 37.0005
R25067 VDD.n832 VDD.n830 37.0005
R25068 VDD.n830 VDD.t612 37.0005
R25069 VDD.n1030 VDD.n831 37.0005
R25070 VDD.n831 VDD.t612 37.0005
R25071 VDD.n845 VDD.n843 37.0005
R25072 VDD.n843 VDD.t434 37.0005
R25073 VDD.n1020 VDD.n844 37.0005
R25074 VDD.n844 VDD.t434 37.0005
R25075 VDD.n856 VDD.n854 37.0005
R25076 VDD.n854 VDD.t168 37.0005
R25077 VDD.n1010 VDD.n855 37.0005
R25078 VDD.n855 VDD.t168 37.0005
R25079 VDD.n866 VDD.n864 37.0005
R25080 VDD.n864 VDD.t138 37.0005
R25081 VDD.n1000 VDD.n865 37.0005
R25082 VDD.n865 VDD.t138 37.0005
R25083 VDD.n882 VDD.n880 37.0005
R25084 VDD.n880 VDD.t136 37.0005
R25085 VDD.n983 VDD.n881 37.0005
R25086 VDD.n881 VDD.t136 37.0005
R25087 VDD.n894 VDD.n892 37.0005
R25088 VDD.n892 VDD.t675 37.0005
R25089 VDD.n973 VDD.n893 37.0005
R25090 VDD.n893 VDD.t675 37.0005
R25091 VDD.n907 VDD.n905 37.0005
R25092 VDD.n905 VDD.t574 37.0005
R25093 VDD.n963 VDD.n906 37.0005
R25094 VDD.n906 VDD.t574 37.0005
R25095 VDD.n918 VDD.n916 37.0005
R25096 VDD.n916 VDD.t313 37.0005
R25097 VDD.n953 VDD.n917 37.0005
R25098 VDD.n917 VDD.t313 37.0005
R25099 VDD.n928 VDD.n926 37.0005
R25100 VDD.n926 VDD.t885 37.0005
R25101 VDD.n943 VDD.n927 37.0005
R25102 VDD.n927 VDD.t885 37.0005
R25103 VDD.n805 VDD.n804 37.0005
R25104 VDD.t941 VDD.n805 37.0005
R25105 VDD.n1058 VDD.n803 37.0005
R25106 VDD.n790 VDD.n789 37.0005
R25107 VDD.n789 VDD.t648 37.0005
R25108 VDD.n557 VDD.n556 37.0005
R25109 VDD.n556 VDD.t648 37.0005
R25110 VDD.n780 VDD.n779 37.0005
R25111 VDD.n779 VDD.t316 37.0005
R25112 VDD.n567 VDD.n566 37.0005
R25113 VDD.n566 VDD.t316 37.0005
R25114 VDD.n770 VDD.n769 37.0005
R25115 VDD.n769 VDD.t514 37.0005
R25116 VDD.n580 VDD.n579 37.0005
R25117 VDD.n579 VDD.t514 37.0005
R25118 VDD.n760 VDD.n759 37.0005
R25119 VDD.n759 VDD.t484 37.0005
R25120 VDD.n591 VDD.n590 37.0005
R25121 VDD.n590 VDD.t484 37.0005
R25122 VDD.n750 VDD.n749 37.0005
R25123 VDD.n749 VDD.t635 37.0005
R25124 VDD.n601 VDD.n600 37.0005
R25125 VDD.n600 VDD.t635 37.0005
R25126 VDD.n740 VDD.n739 37.0005
R25127 VDD.n739 VDD.t176 37.0005
R25128 VDD.n614 VDD.n613 37.0005
R25129 VDD.n613 VDD.t176 37.0005
R25130 VDD.n618 VDD.n616 37.0005
R25131 VDD.n616 VDD.t516 37.0005
R25132 VDD.n731 VDD.n617 37.0005
R25133 VDD.n617 VDD.t516 37.0005
R25134 VDD.n723 VDD.n722 37.0005
R25135 VDD.n722 VDD.t216 37.0005
R25136 VDD.n629 VDD.n628 37.0005
R25137 VDD.n628 VDD.t216 37.0005
R25138 VDD.n713 VDD.n712 37.0005
R25139 VDD.n712 VDD.t266 37.0005
R25140 VDD.n642 VDD.n641 37.0005
R25141 VDD.n641 VDD.t266 37.0005
R25142 VDD.n703 VDD.n702 37.0005
R25143 VDD.n702 VDD.t652 37.0005
R25144 VDD.n653 VDD.n652 37.0005
R25145 VDD.n652 VDD.t652 37.0005
R25146 VDD.n693 VDD.n692 37.0005
R25147 VDD.n692 VDD.t252 37.0005
R25148 VDD.n663 VDD.n662 37.0005
R25149 VDD.n662 VDD.t252 37.0005
R25150 VDD.n683 VDD.n682 37.0005
R25151 VDD.n682 VDD.t240 37.0005
R25152 VDD.n676 VDD.n675 37.0005
R25153 VDD.n675 VDD.t240 37.0005
R25154 VDD.n551 VDD.n549 37.0005
R25155 VDD.n549 VDD.t648 37.0005
R25156 VDD.n790 VDD.n550 37.0005
R25157 VDD.n550 VDD.t648 37.0005
R25158 VDD.n562 VDD.n560 37.0005
R25159 VDD.n560 VDD.t316 37.0005
R25160 VDD.n780 VDD.n561 37.0005
R25161 VDD.n561 VDD.t316 37.0005
R25162 VDD.n572 VDD.n570 37.0005
R25163 VDD.n570 VDD.t514 37.0005
R25164 VDD.n770 VDD.n571 37.0005
R25165 VDD.n571 VDD.t514 37.0005
R25166 VDD.n585 VDD.n583 37.0005
R25167 VDD.n583 VDD.t484 37.0005
R25168 VDD.n760 VDD.n584 37.0005
R25169 VDD.n584 VDD.t484 37.0005
R25170 VDD.n596 VDD.n594 37.0005
R25171 VDD.n594 VDD.t635 37.0005
R25172 VDD.n750 VDD.n595 37.0005
R25173 VDD.n595 VDD.t635 37.0005
R25174 VDD.n606 VDD.n604 37.0005
R25175 VDD.n604 VDD.t176 37.0005
R25176 VDD.n740 VDD.n605 37.0005
R25177 VDD.n605 VDD.t176 37.0005
R25178 VDD.n622 VDD.n620 37.0005
R25179 VDD.n620 VDD.t216 37.0005
R25180 VDD.n723 VDD.n621 37.0005
R25181 VDD.n621 VDD.t216 37.0005
R25182 VDD.n634 VDD.n632 37.0005
R25183 VDD.n632 VDD.t266 37.0005
R25184 VDD.n713 VDD.n633 37.0005
R25185 VDD.n633 VDD.t266 37.0005
R25186 VDD.n647 VDD.n645 37.0005
R25187 VDD.n645 VDD.t652 37.0005
R25188 VDD.n703 VDD.n646 37.0005
R25189 VDD.n646 VDD.t652 37.0005
R25190 VDD.n658 VDD.n656 37.0005
R25191 VDD.n656 VDD.t252 37.0005
R25192 VDD.n693 VDD.n657 37.0005
R25193 VDD.n657 VDD.t252 37.0005
R25194 VDD.n668 VDD.n666 37.0005
R25195 VDD.n666 VDD.t240 37.0005
R25196 VDD.n683 VDD.n667 37.0005
R25197 VDD.n667 VDD.t240 37.0005
R25198 VDD.n545 VDD.n544 37.0005
R25199 VDD.t848 VDD.n545 37.0005
R25200 VDD.n798 VDD.n543 37.0005
R25201 VDD.n530 VDD.n529 37.0005
R25202 VDD.n529 VDD.t933 37.0005
R25203 VDD.n297 VDD.n296 37.0005
R25204 VDD.n296 VDD.t933 37.0005
R25205 VDD.n520 VDD.n519 37.0005
R25206 VDD.n519 VDD.t335 37.0005
R25207 VDD.n307 VDD.n306 37.0005
R25208 VDD.n306 VDD.t335 37.0005
R25209 VDD.n510 VDD.n509 37.0005
R25210 VDD.n509 VDD.t411 37.0005
R25211 VDD.n320 VDD.n319 37.0005
R25212 VDD.n319 VDD.t411 37.0005
R25213 VDD.n500 VDD.n499 37.0005
R25214 VDD.n499 VDD.t394 37.0005
R25215 VDD.n331 VDD.n330 37.0005
R25216 VDD.n330 VDD.t394 37.0005
R25217 VDD.n490 VDD.n489 37.0005
R25218 VDD.n489 VDD.t596 37.0005
R25219 VDD.n341 VDD.n340 37.0005
R25220 VDD.n340 VDD.t596 37.0005
R25221 VDD.n480 VDD.n479 37.0005
R25222 VDD.n479 VDD.t174 37.0005
R25223 VDD.n354 VDD.n353 37.0005
R25224 VDD.n353 VDD.t174 37.0005
R25225 VDD.n358 VDD.n356 37.0005
R25226 VDD.n356 VDD.t414 37.0005
R25227 VDD.n471 VDD.n357 37.0005
R25228 VDD.n357 VDD.t414 37.0005
R25229 VDD.n463 VDD.n462 37.0005
R25230 VDD.n462 VDD.t478 37.0005
R25231 VDD.n369 VDD.n368 37.0005
R25232 VDD.n368 VDD.t478 37.0005
R25233 VDD.n453 VDD.n452 37.0005
R25234 VDD.n452 VDD.t628 37.0005
R25235 VDD.n382 VDD.n381 37.0005
R25236 VDD.n381 VDD.t628 37.0005
R25237 VDD.n443 VDD.n442 37.0005
R25238 VDD.n442 VDD.t466 37.0005
R25239 VDD.n393 VDD.n392 37.0005
R25240 VDD.n392 VDD.t466 37.0005
R25241 VDD.n433 VDD.n432 37.0005
R25242 VDD.n432 VDD.t192 37.0005
R25243 VDD.n403 VDD.n402 37.0005
R25244 VDD.n402 VDD.t192 37.0005
R25245 VDD.n423 VDD.n422 37.0005
R25246 VDD.n422 VDD.t214 37.0005
R25247 VDD.n416 VDD.n415 37.0005
R25248 VDD.n415 VDD.t214 37.0005
R25249 VDD.n291 VDD.n289 37.0005
R25250 VDD.n289 VDD.t933 37.0005
R25251 VDD.n530 VDD.n290 37.0005
R25252 VDD.n290 VDD.t933 37.0005
R25253 VDD.n302 VDD.n300 37.0005
R25254 VDD.n300 VDD.t335 37.0005
R25255 VDD.n520 VDD.n301 37.0005
R25256 VDD.n301 VDD.t335 37.0005
R25257 VDD.n312 VDD.n310 37.0005
R25258 VDD.n310 VDD.t411 37.0005
R25259 VDD.n510 VDD.n311 37.0005
R25260 VDD.n311 VDD.t411 37.0005
R25261 VDD.n325 VDD.n323 37.0005
R25262 VDD.n323 VDD.t394 37.0005
R25263 VDD.n500 VDD.n324 37.0005
R25264 VDD.n324 VDD.t394 37.0005
R25265 VDD.n336 VDD.n334 37.0005
R25266 VDD.n334 VDD.t596 37.0005
R25267 VDD.n490 VDD.n335 37.0005
R25268 VDD.n335 VDD.t596 37.0005
R25269 VDD.n346 VDD.n344 37.0005
R25270 VDD.n344 VDD.t174 37.0005
R25271 VDD.n480 VDD.n345 37.0005
R25272 VDD.n345 VDD.t174 37.0005
R25273 VDD.n362 VDD.n360 37.0005
R25274 VDD.n360 VDD.t478 37.0005
R25275 VDD.n463 VDD.n361 37.0005
R25276 VDD.n361 VDD.t478 37.0005
R25277 VDD.n374 VDD.n372 37.0005
R25278 VDD.n372 VDD.t628 37.0005
R25279 VDD.n453 VDD.n373 37.0005
R25280 VDD.n373 VDD.t628 37.0005
R25281 VDD.n387 VDD.n385 37.0005
R25282 VDD.n385 VDD.t466 37.0005
R25283 VDD.n443 VDD.n386 37.0005
R25284 VDD.n386 VDD.t466 37.0005
R25285 VDD.n398 VDD.n396 37.0005
R25286 VDD.n396 VDD.t192 37.0005
R25287 VDD.n433 VDD.n397 37.0005
R25288 VDD.n397 VDD.t192 37.0005
R25289 VDD.n408 VDD.n406 37.0005
R25290 VDD.n406 VDD.t214 37.0005
R25291 VDD.n423 VDD.n407 37.0005
R25292 VDD.n407 VDD.t214 37.0005
R25293 VDD.n285 VDD.n284 37.0005
R25294 VDD.t978 VDD.n285 37.0005
R25295 VDD.n538 VDD.n283 37.0005
R25296 VDD.n273 VDD.n270 37.0005
R25297 VDD.n277 VDD.n269 37.0005
R25298 VDD.n261 VDD.n260 37.0005
R25299 VDD.n258 VDD.n257 37.0005
R25300 VDD.n257 VDD.t699 37.0005
R25301 VDD.n264 VDD.n263 37.0005
R25302 VDD.n263 VDD.t701 37.0005
R25303 VDD.n255 VDD.n246 37.0005
R25304 VDD.n101 VDD.n98 37.0005
R25305 VDD.n98 VDD.t197 37.0005
R25306 VDD.n105 VDD.n99 37.0005
R25307 VDD.n95 VDD.n94 37.0005
R25308 VDD.t379 VDD.n95 37.0005
R25309 VDD.n112 VDD.n93 37.0005
R25310 VDD.n84 VDD.n82 37.0005
R25311 VDD.n82 VDD.t1071 37.0005
R25312 VDD.n126 VDD.n83 37.0005
R25313 VDD.n83 VDD.t1071 37.0005
R25314 VDD.n115 VDD.n85 37.0005
R25315 VDD.n85 VDD.t250 37.0005
R25316 VDD.n119 VDD.n86 37.0005
R25317 VDD.n79 VDD.n78 37.0005
R25318 VDD.t859 VDD.n79 37.0005
R25319 VDD.n133 VDD.n77 37.0005
R25320 VDD.n136 VDD.n73 37.0005
R25321 VDD.n73 VDD.t827 37.0005
R25322 VDD.n140 VDD.n74 37.0005
R25323 VDD.n70 VDD.n69 37.0005
R25324 VDD.t993 VDD.n70 37.0005
R25325 VDD.n147 VDD.n68 37.0005
R25326 VDD.n59 VDD.n57 37.0005
R25327 VDD.n57 VDD.t1026 37.0005
R25328 VDD.n161 VDD.n58 37.0005
R25329 VDD.n58 VDD.t1026 37.0005
R25330 VDD.n150 VDD.n60 37.0005
R25331 VDD.n60 VDD.t7 37.0005
R25332 VDD.n154 VDD.n61 37.0005
R25333 VDD.n54 VDD.n53 37.0005
R25334 VDD.t326 VDD.n54 37.0005
R25335 VDD.n168 VDD.n52 37.0005
R25336 VDD.n171 VDD.n48 37.0005
R25337 VDD.n48 VDD.t153 37.0005
R25338 VDD.n175 VDD.n49 37.0005
R25339 VDD.n45 VDD.n44 37.0005
R25340 VDD.t568 VDD.n45 37.0005
R25341 VDD.n182 VDD.n43 37.0005
R25342 VDD.n34 VDD.n32 37.0005
R25343 VDD.n32 VDD.t1065 37.0005
R25344 VDD.n196 VDD.n33 37.0005
R25345 VDD.n33 VDD.t1065 37.0005
R25346 VDD.n185 VDD.n35 37.0005
R25347 VDD.n35 VDD.t821 37.0005
R25348 VDD.n189 VDD.n36 37.0005
R25349 VDD.n29 VDD.n28 37.0005
R25350 VDD.t637 VDD.n29 37.0005
R25351 VDD.n203 VDD.n27 37.0005
R25352 VDD.n206 VDD.n23 37.0005
R25353 VDD.n23 VDD.t201 37.0005
R25354 VDD.n210 VDD.n24 37.0005
R25355 VDD.n20 VDD.n19 37.0005
R25356 VDD.t910 VDD.n20 37.0005
R25357 VDD.n217 VDD.n18 37.0005
R25358 VDD.n9 VDD.n7 37.0005
R25359 VDD.n7 VDD.t1092 37.0005
R25360 VDD.n231 VDD.n8 37.0005
R25361 VDD.n8 VDD.t1092 37.0005
R25362 VDD.n220 VDD.n10 37.0005
R25363 VDD.n10 VDD.t539 37.0005
R25364 VDD.n224 VDD.n11 37.0005
R25365 VDD.n4 VDD.n3 37.0005
R25366 VDD.t834 VDD.n4 37.0005
R25367 VDD.n238 VDD.n2 37.0005
R25368 VDD.n7446 VDD.n7445 37.0005
R25369 VDD.n7445 VDD.t650 37.0005
R25370 VDD.n7213 VDD.n7212 37.0005
R25371 VDD.n7212 VDD.t650 37.0005
R25372 VDD.n7436 VDD.n7435 37.0005
R25373 VDD.n7435 VDD.t604 37.0005
R25374 VDD.n7223 VDD.n7222 37.0005
R25375 VDD.n7222 VDD.t604 37.0005
R25376 VDD.n7426 VDD.n7425 37.0005
R25377 VDD.n7425 VDD.t269 37.0005
R25378 VDD.n7236 VDD.n7235 37.0005
R25379 VDD.n7235 VDD.t269 37.0005
R25380 VDD.n7416 VDD.n7415 37.0005
R25381 VDD.n7415 VDD.t985 37.0005
R25382 VDD.n7247 VDD.n7246 37.0005
R25383 VDD.n7246 VDD.t985 37.0005
R25384 VDD.n7406 VDD.n7405 37.0005
R25385 VDD.n7405 VDD.t309 37.0005
R25386 VDD.n7257 VDD.n7256 37.0005
R25387 VDD.n7256 VDD.t309 37.0005
R25388 VDD.n7396 VDD.n7395 37.0005
R25389 VDD.n7395 VDD.t873 37.0005
R25390 VDD.n7270 VDD.n7269 37.0005
R25391 VDD.n7269 VDD.t873 37.0005
R25392 VDD.n7274 VDD.n7272 37.0005
R25393 VDD.n7272 VDD.t271 37.0005
R25394 VDD.n7387 VDD.n7273 37.0005
R25395 VDD.n7273 VDD.t271 37.0005
R25396 VDD.n7379 VDD.n7378 37.0005
R25397 VDD.n7378 VDD.t375 37.0005
R25398 VDD.n7285 VDD.n7284 37.0005
R25399 VDD.n7284 VDD.t375 37.0005
R25400 VDD.n7369 VDD.n7368 37.0005
R25401 VDD.n7368 VDD.t258 37.0005
R25402 VDD.n7298 VDD.n7297 37.0005
R25403 VDD.n7297 VDD.t258 37.0005
R25404 VDD.n7359 VDD.n7358 37.0005
R25405 VDD.n7358 VDD.t331 37.0005
R25406 VDD.n7309 VDD.n7308 37.0005
R25407 VDD.n7308 VDD.t331 37.0005
R25408 VDD.n7349 VDD.n7348 37.0005
R25409 VDD.n7348 VDD.t472 37.0005
R25410 VDD.n7319 VDD.n7318 37.0005
R25411 VDD.n7318 VDD.t472 37.0005
R25412 VDD.n7339 VDD.n7338 37.0005
R25413 VDD.n7338 VDD.t498 37.0005
R25414 VDD.n7332 VDD.n7331 37.0005
R25415 VDD.n7331 VDD.t498 37.0005
R25416 VDD.n7207 VDD.n7205 37.0005
R25417 VDD.n7205 VDD.t650 37.0005
R25418 VDD.n7446 VDD.n7206 37.0005
R25419 VDD.n7206 VDD.t650 37.0005
R25420 VDD.n7218 VDD.n7216 37.0005
R25421 VDD.n7216 VDD.t604 37.0005
R25422 VDD.n7436 VDD.n7217 37.0005
R25423 VDD.n7217 VDD.t604 37.0005
R25424 VDD.n7228 VDD.n7226 37.0005
R25425 VDD.n7226 VDD.t269 37.0005
R25426 VDD.n7426 VDD.n7227 37.0005
R25427 VDD.n7227 VDD.t269 37.0005
R25428 VDD.n7241 VDD.n7239 37.0005
R25429 VDD.n7239 VDD.t985 37.0005
R25430 VDD.n7416 VDD.n7240 37.0005
R25431 VDD.n7240 VDD.t985 37.0005
R25432 VDD.n7252 VDD.n7250 37.0005
R25433 VDD.n7250 VDD.t309 37.0005
R25434 VDD.n7406 VDD.n7251 37.0005
R25435 VDD.n7251 VDD.t309 37.0005
R25436 VDD.n7262 VDD.n7260 37.0005
R25437 VDD.n7260 VDD.t873 37.0005
R25438 VDD.n7396 VDD.n7261 37.0005
R25439 VDD.n7261 VDD.t873 37.0005
R25440 VDD.n7278 VDD.n7276 37.0005
R25441 VDD.n7276 VDD.t375 37.0005
R25442 VDD.n7379 VDD.n7277 37.0005
R25443 VDD.n7277 VDD.t375 37.0005
R25444 VDD.n7290 VDD.n7288 37.0005
R25445 VDD.n7288 VDD.t258 37.0005
R25446 VDD.n7369 VDD.n7289 37.0005
R25447 VDD.n7289 VDD.t258 37.0005
R25448 VDD.n7303 VDD.n7301 37.0005
R25449 VDD.n7301 VDD.t331 37.0005
R25450 VDD.n7359 VDD.n7302 37.0005
R25451 VDD.n7302 VDD.t331 37.0005
R25452 VDD.n7314 VDD.n7312 37.0005
R25453 VDD.n7312 VDD.t472 37.0005
R25454 VDD.n7349 VDD.n7313 37.0005
R25455 VDD.n7313 VDD.t472 37.0005
R25456 VDD.n7324 VDD.n7322 37.0005
R25457 VDD.n7322 VDD.t498 37.0005
R25458 VDD.n7339 VDD.n7323 37.0005
R25459 VDD.n7323 VDD.t498 37.0005
R25460 VDD.n7201 VDD.n7200 37.0005
R25461 VDD.t850 VDD.n7201 37.0005
R25462 VDD.n7454 VDD.n7199 37.0005
R25463 VDD.n7186 VDD.n7185 37.0005
R25464 VDD.n7185 VDD.t29 37.0005
R25465 VDD.n1857 VDD.n1856 37.0005
R25466 VDD.n1856 VDD.t29 37.0005
R25467 VDD.n7176 VDD.n7175 37.0005
R25468 VDD.n7175 VDD.t455 37.0005
R25469 VDD.n1867 VDD.n1866 37.0005
R25470 VDD.n1866 VDD.t455 37.0005
R25471 VDD.n7166 VDD.n7165 37.0005
R25472 VDD.n7165 VDD.t1020 37.0005
R25473 VDD.n1880 VDD.n1879 37.0005
R25474 VDD.n1879 VDD.t1020 37.0005
R25475 VDD.n7156 VDD.n7155 37.0005
R25476 VDD.n7155 VDD.t91 37.0005
R25477 VDD.n1892 VDD.n1891 37.0005
R25478 VDD.n1891 VDD.t91 37.0005
R25479 VDD.n1910 VDD.n1909 37.0005
R25480 VDD.n1909 VDD.t228 37.0005
R25481 VDD.n7142 VDD.n7141 37.0005
R25482 VDD.n7141 VDD.t423 37.0005
R25483 VDD.n1920 VDD.n1919 37.0005
R25484 VDD.t423 VDD.n1920 37.0005
R25485 VDD.n1923 VDD.n1921 37.0005
R25486 VDD.n1921 VDD.t1074 37.0005
R25487 VDD.n7130 VDD.n1922 37.0005
R25488 VDD.n1922 VDD.t1074 37.0005
R25489 VDD.n7122 VDD.n7121 37.0005
R25490 VDD.n7121 VDD.t305 37.0005
R25491 VDD.n1934 VDD.n1933 37.0005
R25492 VDD.n1933 VDD.t305 37.0005
R25493 VDD.n7112 VDD.n7111 37.0005
R25494 VDD.n7111 VDD.t969 37.0005
R25495 VDD.n1947 VDD.n1946 37.0005
R25496 VDD.n1946 VDD.t969 37.0005
R25497 VDD.n7102 VDD.n7101 37.0005
R25498 VDD.n7101 VDD.t113 37.0005
R25499 VDD.n1958 VDD.n1957 37.0005
R25500 VDD.n1957 VDD.t113 37.0005
R25501 VDD.n7092 VDD.n7091 37.0005
R25502 VDD.n7091 VDD.t897 37.0005
R25503 VDD.n1968 VDD.n1967 37.0005
R25504 VDD.n1967 VDD.t897 37.0005
R25505 VDD.n7082 VDD.n7081 37.0005
R25506 VDD.n7081 VDD.t480 37.0005
R25507 VDD.n7075 VDD.n7074 37.0005
R25508 VDD.n7074 VDD.t480 37.0005
R25509 VDD.n1845 VDD.n1844 37.0005
R25510 VDD.t913 VDD.n1845 37.0005
R25511 VDD.n7194 VDD.n1843 37.0005
R25512 VDD.n1851 VDD.n1849 37.0005
R25513 VDD.n1849 VDD.t29 37.0005
R25514 VDD.n7186 VDD.n1850 37.0005
R25515 VDD.n1850 VDD.t29 37.0005
R25516 VDD.n1862 VDD.n1860 37.0005
R25517 VDD.n1860 VDD.t455 37.0005
R25518 VDD.n7176 VDD.n1861 37.0005
R25519 VDD.n1861 VDD.t455 37.0005
R25520 VDD.n1872 VDD.n1870 37.0005
R25521 VDD.n1870 VDD.t1020 37.0005
R25522 VDD.n7166 VDD.n1871 37.0005
R25523 VDD.n1871 VDD.t1020 37.0005
R25524 VDD.n1885 VDD.n1883 37.0005
R25525 VDD.n1883 VDD.t91 37.0005
R25526 VDD.n7156 VDD.n1884 37.0005
R25527 VDD.n1884 VDD.t91 37.0005
R25528 VDD.n7140 VDD.n7139 37.0005
R25529 VDD.t423 VDD.n7140 37.0005
R25530 VDD.n7142 VDD.n1905 37.0005
R25531 VDD.t423 VDD.n1905 37.0005
R25532 VDD.n1927 VDD.n1925 37.0005
R25533 VDD.n1925 VDD.t305 37.0005
R25534 VDD.n7122 VDD.n1926 37.0005
R25535 VDD.n1926 VDD.t305 37.0005
R25536 VDD.n1939 VDD.n1937 37.0005
R25537 VDD.n1937 VDD.t969 37.0005
R25538 VDD.n7112 VDD.n1938 37.0005
R25539 VDD.n1938 VDD.t969 37.0005
R25540 VDD.n1952 VDD.n1950 37.0005
R25541 VDD.n1950 VDD.t113 37.0005
R25542 VDD.n7102 VDD.n1951 37.0005
R25543 VDD.n1951 VDD.t113 37.0005
R25544 VDD.n1963 VDD.n1961 37.0005
R25545 VDD.n1961 VDD.t897 37.0005
R25546 VDD.n7092 VDD.n1962 37.0005
R25547 VDD.n1962 VDD.t897 37.0005
R25548 VDD.n1973 VDD.n1971 37.0005
R25549 VDD.n1971 VDD.t480 37.0005
R25550 VDD.n7082 VDD.n1972 37.0005
R25551 VDD.n1972 VDD.t480 37.0005
R25552 VDD.n1897 VDD.n1895 37.0005
R25553 VDD.n1895 VDD.t228 37.0005
R25554 VDD.n7146 VDD.n1900 37.0005
R25555 VDD.n1900 VDD.t228 37.0005
R25556 VDD.n7146 VDD.n1896 37.0005
R25557 VDD.n1896 VDD.t228 37.0005
R25558 VDD.n6935 VDD.n6932 37.0005
R25559 VDD.n6932 VDD.t694 37.0005
R25560 VDD.n6939 VDD.n6933 37.0005
R25561 VDD.n6929 VDD.n6928 37.0005
R25562 VDD.t329 VDD.n6929 37.0005
R25563 VDD.n6946 VDD.n6927 37.0005
R25564 VDD.n6918 VDD.n6916 37.0005
R25565 VDD.n6916 VDD.t339 37.0005
R25566 VDD.n6960 VDD.n6917 37.0005
R25567 VDD.n6917 VDD.t339 37.0005
R25568 VDD.n6949 VDD.n6919 37.0005
R25569 VDD.n6919 VDD.t1036 37.0005
R25570 VDD.n6953 VDD.n6920 37.0005
R25571 VDD.n6913 VDD.n6912 37.0005
R25572 VDD.t324 VDD.n6913 37.0005
R25573 VDD.n6967 VDD.n6911 37.0005
R25574 VDD.n6970 VDD.n6907 37.0005
R25575 VDD.n6907 VDD.t878 37.0005
R25576 VDD.n6974 VDD.n6908 37.0005
R25577 VDD.n6904 VDD.n6903 37.0005
R25578 VDD.t357 VDD.n6904 37.0005
R25579 VDD.n6981 VDD.n6902 37.0005
R25580 VDD.n6893 VDD.n6891 37.0005
R25581 VDD.n6891 VDD.t620 37.0005
R25582 VDD.n6995 VDD.n6892 37.0005
R25583 VDD.n6892 VDD.t620 37.0005
R25584 VDD.n6984 VDD.n6894 37.0005
R25585 VDD.n6894 VDD.t1012 37.0005
R25586 VDD.n6988 VDD.n6895 37.0005
R25587 VDD.n6888 VDD.n6887 37.0005
R25588 VDD.t576 VDD.n6888 37.0005
R25589 VDD.n7002 VDD.n6886 37.0005
R25590 VDD.n7005 VDD.n6882 37.0005
R25591 VDD.n6882 VDD.t905 37.0005
R25592 VDD.n7009 VDD.n6883 37.0005
R25593 VDD.n6879 VDD.n6878 37.0005
R25594 VDD.t582 VDD.n6879 37.0005
R25595 VDD.n7016 VDD.n6877 37.0005
R25596 VDD.n6868 VDD.n6866 37.0005
R25597 VDD.n6866 VDD.t958 37.0005
R25598 VDD.n7030 VDD.n6867 37.0005
R25599 VDD.n6867 VDD.t958 37.0005
R25600 VDD.n7019 VDD.n6869 37.0005
R25601 VDD.n6869 VDD.t1040 37.0005
R25602 VDD.n7023 VDD.n6870 37.0005
R25603 VDD.n6863 VDD.n6862 37.0005
R25604 VDD.t600 VDD.n6863 37.0005
R25605 VDD.n7037 VDD.n6861 37.0005
R25606 VDD.n7040 VDD.n6857 37.0005
R25607 VDD.n6857 VDD.t870 37.0005
R25608 VDD.n7044 VDD.n6858 37.0005
R25609 VDD.n6854 VDD.n6853 37.0005
R25610 VDD.t367 VDD.n6854 37.0005
R25611 VDD.n7051 VDD.n6852 37.0005
R25612 VDD.n7066 VDD.n7065 37.0005
R25613 VDD.n7065 VDD.t409 37.0005
R25614 VDD.n7064 VDD.n7063 37.0005
R25615 VDD.t409 VDD.n7064 37.0005
R25616 VDD.n7054 VDD.n6847 37.0005
R25617 VDD.n6847 VDD.t1008 37.0005
R25618 VDD.n7058 VDD.n6848 37.0005
R25619 VDD.n6842 VDD.n6836 37.0005
R25620 VDD.n6836 VDD.t589 37.0005
R25621 VDD.n6838 VDD.n6835 37.0005
R25622 VDD.n5842 VDD.n5841 37.0005
R25623 VDD.t390 VDD.n5842 37.0005
R25624 VDD.n6074 VDD.n6073 37.0005
R25625 VDD.n6073 VDD.t706 37.0005
R25626 VDD.n5851 VDD.n5850 37.0005
R25627 VDD.n5850 VDD.t706 37.0005
R25628 VDD.n6064 VDD.n6063 37.0005
R25629 VDD.n6063 VDD.t121 37.0005
R25630 VDD.n5861 VDD.n5860 37.0005
R25631 VDD.n5860 VDD.t121 37.0005
R25632 VDD.n6054 VDD.n6053 37.0005
R25633 VDD.n6053 VDD.t297 37.0005
R25634 VDD.n5872 VDD.n5871 37.0005
R25635 VDD.n5871 VDD.t297 37.0005
R25636 VDD.n6044 VDD.n6043 37.0005
R25637 VDD.n6043 VDD.t274 37.0005
R25638 VDD.n5885 VDD.n5884 37.0005
R25639 VDD.n5884 VDD.t274 37.0005
R25640 VDD.n5889 VDD.n5887 37.0005
R25641 VDD.n5887 VDD.t1024 37.0005
R25642 VDD.n6035 VDD.n5888 37.0005
R25643 VDD.n5888 VDD.t1024 37.0005
R25644 VDD.n6027 VDD.n6026 37.0005
R25645 VDD.n6026 VDD.t276 37.0005
R25646 VDD.n5900 VDD.n5899 37.0005
R25647 VDD.n5899 VDD.t276 37.0005
R25648 VDD.n6017 VDD.n6016 37.0005
R25649 VDD.n6016 VDD.t219 37.0005
R25650 VDD.n5913 VDD.n5912 37.0005
R25651 VDD.n5912 VDD.t219 37.0005
R25652 VDD.n6007 VDD.n6006 37.0005
R25653 VDD.n6006 VDD.t125 37.0005
R25654 VDD.n5923 VDD.n5922 37.0005
R25655 VDD.n5922 VDD.t125 37.0005
R25656 VDD.n5997 VDD.n5996 37.0005
R25657 VDD.n5996 VDD.t1000 37.0005
R25658 VDD.n5934 VDD.n5933 37.0005
R25659 VDD.n5933 VDD.t1000 37.0005
R25660 VDD.n5987 VDD.n5986 37.0005
R25661 VDD.n5986 VDD.t343 37.0005
R25662 VDD.n5947 VDD.n5946 37.0005
R25663 VDD.n5946 VDD.t343 37.0005
R25664 VDD.n5977 VDD.n5976 37.0005
R25665 VDD.n5976 VDD.t85 37.0005
R25666 VDD.n5957 VDD.n5956 37.0005
R25667 VDD.n5956 VDD.t85 37.0005
R25668 VDD.n5846 VDD.n5844 37.0005
R25669 VDD.n5844 VDD.t706 37.0005
R25670 VDD.n6074 VDD.n5845 37.0005
R25671 VDD.n5845 VDD.t706 37.0005
R25672 VDD.n5856 VDD.n5854 37.0005
R25673 VDD.n5854 VDD.t121 37.0005
R25674 VDD.n6064 VDD.n5855 37.0005
R25675 VDD.n5855 VDD.t121 37.0005
R25676 VDD.n5866 VDD.n5864 37.0005
R25677 VDD.n5864 VDD.t297 37.0005
R25678 VDD.n6054 VDD.n5865 37.0005
R25679 VDD.n5865 VDD.t297 37.0005
R25680 VDD.n5877 VDD.n5875 37.0005
R25681 VDD.n5875 VDD.t274 37.0005
R25682 VDD.n6044 VDD.n5876 37.0005
R25683 VDD.n5876 VDD.t274 37.0005
R25684 VDD.n5893 VDD.n5891 37.0005
R25685 VDD.n5891 VDD.t276 37.0005
R25686 VDD.n6027 VDD.n5892 37.0005
R25687 VDD.n5892 VDD.t276 37.0005
R25688 VDD.n5905 VDD.n5903 37.0005
R25689 VDD.n5903 VDD.t219 37.0005
R25690 VDD.n6017 VDD.n5904 37.0005
R25691 VDD.n5904 VDD.t219 37.0005
R25692 VDD.n5918 VDD.n5916 37.0005
R25693 VDD.n5916 VDD.t125 37.0005
R25694 VDD.n6007 VDD.n5917 37.0005
R25695 VDD.n5917 VDD.t125 37.0005
R25696 VDD.n5928 VDD.n5926 37.0005
R25697 VDD.n5926 VDD.t1000 37.0005
R25698 VDD.n5997 VDD.n5927 37.0005
R25699 VDD.n5927 VDD.t1000 37.0005
R25700 VDD.n5939 VDD.n5937 37.0005
R25701 VDD.n5937 VDD.t343 37.0005
R25702 VDD.n5987 VDD.n5938 37.0005
R25703 VDD.n5938 VDD.t343 37.0005
R25704 VDD.n5952 VDD.n5950 37.0005
R25705 VDD.n5950 VDD.t85 37.0005
R25706 VDD.n5977 VDD.n5951 37.0005
R25707 VDD.n5951 VDD.t85 37.0005
R25708 VDD.n5961 VDD.n5959 37.0005
R25709 VDD.n5959 VDD.t345 37.0005
R25710 VDD.n5968 VDD.n5960 37.0005
R25711 VDD.n6085 VDD.n6084 37.0005
R25712 VDD.t390 VDD.n6085 37.0005
R25713 VDD.n6087 VDD.n6086 37.0005
R25714 VDD.n6086 VDD.t390 37.0005
R25715 VDD.n6087 VDD.n5834 37.0005
R25716 VDD.t390 VDD.n5834 37.0005
R25717 VDD.n5706 VDD.n5705 37.0005
R25718 VDD.t207 VDD.n5706 37.0005
R25719 VDD.n6197 VDD.n6196 37.0005
R25720 VDD.n6196 VDD.t351 37.0005
R25721 VDD.n5715 VDD.n5714 37.0005
R25722 VDD.n5714 VDD.t351 37.0005
R25723 VDD.n6187 VDD.n6186 37.0005
R25724 VDD.n6186 VDD.t25 37.0005
R25725 VDD.n5725 VDD.n5724 37.0005
R25726 VDD.n5724 VDD.t25 37.0005
R25727 VDD.n6177 VDD.n6176 37.0005
R25728 VDD.n6176 VDD.t529 37.0005
R25729 VDD.n5736 VDD.n5735 37.0005
R25730 VDD.n5735 VDD.t529 37.0005
R25731 VDD.n6167 VDD.n6166 37.0005
R25732 VDD.n6166 VDD.t490 37.0005
R25733 VDD.n5749 VDD.n5748 37.0005
R25734 VDD.n5748 VDD.t490 37.0005
R25735 VDD.n5753 VDD.n5751 37.0005
R25736 VDD.n5751 VDD.t1079 37.0005
R25737 VDD.n6158 VDD.n5752 37.0005
R25738 VDD.n5752 VDD.t1079 37.0005
R25739 VDD.n6150 VDD.n6149 37.0005
R25740 VDD.n6149 VDD.t501 37.0005
R25741 VDD.n5764 VDD.n5763 37.0005
R25742 VDD.n5763 VDD.t501 37.0005
R25743 VDD.n6140 VDD.n6139 37.0005
R25744 VDD.n6139 VDD.t299 37.0005
R25745 VDD.n5777 VDD.n5776 37.0005
R25746 VDD.n5776 VDD.t299 37.0005
R25747 VDD.n6130 VDD.n6129 37.0005
R25748 VDD.n6129 VDD.t61 37.0005
R25749 VDD.n5787 VDD.n5786 37.0005
R25750 VDD.n5786 VDD.t61 37.0005
R25751 VDD.n6120 VDD.n6119 37.0005
R25752 VDD.n6119 VDD.t1056 37.0005
R25753 VDD.n5798 VDD.n5797 37.0005
R25754 VDD.n5797 VDD.t1056 37.0005
R25755 VDD.n6110 VDD.n6109 37.0005
R25756 VDD.n6109 VDD.t468 37.0005
R25757 VDD.n5811 VDD.n5810 37.0005
R25758 VDD.n5810 VDD.t468 37.0005
R25759 VDD.n6100 VDD.n6099 37.0005
R25760 VDD.n6099 VDD.t107 37.0005
R25761 VDD.n5821 VDD.n5820 37.0005
R25762 VDD.n5820 VDD.t107 37.0005
R25763 VDD.n5710 VDD.n5708 37.0005
R25764 VDD.n5708 VDD.t351 37.0005
R25765 VDD.n6197 VDD.n5709 37.0005
R25766 VDD.n5709 VDD.t351 37.0005
R25767 VDD.n5720 VDD.n5718 37.0005
R25768 VDD.n5718 VDD.t25 37.0005
R25769 VDD.n6187 VDD.n5719 37.0005
R25770 VDD.n5719 VDD.t25 37.0005
R25771 VDD.n5730 VDD.n5728 37.0005
R25772 VDD.n5728 VDD.t529 37.0005
R25773 VDD.n6177 VDD.n5729 37.0005
R25774 VDD.n5729 VDD.t529 37.0005
R25775 VDD.n5741 VDD.n5739 37.0005
R25776 VDD.n5739 VDD.t490 37.0005
R25777 VDD.n6167 VDD.n5740 37.0005
R25778 VDD.n5740 VDD.t490 37.0005
R25779 VDD.n5757 VDD.n5755 37.0005
R25780 VDD.n5755 VDD.t501 37.0005
R25781 VDD.n6150 VDD.n5756 37.0005
R25782 VDD.n5756 VDD.t501 37.0005
R25783 VDD.n5769 VDD.n5767 37.0005
R25784 VDD.n5767 VDD.t299 37.0005
R25785 VDD.n6140 VDD.n5768 37.0005
R25786 VDD.n5768 VDD.t299 37.0005
R25787 VDD.n5782 VDD.n5780 37.0005
R25788 VDD.n5780 VDD.t61 37.0005
R25789 VDD.n6130 VDD.n5781 37.0005
R25790 VDD.n5781 VDD.t61 37.0005
R25791 VDD.n5792 VDD.n5790 37.0005
R25792 VDD.n5790 VDD.t1056 37.0005
R25793 VDD.n6120 VDD.n5791 37.0005
R25794 VDD.n5791 VDD.t1056 37.0005
R25795 VDD.n5803 VDD.n5801 37.0005
R25796 VDD.n5801 VDD.t468 37.0005
R25797 VDD.n6110 VDD.n5802 37.0005
R25798 VDD.n5802 VDD.t468 37.0005
R25799 VDD.n5816 VDD.n5814 37.0005
R25800 VDD.n5814 VDD.t107 37.0005
R25801 VDD.n6100 VDD.n5815 37.0005
R25802 VDD.n5815 VDD.t107 37.0005
R25803 VDD.n5825 VDD.n5823 37.0005
R25804 VDD.n5823 VDD.t946 37.0005
R25805 VDD.n6091 VDD.n5824 37.0005
R25806 VDD.n6208 VDD.n6207 37.0005
R25807 VDD.t207 VDD.n6208 37.0005
R25808 VDD.n6210 VDD.n6209 37.0005
R25809 VDD.n6209 VDD.t207 37.0005
R25810 VDD.n6210 VDD.n5698 37.0005
R25811 VDD.t207 VDD.n5698 37.0005
R25812 VDD.n5570 VDD.n5569 37.0005
R25813 VDD.t311 VDD.n5570 37.0005
R25814 VDD.n6320 VDD.n6319 37.0005
R25815 VDD.n6319 VDD.t184 37.0005
R25816 VDD.n5579 VDD.n5578 37.0005
R25817 VDD.n5578 VDD.t184 37.0005
R25818 VDD.n6310 VDD.n6309 37.0005
R25819 VDD.n6309 VDD.t103 37.0005
R25820 VDD.n5589 VDD.n5588 37.0005
R25821 VDD.n5588 VDD.t103 37.0005
R25822 VDD.n6300 VDD.n6299 37.0005
R25823 VDD.n6299 VDD.t855 37.0005
R25824 VDD.n5600 VDD.n5599 37.0005
R25825 VDD.n5599 VDD.t855 37.0005
R25826 VDD.n6290 VDD.n6289 37.0005
R25827 VDD.n6289 VDD.t301 37.0005
R25828 VDD.n5613 VDD.n5612 37.0005
R25829 VDD.n5612 VDD.t301 37.0005
R25830 VDD.n5617 VDD.n5615 37.0005
R25831 VDD.n5615 VDD.t1054 37.0005
R25832 VDD.n6281 VDD.n5616 37.0005
R25833 VDD.n5616 VDD.t1054 37.0005
R25834 VDD.n6273 VDD.n6272 37.0005
R25835 VDD.n6272 VDD.t303 37.0005
R25836 VDD.n5628 VDD.n5627 37.0005
R25837 VDD.n5627 VDD.t303 37.0005
R25838 VDD.n6263 VDD.n6262 37.0005
R25839 VDD.n6262 VDD.t548 37.0005
R25840 VDD.n5641 VDD.n5640 37.0005
R25841 VDD.n5640 VDD.t548 37.0005
R25842 VDD.n6253 VDD.n6252 37.0005
R25843 VDD.n6252 VDD.t43 37.0005
R25844 VDD.n5651 VDD.n5650 37.0005
R25845 VDD.n5650 VDD.t43 37.0005
R25846 VDD.n6243 VDD.n6242 37.0005
R25847 VDD.n6242 VDD.t1028 37.0005
R25848 VDD.n5662 VDD.n5661 37.0005
R25849 VDD.n5661 VDD.t1028 37.0005
R25850 VDD.n6233 VDD.n6232 37.0005
R25851 VDD.n6232 VDD.t377 37.0005
R25852 VDD.n5675 VDD.n5674 37.0005
R25853 VDD.n5674 VDD.t377 37.0005
R25854 VDD.n6223 VDD.n6222 37.0005
R25855 VDD.n6222 VDD.t53 37.0005
R25856 VDD.n5685 VDD.n5684 37.0005
R25857 VDD.n5684 VDD.t53 37.0005
R25858 VDD.n5574 VDD.n5572 37.0005
R25859 VDD.n5572 VDD.t184 37.0005
R25860 VDD.n6320 VDD.n5573 37.0005
R25861 VDD.n5573 VDD.t184 37.0005
R25862 VDD.n5584 VDD.n5582 37.0005
R25863 VDD.n5582 VDD.t103 37.0005
R25864 VDD.n6310 VDD.n5583 37.0005
R25865 VDD.n5583 VDD.t103 37.0005
R25866 VDD.n5594 VDD.n5592 37.0005
R25867 VDD.n5592 VDD.t855 37.0005
R25868 VDD.n6300 VDD.n5593 37.0005
R25869 VDD.n5593 VDD.t855 37.0005
R25870 VDD.n5605 VDD.n5603 37.0005
R25871 VDD.n5603 VDD.t301 37.0005
R25872 VDD.n6290 VDD.n5604 37.0005
R25873 VDD.n5604 VDD.t301 37.0005
R25874 VDD.n5621 VDD.n5619 37.0005
R25875 VDD.n5619 VDD.t303 37.0005
R25876 VDD.n6273 VDD.n5620 37.0005
R25877 VDD.n5620 VDD.t303 37.0005
R25878 VDD.n5633 VDD.n5631 37.0005
R25879 VDD.n5631 VDD.t548 37.0005
R25880 VDD.n6263 VDD.n5632 37.0005
R25881 VDD.n5632 VDD.t548 37.0005
R25882 VDD.n5646 VDD.n5644 37.0005
R25883 VDD.n5644 VDD.t43 37.0005
R25884 VDD.n6253 VDD.n5645 37.0005
R25885 VDD.n5645 VDD.t43 37.0005
R25886 VDD.n5656 VDD.n5654 37.0005
R25887 VDD.n5654 VDD.t1028 37.0005
R25888 VDD.n6243 VDD.n5655 37.0005
R25889 VDD.n5655 VDD.t1028 37.0005
R25890 VDD.n5667 VDD.n5665 37.0005
R25891 VDD.n5665 VDD.t377 37.0005
R25892 VDD.n6233 VDD.n5666 37.0005
R25893 VDD.n5666 VDD.t377 37.0005
R25894 VDD.n5680 VDD.n5678 37.0005
R25895 VDD.n5678 VDD.t53 37.0005
R25896 VDD.n6223 VDD.n5679 37.0005
R25897 VDD.n5679 VDD.t53 37.0005
R25898 VDD.n5689 VDD.n5687 37.0005
R25899 VDD.n5687 VDD.t209 37.0005
R25900 VDD.n6214 VDD.n5688 37.0005
R25901 VDD.n6331 VDD.n6330 37.0005
R25902 VDD.t311 VDD.n6331 37.0005
R25903 VDD.n6333 VDD.n6332 37.0005
R25904 VDD.n6332 VDD.t311 37.0005
R25905 VDD.n6333 VDD.n5562 37.0005
R25906 VDD.t311 VDD.n5562 37.0005
R25907 VDD.n5434 VDD.n5433 37.0005
R25908 VDD.t658 VDD.n5434 37.0005
R25909 VDD.n6443 VDD.n6442 37.0005
R25910 VDD.n6442 VDD.t199 37.0005
R25911 VDD.n5443 VDD.n5442 37.0005
R25912 VDD.n5442 VDD.t199 37.0005
R25913 VDD.n6433 VDD.n6432 37.0005
R25914 VDD.n6432 VDD.t49 37.0005
R25915 VDD.n5453 VDD.n5452 37.0005
R25916 VDD.n5452 VDD.t49 37.0005
R25917 VDD.n6423 VDD.n6422 37.0005
R25918 VDD.n6422 VDD.t428 37.0005
R25919 VDD.n5464 VDD.n5463 37.0005
R25920 VDD.n5463 VDD.t428 37.0005
R25921 VDD.n6413 VDD.n6412 37.0005
R25922 VDD.n6412 VDD.t170 37.0005
R25923 VDD.n5477 VDD.n5476 37.0005
R25924 VDD.n5476 VDD.t170 37.0005
R25925 VDD.n5481 VDD.n5479 37.0005
R25926 VDD.n5479 VDD.t1089 37.0005
R25927 VDD.n6404 VDD.n5480 37.0005
R25928 VDD.n5480 VDD.t1089 37.0005
R25929 VDD.n6396 VDD.n6395 37.0005
R25930 VDD.n6395 VDD.t280 37.0005
R25931 VDD.n5492 VDD.n5491 37.0005
R25932 VDD.n5491 VDD.t280 37.0005
R25933 VDD.n6386 VDD.n6385 37.0005
R25934 VDD.n6385 VDD.t365 37.0005
R25935 VDD.n5505 VDD.n5504 37.0005
R25936 VDD.n5504 VDD.t365 37.0005
R25937 VDD.n6376 VDD.n6375 37.0005
R25938 VDD.n6375 VDD.t81 37.0005
R25939 VDD.n5515 VDD.n5514 37.0005
R25940 VDD.n5514 VDD.t81 37.0005
R25941 VDD.n6366 VDD.n6365 37.0005
R25942 VDD.n6365 VDD.t1002 37.0005
R25943 VDD.n5526 VDD.n5525 37.0005
R25944 VDD.n5525 VDD.t1002 37.0005
R25945 VDD.n6356 VDD.n6355 37.0005
R25946 VDD.n6355 VDD.t254 37.0005
R25947 VDD.n5539 VDD.n5538 37.0005
R25948 VDD.n5538 VDD.t254 37.0005
R25949 VDD.n6346 VDD.n6345 37.0005
R25950 VDD.n6345 VDD.t33 37.0005
R25951 VDD.n5549 VDD.n5548 37.0005
R25952 VDD.n5548 VDD.t33 37.0005
R25953 VDD.n5438 VDD.n5436 37.0005
R25954 VDD.n5436 VDD.t199 37.0005
R25955 VDD.n6443 VDD.n5437 37.0005
R25956 VDD.n5437 VDD.t199 37.0005
R25957 VDD.n5448 VDD.n5446 37.0005
R25958 VDD.n5446 VDD.t49 37.0005
R25959 VDD.n6433 VDD.n5447 37.0005
R25960 VDD.n5447 VDD.t49 37.0005
R25961 VDD.n5458 VDD.n5456 37.0005
R25962 VDD.n5456 VDD.t428 37.0005
R25963 VDD.n6423 VDD.n5457 37.0005
R25964 VDD.n5457 VDD.t428 37.0005
R25965 VDD.n5469 VDD.n5467 37.0005
R25966 VDD.n5467 VDD.t170 37.0005
R25967 VDD.n6413 VDD.n5468 37.0005
R25968 VDD.n5468 VDD.t170 37.0005
R25969 VDD.n5485 VDD.n5483 37.0005
R25970 VDD.n5483 VDD.t280 37.0005
R25971 VDD.n6396 VDD.n5484 37.0005
R25972 VDD.n5484 VDD.t280 37.0005
R25973 VDD.n5497 VDD.n5495 37.0005
R25974 VDD.n5495 VDD.t365 37.0005
R25975 VDD.n6386 VDD.n5496 37.0005
R25976 VDD.n5496 VDD.t365 37.0005
R25977 VDD.n5510 VDD.n5508 37.0005
R25978 VDD.n5508 VDD.t81 37.0005
R25979 VDD.n6376 VDD.n5509 37.0005
R25980 VDD.n5509 VDD.t81 37.0005
R25981 VDD.n5520 VDD.n5518 37.0005
R25982 VDD.n5518 VDD.t1002 37.0005
R25983 VDD.n6366 VDD.n5519 37.0005
R25984 VDD.n5519 VDD.t1002 37.0005
R25985 VDD.n5531 VDD.n5529 37.0005
R25986 VDD.n5529 VDD.t254 37.0005
R25987 VDD.n6356 VDD.n5530 37.0005
R25988 VDD.n5530 VDD.t254 37.0005
R25989 VDD.n5544 VDD.n5542 37.0005
R25990 VDD.n5542 VDD.t33 37.0005
R25991 VDD.n6346 VDD.n5543 37.0005
R25992 VDD.n5543 VDD.t33 37.0005
R25993 VDD.n5553 VDD.n5551 37.0005
R25994 VDD.n5551 VDD.t829 37.0005
R25995 VDD.n6337 VDD.n5552 37.0005
R25996 VDD.n6454 VDD.n6453 37.0005
R25997 VDD.t658 VDD.n6454 37.0005
R25998 VDD.n6456 VDD.n6455 37.0005
R25999 VDD.n6455 VDD.t658 37.0005
R26000 VDD.n6456 VDD.n5426 37.0005
R26001 VDD.t658 VDD.n5426 37.0005
R26002 VDD.n5298 VDD.n5297 37.0005
R26003 VDD.t151 VDD.n5298 37.0005
R26004 VDD.n6566 VDD.n6565 37.0005
R26005 VDD.n6565 VDD.t447 37.0005
R26006 VDD.n5307 VDD.n5306 37.0005
R26007 VDD.n5306 VDD.t447 37.0005
R26008 VDD.n6556 VDD.n6555 37.0005
R26009 VDD.n6555 VDD.t83 37.0005
R26010 VDD.n5317 VDD.n5316 37.0005
R26011 VDD.n5316 VDD.t83 37.0005
R26012 VDD.n6546 VDD.n6545 37.0005
R26013 VDD.n6545 VDD.t363 37.0005
R26014 VDD.n5328 VDD.n5327 37.0005
R26015 VDD.n5327 VDD.t363 37.0005
R26016 VDD.n6536 VDD.n6535 37.0005
R26017 VDD.n6535 VDD.t15 37.0005
R26018 VDD.n5341 VDD.n5340 37.0005
R26019 VDD.n5340 VDD.t15 37.0005
R26020 VDD.n5345 VDD.n5343 37.0005
R26021 VDD.n5343 VDD.t1084 37.0005
R26022 VDD.n6527 VDD.n5344 37.0005
R26023 VDD.n5344 VDD.t1084 37.0005
R26024 VDD.n6519 VDD.n6518 37.0005
R26025 VDD.n6518 VDD.t21 37.0005
R26026 VDD.n5356 VDD.n5355 37.0005
R26027 VDD.n5355 VDD.t21 37.0005
R26028 VDD.n6509 VDD.n6508 37.0005
R26029 VDD.n6508 VDD.t615 37.0005
R26030 VDD.n5369 VDD.n5368 37.0005
R26031 VDD.n5368 VDD.t615 37.0005
R26032 VDD.n6499 VDD.n6498 37.0005
R26033 VDD.n6498 VDD.t65 37.0005
R26034 VDD.n5379 VDD.n5378 37.0005
R26035 VDD.n5378 VDD.t65 37.0005
R26036 VDD.n6489 VDD.n6488 37.0005
R26037 VDD.n6488 VDD.t1060 37.0005
R26038 VDD.n5390 VDD.n5389 37.0005
R26039 VDD.n5389 VDD.t1060 37.0005
R26040 VDD.n6479 VDD.n6478 37.0005
R26041 VDD.n6478 VDD.t172 37.0005
R26042 VDD.n5403 VDD.n5402 37.0005
R26043 VDD.n5402 VDD.t172 37.0005
R26044 VDD.n6469 VDD.n6468 37.0005
R26045 VDD.n6468 VDD.t69 37.0005
R26046 VDD.n5413 VDD.n5412 37.0005
R26047 VDD.n5412 VDD.t69 37.0005
R26048 VDD.n5302 VDD.n5300 37.0005
R26049 VDD.n5300 VDD.t447 37.0005
R26050 VDD.n6566 VDD.n5301 37.0005
R26051 VDD.n5301 VDD.t447 37.0005
R26052 VDD.n5312 VDD.n5310 37.0005
R26053 VDD.n5310 VDD.t83 37.0005
R26054 VDD.n6556 VDD.n5311 37.0005
R26055 VDD.n5311 VDD.t83 37.0005
R26056 VDD.n5322 VDD.n5320 37.0005
R26057 VDD.n5320 VDD.t363 37.0005
R26058 VDD.n6546 VDD.n5321 37.0005
R26059 VDD.n5321 VDD.t363 37.0005
R26060 VDD.n5333 VDD.n5331 37.0005
R26061 VDD.n5331 VDD.t15 37.0005
R26062 VDD.n6536 VDD.n5332 37.0005
R26063 VDD.n5332 VDD.t15 37.0005
R26064 VDD.n5349 VDD.n5347 37.0005
R26065 VDD.n5347 VDD.t21 37.0005
R26066 VDD.n6519 VDD.n5348 37.0005
R26067 VDD.n5348 VDD.t21 37.0005
R26068 VDD.n5361 VDD.n5359 37.0005
R26069 VDD.n5359 VDD.t615 37.0005
R26070 VDD.n6509 VDD.n5360 37.0005
R26071 VDD.n5360 VDD.t615 37.0005
R26072 VDD.n5374 VDD.n5372 37.0005
R26073 VDD.n5372 VDD.t65 37.0005
R26074 VDD.n6499 VDD.n5373 37.0005
R26075 VDD.n5373 VDD.t65 37.0005
R26076 VDD.n5384 VDD.n5382 37.0005
R26077 VDD.n5382 VDD.t1060 37.0005
R26078 VDD.n6489 VDD.n5383 37.0005
R26079 VDD.n5383 VDD.t1060 37.0005
R26080 VDD.n5395 VDD.n5393 37.0005
R26081 VDD.n5393 VDD.t172 37.0005
R26082 VDD.n6479 VDD.n5394 37.0005
R26083 VDD.n5394 VDD.t172 37.0005
R26084 VDD.n5408 VDD.n5406 37.0005
R26085 VDD.n5406 VDD.t69 37.0005
R26086 VDD.n6469 VDD.n5407 37.0005
R26087 VDD.n5407 VDD.t69 37.0005
R26088 VDD.n5417 VDD.n5415 37.0005
R26089 VDD.n5415 VDD.t837 37.0005
R26090 VDD.n6460 VDD.n5416 37.0005
R26091 VDD.n6577 VDD.n6576 37.0005
R26092 VDD.t151 VDD.n6577 37.0005
R26093 VDD.n6579 VDD.n6578 37.0005
R26094 VDD.n6578 VDD.t151 37.0005
R26095 VDD.n6579 VDD.n5290 37.0005
R26096 VDD.t151 VDD.n5290 37.0005
R26097 VDD.n5162 VDD.n5161 37.0005
R26098 VDD.t862 VDD.n5162 37.0005
R26099 VDD.n6689 VDD.n6688 37.0005
R26100 VDD.n6688 VDD.t285 37.0005
R26101 VDD.n5171 VDD.n5170 37.0005
R26102 VDD.n5170 VDD.t285 37.0005
R26103 VDD.n6679 VDD.n6678 37.0005
R26104 VDD.n6678 VDD.t73 37.0005
R26105 VDD.n5181 VDD.n5180 37.0005
R26106 VDD.n5180 VDD.t73 37.0005
R26107 VDD.n6669 VDD.n6668 37.0005
R26108 VDD.n6668 VDD.t341 37.0005
R26109 VDD.n5192 VDD.n5191 37.0005
R26110 VDD.n5191 VDD.t341 37.0005
R26111 VDD.n6659 VDD.n6658 37.0005
R26112 VDD.n6658 VDD.t665 37.0005
R26113 VDD.n5205 VDD.n5204 37.0005
R26114 VDD.n5204 VDD.t665 37.0005
R26115 VDD.n5209 VDD.n5207 37.0005
R26116 VDD.n5207 VDD.t1058 37.0005
R26117 VDD.n6650 VDD.n5208 37.0005
R26118 VDD.n5208 VDD.t1058 37.0005
R26119 VDD.n6642 VDD.n6641 37.0005
R26120 VDD.n6641 VDD.t643 37.0005
R26121 VDD.n5220 VDD.n5219 37.0005
R26122 VDD.n5219 VDD.t643 37.0005
R26123 VDD.n6632 VDD.n6631 37.0005
R26124 VDD.n6631 VDD.t486 37.0005
R26125 VDD.n5233 VDD.n5232 37.0005
R26126 VDD.n5232 VDD.t486 37.0005
R26127 VDD.n6622 VDD.n6621 37.0005
R26128 VDD.n6621 VDD.t111 37.0005
R26129 VDD.n5243 VDD.n5242 37.0005
R26130 VDD.n5242 VDD.t111 37.0005
R26131 VDD.n6612 VDD.n6611 37.0005
R26132 VDD.n6611 VDD.t1032 37.0005
R26133 VDD.n5254 VDD.n5253 37.0005
R26134 VDD.n5253 VDD.t1032 37.0005
R26135 VDD.n6602 VDD.n6601 37.0005
R26136 VDD.n6601 VDD.t398 37.0005
R26137 VDD.n5267 VDD.n5266 37.0005
R26138 VDD.n5266 VDD.t398 37.0005
R26139 VDD.n6592 VDD.n6591 37.0005
R26140 VDD.n6591 VDD.t55 37.0005
R26141 VDD.n5277 VDD.n5276 37.0005
R26142 VDD.n5276 VDD.t55 37.0005
R26143 VDD.n5166 VDD.n5164 37.0005
R26144 VDD.n5164 VDD.t285 37.0005
R26145 VDD.n6689 VDD.n5165 37.0005
R26146 VDD.n5165 VDD.t285 37.0005
R26147 VDD.n5176 VDD.n5174 37.0005
R26148 VDD.n5174 VDD.t73 37.0005
R26149 VDD.n6679 VDD.n5175 37.0005
R26150 VDD.n5175 VDD.t73 37.0005
R26151 VDD.n5186 VDD.n5184 37.0005
R26152 VDD.n5184 VDD.t341 37.0005
R26153 VDD.n6669 VDD.n5185 37.0005
R26154 VDD.n5185 VDD.t341 37.0005
R26155 VDD.n5197 VDD.n5195 37.0005
R26156 VDD.n5195 VDD.t665 37.0005
R26157 VDD.n6659 VDD.n5196 37.0005
R26158 VDD.n5196 VDD.t665 37.0005
R26159 VDD.n5213 VDD.n5211 37.0005
R26160 VDD.n5211 VDD.t643 37.0005
R26161 VDD.n6642 VDD.n5212 37.0005
R26162 VDD.n5212 VDD.t643 37.0005
R26163 VDD.n5225 VDD.n5223 37.0005
R26164 VDD.n5223 VDD.t486 37.0005
R26165 VDD.n6632 VDD.n5224 37.0005
R26166 VDD.n5224 VDD.t486 37.0005
R26167 VDD.n5238 VDD.n5236 37.0005
R26168 VDD.n5236 VDD.t111 37.0005
R26169 VDD.n6622 VDD.n5237 37.0005
R26170 VDD.n5237 VDD.t111 37.0005
R26171 VDD.n5248 VDD.n5246 37.0005
R26172 VDD.n5246 VDD.t1032 37.0005
R26173 VDD.n6612 VDD.n5247 37.0005
R26174 VDD.n5247 VDD.t1032 37.0005
R26175 VDD.n5259 VDD.n5257 37.0005
R26176 VDD.n5257 VDD.t398 37.0005
R26177 VDD.n6602 VDD.n5258 37.0005
R26178 VDD.n5258 VDD.t398 37.0005
R26179 VDD.n5272 VDD.n5270 37.0005
R26180 VDD.n5270 VDD.t55 37.0005
R26181 VDD.n6592 VDD.n5271 37.0005
R26182 VDD.n5271 VDD.t55 37.0005
R26183 VDD.n5281 VDD.n5279 37.0005
R26184 VDD.n5279 VDD.t155 37.0005
R26185 VDD.n6583 VDD.n5280 37.0005
R26186 VDD.n6700 VDD.n6699 37.0005
R26187 VDD.t862 VDD.n6700 37.0005
R26188 VDD.n6702 VDD.n6701 37.0005
R26189 VDD.n6701 VDD.t862 37.0005
R26190 VDD.n6702 VDD.n5154 37.0005
R26191 VDD.t862 VDD.n5154 37.0005
R26192 VDD.n5026 VDD.n5025 37.0005
R26193 VDD.t937 VDD.n5026 37.0005
R26194 VDD.n6812 VDD.n6811 37.0005
R26195 VDD.n6811 VDD.t144 37.0005
R26196 VDD.n5035 VDD.n5034 37.0005
R26197 VDD.n5034 VDD.t144 37.0005
R26198 VDD.n6802 VDD.n6801 37.0005
R26199 VDD.n6801 VDD.t23 37.0005
R26200 VDD.n5045 VDD.n5044 37.0005
R26201 VDD.n5044 VDD.t23 37.0005
R26202 VDD.n6792 VDD.n6791 37.0005
R26203 VDD.n6791 VDD.t507 37.0005
R26204 VDD.n5056 VDD.n5055 37.0005
R26205 VDD.n5055 VDD.t507 37.0005
R26206 VDD.n6782 VDD.n6781 37.0005
R26207 VDD.n6781 VDD.t9 37.0005
R26208 VDD.n5069 VDD.n5068 37.0005
R26209 VDD.n5068 VDD.t9 37.0005
R26210 VDD.n5073 VDD.n5071 37.0005
R26211 VDD.n5071 VDD.t1076 37.0005
R26212 VDD.n6773 VDD.n5072 37.0005
R26213 VDD.n5072 VDD.t1076 37.0005
R26214 VDD.n6765 VDD.n6764 37.0005
R26215 VDD.n6764 VDD.t11 37.0005
R26216 VDD.n5084 VDD.n5083 37.0005
R26217 VDD.n5083 VDD.t11 37.0005
R26218 VDD.n6755 VDD.n6754 37.0005
R26219 VDD.n6754 VDD.t561 37.0005
R26220 VDD.n5097 VDD.n5096 37.0005
R26221 VDD.n5096 VDD.t561 37.0005
R26222 VDD.n6745 VDD.n6744 37.0005
R26223 VDD.n6744 VDD.t99 37.0005
R26224 VDD.n5107 VDD.n5106 37.0005
R26225 VDD.n5106 VDD.t99 37.0005
R26226 VDD.n6735 VDD.n6734 37.0005
R26227 VDD.n6734 VDD.t1030 37.0005
R26228 VDD.n5118 VDD.n5117 37.0005
R26229 VDD.n5117 VDD.t1030 37.0005
R26230 VDD.n6725 VDD.n6724 37.0005
R26231 VDD.n6724 VDD.t598 37.0005
R26232 VDD.n5131 VDD.n5130 37.0005
R26233 VDD.n5130 VDD.t598 37.0005
R26234 VDD.n6715 VDD.n6714 37.0005
R26235 VDD.n6714 VDD.t47 37.0005
R26236 VDD.n5141 VDD.n5140 37.0005
R26237 VDD.n5140 VDD.t47 37.0005
R26238 VDD.n5030 VDD.n5028 37.0005
R26239 VDD.n5028 VDD.t144 37.0005
R26240 VDD.n6812 VDD.n5029 37.0005
R26241 VDD.n5029 VDD.t144 37.0005
R26242 VDD.n5040 VDD.n5038 37.0005
R26243 VDD.n5038 VDD.t23 37.0005
R26244 VDD.n6802 VDD.n5039 37.0005
R26245 VDD.n5039 VDD.t23 37.0005
R26246 VDD.n5050 VDD.n5048 37.0005
R26247 VDD.n5048 VDD.t507 37.0005
R26248 VDD.n6792 VDD.n5049 37.0005
R26249 VDD.n5049 VDD.t507 37.0005
R26250 VDD.n5061 VDD.n5059 37.0005
R26251 VDD.n5059 VDD.t9 37.0005
R26252 VDD.n6782 VDD.n5060 37.0005
R26253 VDD.n5060 VDD.t9 37.0005
R26254 VDD.n5077 VDD.n5075 37.0005
R26255 VDD.n5075 VDD.t11 37.0005
R26256 VDD.n6765 VDD.n5076 37.0005
R26257 VDD.n5076 VDD.t11 37.0005
R26258 VDD.n5089 VDD.n5087 37.0005
R26259 VDD.n5087 VDD.t561 37.0005
R26260 VDD.n6755 VDD.n5088 37.0005
R26261 VDD.n5088 VDD.t561 37.0005
R26262 VDD.n5102 VDD.n5100 37.0005
R26263 VDD.n5100 VDD.t99 37.0005
R26264 VDD.n6745 VDD.n5101 37.0005
R26265 VDD.n5101 VDD.t99 37.0005
R26266 VDD.n5112 VDD.n5110 37.0005
R26267 VDD.n5110 VDD.t1030 37.0005
R26268 VDD.n6735 VDD.n5111 37.0005
R26269 VDD.n5111 VDD.t1030 37.0005
R26270 VDD.n5123 VDD.n5121 37.0005
R26271 VDD.n5121 VDD.t598 37.0005
R26272 VDD.n6725 VDD.n5122 37.0005
R26273 VDD.n5122 VDD.t598 37.0005
R26274 VDD.n5136 VDD.n5134 37.0005
R26275 VDD.n5134 VDD.t47 37.0005
R26276 VDD.n6715 VDD.n5135 37.0005
R26277 VDD.n5135 VDD.t47 37.0005
R26278 VDD.n5145 VDD.n5143 37.0005
R26279 VDD.n5143 VDD.t566 37.0005
R26280 VDD.n6706 VDD.n5144 37.0005
R26281 VDD.n6823 VDD.n6822 37.0005
R26282 VDD.t937 VDD.n6823 37.0005
R26283 VDD.n6825 VDD.n6824 37.0005
R26284 VDD.n6824 VDD.t937 37.0005
R26285 VDD.n6825 VDD.n5018 37.0005
R26286 VDD.t937 VDD.n5018 37.0005
R26287 VDD.n4884 VDD.n4883 37.0005
R26288 VDD.n4883 VDD.t492 37.0005
R26289 VDD.n4904 VDD.n4903 37.0005
R26290 VDD.n4903 VDD.t248 37.0005
R26291 VDD.n4875 VDD.n4874 37.0005
R26292 VDD.n4874 VDD.t248 37.0005
R26293 VDD.n4914 VDD.n4913 37.0005
R26294 VDD.n4913 VDD.t101 37.0005
R26295 VDD.n4865 VDD.n4864 37.0005
R26296 VDD.n4864 VDD.t101 37.0005
R26297 VDD.n4924 VDD.n4923 37.0005
R26298 VDD.n4923 VDD.t655 37.0005
R26299 VDD.n4854 VDD.n4853 37.0005
R26300 VDD.n4853 VDD.t655 37.0005
R26301 VDD.n4934 VDD.n4933 37.0005
R26302 VDD.n4933 VDD.t242 37.0005
R26303 VDD.n4841 VDD.n4840 37.0005
R26304 VDD.n4840 VDD.t242 37.0005
R26305 VDD.n4830 VDD.n4828 37.0005
R26306 VDD.n4828 VDD.t1052 37.0005
R26307 VDD.n4942 VDD.n4829 37.0005
R26308 VDD.n4829 VDD.t1052 37.0005
R26309 VDD.n4951 VDD.n4950 37.0005
R26310 VDD.n4950 VDD.t244 37.0005
R26311 VDD.n4826 VDD.n4825 37.0005
R26312 VDD.n4825 VDD.t244 37.0005
R26313 VDD.n4961 VDD.n4960 37.0005
R26314 VDD.n4960 VDD.t445 37.0005
R26315 VDD.n4813 VDD.n4812 37.0005
R26316 VDD.n4812 VDD.t445 37.0005
R26317 VDD.n4971 VDD.n4970 37.0005
R26318 VDD.n4970 VDD.t77 37.0005
R26319 VDD.n4803 VDD.n4802 37.0005
R26320 VDD.n4802 VDD.t77 37.0005
R26321 VDD.n4981 VDD.n4980 37.0005
R26322 VDD.n4980 VDD.t1004 37.0005
R26323 VDD.n4792 VDD.n4791 37.0005
R26324 VDD.n4791 VDD.t1004 37.0005
R26325 VDD.n4991 VDD.n4990 37.0005
R26326 VDD.n4990 VDD.t205 37.0005
R26327 VDD.n4779 VDD.n4778 37.0005
R26328 VDD.n4778 VDD.t205 37.0005
R26329 VDD.n5001 VDD.n5000 37.0005
R26330 VDD.n5000 VDD.t87 37.0005
R26331 VDD.n4769 VDD.n4768 37.0005
R26332 VDD.n4768 VDD.t87 37.0005
R26333 VDD.n4870 VDD.n4868 37.0005
R26334 VDD.n4868 VDD.t248 37.0005
R26335 VDD.n4904 VDD.n4869 37.0005
R26336 VDD.n4869 VDD.t248 37.0005
R26337 VDD.n4859 VDD.n4857 37.0005
R26338 VDD.n4857 VDD.t101 37.0005
R26339 VDD.n4914 VDD.n4858 37.0005
R26340 VDD.n4858 VDD.t101 37.0005
R26341 VDD.n4846 VDD.n4844 37.0005
R26342 VDD.n4844 VDD.t655 37.0005
R26343 VDD.n4924 VDD.n4845 37.0005
R26344 VDD.n4845 VDD.t655 37.0005
R26345 VDD.n4834 VDD.n4832 37.0005
R26346 VDD.n4832 VDD.t242 37.0005
R26347 VDD.n4934 VDD.n4833 37.0005
R26348 VDD.n4833 VDD.t242 37.0005
R26349 VDD.n4818 VDD.n4816 37.0005
R26350 VDD.n4816 VDD.t244 37.0005
R26351 VDD.n4951 VDD.n4817 37.0005
R26352 VDD.n4817 VDD.t244 37.0005
R26353 VDD.n4808 VDD.n4806 37.0005
R26354 VDD.n4806 VDD.t445 37.0005
R26355 VDD.n4961 VDD.n4807 37.0005
R26356 VDD.n4807 VDD.t445 37.0005
R26357 VDD.n4797 VDD.n4795 37.0005
R26358 VDD.n4795 VDD.t77 37.0005
R26359 VDD.n4971 VDD.n4796 37.0005
R26360 VDD.n4796 VDD.t77 37.0005
R26361 VDD.n4784 VDD.n4782 37.0005
R26362 VDD.n4782 VDD.t1004 37.0005
R26363 VDD.n4981 VDD.n4783 37.0005
R26364 VDD.n4783 VDD.t1004 37.0005
R26365 VDD.n4774 VDD.n4772 37.0005
R26366 VDD.n4772 VDD.t205 37.0005
R26367 VDD.n4991 VDD.n4773 37.0005
R26368 VDD.n4773 VDD.t205 37.0005
R26369 VDD.n4763 VDD.n4761 37.0005
R26370 VDD.n4761 VDD.t87 37.0005
R26371 VDD.n5001 VDD.n4762 37.0005
R26372 VDD.n4762 VDD.t87 37.0005
R26373 VDD.n4759 VDD.n4758 37.0005
R26374 VDD.t203 VDD.n4759 37.0005
R26375 VDD.n5011 VDD.n4757 37.0005
R26376 VDD.n4880 VDD.n4878 37.0005
R26377 VDD.n4878 VDD.t492 37.0005
R26378 VDD.n4894 VDD.n4890 37.0005
R26379 VDD.n4890 VDD.t492 37.0005
R26380 VDD.n4894 VDD.n4879 37.0005
R26381 VDD.n4879 VDD.t492 37.0005
R26382 VDD.n4745 VDD.n4744 37.0005
R26383 VDD.n4744 VDD.t51 37.0005
R26384 VDD.n1993 VDD.n1992 37.0005
R26385 VDD.n1992 VDD.t51 37.0005
R26386 VDD.n4735 VDD.n4734 37.0005
R26387 VDD.n4734 VDD.t646 37.0005
R26388 VDD.n2003 VDD.n2002 37.0005
R26389 VDD.n2002 VDD.t646 37.0005
R26390 VDD.n4725 VDD.n4724 37.0005
R26391 VDD.n4724 VDD.t1016 37.0005
R26392 VDD.n2016 VDD.n2015 37.0005
R26393 VDD.n2015 VDD.t1016 37.0005
R26394 VDD.n4715 VDD.n4714 37.0005
R26395 VDD.n4714 VDD.t117 37.0005
R26396 VDD.n2028 VDD.n2027 37.0005
R26397 VDD.n2027 VDD.t117 37.0005
R26398 VDD.n2046 VDD.n2045 37.0005
R26399 VDD.n2045 VDD.t256 37.0005
R26400 VDD.n4701 VDD.n4700 37.0005
R26401 VDD.n4700 VDD.t17 37.0005
R26402 VDD.n2056 VDD.n2055 37.0005
R26403 VDD.t17 VDD.n2056 37.0005
R26404 VDD.n2059 VDD.n2057 37.0005
R26405 VDD.n2057 VDD.t1068 37.0005
R26406 VDD.n4689 VDD.n2058 37.0005
R26407 VDD.n2058 VDD.t1068 37.0005
R26408 VDD.n4681 VDD.n4680 37.0005
R26409 VDD.n4680 VDD.t19 37.0005
R26410 VDD.n2070 VDD.n2069 37.0005
R26411 VDD.n2069 VDD.t19 37.0005
R26412 VDD.n4671 VDD.n4670 37.0005
R26413 VDD.n4670 VDD.t607 37.0005
R26414 VDD.n2083 VDD.n2082 37.0005
R26415 VDD.n2082 VDD.t607 37.0005
R26416 VDD.n4661 VDD.n4660 37.0005
R26417 VDD.n4660 VDD.t57 37.0005
R26418 VDD.n2094 VDD.n2093 37.0005
R26419 VDD.n2093 VDD.t57 37.0005
R26420 VDD.n4651 VDD.n4650 37.0005
R26421 VDD.n4650 VDD.t232 37.0005
R26422 VDD.n2104 VDD.n2103 37.0005
R26423 VDD.n2103 VDD.t232 37.0005
R26424 VDD.n4641 VDD.n4640 37.0005
R26425 VDD.n4640 VDD.t602 37.0005
R26426 VDD.n4634 VDD.n4633 37.0005
R26427 VDD.n4633 VDD.t602 37.0005
R26428 VDD.n1981 VDD.n1980 37.0005
R26429 VDD.t2 VDD.n1981 37.0005
R26430 VDD.n4753 VDD.n1979 37.0005
R26431 VDD.n1987 VDD.n1985 37.0005
R26432 VDD.n1985 VDD.t51 37.0005
R26433 VDD.n4745 VDD.n1986 37.0005
R26434 VDD.n1986 VDD.t51 37.0005
R26435 VDD.n1998 VDD.n1996 37.0005
R26436 VDD.n1996 VDD.t646 37.0005
R26437 VDD.n4735 VDD.n1997 37.0005
R26438 VDD.n1997 VDD.t646 37.0005
R26439 VDD.n2008 VDD.n2006 37.0005
R26440 VDD.n2006 VDD.t1016 37.0005
R26441 VDD.n4725 VDD.n2007 37.0005
R26442 VDD.n2007 VDD.t1016 37.0005
R26443 VDD.n2021 VDD.n2019 37.0005
R26444 VDD.n2019 VDD.t117 37.0005
R26445 VDD.n4715 VDD.n2020 37.0005
R26446 VDD.n2020 VDD.t117 37.0005
R26447 VDD.n4699 VDD.n4698 37.0005
R26448 VDD.t17 VDD.n4699 37.0005
R26449 VDD.n4701 VDD.n2041 37.0005
R26450 VDD.t17 VDD.n2041 37.0005
R26451 VDD.n2063 VDD.n2061 37.0005
R26452 VDD.n2061 VDD.t19 37.0005
R26453 VDD.n4681 VDD.n2062 37.0005
R26454 VDD.n2062 VDD.t19 37.0005
R26455 VDD.n2075 VDD.n2073 37.0005
R26456 VDD.n2073 VDD.t607 37.0005
R26457 VDD.n4671 VDD.n2074 37.0005
R26458 VDD.n2074 VDD.t607 37.0005
R26459 VDD.n2088 VDD.n2086 37.0005
R26460 VDD.n2086 VDD.t57 37.0005
R26461 VDD.n4661 VDD.n2087 37.0005
R26462 VDD.n2087 VDD.t57 37.0005
R26463 VDD.n2099 VDD.n2097 37.0005
R26464 VDD.n2097 VDD.t232 37.0005
R26465 VDD.n4651 VDD.n2098 37.0005
R26466 VDD.n2098 VDD.t232 37.0005
R26467 VDD.n2109 VDD.n2107 37.0005
R26468 VDD.n2107 VDD.t602 37.0005
R26469 VDD.n4641 VDD.n2108 37.0005
R26470 VDD.n2108 VDD.t602 37.0005
R26471 VDD.n2033 VDD.n2031 37.0005
R26472 VDD.n2031 VDD.t256 37.0005
R26473 VDD.n4705 VDD.n2036 37.0005
R26474 VDD.n2036 VDD.t256 37.0005
R26475 VDD.n4705 VDD.n2032 37.0005
R26476 VDD.n2032 VDD.t256 37.0005
R26477 VDD.n4620 VDD.n4619 37.0005
R26478 VDD.n4619 VDD.t89 37.0005
R26479 VDD.n2129 VDD.n2128 37.0005
R26480 VDD.n2128 VDD.t89 37.0005
R26481 VDD.n4610 VDD.n4609 37.0005
R26482 VDD.n4609 VDD.t186 37.0005
R26483 VDD.n2139 VDD.n2138 37.0005
R26484 VDD.n2138 VDD.t186 37.0005
R26485 VDD.n4600 VDD.n4599 37.0005
R26486 VDD.n4599 VDD.t1042 37.0005
R26487 VDD.n2152 VDD.n2151 37.0005
R26488 VDD.n2151 VDD.t1042 37.0005
R26489 VDD.n4590 VDD.n4589 37.0005
R26490 VDD.n4589 VDD.t39 37.0005
R26491 VDD.n2164 VDD.n2163 37.0005
R26492 VDD.n2163 VDD.t39 37.0005
R26493 VDD.n2182 VDD.n2181 37.0005
R26494 VDD.n2181 VDD.t512 37.0005
R26495 VDD.n4576 VDD.n4575 37.0005
R26496 VDD.n4575 VDD.t221 37.0005
R26497 VDD.n2192 VDD.n2191 37.0005
R26498 VDD.t221 VDD.n2192 37.0005
R26499 VDD.n2195 VDD.n2193 37.0005
R26500 VDD.n2193 VDD.t1082 37.0005
R26501 VDD.n4564 VDD.n2194 37.0005
R26502 VDD.n2194 VDD.t1082 37.0005
R26503 VDD.n4556 VDD.n4555 37.0005
R26504 VDD.n4555 VDD.t223 37.0005
R26505 VDD.n2206 VDD.n2205 37.0005
R26506 VDD.n2205 VDD.t223 37.0005
R26507 VDD.n4546 VDD.n4545 37.0005
R26508 VDD.n4545 VDD.t685 37.0005
R26509 VDD.n2219 VDD.n2218 37.0005
R26510 VDD.n2218 VDD.t685 37.0005
R26511 VDD.n4536 VDD.n4535 37.0005
R26512 VDD.n4535 VDD.t63 37.0005
R26513 VDD.n2230 VDD.n2229 37.0005
R26514 VDD.n2229 VDD.t63 37.0005
R26515 VDD.n4526 VDD.n4525 37.0005
R26516 VDD.n4525 VDD.t460 37.0005
R26517 VDD.n2240 VDD.n2239 37.0005
R26518 VDD.n2239 VDD.t460 37.0005
R26519 VDD.n4516 VDD.n4515 37.0005
R26520 VDD.n4515 VDD.t578 37.0005
R26521 VDD.n4509 VDD.n4508 37.0005
R26522 VDD.n4508 VDD.t578 37.0005
R26523 VDD.n2117 VDD.n2116 37.0005
R26524 VDD.t920 VDD.n2117 37.0005
R26525 VDD.n4628 VDD.n2115 37.0005
R26526 VDD.n2123 VDD.n2121 37.0005
R26527 VDD.n2121 VDD.t89 37.0005
R26528 VDD.n4620 VDD.n2122 37.0005
R26529 VDD.n2122 VDD.t89 37.0005
R26530 VDD.n2134 VDD.n2132 37.0005
R26531 VDD.n2132 VDD.t186 37.0005
R26532 VDD.n4610 VDD.n2133 37.0005
R26533 VDD.n2133 VDD.t186 37.0005
R26534 VDD.n2144 VDD.n2142 37.0005
R26535 VDD.n2142 VDD.t1042 37.0005
R26536 VDD.n4600 VDD.n2143 37.0005
R26537 VDD.n2143 VDD.t1042 37.0005
R26538 VDD.n2157 VDD.n2155 37.0005
R26539 VDD.n2155 VDD.t39 37.0005
R26540 VDD.n4590 VDD.n2156 37.0005
R26541 VDD.n2156 VDD.t39 37.0005
R26542 VDD.n4574 VDD.n4573 37.0005
R26543 VDD.t221 VDD.n4574 37.0005
R26544 VDD.n4576 VDD.n2177 37.0005
R26545 VDD.t221 VDD.n2177 37.0005
R26546 VDD.n2199 VDD.n2197 37.0005
R26547 VDD.n2197 VDD.t223 37.0005
R26548 VDD.n4556 VDD.n2198 37.0005
R26549 VDD.n2198 VDD.t223 37.0005
R26550 VDD.n2211 VDD.n2209 37.0005
R26551 VDD.n2209 VDD.t685 37.0005
R26552 VDD.n4546 VDD.n2210 37.0005
R26553 VDD.n2210 VDD.t685 37.0005
R26554 VDD.n2224 VDD.n2222 37.0005
R26555 VDD.n2222 VDD.t63 37.0005
R26556 VDD.n4536 VDD.n2223 37.0005
R26557 VDD.n2223 VDD.t63 37.0005
R26558 VDD.n2235 VDD.n2233 37.0005
R26559 VDD.n2233 VDD.t460 37.0005
R26560 VDD.n4526 VDD.n2234 37.0005
R26561 VDD.n2234 VDD.t460 37.0005
R26562 VDD.n2245 VDD.n2243 37.0005
R26563 VDD.n2243 VDD.t578 37.0005
R26564 VDD.n4516 VDD.n2244 37.0005
R26565 VDD.n2244 VDD.t578 37.0005
R26566 VDD.n2169 VDD.n2167 37.0005
R26567 VDD.n2167 VDD.t512 37.0005
R26568 VDD.n4580 VDD.n2172 37.0005
R26569 VDD.n2172 VDD.t512 37.0005
R26570 VDD.n4580 VDD.n2168 37.0005
R26571 VDD.n2168 VDD.t512 37.0005
R26572 VDD.n4495 VDD.n4494 37.0005
R26573 VDD.n4494 VDD.t97 37.0005
R26574 VDD.n2265 VDD.n2264 37.0005
R26575 VDD.n2264 VDD.t97 37.0005
R26576 VDD.n4485 VDD.n4484 37.0005
R26577 VDD.n4484 VDD.t564 37.0005
R26578 VDD.n2275 VDD.n2274 37.0005
R26579 VDD.n2274 VDD.t564 37.0005
R26580 VDD.n4475 VDD.n4474 37.0005
R26581 VDD.n4474 VDD.t1050 37.0005
R26582 VDD.n2288 VDD.n2287 37.0005
R26583 VDD.n2287 VDD.t1050 37.0005
R26584 VDD.n4465 VDD.n4464 37.0005
R26585 VDD.n4464 VDD.t109 37.0005
R26586 VDD.n2300 VDD.n2299 37.0005
R26587 VDD.n2299 VDD.t109 37.0005
R26588 VDD.n2318 VDD.n2317 37.0005
R26589 VDD.n2317 VDD.t451 37.0005
R26590 VDD.n4451 VDD.n4450 37.0005
R26591 VDD.n4450 VDD.t954 37.0005
R26592 VDD.n2328 VDD.n2327 37.0005
R26593 VDD.t954 VDD.n2328 37.0005
R26594 VDD.n2331 VDD.n2329 37.0005
R26595 VDD.n2329 VDD.t1010 37.0005
R26596 VDD.n4439 VDD.n2330 37.0005
R26597 VDD.n2330 VDD.t1010 37.0005
R26598 VDD.n4431 VDD.n4430 37.0005
R26599 VDD.n4430 VDD.t660 37.0005
R26600 VDD.n2342 VDD.n2341 37.0005
R26601 VDD.n2341 VDD.t660 37.0005
R26602 VDD.n4421 VDD.n4420 37.0005
R26603 VDD.n4420 VDD.t337 37.0005
R26604 VDD.n2355 VDD.n2354 37.0005
R26605 VDD.n2354 VDD.t337 37.0005
R26606 VDD.n4411 VDD.n4410 37.0005
R26607 VDD.n4410 VDD.t123 37.0005
R26608 VDD.n2366 VDD.n2365 37.0005
R26609 VDD.n2365 VDD.t123 37.0005
R26610 VDD.n4401 VDD.n4400 37.0005
R26611 VDD.n4400 VDD.t625 37.0005
R26612 VDD.n2376 VDD.n2375 37.0005
R26613 VDD.n2375 VDD.t625 37.0005
R26614 VDD.n4391 VDD.n4390 37.0005
R26615 VDD.n4390 VDD.t453 37.0005
R26616 VDD.n4384 VDD.n4383 37.0005
R26617 VDD.n4383 VDD.t453 37.0005
R26618 VDD.n2253 VDD.n2252 37.0005
R26619 VDD.t291 VDD.n2253 37.0005
R26620 VDD.n4503 VDD.n2251 37.0005
R26621 VDD.n2259 VDD.n2257 37.0005
R26622 VDD.n2257 VDD.t97 37.0005
R26623 VDD.n4495 VDD.n2258 37.0005
R26624 VDD.n2258 VDD.t97 37.0005
R26625 VDD.n2270 VDD.n2268 37.0005
R26626 VDD.n2268 VDD.t564 37.0005
R26627 VDD.n4485 VDD.n2269 37.0005
R26628 VDD.n2269 VDD.t564 37.0005
R26629 VDD.n2280 VDD.n2278 37.0005
R26630 VDD.n2278 VDD.t1050 37.0005
R26631 VDD.n4475 VDD.n2279 37.0005
R26632 VDD.n2279 VDD.t1050 37.0005
R26633 VDD.n2293 VDD.n2291 37.0005
R26634 VDD.n2291 VDD.t109 37.0005
R26635 VDD.n4465 VDD.n2292 37.0005
R26636 VDD.n2292 VDD.t109 37.0005
R26637 VDD.n4449 VDD.n4448 37.0005
R26638 VDD.t954 VDD.n4449 37.0005
R26639 VDD.n4451 VDD.n2313 37.0005
R26640 VDD.t954 VDD.n2313 37.0005
R26641 VDD.n2335 VDD.n2333 37.0005
R26642 VDD.n2333 VDD.t660 37.0005
R26643 VDD.n4431 VDD.n2334 37.0005
R26644 VDD.n2334 VDD.t660 37.0005
R26645 VDD.n2347 VDD.n2345 37.0005
R26646 VDD.n2345 VDD.t337 37.0005
R26647 VDD.n4421 VDD.n2346 37.0005
R26648 VDD.n2346 VDD.t337 37.0005
R26649 VDD.n2360 VDD.n2358 37.0005
R26650 VDD.n2358 VDD.t123 37.0005
R26651 VDD.n4411 VDD.n2359 37.0005
R26652 VDD.n2359 VDD.t123 37.0005
R26653 VDD.n2371 VDD.n2369 37.0005
R26654 VDD.n2369 VDD.t625 37.0005
R26655 VDD.n4401 VDD.n2370 37.0005
R26656 VDD.n2370 VDD.t625 37.0005
R26657 VDD.n2381 VDD.n2379 37.0005
R26658 VDD.n2379 VDD.t453 37.0005
R26659 VDD.n4391 VDD.n2380 37.0005
R26660 VDD.n2380 VDD.t453 37.0005
R26661 VDD.n2305 VDD.n2303 37.0005
R26662 VDD.n2303 VDD.t451 37.0005
R26663 VDD.n4455 VDD.n2308 37.0005
R26664 VDD.n2308 VDD.t451 37.0005
R26665 VDD.n4455 VDD.n2304 37.0005
R26666 VDD.n2304 VDD.t451 37.0005
R26667 VDD.n4370 VDD.n4369 37.0005
R26668 VDD.n4369 VDD.t95 37.0005
R26669 VDD.n2401 VDD.n2400 37.0005
R26670 VDD.n2400 VDD.t95 37.0005
R26671 VDD.n4360 VDD.n4359 37.0005
R26672 VDD.n4359 VDD.t591 37.0005
R26673 VDD.n2411 VDD.n2410 37.0005
R26674 VDD.n2410 VDD.t591 37.0005
R26675 VDD.n4350 VDD.n4349 37.0005
R26676 VDD.n4349 VDD.t1048 37.0005
R26677 VDD.n2424 VDD.n2423 37.0005
R26678 VDD.n2423 VDD.t1048 37.0005
R26679 VDD.n4340 VDD.n4339 37.0005
R26680 VDD.n4339 VDD.t31 37.0005
R26681 VDD.n2436 VDD.n2435 37.0005
R26682 VDD.n2435 VDD.t31 37.0005
R26683 VDD.n2454 VDD.n2453 37.0005
R26684 VDD.n2453 VDD.t426 37.0005
R26685 VDD.n4326 VDD.n4325 37.0005
R26686 VDD.n4325 VDD.t236 37.0005
R26687 VDD.n2464 VDD.n2463 37.0005
R26688 VDD.t236 VDD.n2464 37.0005
R26689 VDD.n2467 VDD.n2465 37.0005
R26690 VDD.n2465 VDD.t1038 37.0005
R26691 VDD.n4314 VDD.n2466 37.0005
R26692 VDD.n2466 VDD.t1038 37.0005
R26693 VDD.n4306 VDD.n4305 37.0005
R26694 VDD.n4305 VDD.t234 37.0005
R26695 VDD.n2478 VDD.n2477 37.0005
R26696 VDD.n2477 VDD.t234 37.0005
R26697 VDD.n4296 VDD.n4295 37.0005
R26698 VDD.n4295 VDD.t262 37.0005
R26699 VDD.n2491 VDD.n2490 37.0005
R26700 VDD.n2490 VDD.t262 37.0005
R26701 VDD.n4286 VDD.n4285 37.0005
R26702 VDD.n4285 VDD.t41 37.0005
R26703 VDD.n2502 VDD.n2501 37.0005
R26704 VDD.n2501 VDD.t41 37.0005
R26705 VDD.n4276 VDD.n4275 37.0005
R26706 VDD.n4275 VDD.t322 37.0005
R26707 VDD.n2512 VDD.n2511 37.0005
R26708 VDD.n2511 VDD.t322 37.0005
R26709 VDD.n4266 VDD.n4265 37.0005
R26710 VDD.n4265 VDD.t355 37.0005
R26711 VDD.n4259 VDD.n4258 37.0005
R26712 VDD.n4258 VDD.t355 37.0005
R26713 VDD.n2389 VDD.n2388 37.0005
R26714 VDD.t903 VDD.n2389 37.0005
R26715 VDD.n4378 VDD.n2387 37.0005
R26716 VDD.n2395 VDD.n2393 37.0005
R26717 VDD.n2393 VDD.t95 37.0005
R26718 VDD.n4370 VDD.n2394 37.0005
R26719 VDD.n2394 VDD.t95 37.0005
R26720 VDD.n2406 VDD.n2404 37.0005
R26721 VDD.n2404 VDD.t591 37.0005
R26722 VDD.n4360 VDD.n2405 37.0005
R26723 VDD.n2405 VDD.t591 37.0005
R26724 VDD.n2416 VDD.n2414 37.0005
R26725 VDD.n2414 VDD.t1048 37.0005
R26726 VDD.n4350 VDD.n2415 37.0005
R26727 VDD.n2415 VDD.t1048 37.0005
R26728 VDD.n2429 VDD.n2427 37.0005
R26729 VDD.n2427 VDD.t31 37.0005
R26730 VDD.n4340 VDD.n2428 37.0005
R26731 VDD.n2428 VDD.t31 37.0005
R26732 VDD.n4324 VDD.n4323 37.0005
R26733 VDD.t236 VDD.n4324 37.0005
R26734 VDD.n4326 VDD.n2449 37.0005
R26735 VDD.t236 VDD.n2449 37.0005
R26736 VDD.n2471 VDD.n2469 37.0005
R26737 VDD.n2469 VDD.t234 37.0005
R26738 VDD.n4306 VDD.n2470 37.0005
R26739 VDD.n2470 VDD.t234 37.0005
R26740 VDD.n2483 VDD.n2481 37.0005
R26741 VDD.n2481 VDD.t262 37.0005
R26742 VDD.n4296 VDD.n2482 37.0005
R26743 VDD.n2482 VDD.t262 37.0005
R26744 VDD.n2496 VDD.n2494 37.0005
R26745 VDD.n2494 VDD.t41 37.0005
R26746 VDD.n4286 VDD.n2495 37.0005
R26747 VDD.n2495 VDD.t41 37.0005
R26748 VDD.n2507 VDD.n2505 37.0005
R26749 VDD.n2505 VDD.t322 37.0005
R26750 VDD.n4276 VDD.n2506 37.0005
R26751 VDD.n2506 VDD.t322 37.0005
R26752 VDD.n2517 VDD.n2515 37.0005
R26753 VDD.n2515 VDD.t355 37.0005
R26754 VDD.n4266 VDD.n2516 37.0005
R26755 VDD.n2516 VDD.t355 37.0005
R26756 VDD.n2441 VDD.n2439 37.0005
R26757 VDD.n2439 VDD.t426 37.0005
R26758 VDD.n4330 VDD.n2444 37.0005
R26759 VDD.n2444 VDD.t426 37.0005
R26760 VDD.n4330 VDD.n2440 37.0005
R26761 VDD.n2440 VDD.t426 37.0005
R26762 VDD.n4245 VDD.n4244 37.0005
R26763 VDD.n4244 VDD.t127 37.0005
R26764 VDD.n2537 VDD.n2536 37.0005
R26765 VDD.n2536 VDD.t127 37.0005
R26766 VDD.n4235 VDD.n4234 37.0005
R26767 VDD.n4234 VDD.t353 37.0005
R26768 VDD.n2547 VDD.n2546 37.0005
R26769 VDD.n2546 VDD.t353 37.0005
R26770 VDD.n4225 VDD.n4224 37.0005
R26771 VDD.n4224 VDD.t1022 37.0005
R26772 VDD.n2560 VDD.n2559 37.0005
R26773 VDD.n2559 VDD.t1022 37.0005
R26774 VDD.n4215 VDD.n4214 37.0005
R26775 VDD.n4214 VDD.t79 37.0005
R26776 VDD.n2572 VDD.n2571 37.0005
R26777 VDD.n2571 VDD.t79 37.0005
R26778 VDD.n2590 VDD.n2589 37.0005
R26779 VDD.n2589 VDD.t476 37.0005
R26780 VDD.n4201 VDD.n4200 37.0005
R26781 VDD.n4200 VDD.t438 37.0005
R26782 VDD.n2600 VDD.n2599 37.0005
R26783 VDD.t438 VDD.n2600 37.0005
R26784 VDD.n2603 VDD.n2601 37.0005
R26785 VDD.n2601 VDD.t1062 37.0005
R26786 VDD.n4189 VDD.n2602 37.0005
R26787 VDD.n2602 VDD.t1062 37.0005
R26788 VDD.n4181 VDD.n4180 37.0005
R26789 VDD.n4180 VDD.t440 37.0005
R26790 VDD.n2614 VDD.n2613 37.0005
R26791 VDD.n2613 VDD.t440 37.0005
R26792 VDD.n4171 VDD.n4170 37.0005
R26793 VDD.n4170 VDD.t817 37.0005
R26794 VDD.n2627 VDD.n2626 37.0005
R26795 VDD.n2626 VDD.t817 37.0005
R26796 VDD.n4161 VDD.n4160 37.0005
R26797 VDD.n4160 VDD.t59 37.0005
R26798 VDD.n2638 VDD.n2637 37.0005
R26799 VDD.n2637 VDD.t59 37.0005
R26800 VDD.n4151 VDD.n4150 37.0005
R26801 VDD.n4150 VDD.t474 37.0005
R26802 VDD.n2648 VDD.n2647 37.0005
R26803 VDD.n2647 VDD.t474 37.0005
R26804 VDD.n4141 VDD.n4140 37.0005
R26805 VDD.n4140 VDD.t320 37.0005
R26806 VDD.n4134 VDD.n4133 37.0005
R26807 VDD.n4133 VDD.t320 37.0005
R26808 VDD.n2525 VDD.n2524 37.0005
R26809 VDD.t571 VDD.n2525 37.0005
R26810 VDD.n4253 VDD.n2523 37.0005
R26811 VDD.n2531 VDD.n2529 37.0005
R26812 VDD.n2529 VDD.t127 37.0005
R26813 VDD.n4245 VDD.n2530 37.0005
R26814 VDD.n2530 VDD.t127 37.0005
R26815 VDD.n2542 VDD.n2540 37.0005
R26816 VDD.n2540 VDD.t353 37.0005
R26817 VDD.n4235 VDD.n2541 37.0005
R26818 VDD.n2541 VDD.t353 37.0005
R26819 VDD.n2552 VDD.n2550 37.0005
R26820 VDD.n2550 VDD.t1022 37.0005
R26821 VDD.n4225 VDD.n2551 37.0005
R26822 VDD.n2551 VDD.t1022 37.0005
R26823 VDD.n2565 VDD.n2563 37.0005
R26824 VDD.n2563 VDD.t79 37.0005
R26825 VDD.n4215 VDD.n2564 37.0005
R26826 VDD.n2564 VDD.t79 37.0005
R26827 VDD.n4199 VDD.n4198 37.0005
R26828 VDD.t438 VDD.n4199 37.0005
R26829 VDD.n4201 VDD.n2585 37.0005
R26830 VDD.t438 VDD.n2585 37.0005
R26831 VDD.n2607 VDD.n2605 37.0005
R26832 VDD.n2605 VDD.t440 37.0005
R26833 VDD.n4181 VDD.n2606 37.0005
R26834 VDD.n2606 VDD.t440 37.0005
R26835 VDD.n2619 VDD.n2617 37.0005
R26836 VDD.n2617 VDD.t817 37.0005
R26837 VDD.n4171 VDD.n2618 37.0005
R26838 VDD.n2618 VDD.t817 37.0005
R26839 VDD.n2632 VDD.n2630 37.0005
R26840 VDD.n2630 VDD.t59 37.0005
R26841 VDD.n4161 VDD.n2631 37.0005
R26842 VDD.n2631 VDD.t59 37.0005
R26843 VDD.n2643 VDD.n2641 37.0005
R26844 VDD.n2641 VDD.t474 37.0005
R26845 VDD.n4151 VDD.n2642 37.0005
R26846 VDD.n2642 VDD.t474 37.0005
R26847 VDD.n2653 VDD.n2651 37.0005
R26848 VDD.n2651 VDD.t320 37.0005
R26849 VDD.n4141 VDD.n2652 37.0005
R26850 VDD.n2652 VDD.t320 37.0005
R26851 VDD.n2577 VDD.n2575 37.0005
R26852 VDD.n2575 VDD.t476 37.0005
R26853 VDD.n4205 VDD.n2580 37.0005
R26854 VDD.n2580 VDD.t476 37.0005
R26855 VDD.n4205 VDD.n2576 37.0005
R26856 VDD.n2576 VDD.t476 37.0005
R26857 VDD.n4120 VDD.n4119 37.0005
R26858 VDD.n4119 VDD.t45 37.0005
R26859 VDD.n2673 VDD.n2672 37.0005
R26860 VDD.n2672 VDD.t45 37.0005
R26861 VDD.n4110 VDD.n4109 37.0005
R26862 VDD.n4109 VDD.t318 37.0005
R26863 VDD.n2683 VDD.n2682 37.0005
R26864 VDD.n2682 VDD.t318 37.0005
R26865 VDD.n4100 VDD.n4099 37.0005
R26866 VDD.n4099 VDD.t1018 37.0005
R26867 VDD.n2696 VDD.n2695 37.0005
R26868 VDD.n2695 VDD.t1018 37.0005
R26869 VDD.n4090 VDD.n4089 37.0005
R26870 VDD.n4089 VDD.t105 37.0005
R26871 VDD.n2708 VDD.n2707 37.0005
R26872 VDD.n2707 VDD.t105 37.0005
R26873 VDD.n2726 VDD.n2725 37.0005
R26874 VDD.n2725 VDD.t925 37.0005
R26875 VDD.n4076 VDD.n4075 37.0005
R26876 VDD.n4075 VDD.t525 37.0005
R26877 VDD.n2736 VDD.n2735 37.0005
R26878 VDD.t525 VDD.n2736 37.0005
R26879 VDD.n2739 VDD.n2737 37.0005
R26880 VDD.n2737 VDD.t1006 37.0005
R26881 VDD.n4064 VDD.n2738 37.0005
R26882 VDD.n2738 VDD.t1006 37.0005
R26883 VDD.n4056 VDD.n4055 37.0005
R26884 VDD.n4055 VDD.t527 37.0005
R26885 VDD.n2750 VDD.n2749 37.0005
R26886 VDD.n2749 VDD.t527 37.0005
R26887 VDD.n4046 VDD.n4045 37.0005
R26888 VDD.n4045 VDD.t295 37.0005
R26889 VDD.n2763 VDD.n2762 37.0005
R26890 VDD.n2762 VDD.t295 37.0005
R26891 VDD.n4036 VDD.n4035 37.0005
R26892 VDD.n4035 VDD.t115 37.0005
R26893 VDD.n2774 VDD.n2773 37.0005
R26894 VDD.n2773 VDD.t115 37.0005
R26895 VDD.n4026 VDD.n4025 37.0005
R26896 VDD.n4025 VDD.t0 37.0005
R26897 VDD.n2784 VDD.n2783 37.0005
R26898 VDD.n2783 VDD.t0 37.0005
R26899 VDD.n4016 VDD.n4015 37.0005
R26900 VDD.n4015 VDD.t182 37.0005
R26901 VDD.n4009 VDD.n4008 37.0005
R26902 VDD.n4008 VDD.t182 37.0005
R26903 VDD.n2661 VDD.n2660 37.0005
R26904 VDD.t876 VDD.n2661 37.0005
R26905 VDD.n4128 VDD.n2659 37.0005
R26906 VDD.n2667 VDD.n2665 37.0005
R26907 VDD.n2665 VDD.t45 37.0005
R26908 VDD.n4120 VDD.n2666 37.0005
R26909 VDD.n2666 VDD.t45 37.0005
R26910 VDD.n2678 VDD.n2676 37.0005
R26911 VDD.n2676 VDD.t318 37.0005
R26912 VDD.n4110 VDD.n2677 37.0005
R26913 VDD.n2677 VDD.t318 37.0005
R26914 VDD.n2688 VDD.n2686 37.0005
R26915 VDD.n2686 VDD.t1018 37.0005
R26916 VDD.n4100 VDD.n2687 37.0005
R26917 VDD.n2687 VDD.t1018 37.0005
R26918 VDD.n2701 VDD.n2699 37.0005
R26919 VDD.n2699 VDD.t105 37.0005
R26920 VDD.n4090 VDD.n2700 37.0005
R26921 VDD.n2700 VDD.t105 37.0005
R26922 VDD.n4074 VDD.n4073 37.0005
R26923 VDD.t525 VDD.n4074 37.0005
R26924 VDD.n4076 VDD.n2721 37.0005
R26925 VDD.t525 VDD.n2721 37.0005
R26926 VDD.n2743 VDD.n2741 37.0005
R26927 VDD.n2741 VDD.t527 37.0005
R26928 VDD.n4056 VDD.n2742 37.0005
R26929 VDD.n2742 VDD.t527 37.0005
R26930 VDD.n2755 VDD.n2753 37.0005
R26931 VDD.n2753 VDD.t295 37.0005
R26932 VDD.n4046 VDD.n2754 37.0005
R26933 VDD.n2754 VDD.t295 37.0005
R26934 VDD.n2768 VDD.n2766 37.0005
R26935 VDD.n2766 VDD.t115 37.0005
R26936 VDD.n4036 VDD.n2767 37.0005
R26937 VDD.n2767 VDD.t115 37.0005
R26938 VDD.n2779 VDD.n2777 37.0005
R26939 VDD.n2777 VDD.t0 37.0005
R26940 VDD.n4026 VDD.n2778 37.0005
R26941 VDD.n2778 VDD.t0 37.0005
R26942 VDD.n2789 VDD.n2787 37.0005
R26943 VDD.n2787 VDD.t182 37.0005
R26944 VDD.n4016 VDD.n2788 37.0005
R26945 VDD.n2788 VDD.t182 37.0005
R26946 VDD.n2713 VDD.n2711 37.0005
R26947 VDD.n2711 VDD.t925 37.0005
R26948 VDD.n4080 VDD.n2716 37.0005
R26949 VDD.n2716 VDD.t925 37.0005
R26950 VDD.n4080 VDD.n2712 37.0005
R26951 VDD.n2712 VDD.t925 37.0005
R26952 VDD.n3995 VDD.n3994 37.0005
R26953 VDD.n3994 VDD.t93 37.0005
R26954 VDD.n2809 VDD.n2808 37.0005
R26955 VDD.n2808 VDD.t93 37.0005
R26956 VDD.n3985 VDD.n3984 37.0005
R26957 VDD.n3984 VDD.t180 37.0005
R26958 VDD.n2819 VDD.n2818 37.0005
R26959 VDD.n2818 VDD.t180 37.0005
R26960 VDD.n3975 VDD.n3974 37.0005
R26961 VDD.n3974 VDD.t1045 37.0005
R26962 VDD.n2832 VDD.n2831 37.0005
R26963 VDD.n2831 VDD.t1045 37.0005
R26964 VDD.n3965 VDD.n3964 37.0005
R26965 VDD.n3964 VDD.t27 37.0005
R26966 VDD.n2844 VDD.n2843 37.0005
R26967 VDD.n2843 VDD.t27 37.0005
R26968 VDD.n2862 VDD.n2861 37.0005
R26969 VDD.n2861 VDD.t373 37.0005
R26970 VDD.n3951 VDD.n3950 37.0005
R26971 VDD.n3950 VDD.t510 37.0005
R26972 VDD.n2872 VDD.n2871 37.0005
R26973 VDD.t510 VDD.n2872 37.0005
R26974 VDD.n2875 VDD.n2873 37.0005
R26975 VDD.n2873 VDD.t1034 37.0005
R26976 VDD.n3939 VDD.n2874 37.0005
R26977 VDD.n2874 VDD.t1034 37.0005
R26978 VDD.n3931 VDD.n3930 37.0005
R26979 VDD.n3930 VDD.t543 37.0005
R26980 VDD.n2886 VDD.n2885 37.0005
R26981 VDD.n2885 VDD.t543 37.0005
R26982 VDD.n3921 VDD.n3920 37.0005
R26983 VDD.n3920 VDD.t166 37.0005
R26984 VDD.n2899 VDD.n2898 37.0005
R26985 VDD.n2898 VDD.t166 37.0005
R26986 VDD.n3911 VDD.n3910 37.0005
R26987 VDD.n3910 VDD.t37 37.0005
R26988 VDD.n2910 VDD.n2909 37.0005
R26989 VDD.n2909 VDD.t37 37.0005
R26990 VDD.n3901 VDD.n3900 37.0005
R26991 VDD.n3900 VDD.t704 37.0005
R26992 VDD.n2920 VDD.n2919 37.0005
R26993 VDD.n2919 VDD.t704 37.0005
R26994 VDD.n3891 VDD.n3890 37.0005
R26995 VDD.n3890 VDD.t689 37.0005
R26996 VDD.n3884 VDD.n3883 37.0005
R26997 VDD.n3883 VDD.t689 37.0005
R26998 VDD.n2797 VDD.n2796 37.0005
R26999 VDD.t1102 VDD.n2797 37.0005
R27000 VDD.n4003 VDD.n2795 37.0005
R27001 VDD.n2803 VDD.n2801 37.0005
R27002 VDD.n2801 VDD.t93 37.0005
R27003 VDD.n3995 VDD.n2802 37.0005
R27004 VDD.n2802 VDD.t93 37.0005
R27005 VDD.n2814 VDD.n2812 37.0005
R27006 VDD.n2812 VDD.t180 37.0005
R27007 VDD.n3985 VDD.n2813 37.0005
R27008 VDD.n2813 VDD.t180 37.0005
R27009 VDD.n2824 VDD.n2822 37.0005
R27010 VDD.n2822 VDD.t1045 37.0005
R27011 VDD.n3975 VDD.n2823 37.0005
R27012 VDD.n2823 VDD.t1045 37.0005
R27013 VDD.n2837 VDD.n2835 37.0005
R27014 VDD.n2835 VDD.t27 37.0005
R27015 VDD.n3965 VDD.n2836 37.0005
R27016 VDD.n2836 VDD.t27 37.0005
R27017 VDD.n3949 VDD.n3948 37.0005
R27018 VDD.t510 VDD.n3949 37.0005
R27019 VDD.n3951 VDD.n2857 37.0005
R27020 VDD.t510 VDD.n2857 37.0005
R27021 VDD.n2879 VDD.n2877 37.0005
R27022 VDD.n2877 VDD.t543 37.0005
R27023 VDD.n3931 VDD.n2878 37.0005
R27024 VDD.n2878 VDD.t543 37.0005
R27025 VDD.n2891 VDD.n2889 37.0005
R27026 VDD.n2889 VDD.t166 37.0005
R27027 VDD.n3921 VDD.n2890 37.0005
R27028 VDD.n2890 VDD.t166 37.0005
R27029 VDD.n2904 VDD.n2902 37.0005
R27030 VDD.n2902 VDD.t37 37.0005
R27031 VDD.n3911 VDD.n2903 37.0005
R27032 VDD.n2903 VDD.t37 37.0005
R27033 VDD.n2915 VDD.n2913 37.0005
R27034 VDD.n2913 VDD.t704 37.0005
R27035 VDD.n3901 VDD.n2914 37.0005
R27036 VDD.n2914 VDD.t704 37.0005
R27037 VDD.n2925 VDD.n2923 37.0005
R27038 VDD.n2923 VDD.t689 37.0005
R27039 VDD.n3891 VDD.n2924 37.0005
R27040 VDD.n2924 VDD.t689 37.0005
R27041 VDD.n2849 VDD.n2847 37.0005
R27042 VDD.n2847 VDD.t373 37.0005
R27043 VDD.n3955 VDD.n2852 37.0005
R27044 VDD.n2852 VDD.t373 37.0005
R27045 VDD.n3955 VDD.n2848 37.0005
R27046 VDD.n2848 VDD.t373 37.0005
R27047 VDD.n3556 VDD.n3555 37.0005
R27048 VDD.n3555 VDD.t160 37.0005
R27049 VDD.n3215 VDD.n3214 37.0005
R27050 VDD.t160 VDD.n3215 37.0005
R27051 VDD.n3543 VDD.n3542 37.0005
R27052 VDD.n3542 VDD.t315 37.0005
R27053 VDD.n3224 VDD.n3223 37.0005
R27054 VDD.n3223 VDD.t315 37.0005
R27055 VDD.n3233 VDD.n3232 37.0005
R27056 VDD.n3232 VDD.t282 37.0005
R27057 VDD.n3554 VDD.n3553 37.0005
R27058 VDD.t160 VDD.n3554 37.0005
R27059 VDD.n3556 VDD.n3207 37.0005
R27060 VDD.t160 VDD.n3207 37.0005
R27061 VDD.n3219 VDD.n3217 37.0005
R27062 VDD.n3217 VDD.t315 37.0005
R27063 VDD.n3543 VDD.n3218 37.0005
R27064 VDD.n3218 VDD.t315 37.0005
R27065 VDD.n3229 VDD.n3227 37.0005
R27066 VDD.n3227 VDD.t282 37.0005
R27067 VDD.n3533 VDD.n3239 37.0005
R27068 VDD.n3239 VDD.t282 37.0005
R27069 VDD.n3533 VDD.n3228 37.0005
R27070 VDD.n3228 VDD.t282 37.0005
R27071 VDD.n3289 VDD.n3287 37.0005
R27072 VDD.n3287 VDD.t386 37.0005
R27073 VDD.n3379 VDD.n3288 37.0005
R27074 VDD.n3288 VDD.t386 37.0005
R27075 VDD.n3286 VDD.n3285 37.0005
R27076 VDD.t307 VDD.n3286 37.0005
R27077 VDD.n3388 VDD.n3284 37.0005
R27078 VDD.n3366 VDD.n3365 37.0005
R27079 VDD.t384 VDD.n3366 37.0005
R27080 VDD.n3374 VDD.n3364 37.0005
R27081 VDD.n3398 VDD.n3396 37.0005
R27082 VDD.n3396 VDD.t992 37.0005
R27083 VDD.n3416 VDD.n3397 37.0005
R27084 VDD.n3397 VDD.t992 37.0005
R27085 VDD.n3395 VDD.n3394 37.0005
R27086 VDD.t618 VDD.n3395 37.0005
R27087 VDD.n3425 VDD.n3393 37.0005
R27088 VDD.n3404 VDD.n3403 37.0005
R27089 VDD.t990 VDD.n3404 37.0005
R27090 VDD.n3412 VDD.n3402 37.0005
R27091 VDD.n3264 VDD.n3262 37.0005
R27092 VDD.n3262 VDD.t225 37.0005
R27093 VDD.n3445 VDD.n3263 37.0005
R27094 VDD.n3263 VDD.t225 37.0005
R27095 VDD.n3269 VDD.n3268 37.0005
R27096 VDD.t381 VDD.n3269 37.0005
R27097 VDD.n3277 VDD.n3267 37.0005
R27098 VDD.n3259 VDD.n3258 37.0005
R27099 VDD.t464 VDD.n3259 37.0005
R27100 VDD.n3452 VDD.n3257 37.0005
R27101 VDD.n3252 VDD.n3250 37.0005
R27102 VDD.n3250 VDD.t407 37.0005
R27103 VDD.n3474 VDD.n3251 37.0005
R27104 VDD.n3251 VDD.t407 37.0005
R27105 VDD.n3249 VDD.n3248 37.0005
R27106 VDD.t867 VDD.n3249 37.0005
R27107 VDD.n3483 VDD.n3247 37.0005
R27108 VDD.n3461 VDD.n3460 37.0005
R27109 VDD.t405 VDD.n3461 37.0005
R27110 VDD.n3469 VDD.n3459 37.0005
R27111 VDD.n3492 VDD.n3490 37.0005
R27112 VDD.n3490 VDD.t642 37.0005
R27113 VDD.n3510 VDD.n3491 37.0005
R27114 VDD.n3491 VDD.t642 37.0005
R27115 VDD.n3489 VDD.n3488 37.0005
R27116 VDD.t966 VDD.n3489 37.0005
R27117 VDD.n3519 VDD.n3487 37.0005
R27118 VDD.n3498 VDD.n3497 37.0005
R27119 VDD.t640 VDD.n3498 37.0005
R27120 VDD.n3506 VDD.n3496 37.0005
R27121 VDD.n3320 VDD.n3318 37.0005
R27122 VDD.n3318 VDD.t213 37.0005
R27123 VDD.n3350 VDD.n3319 37.0005
R27124 VDD.n3319 VDD.t213 37.0005
R27125 VDD.n3325 VDD.n3324 37.0005
R27126 VDD.t533 VDD.n3325 37.0005
R27127 VDD.n3333 VDD.n3323 37.0005
R27128 VDD.n3315 VDD.n3314 37.0005
R27129 VDD.t211 VDD.n3315 37.0005
R27130 VDD.n3357 VDD.n3313 37.0005
R27131 VDD.n3870 VDD.n3869 37.0005
R27132 VDD.n3869 VDD.t119 37.0005
R27133 VDD.n2945 VDD.n2944 37.0005
R27134 VDD.n2944 VDD.t119 37.0005
R27135 VDD.n3860 VDD.n3859 37.0005
R27136 VDD.n3859 VDD.t692 37.0005
R27137 VDD.n2955 VDD.n2954 37.0005
R27138 VDD.n2954 VDD.t692 37.0005
R27139 VDD.n3850 VDD.n3849 37.0005
R27140 VDD.n3849 VDD.t1014 37.0005
R27141 VDD.n2968 VDD.n2967 37.0005
R27142 VDD.n2967 VDD.t1014 37.0005
R27143 VDD.n3840 VDD.n3839 37.0005
R27144 VDD.n3839 VDD.t75 37.0005
R27145 VDD.n3670 VDD.n3669 37.0005
R27146 VDD.n3669 VDD.t75 37.0005
R27147 VDD.n3688 VDD.n3687 37.0005
R27148 VDD.n3687 VDD.t164 37.0005
R27149 VDD.n3826 VDD.n3825 37.0005
R27150 VDD.n3825 VDD.t162 37.0005
R27151 VDD.n3698 VDD.n3697 37.0005
R27152 VDD.t162 VDD.n3698 37.0005
R27153 VDD.n3701 VDD.n3699 37.0005
R27154 VDD.n3699 VDD.t1094 37.0005
R27155 VDD.n3814 VDD.n3700 37.0005
R27156 VDD.n3700 VDD.t1094 37.0005
R27157 VDD.n3806 VDD.n3805 37.0005
R27158 VDD.n3805 VDD.t246 37.0005
R27159 VDD.n3712 VDD.n3711 37.0005
R27160 VDD.n3711 VDD.t246 37.0005
R27161 VDD.n3796 VDD.n3795 37.0005
R27162 VDD.n3795 VDD.t550 37.0005
R27163 VDD.n3725 VDD.n3724 37.0005
R27164 VDD.n3724 VDD.t550 37.0005
R27165 VDD.n3786 VDD.n3785 37.0005
R27166 VDD.n3785 VDD.t35 37.0005
R27167 VDD.n3736 VDD.n3735 37.0005
R27168 VDD.n3735 VDD.t35 37.0005
R27169 VDD.n3776 VDD.n3775 37.0005
R27170 VDD.n3775 VDD.t633 37.0005
R27171 VDD.n3746 VDD.n3745 37.0005
R27172 VDD.n3745 VDD.t633 37.0005
R27173 VDD.n3766 VDD.n3765 37.0005
R27174 VDD.n3765 VDD.t347 37.0005
R27175 VDD.n3759 VDD.n3758 37.0005
R27176 VDD.n3758 VDD.t347 37.0005
R27177 VDD.n2933 VDD.n2932 37.0005
R27178 VDD.t696 VDD.n2933 37.0005
R27179 VDD.n3878 VDD.n2931 37.0005
R27180 VDD.n2939 VDD.n2937 37.0005
R27181 VDD.n2937 VDD.t119 37.0005
R27182 VDD.n3870 VDD.n2938 37.0005
R27183 VDD.n2938 VDD.t119 37.0005
R27184 VDD.n2950 VDD.n2948 37.0005
R27185 VDD.n2948 VDD.t692 37.0005
R27186 VDD.n3860 VDD.n2949 37.0005
R27187 VDD.n2949 VDD.t692 37.0005
R27188 VDD.n2960 VDD.n2958 37.0005
R27189 VDD.n2958 VDD.t1014 37.0005
R27190 VDD.n3850 VDD.n2959 37.0005
R27191 VDD.n2959 VDD.t1014 37.0005
R27192 VDD.n2973 VDD.n2971 37.0005
R27193 VDD.n2971 VDD.t75 37.0005
R27194 VDD.n3840 VDD.n2972 37.0005
R27195 VDD.n2972 VDD.t75 37.0005
R27196 VDD.n3824 VDD.n3823 37.0005
R27197 VDD.t162 VDD.n3824 37.0005
R27198 VDD.n3826 VDD.n3683 37.0005
R27199 VDD.t162 VDD.n3683 37.0005
R27200 VDD.n3705 VDD.n3703 37.0005
R27201 VDD.n3703 VDD.t246 37.0005
R27202 VDD.n3806 VDD.n3704 37.0005
R27203 VDD.n3704 VDD.t246 37.0005
R27204 VDD.n3717 VDD.n3715 37.0005
R27205 VDD.n3715 VDD.t550 37.0005
R27206 VDD.n3796 VDD.n3716 37.0005
R27207 VDD.n3716 VDD.t550 37.0005
R27208 VDD.n3730 VDD.n3728 37.0005
R27209 VDD.n3728 VDD.t35 37.0005
R27210 VDD.n3786 VDD.n3729 37.0005
R27211 VDD.n3729 VDD.t35 37.0005
R27212 VDD.n3741 VDD.n3739 37.0005
R27213 VDD.n3739 VDD.t633 37.0005
R27214 VDD.n3776 VDD.n3740 37.0005
R27215 VDD.n3740 VDD.t633 37.0005
R27216 VDD.n3751 VDD.n3749 37.0005
R27217 VDD.n3749 VDD.t347 37.0005
R27218 VDD.n3766 VDD.n3750 37.0005
R27219 VDD.n3750 VDD.t347 37.0005
R27220 VDD.n3675 VDD.n3673 37.0005
R27221 VDD.n3673 VDD.t164 37.0005
R27222 VDD.n3830 VDD.n3678 37.0005
R27223 VDD.n3678 VDD.t164 37.0005
R27224 VDD.n3830 VDD.n3674 37.0005
R27225 VDD.n3674 VDD.t164 37.0005
R27226 VDD.n271 VDD.n269 36.8325
R27227 VDD.n274 VDD.n273 36.8325
R27228 VDD.n256 VDD.n255 36.7882
R27229 VDD.n262 VDD.n261 36.7882
R27230 VDD.n3666 VDD.n3647 34.7977
R27231 VDD.n281 VDD.n240 34.146
R27232 VDD.n7070 VDD.n6827 33.6641
R27233 VDD.n3626 VDD.n3625 33.3344
R27234 VDD.n3139 VDD.n3075 33.3344
R27235 VDD.n7470 VDD.n7468 31.6493
R27236 VDD.n1587 VDD.n1583 31.6493
R27237 VDD.n1327 VDD.n1323 31.6493
R27238 VDD.n1067 VDD.n1063 31.6493
R27239 VDD.n807 VDD.n803 31.6493
R27240 VDD.n547 VDD.n543 31.6493
R27241 VDD.n287 VDD.n283 31.6493
R27242 VDD.n7203 VDD.n7199 31.6493
R27243 VDD.n1847 VDD.n1843 31.6493
R27244 VDD.n5962 VDD.n5960 31.6493
R27245 VDD.n5826 VDD.n5824 31.6493
R27246 VDD.n5690 VDD.n5688 31.6493
R27247 VDD.n5554 VDD.n5552 31.6493
R27248 VDD.n5418 VDD.n5416 31.6493
R27249 VDD.n5282 VDD.n5280 31.6493
R27250 VDD.n5146 VDD.n5144 31.6493
R27251 VDD.n5008 VDD.n4757 31.6493
R27252 VDD.n1983 VDD.n1979 31.6493
R27253 VDD.n2119 VDD.n2115 31.6493
R27254 VDD.n2255 VDD.n2251 31.6493
R27255 VDD.n2391 VDD.n2387 31.6493
R27256 VDD.n2527 VDD.n2523 31.6493
R27257 VDD.n2663 VDD.n2659 31.6493
R27258 VDD.n2799 VDD.n2795 31.6493
R27259 VDD.n2935 VDD.n2931 31.6493
R27260 VDD.n3625 VDD.n3584 29.9244
R27261 VDD.n3584 VDD.n2997 29.9244
R27262 VDD.n3181 VDD.n2997 29.9244
R27263 VDD.n3181 VDD.n3180 29.9244
R27264 VDD.n3180 VDD.n3139 29.9244
R27265 VDD.n3136 VDD.n3036 29.9244
R27266 VDD.n3203 VDD.n3036 29.9244
R27267 VDD.n3580 VDD.n3203 29.9244
R27268 VDD.n3581 VDD.n3580 29.9244
R27269 VDD.n3581 VDD.n2977 29.9244
R27270 VDD.n3647 VDD.n2977 29.9244
R27271 VDD.n3135 VDD.n3134 29.7994
R27272 VDD.n102 VDD.n99 28.7118
R27273 VDD.n97 VDD.n93 28.7118
R27274 VDD.n116 VDD.n86 28.7118
R27275 VDD.n81 VDD.n77 28.7118
R27276 VDD.n137 VDD.n74 28.7118
R27277 VDD.n72 VDD.n68 28.7118
R27278 VDD.n151 VDD.n61 28.7118
R27279 VDD.n56 VDD.n52 28.7118
R27280 VDD.n172 VDD.n49 28.7118
R27281 VDD.n47 VDD.n43 28.7118
R27282 VDD.n186 VDD.n36 28.7118
R27283 VDD.n31 VDD.n27 28.7118
R27284 VDD.n207 VDD.n24 28.7118
R27285 VDD.n22 VDD.n18 28.7118
R27286 VDD.n221 VDD.n11 28.7118
R27287 VDD.n6 VDD.n2 28.7118
R27288 VDD.n6936 VDD.n6933 28.7118
R27289 VDD.n6931 VDD.n6927 28.7118
R27290 VDD.n6950 VDD.n6920 28.7118
R27291 VDD.n6915 VDD.n6911 28.7118
R27292 VDD.n6971 VDD.n6908 28.7118
R27293 VDD.n6906 VDD.n6902 28.7118
R27294 VDD.n6985 VDD.n6895 28.7118
R27295 VDD.n6890 VDD.n6886 28.7118
R27296 VDD.n7006 VDD.n6883 28.7118
R27297 VDD.n6881 VDD.n6877 28.7118
R27298 VDD.n7020 VDD.n6870 28.7118
R27299 VDD.n6865 VDD.n6861 28.7118
R27300 VDD.n7041 VDD.n6858 28.7118
R27301 VDD.n6856 VDD.n6852 28.7118
R27302 VDD.n7055 VDD.n6848 28.7118
R27303 VDD.n6839 VDD.n6835 28.7118
R27304 VDD.n3385 VDD.n3284 28.7118
R27305 VDD.n3368 VDD.n3364 28.7118
R27306 VDD.n3422 VDD.n3393 28.7118
R27307 VDD.n3406 VDD.n3402 28.7118
R27308 VDD.n3274 VDD.n3267 28.7118
R27309 VDD.n3261 VDD.n3257 28.7118
R27310 VDD.n3480 VDD.n3247 28.7118
R27311 VDD.n3463 VDD.n3459 28.7118
R27312 VDD.n3516 VDD.n3487 28.7118
R27313 VDD.n3500 VDD.n3496 28.7118
R27314 VDD.n3330 VDD.n3323 28.7118
R27315 VDD.n3317 VDD.n3313 28.7118
R27316 VDD VDD.n218 26.3103
R27317 VDD VDD.n204 26.3103
R27318 VDD VDD.n183 26.3103
R27319 VDD VDD.n169 26.3103
R27320 VDD VDD.n148 26.3103
R27321 VDD VDD.n134 26.3103
R27322 VDD VDD.n113 26.3103
R27323 VDD VDD.n7052 26.3103
R27324 VDD VDD.n7038 26.3103
R27325 VDD VDD.n7017 26.3103
R27326 VDD VDD.n7003 26.3103
R27327 VDD VDD.n6982 26.3103
R27328 VDD VDD.n6968 26.3103
R27329 VDD VDD.n6947 26.3103
R27330 VDD.n3138 VDD.n3137 25.8669
R27331 VDD.n3179 VDD.n3178 25.8669
R27332 VDD.n3202 VDD.n3182 25.8669
R27333 VDD.n3583 VDD.n3582 25.8669
R27334 VDD.n3624 VDD.n3623 25.8669
R27335 VDD.n3646 VDD.n3626 25.8669
R27336 VDD.n3133 VDD.n3075 25.8669
R27337 VDD.n256 VDD.n254 24.6676
R27338 VDD.n262 VDD.n249 24.6676
R27339 VDD.n3245 VDD 24.3918
R27340 VDD.t699 VDD.n250 23.5846
R27341 VDD.t701 VDD.n250 23.5846
R27342 VDD.n7478 VDD.n7465 23.1255
R27343 VDD.n7477 VDD.n7465 23.1255
R27344 VDD.n7479 VDD.n7466 23.1255
R27345 VDD.n7707 VDD.n7466 23.1255
R27346 VDD.n7486 VDD.n7482 23.1255
R27347 VDD.n7706 VDD.n7482 23.1255
R27348 VDD.n7700 VDD.n7490 23.1255
R27349 VDD.n7700 VDD.n7699 23.1255
R27350 VDD.n7495 VDD.n7491 23.1255
R27351 VDD.n7696 VDD.n7491 23.1255
R27352 VDD.n7690 VDD.n7503 23.1255
R27353 VDD.n7690 VDD.n7689 23.1255
R27354 VDD.n7508 VDD.n7504 23.1255
R27355 VDD.n7686 VDD.n7504 23.1255
R27356 VDD.n7680 VDD.n7514 23.1255
R27357 VDD.n7680 VDD.n7679 23.1255
R27358 VDD.n7519 VDD.n7515 23.1255
R27359 VDD.n7676 VDD.n7515 23.1255
R27360 VDD.n7670 VDD.n7524 23.1255
R27361 VDD.n7670 VDD.n7669 23.1255
R27362 VDD.n7529 VDD.n7525 23.1255
R27363 VDD.n7666 VDD.n7525 23.1255
R27364 VDD.n7660 VDD.n7537 23.1255
R27365 VDD.n7660 VDD.n7659 23.1255
R27366 VDD.n7655 VDD.n7654 23.1255
R27367 VDD.n7656 VDD.n7655 23.1255
R27368 VDD.n7652 VDD.n7651 23.1255
R27369 VDD.n7651 VDD.n7650 23.1255
R27370 VDD.n7545 VDD.n7541 23.1255
R27371 VDD.n7649 VDD.n7541 23.1255
R27372 VDD.n7643 VDD.n7552 23.1255
R27373 VDD.n7643 VDD.n7642 23.1255
R27374 VDD.n7557 VDD.n7553 23.1255
R27375 VDD.n7639 VDD.n7553 23.1255
R27376 VDD.n7633 VDD.n7565 23.1255
R27377 VDD.n7633 VDD.n7632 23.1255
R27378 VDD.n7570 VDD.n7566 23.1255
R27379 VDD.n7629 VDD.n7566 23.1255
R27380 VDD.n7623 VDD.n7576 23.1255
R27381 VDD.n7623 VDD.n7622 23.1255
R27382 VDD.n7581 VDD.n7577 23.1255
R27383 VDD.n7619 VDD.n7577 23.1255
R27384 VDD.n7613 VDD.n7586 23.1255
R27385 VDD.n7613 VDD.n7612 23.1255
R27386 VDD.n7591 VDD.n7587 23.1255
R27387 VDD.n7609 VDD.n7587 23.1255
R27388 VDD.n7603 VDD.n7599 23.1255
R27389 VDD.n7603 VDD.n7602 23.1255
R27390 VDD.n7710 VDD.n7708 23.1255
R27391 VDD.n7708 VDD.n7477 23.1255
R27392 VDD.n7711 VDD.n7709 23.1255
R27393 VDD.n7709 VDD.n7707 23.1255
R27394 VDD.n7705 VDD.n7704 23.1255
R27395 VDD.n7706 VDD.n7705 23.1255
R27396 VDD.n7698 VDD.n7697 23.1255
R27397 VDD.n7699 VDD.n7698 23.1255
R27398 VDD.n7695 VDD.n7694 23.1255
R27399 VDD.n7696 VDD.n7695 23.1255
R27400 VDD.n7688 VDD.n7687 23.1255
R27401 VDD.n7689 VDD.n7688 23.1255
R27402 VDD.n7685 VDD.n7684 23.1255
R27403 VDD.n7686 VDD.n7685 23.1255
R27404 VDD.n7678 VDD.n7677 23.1255
R27405 VDD.n7679 VDD.n7678 23.1255
R27406 VDD.n7675 VDD.n7674 23.1255
R27407 VDD.n7676 VDD.n7675 23.1255
R27408 VDD.n7668 VDD.n7667 23.1255
R27409 VDD.n7669 VDD.n7668 23.1255
R27410 VDD.n7665 VDD.n7664 23.1255
R27411 VDD.n7666 VDD.n7665 23.1255
R27412 VDD.n7658 VDD.n7657 23.1255
R27413 VDD.n7659 VDD.n7658 23.1255
R27414 VDD.n7648 VDD.n7647 23.1255
R27415 VDD.n7649 VDD.n7648 23.1255
R27416 VDD.n7641 VDD.n7640 23.1255
R27417 VDD.n7642 VDD.n7641 23.1255
R27418 VDD.n7638 VDD.n7637 23.1255
R27419 VDD.n7639 VDD.n7638 23.1255
R27420 VDD.n7631 VDD.n7630 23.1255
R27421 VDD.n7632 VDD.n7631 23.1255
R27422 VDD.n7628 VDD.n7627 23.1255
R27423 VDD.n7629 VDD.n7628 23.1255
R27424 VDD.n7621 VDD.n7620 23.1255
R27425 VDD.n7622 VDD.n7621 23.1255
R27426 VDD.n7618 VDD.n7617 23.1255
R27427 VDD.n7619 VDD.n7618 23.1255
R27428 VDD.n7611 VDD.n7610 23.1255
R27429 VDD.n7612 VDD.n7611 23.1255
R27430 VDD.n7608 VDD.n7607 23.1255
R27431 VDD.n7609 VDD.n7608 23.1255
R27432 VDD.n7601 VDD.n7600 23.1255
R27433 VDD.n7602 VDD.n7601 23.1255
R27434 VDD.n7475 VDD.n7474 23.1255
R27435 VDD.n7476 VDD.n7475 23.1255
R27436 VDD.n7472 VDD.n7471 23.1255
R27437 VDD.n1592 VDD.n1588 23.1255
R27438 VDD.n1834 VDD.n1588 23.1255
R27439 VDD.n1828 VDD.n1598 23.1255
R27440 VDD.n1828 VDD.n1827 23.1255
R27441 VDD.n1603 VDD.n1599 23.1255
R27442 VDD.n1824 VDD.n1599 23.1255
R27443 VDD.n1818 VDD.n1608 23.1255
R27444 VDD.n1818 VDD.n1817 23.1255
R27445 VDD.n1613 VDD.n1609 23.1255
R27446 VDD.n1814 VDD.n1609 23.1255
R27447 VDD.n1808 VDD.n1621 23.1255
R27448 VDD.n1808 VDD.n1807 23.1255
R27449 VDD.n1626 VDD.n1622 23.1255
R27450 VDD.n1804 VDD.n1622 23.1255
R27451 VDD.n1798 VDD.n1632 23.1255
R27452 VDD.n1798 VDD.n1797 23.1255
R27453 VDD.n1637 VDD.n1633 23.1255
R27454 VDD.n1794 VDD.n1633 23.1255
R27455 VDD.n1788 VDD.n1642 23.1255
R27456 VDD.n1788 VDD.n1787 23.1255
R27457 VDD.n1647 VDD.n1643 23.1255
R27458 VDD.n1784 VDD.n1643 23.1255
R27459 VDD.n1778 VDD.n1655 23.1255
R27460 VDD.n1778 VDD.n1777 23.1255
R27461 VDD.n1773 VDD.n1772 23.1255
R27462 VDD.n1774 VDD.n1773 23.1255
R27463 VDD.n1770 VDD.n1769 23.1255
R27464 VDD.n1769 VDD.n1768 23.1255
R27465 VDD.n1663 VDD.n1659 23.1255
R27466 VDD.n1767 VDD.n1659 23.1255
R27467 VDD.n1761 VDD.n1670 23.1255
R27468 VDD.n1761 VDD.n1760 23.1255
R27469 VDD.n1675 VDD.n1671 23.1255
R27470 VDD.n1757 VDD.n1671 23.1255
R27471 VDD.n1751 VDD.n1683 23.1255
R27472 VDD.n1751 VDD.n1750 23.1255
R27473 VDD.n1688 VDD.n1684 23.1255
R27474 VDD.n1747 VDD.n1684 23.1255
R27475 VDD.n1741 VDD.n1694 23.1255
R27476 VDD.n1741 VDD.n1740 23.1255
R27477 VDD.n1699 VDD.n1695 23.1255
R27478 VDD.n1737 VDD.n1695 23.1255
R27479 VDD.n1731 VDD.n1704 23.1255
R27480 VDD.n1731 VDD.n1730 23.1255
R27481 VDD.n1709 VDD.n1705 23.1255
R27482 VDD.n1727 VDD.n1705 23.1255
R27483 VDD.n1721 VDD.n1717 23.1255
R27484 VDD.n1721 VDD.n1720 23.1255
R27485 VDD.n1833 VDD.n1832 23.1255
R27486 VDD.n1834 VDD.n1833 23.1255
R27487 VDD.n1826 VDD.n1825 23.1255
R27488 VDD.n1827 VDD.n1826 23.1255
R27489 VDD.n1823 VDD.n1822 23.1255
R27490 VDD.n1824 VDD.n1823 23.1255
R27491 VDD.n1816 VDD.n1815 23.1255
R27492 VDD.n1817 VDD.n1816 23.1255
R27493 VDD.n1813 VDD.n1812 23.1255
R27494 VDD.n1814 VDD.n1813 23.1255
R27495 VDD.n1806 VDD.n1805 23.1255
R27496 VDD.n1807 VDD.n1806 23.1255
R27497 VDD.n1803 VDD.n1802 23.1255
R27498 VDD.n1804 VDD.n1803 23.1255
R27499 VDD.n1796 VDD.n1795 23.1255
R27500 VDD.n1797 VDD.n1796 23.1255
R27501 VDD.n1793 VDD.n1792 23.1255
R27502 VDD.n1794 VDD.n1793 23.1255
R27503 VDD.n1786 VDD.n1785 23.1255
R27504 VDD.n1787 VDD.n1786 23.1255
R27505 VDD.n1783 VDD.n1782 23.1255
R27506 VDD.n1784 VDD.n1783 23.1255
R27507 VDD.n1776 VDD.n1775 23.1255
R27508 VDD.n1777 VDD.n1776 23.1255
R27509 VDD.n1766 VDD.n1765 23.1255
R27510 VDD.n1767 VDD.n1766 23.1255
R27511 VDD.n1759 VDD.n1758 23.1255
R27512 VDD.n1760 VDD.n1759 23.1255
R27513 VDD.n1756 VDD.n1755 23.1255
R27514 VDD.n1757 VDD.n1756 23.1255
R27515 VDD.n1749 VDD.n1748 23.1255
R27516 VDD.n1750 VDD.n1749 23.1255
R27517 VDD.n1746 VDD.n1745 23.1255
R27518 VDD.n1747 VDD.n1746 23.1255
R27519 VDD.n1739 VDD.n1738 23.1255
R27520 VDD.n1740 VDD.n1739 23.1255
R27521 VDD.n1736 VDD.n1735 23.1255
R27522 VDD.n1737 VDD.n1736 23.1255
R27523 VDD.n1729 VDD.n1728 23.1255
R27524 VDD.n1730 VDD.n1729 23.1255
R27525 VDD.n1726 VDD.n1725 23.1255
R27526 VDD.n1727 VDD.n1726 23.1255
R27527 VDD.n1719 VDD.n1718 23.1255
R27528 VDD.n1720 VDD.n1719 23.1255
R27529 VDD.n1837 VDD.n1836 23.1255
R27530 VDD.n1836 VDD.n1835 23.1255
R27531 VDD.n1586 VDD.n1582 23.1255
R27532 VDD.n1332 VDD.n1328 23.1255
R27533 VDD.n1574 VDD.n1328 23.1255
R27534 VDD.n1568 VDD.n1338 23.1255
R27535 VDD.n1568 VDD.n1567 23.1255
R27536 VDD.n1343 VDD.n1339 23.1255
R27537 VDD.n1564 VDD.n1339 23.1255
R27538 VDD.n1558 VDD.n1348 23.1255
R27539 VDD.n1558 VDD.n1557 23.1255
R27540 VDD.n1353 VDD.n1349 23.1255
R27541 VDD.n1554 VDD.n1349 23.1255
R27542 VDD.n1548 VDD.n1361 23.1255
R27543 VDD.n1548 VDD.n1547 23.1255
R27544 VDD.n1366 VDD.n1362 23.1255
R27545 VDD.n1544 VDD.n1362 23.1255
R27546 VDD.n1538 VDD.n1372 23.1255
R27547 VDD.n1538 VDD.n1537 23.1255
R27548 VDD.n1377 VDD.n1373 23.1255
R27549 VDD.n1534 VDD.n1373 23.1255
R27550 VDD.n1528 VDD.n1382 23.1255
R27551 VDD.n1528 VDD.n1527 23.1255
R27552 VDD.n1387 VDD.n1383 23.1255
R27553 VDD.n1524 VDD.n1383 23.1255
R27554 VDD.n1518 VDD.n1395 23.1255
R27555 VDD.n1518 VDD.n1517 23.1255
R27556 VDD.n1513 VDD.n1512 23.1255
R27557 VDD.n1514 VDD.n1513 23.1255
R27558 VDD.n1510 VDD.n1509 23.1255
R27559 VDD.n1509 VDD.n1508 23.1255
R27560 VDD.n1403 VDD.n1399 23.1255
R27561 VDD.n1507 VDD.n1399 23.1255
R27562 VDD.n1501 VDD.n1410 23.1255
R27563 VDD.n1501 VDD.n1500 23.1255
R27564 VDD.n1415 VDD.n1411 23.1255
R27565 VDD.n1497 VDD.n1411 23.1255
R27566 VDD.n1491 VDD.n1423 23.1255
R27567 VDD.n1491 VDD.n1490 23.1255
R27568 VDD.n1428 VDD.n1424 23.1255
R27569 VDD.n1487 VDD.n1424 23.1255
R27570 VDD.n1481 VDD.n1434 23.1255
R27571 VDD.n1481 VDD.n1480 23.1255
R27572 VDD.n1439 VDD.n1435 23.1255
R27573 VDD.n1477 VDD.n1435 23.1255
R27574 VDD.n1471 VDD.n1444 23.1255
R27575 VDD.n1471 VDD.n1470 23.1255
R27576 VDD.n1449 VDD.n1445 23.1255
R27577 VDD.n1467 VDD.n1445 23.1255
R27578 VDD.n1461 VDD.n1457 23.1255
R27579 VDD.n1461 VDD.n1460 23.1255
R27580 VDD.n1573 VDD.n1572 23.1255
R27581 VDD.n1574 VDD.n1573 23.1255
R27582 VDD.n1566 VDD.n1565 23.1255
R27583 VDD.n1567 VDD.n1566 23.1255
R27584 VDD.n1563 VDD.n1562 23.1255
R27585 VDD.n1564 VDD.n1563 23.1255
R27586 VDD.n1556 VDD.n1555 23.1255
R27587 VDD.n1557 VDD.n1556 23.1255
R27588 VDD.n1553 VDD.n1552 23.1255
R27589 VDD.n1554 VDD.n1553 23.1255
R27590 VDD.n1546 VDD.n1545 23.1255
R27591 VDD.n1547 VDD.n1546 23.1255
R27592 VDD.n1543 VDD.n1542 23.1255
R27593 VDD.n1544 VDD.n1543 23.1255
R27594 VDD.n1536 VDD.n1535 23.1255
R27595 VDD.n1537 VDD.n1536 23.1255
R27596 VDD.n1533 VDD.n1532 23.1255
R27597 VDD.n1534 VDD.n1533 23.1255
R27598 VDD.n1526 VDD.n1525 23.1255
R27599 VDD.n1527 VDD.n1526 23.1255
R27600 VDD.n1523 VDD.n1522 23.1255
R27601 VDD.n1524 VDD.n1523 23.1255
R27602 VDD.n1516 VDD.n1515 23.1255
R27603 VDD.n1517 VDD.n1516 23.1255
R27604 VDD.n1506 VDD.n1505 23.1255
R27605 VDD.n1507 VDD.n1506 23.1255
R27606 VDD.n1499 VDD.n1498 23.1255
R27607 VDD.n1500 VDD.n1499 23.1255
R27608 VDD.n1496 VDD.n1495 23.1255
R27609 VDD.n1497 VDD.n1496 23.1255
R27610 VDD.n1489 VDD.n1488 23.1255
R27611 VDD.n1490 VDD.n1489 23.1255
R27612 VDD.n1486 VDD.n1485 23.1255
R27613 VDD.n1487 VDD.n1486 23.1255
R27614 VDD.n1479 VDD.n1478 23.1255
R27615 VDD.n1480 VDD.n1479 23.1255
R27616 VDD.n1476 VDD.n1475 23.1255
R27617 VDD.n1477 VDD.n1476 23.1255
R27618 VDD.n1469 VDD.n1468 23.1255
R27619 VDD.n1470 VDD.n1469 23.1255
R27620 VDD.n1466 VDD.n1465 23.1255
R27621 VDD.n1467 VDD.n1466 23.1255
R27622 VDD.n1459 VDD.n1458 23.1255
R27623 VDD.n1460 VDD.n1459 23.1255
R27624 VDD.n1577 VDD.n1576 23.1255
R27625 VDD.n1576 VDD.n1575 23.1255
R27626 VDD.n1326 VDD.n1322 23.1255
R27627 VDD.n1072 VDD.n1068 23.1255
R27628 VDD.n1314 VDD.n1068 23.1255
R27629 VDD.n1308 VDD.n1078 23.1255
R27630 VDD.n1308 VDD.n1307 23.1255
R27631 VDD.n1083 VDD.n1079 23.1255
R27632 VDD.n1304 VDD.n1079 23.1255
R27633 VDD.n1298 VDD.n1088 23.1255
R27634 VDD.n1298 VDD.n1297 23.1255
R27635 VDD.n1093 VDD.n1089 23.1255
R27636 VDD.n1294 VDD.n1089 23.1255
R27637 VDD.n1288 VDD.n1101 23.1255
R27638 VDD.n1288 VDD.n1287 23.1255
R27639 VDD.n1106 VDD.n1102 23.1255
R27640 VDD.n1284 VDD.n1102 23.1255
R27641 VDD.n1278 VDD.n1112 23.1255
R27642 VDD.n1278 VDD.n1277 23.1255
R27643 VDD.n1117 VDD.n1113 23.1255
R27644 VDD.n1274 VDD.n1113 23.1255
R27645 VDD.n1268 VDD.n1122 23.1255
R27646 VDD.n1268 VDD.n1267 23.1255
R27647 VDD.n1127 VDD.n1123 23.1255
R27648 VDD.n1264 VDD.n1123 23.1255
R27649 VDD.n1258 VDD.n1135 23.1255
R27650 VDD.n1258 VDD.n1257 23.1255
R27651 VDD.n1253 VDD.n1252 23.1255
R27652 VDD.n1254 VDD.n1253 23.1255
R27653 VDD.n1250 VDD.n1249 23.1255
R27654 VDD.n1249 VDD.n1248 23.1255
R27655 VDD.n1143 VDD.n1139 23.1255
R27656 VDD.n1247 VDD.n1139 23.1255
R27657 VDD.n1241 VDD.n1150 23.1255
R27658 VDD.n1241 VDD.n1240 23.1255
R27659 VDD.n1155 VDD.n1151 23.1255
R27660 VDD.n1237 VDD.n1151 23.1255
R27661 VDD.n1231 VDD.n1163 23.1255
R27662 VDD.n1231 VDD.n1230 23.1255
R27663 VDD.n1168 VDD.n1164 23.1255
R27664 VDD.n1227 VDD.n1164 23.1255
R27665 VDD.n1221 VDD.n1174 23.1255
R27666 VDD.n1221 VDD.n1220 23.1255
R27667 VDD.n1179 VDD.n1175 23.1255
R27668 VDD.n1217 VDD.n1175 23.1255
R27669 VDD.n1211 VDD.n1184 23.1255
R27670 VDD.n1211 VDD.n1210 23.1255
R27671 VDD.n1189 VDD.n1185 23.1255
R27672 VDD.n1207 VDD.n1185 23.1255
R27673 VDD.n1201 VDD.n1197 23.1255
R27674 VDD.n1201 VDD.n1200 23.1255
R27675 VDD.n1313 VDD.n1312 23.1255
R27676 VDD.n1314 VDD.n1313 23.1255
R27677 VDD.n1306 VDD.n1305 23.1255
R27678 VDD.n1307 VDD.n1306 23.1255
R27679 VDD.n1303 VDD.n1302 23.1255
R27680 VDD.n1304 VDD.n1303 23.1255
R27681 VDD.n1296 VDD.n1295 23.1255
R27682 VDD.n1297 VDD.n1296 23.1255
R27683 VDD.n1293 VDD.n1292 23.1255
R27684 VDD.n1294 VDD.n1293 23.1255
R27685 VDD.n1286 VDD.n1285 23.1255
R27686 VDD.n1287 VDD.n1286 23.1255
R27687 VDD.n1283 VDD.n1282 23.1255
R27688 VDD.n1284 VDD.n1283 23.1255
R27689 VDD.n1276 VDD.n1275 23.1255
R27690 VDD.n1277 VDD.n1276 23.1255
R27691 VDD.n1273 VDD.n1272 23.1255
R27692 VDD.n1274 VDD.n1273 23.1255
R27693 VDD.n1266 VDD.n1265 23.1255
R27694 VDD.n1267 VDD.n1266 23.1255
R27695 VDD.n1263 VDD.n1262 23.1255
R27696 VDD.n1264 VDD.n1263 23.1255
R27697 VDD.n1256 VDD.n1255 23.1255
R27698 VDD.n1257 VDD.n1256 23.1255
R27699 VDD.n1246 VDD.n1245 23.1255
R27700 VDD.n1247 VDD.n1246 23.1255
R27701 VDD.n1239 VDD.n1238 23.1255
R27702 VDD.n1240 VDD.n1239 23.1255
R27703 VDD.n1236 VDD.n1235 23.1255
R27704 VDD.n1237 VDD.n1236 23.1255
R27705 VDD.n1229 VDD.n1228 23.1255
R27706 VDD.n1230 VDD.n1229 23.1255
R27707 VDD.n1226 VDD.n1225 23.1255
R27708 VDD.n1227 VDD.n1226 23.1255
R27709 VDD.n1219 VDD.n1218 23.1255
R27710 VDD.n1220 VDD.n1219 23.1255
R27711 VDD.n1216 VDD.n1215 23.1255
R27712 VDD.n1217 VDD.n1216 23.1255
R27713 VDD.n1209 VDD.n1208 23.1255
R27714 VDD.n1210 VDD.n1209 23.1255
R27715 VDD.n1206 VDD.n1205 23.1255
R27716 VDD.n1207 VDD.n1206 23.1255
R27717 VDD.n1199 VDD.n1198 23.1255
R27718 VDD.n1200 VDD.n1199 23.1255
R27719 VDD.n1317 VDD.n1316 23.1255
R27720 VDD.n1316 VDD.n1315 23.1255
R27721 VDD.n1066 VDD.n1062 23.1255
R27722 VDD.n812 VDD.n808 23.1255
R27723 VDD.n1054 VDD.n808 23.1255
R27724 VDD.n1048 VDD.n818 23.1255
R27725 VDD.n1048 VDD.n1047 23.1255
R27726 VDD.n823 VDD.n819 23.1255
R27727 VDD.n1044 VDD.n819 23.1255
R27728 VDD.n1038 VDD.n828 23.1255
R27729 VDD.n1038 VDD.n1037 23.1255
R27730 VDD.n833 VDD.n829 23.1255
R27731 VDD.n1034 VDD.n829 23.1255
R27732 VDD.n1028 VDD.n841 23.1255
R27733 VDD.n1028 VDD.n1027 23.1255
R27734 VDD.n846 VDD.n842 23.1255
R27735 VDD.n1024 VDD.n842 23.1255
R27736 VDD.n1018 VDD.n852 23.1255
R27737 VDD.n1018 VDD.n1017 23.1255
R27738 VDD.n857 VDD.n853 23.1255
R27739 VDD.n1014 VDD.n853 23.1255
R27740 VDD.n1008 VDD.n862 23.1255
R27741 VDD.n1008 VDD.n1007 23.1255
R27742 VDD.n867 VDD.n863 23.1255
R27743 VDD.n1004 VDD.n863 23.1255
R27744 VDD.n998 VDD.n875 23.1255
R27745 VDD.n998 VDD.n997 23.1255
R27746 VDD.n993 VDD.n992 23.1255
R27747 VDD.n994 VDD.n993 23.1255
R27748 VDD.n990 VDD.n989 23.1255
R27749 VDD.n989 VDD.n988 23.1255
R27750 VDD.n883 VDD.n879 23.1255
R27751 VDD.n987 VDD.n879 23.1255
R27752 VDD.n981 VDD.n890 23.1255
R27753 VDD.n981 VDD.n980 23.1255
R27754 VDD.n895 VDD.n891 23.1255
R27755 VDD.n977 VDD.n891 23.1255
R27756 VDD.n971 VDD.n903 23.1255
R27757 VDD.n971 VDD.n970 23.1255
R27758 VDD.n908 VDD.n904 23.1255
R27759 VDD.n967 VDD.n904 23.1255
R27760 VDD.n961 VDD.n914 23.1255
R27761 VDD.n961 VDD.n960 23.1255
R27762 VDD.n919 VDD.n915 23.1255
R27763 VDD.n957 VDD.n915 23.1255
R27764 VDD.n951 VDD.n924 23.1255
R27765 VDD.n951 VDD.n950 23.1255
R27766 VDD.n929 VDD.n925 23.1255
R27767 VDD.n947 VDD.n925 23.1255
R27768 VDD.n941 VDD.n937 23.1255
R27769 VDD.n941 VDD.n940 23.1255
R27770 VDD.n1053 VDD.n1052 23.1255
R27771 VDD.n1054 VDD.n1053 23.1255
R27772 VDD.n1046 VDD.n1045 23.1255
R27773 VDD.n1047 VDD.n1046 23.1255
R27774 VDD.n1043 VDD.n1042 23.1255
R27775 VDD.n1044 VDD.n1043 23.1255
R27776 VDD.n1036 VDD.n1035 23.1255
R27777 VDD.n1037 VDD.n1036 23.1255
R27778 VDD.n1033 VDD.n1032 23.1255
R27779 VDD.n1034 VDD.n1033 23.1255
R27780 VDD.n1026 VDD.n1025 23.1255
R27781 VDD.n1027 VDD.n1026 23.1255
R27782 VDD.n1023 VDD.n1022 23.1255
R27783 VDD.n1024 VDD.n1023 23.1255
R27784 VDD.n1016 VDD.n1015 23.1255
R27785 VDD.n1017 VDD.n1016 23.1255
R27786 VDD.n1013 VDD.n1012 23.1255
R27787 VDD.n1014 VDD.n1013 23.1255
R27788 VDD.n1006 VDD.n1005 23.1255
R27789 VDD.n1007 VDD.n1006 23.1255
R27790 VDD.n1003 VDD.n1002 23.1255
R27791 VDD.n1004 VDD.n1003 23.1255
R27792 VDD.n996 VDD.n995 23.1255
R27793 VDD.n997 VDD.n996 23.1255
R27794 VDD.n986 VDD.n985 23.1255
R27795 VDD.n987 VDD.n986 23.1255
R27796 VDD.n979 VDD.n978 23.1255
R27797 VDD.n980 VDD.n979 23.1255
R27798 VDD.n976 VDD.n975 23.1255
R27799 VDD.n977 VDD.n976 23.1255
R27800 VDD.n969 VDD.n968 23.1255
R27801 VDD.n970 VDD.n969 23.1255
R27802 VDD.n966 VDD.n965 23.1255
R27803 VDD.n967 VDD.n966 23.1255
R27804 VDD.n959 VDD.n958 23.1255
R27805 VDD.n960 VDD.n959 23.1255
R27806 VDD.n956 VDD.n955 23.1255
R27807 VDD.n957 VDD.n956 23.1255
R27808 VDD.n949 VDD.n948 23.1255
R27809 VDD.n950 VDD.n949 23.1255
R27810 VDD.n946 VDD.n945 23.1255
R27811 VDD.n947 VDD.n946 23.1255
R27812 VDD.n939 VDD.n938 23.1255
R27813 VDD.n940 VDD.n939 23.1255
R27814 VDD.n1057 VDD.n1056 23.1255
R27815 VDD.n1056 VDD.n1055 23.1255
R27816 VDD.n806 VDD.n802 23.1255
R27817 VDD.n552 VDD.n548 23.1255
R27818 VDD.n794 VDD.n548 23.1255
R27819 VDD.n788 VDD.n558 23.1255
R27820 VDD.n788 VDD.n787 23.1255
R27821 VDD.n563 VDD.n559 23.1255
R27822 VDD.n784 VDD.n559 23.1255
R27823 VDD.n778 VDD.n568 23.1255
R27824 VDD.n778 VDD.n777 23.1255
R27825 VDD.n573 VDD.n569 23.1255
R27826 VDD.n774 VDD.n569 23.1255
R27827 VDD.n768 VDD.n581 23.1255
R27828 VDD.n768 VDD.n767 23.1255
R27829 VDD.n586 VDD.n582 23.1255
R27830 VDD.n764 VDD.n582 23.1255
R27831 VDD.n758 VDD.n592 23.1255
R27832 VDD.n758 VDD.n757 23.1255
R27833 VDD.n597 VDD.n593 23.1255
R27834 VDD.n754 VDD.n593 23.1255
R27835 VDD.n748 VDD.n602 23.1255
R27836 VDD.n748 VDD.n747 23.1255
R27837 VDD.n607 VDD.n603 23.1255
R27838 VDD.n744 VDD.n603 23.1255
R27839 VDD.n738 VDD.n615 23.1255
R27840 VDD.n738 VDD.n737 23.1255
R27841 VDD.n733 VDD.n732 23.1255
R27842 VDD.n734 VDD.n733 23.1255
R27843 VDD.n730 VDD.n729 23.1255
R27844 VDD.n729 VDD.n728 23.1255
R27845 VDD.n623 VDD.n619 23.1255
R27846 VDD.n727 VDD.n619 23.1255
R27847 VDD.n721 VDD.n630 23.1255
R27848 VDD.n721 VDD.n720 23.1255
R27849 VDD.n635 VDD.n631 23.1255
R27850 VDD.n717 VDD.n631 23.1255
R27851 VDD.n711 VDD.n643 23.1255
R27852 VDD.n711 VDD.n710 23.1255
R27853 VDD.n648 VDD.n644 23.1255
R27854 VDD.n707 VDD.n644 23.1255
R27855 VDD.n701 VDD.n654 23.1255
R27856 VDD.n701 VDD.n700 23.1255
R27857 VDD.n659 VDD.n655 23.1255
R27858 VDD.n697 VDD.n655 23.1255
R27859 VDD.n691 VDD.n664 23.1255
R27860 VDD.n691 VDD.n690 23.1255
R27861 VDD.n669 VDD.n665 23.1255
R27862 VDD.n687 VDD.n665 23.1255
R27863 VDD.n681 VDD.n677 23.1255
R27864 VDD.n681 VDD.n680 23.1255
R27865 VDD.n793 VDD.n792 23.1255
R27866 VDD.n794 VDD.n793 23.1255
R27867 VDD.n786 VDD.n785 23.1255
R27868 VDD.n787 VDD.n786 23.1255
R27869 VDD.n783 VDD.n782 23.1255
R27870 VDD.n784 VDD.n783 23.1255
R27871 VDD.n776 VDD.n775 23.1255
R27872 VDD.n777 VDD.n776 23.1255
R27873 VDD.n773 VDD.n772 23.1255
R27874 VDD.n774 VDD.n773 23.1255
R27875 VDD.n766 VDD.n765 23.1255
R27876 VDD.n767 VDD.n766 23.1255
R27877 VDD.n763 VDD.n762 23.1255
R27878 VDD.n764 VDD.n763 23.1255
R27879 VDD.n756 VDD.n755 23.1255
R27880 VDD.n757 VDD.n756 23.1255
R27881 VDD.n753 VDD.n752 23.1255
R27882 VDD.n754 VDD.n753 23.1255
R27883 VDD.n746 VDD.n745 23.1255
R27884 VDD.n747 VDD.n746 23.1255
R27885 VDD.n743 VDD.n742 23.1255
R27886 VDD.n744 VDD.n743 23.1255
R27887 VDD.n736 VDD.n735 23.1255
R27888 VDD.n737 VDD.n736 23.1255
R27889 VDD.n726 VDD.n725 23.1255
R27890 VDD.n727 VDD.n726 23.1255
R27891 VDD.n719 VDD.n718 23.1255
R27892 VDD.n720 VDD.n719 23.1255
R27893 VDD.n716 VDD.n715 23.1255
R27894 VDD.n717 VDD.n716 23.1255
R27895 VDD.n709 VDD.n708 23.1255
R27896 VDD.n710 VDD.n709 23.1255
R27897 VDD.n706 VDD.n705 23.1255
R27898 VDD.n707 VDD.n706 23.1255
R27899 VDD.n699 VDD.n698 23.1255
R27900 VDD.n700 VDD.n699 23.1255
R27901 VDD.n696 VDD.n695 23.1255
R27902 VDD.n697 VDD.n696 23.1255
R27903 VDD.n689 VDD.n688 23.1255
R27904 VDD.n690 VDD.n689 23.1255
R27905 VDD.n686 VDD.n685 23.1255
R27906 VDD.n687 VDD.n686 23.1255
R27907 VDD.n679 VDD.n678 23.1255
R27908 VDD.n680 VDD.n679 23.1255
R27909 VDD.n797 VDD.n796 23.1255
R27910 VDD.n796 VDD.n795 23.1255
R27911 VDD.n546 VDD.n542 23.1255
R27912 VDD.n292 VDD.n288 23.1255
R27913 VDD.n534 VDD.n288 23.1255
R27914 VDD.n528 VDD.n298 23.1255
R27915 VDD.n528 VDD.n527 23.1255
R27916 VDD.n303 VDD.n299 23.1255
R27917 VDD.n524 VDD.n299 23.1255
R27918 VDD.n518 VDD.n308 23.1255
R27919 VDD.n518 VDD.n517 23.1255
R27920 VDD.n313 VDD.n309 23.1255
R27921 VDD.n514 VDD.n309 23.1255
R27922 VDD.n508 VDD.n321 23.1255
R27923 VDD.n508 VDD.n507 23.1255
R27924 VDD.n326 VDD.n322 23.1255
R27925 VDD.n504 VDD.n322 23.1255
R27926 VDD.n498 VDD.n332 23.1255
R27927 VDD.n498 VDD.n497 23.1255
R27928 VDD.n337 VDD.n333 23.1255
R27929 VDD.n494 VDD.n333 23.1255
R27930 VDD.n488 VDD.n342 23.1255
R27931 VDD.n488 VDD.n487 23.1255
R27932 VDD.n347 VDD.n343 23.1255
R27933 VDD.n484 VDD.n343 23.1255
R27934 VDD.n478 VDD.n355 23.1255
R27935 VDD.n478 VDD.n477 23.1255
R27936 VDD.n473 VDD.n472 23.1255
R27937 VDD.n474 VDD.n473 23.1255
R27938 VDD.n470 VDD.n469 23.1255
R27939 VDD.n469 VDD.n468 23.1255
R27940 VDD.n363 VDD.n359 23.1255
R27941 VDD.n467 VDD.n359 23.1255
R27942 VDD.n461 VDD.n370 23.1255
R27943 VDD.n461 VDD.n460 23.1255
R27944 VDD.n375 VDD.n371 23.1255
R27945 VDD.n457 VDD.n371 23.1255
R27946 VDD.n451 VDD.n383 23.1255
R27947 VDD.n451 VDD.n450 23.1255
R27948 VDD.n388 VDD.n384 23.1255
R27949 VDD.n447 VDD.n384 23.1255
R27950 VDD.n441 VDD.n394 23.1255
R27951 VDD.n441 VDD.n440 23.1255
R27952 VDD.n399 VDD.n395 23.1255
R27953 VDD.n437 VDD.n395 23.1255
R27954 VDD.n431 VDD.n404 23.1255
R27955 VDD.n431 VDD.n430 23.1255
R27956 VDD.n409 VDD.n405 23.1255
R27957 VDD.n427 VDD.n405 23.1255
R27958 VDD.n421 VDD.n417 23.1255
R27959 VDD.n421 VDD.n420 23.1255
R27960 VDD.n533 VDD.n532 23.1255
R27961 VDD.n534 VDD.n533 23.1255
R27962 VDD.n526 VDD.n525 23.1255
R27963 VDD.n527 VDD.n526 23.1255
R27964 VDD.n523 VDD.n522 23.1255
R27965 VDD.n524 VDD.n523 23.1255
R27966 VDD.n516 VDD.n515 23.1255
R27967 VDD.n517 VDD.n516 23.1255
R27968 VDD.n513 VDD.n512 23.1255
R27969 VDD.n514 VDD.n513 23.1255
R27970 VDD.n506 VDD.n505 23.1255
R27971 VDD.n507 VDD.n506 23.1255
R27972 VDD.n503 VDD.n502 23.1255
R27973 VDD.n504 VDD.n503 23.1255
R27974 VDD.n496 VDD.n495 23.1255
R27975 VDD.n497 VDD.n496 23.1255
R27976 VDD.n493 VDD.n492 23.1255
R27977 VDD.n494 VDD.n493 23.1255
R27978 VDD.n486 VDD.n485 23.1255
R27979 VDD.n487 VDD.n486 23.1255
R27980 VDD.n483 VDD.n482 23.1255
R27981 VDD.n484 VDD.n483 23.1255
R27982 VDD.n476 VDD.n475 23.1255
R27983 VDD.n477 VDD.n476 23.1255
R27984 VDD.n466 VDD.n465 23.1255
R27985 VDD.n467 VDD.n466 23.1255
R27986 VDD.n459 VDD.n458 23.1255
R27987 VDD.n460 VDD.n459 23.1255
R27988 VDD.n456 VDD.n455 23.1255
R27989 VDD.n457 VDD.n456 23.1255
R27990 VDD.n449 VDD.n448 23.1255
R27991 VDD.n450 VDD.n449 23.1255
R27992 VDD.n446 VDD.n445 23.1255
R27993 VDD.n447 VDD.n446 23.1255
R27994 VDD.n439 VDD.n438 23.1255
R27995 VDD.n440 VDD.n439 23.1255
R27996 VDD.n436 VDD.n435 23.1255
R27997 VDD.n437 VDD.n436 23.1255
R27998 VDD.n429 VDD.n428 23.1255
R27999 VDD.n430 VDD.n429 23.1255
R28000 VDD.n426 VDD.n425 23.1255
R28001 VDD.n427 VDD.n426 23.1255
R28002 VDD.n419 VDD.n418 23.1255
R28003 VDD.n420 VDD.n419 23.1255
R28004 VDD.n537 VDD.n536 23.1255
R28005 VDD.n536 VDD.n535 23.1255
R28006 VDD.n286 VDD.n282 23.1255
R28007 VDD.n107 VDD.n106 23.1255
R28008 VDD.n108 VDD.n107 23.1255
R28009 VDD.n104 VDD.n103 23.1255
R28010 VDD.n111 VDD.n110 23.1255
R28011 VDD.n110 VDD.n109 23.1255
R28012 VDD.n96 VDD.n92 23.1255
R28013 VDD.n128 VDD.n127 23.1255
R28014 VDD.n129 VDD.n128 23.1255
R28015 VDD.n125 VDD.n124 23.1255
R28016 VDD.n124 VDD.n123 23.1255
R28017 VDD.n121 VDD.n120 23.1255
R28018 VDD.n122 VDD.n121 23.1255
R28019 VDD.n118 VDD.n117 23.1255
R28020 VDD.n132 VDD.n131 23.1255
R28021 VDD.n131 VDD.n130 23.1255
R28022 VDD.n80 VDD.n76 23.1255
R28023 VDD.n142 VDD.n141 23.1255
R28024 VDD.n143 VDD.n142 23.1255
R28025 VDD.n139 VDD.n138 23.1255
R28026 VDD.n146 VDD.n145 23.1255
R28027 VDD.n145 VDD.n144 23.1255
R28028 VDD.n71 VDD.n67 23.1255
R28029 VDD.n163 VDD.n162 23.1255
R28030 VDD.n164 VDD.n163 23.1255
R28031 VDD.n160 VDD.n159 23.1255
R28032 VDD.n159 VDD.n158 23.1255
R28033 VDD.n156 VDD.n155 23.1255
R28034 VDD.n157 VDD.n156 23.1255
R28035 VDD.n153 VDD.n152 23.1255
R28036 VDD.n167 VDD.n166 23.1255
R28037 VDD.n166 VDD.n165 23.1255
R28038 VDD.n55 VDD.n51 23.1255
R28039 VDD.n177 VDD.n176 23.1255
R28040 VDD.n178 VDD.n177 23.1255
R28041 VDD.n174 VDD.n173 23.1255
R28042 VDD.n181 VDD.n180 23.1255
R28043 VDD.n180 VDD.n179 23.1255
R28044 VDD.n46 VDD.n42 23.1255
R28045 VDD.n198 VDD.n197 23.1255
R28046 VDD.n199 VDD.n198 23.1255
R28047 VDD.n195 VDD.n194 23.1255
R28048 VDD.n194 VDD.n193 23.1255
R28049 VDD.n191 VDD.n190 23.1255
R28050 VDD.n192 VDD.n191 23.1255
R28051 VDD.n188 VDD.n187 23.1255
R28052 VDD.n202 VDD.n201 23.1255
R28053 VDD.n201 VDD.n200 23.1255
R28054 VDD.n30 VDD.n26 23.1255
R28055 VDD.n212 VDD.n211 23.1255
R28056 VDD.n213 VDD.n212 23.1255
R28057 VDD.n209 VDD.n208 23.1255
R28058 VDD.n216 VDD.n215 23.1255
R28059 VDD.n215 VDD.n214 23.1255
R28060 VDD.n21 VDD.n17 23.1255
R28061 VDD.n233 VDD.n232 23.1255
R28062 VDD.n234 VDD.n233 23.1255
R28063 VDD.n230 VDD.n229 23.1255
R28064 VDD.n229 VDD.n228 23.1255
R28065 VDD.n226 VDD.n225 23.1255
R28066 VDD.n227 VDD.n226 23.1255
R28067 VDD.n223 VDD.n222 23.1255
R28068 VDD.n237 VDD.n236 23.1255
R28069 VDD.n236 VDD.n235 23.1255
R28070 VDD.n5 VDD.n1 23.1255
R28071 VDD.n7208 VDD.n7204 23.1255
R28072 VDD.n7450 VDD.n7204 23.1255
R28073 VDD.n7444 VDD.n7214 23.1255
R28074 VDD.n7444 VDD.n7443 23.1255
R28075 VDD.n7219 VDD.n7215 23.1255
R28076 VDD.n7440 VDD.n7215 23.1255
R28077 VDD.n7434 VDD.n7224 23.1255
R28078 VDD.n7434 VDD.n7433 23.1255
R28079 VDD.n7229 VDD.n7225 23.1255
R28080 VDD.n7430 VDD.n7225 23.1255
R28081 VDD.n7424 VDD.n7237 23.1255
R28082 VDD.n7424 VDD.n7423 23.1255
R28083 VDD.n7242 VDD.n7238 23.1255
R28084 VDD.n7420 VDD.n7238 23.1255
R28085 VDD.n7414 VDD.n7248 23.1255
R28086 VDD.n7414 VDD.n7413 23.1255
R28087 VDD.n7253 VDD.n7249 23.1255
R28088 VDD.n7410 VDD.n7249 23.1255
R28089 VDD.n7404 VDD.n7258 23.1255
R28090 VDD.n7404 VDD.n7403 23.1255
R28091 VDD.n7263 VDD.n7259 23.1255
R28092 VDD.n7400 VDD.n7259 23.1255
R28093 VDD.n7394 VDD.n7271 23.1255
R28094 VDD.n7394 VDD.n7393 23.1255
R28095 VDD.n7389 VDD.n7388 23.1255
R28096 VDD.n7390 VDD.n7389 23.1255
R28097 VDD.n7386 VDD.n7385 23.1255
R28098 VDD.n7385 VDD.n7384 23.1255
R28099 VDD.n7279 VDD.n7275 23.1255
R28100 VDD.n7383 VDD.n7275 23.1255
R28101 VDD.n7377 VDD.n7286 23.1255
R28102 VDD.n7377 VDD.n7376 23.1255
R28103 VDD.n7291 VDD.n7287 23.1255
R28104 VDD.n7373 VDD.n7287 23.1255
R28105 VDD.n7367 VDD.n7299 23.1255
R28106 VDD.n7367 VDD.n7366 23.1255
R28107 VDD.n7304 VDD.n7300 23.1255
R28108 VDD.n7363 VDD.n7300 23.1255
R28109 VDD.n7357 VDD.n7310 23.1255
R28110 VDD.n7357 VDD.n7356 23.1255
R28111 VDD.n7315 VDD.n7311 23.1255
R28112 VDD.n7353 VDD.n7311 23.1255
R28113 VDD.n7347 VDD.n7320 23.1255
R28114 VDD.n7347 VDD.n7346 23.1255
R28115 VDD.n7325 VDD.n7321 23.1255
R28116 VDD.n7343 VDD.n7321 23.1255
R28117 VDD.n7337 VDD.n7333 23.1255
R28118 VDD.n7337 VDD.n7336 23.1255
R28119 VDD.n7449 VDD.n7448 23.1255
R28120 VDD.n7450 VDD.n7449 23.1255
R28121 VDD.n7442 VDD.n7441 23.1255
R28122 VDD.n7443 VDD.n7442 23.1255
R28123 VDD.n7439 VDD.n7438 23.1255
R28124 VDD.n7440 VDD.n7439 23.1255
R28125 VDD.n7432 VDD.n7431 23.1255
R28126 VDD.n7433 VDD.n7432 23.1255
R28127 VDD.n7429 VDD.n7428 23.1255
R28128 VDD.n7430 VDD.n7429 23.1255
R28129 VDD.n7422 VDD.n7421 23.1255
R28130 VDD.n7423 VDD.n7422 23.1255
R28131 VDD.n7419 VDD.n7418 23.1255
R28132 VDD.n7420 VDD.n7419 23.1255
R28133 VDD.n7412 VDD.n7411 23.1255
R28134 VDD.n7413 VDD.n7412 23.1255
R28135 VDD.n7409 VDD.n7408 23.1255
R28136 VDD.n7410 VDD.n7409 23.1255
R28137 VDD.n7402 VDD.n7401 23.1255
R28138 VDD.n7403 VDD.n7402 23.1255
R28139 VDD.n7399 VDD.n7398 23.1255
R28140 VDD.n7400 VDD.n7399 23.1255
R28141 VDD.n7392 VDD.n7391 23.1255
R28142 VDD.n7393 VDD.n7392 23.1255
R28143 VDD.n7382 VDD.n7381 23.1255
R28144 VDD.n7383 VDD.n7382 23.1255
R28145 VDD.n7375 VDD.n7374 23.1255
R28146 VDD.n7376 VDD.n7375 23.1255
R28147 VDD.n7372 VDD.n7371 23.1255
R28148 VDD.n7373 VDD.n7372 23.1255
R28149 VDD.n7365 VDD.n7364 23.1255
R28150 VDD.n7366 VDD.n7365 23.1255
R28151 VDD.n7362 VDD.n7361 23.1255
R28152 VDD.n7363 VDD.n7362 23.1255
R28153 VDD.n7355 VDD.n7354 23.1255
R28154 VDD.n7356 VDD.n7355 23.1255
R28155 VDD.n7352 VDD.n7351 23.1255
R28156 VDD.n7353 VDD.n7352 23.1255
R28157 VDD.n7345 VDD.n7344 23.1255
R28158 VDD.n7346 VDD.n7345 23.1255
R28159 VDD.n7342 VDD.n7341 23.1255
R28160 VDD.n7343 VDD.n7342 23.1255
R28161 VDD.n7335 VDD.n7334 23.1255
R28162 VDD.n7336 VDD.n7335 23.1255
R28163 VDD.n7453 VDD.n7452 23.1255
R28164 VDD.n7452 VDD.n7451 23.1255
R28165 VDD.n7202 VDD.n7198 23.1255
R28166 VDD.n1852 VDD.n1848 23.1255
R28167 VDD.n7190 VDD.n1848 23.1255
R28168 VDD.n7184 VDD.n1858 23.1255
R28169 VDD.n7184 VDD.n7183 23.1255
R28170 VDD.n1863 VDD.n1859 23.1255
R28171 VDD.n7180 VDD.n1859 23.1255
R28172 VDD.n7174 VDD.n1868 23.1255
R28173 VDD.n7174 VDD.n7173 23.1255
R28174 VDD.n1873 VDD.n1869 23.1255
R28175 VDD.n7170 VDD.n1869 23.1255
R28176 VDD.n7164 VDD.n1881 23.1255
R28177 VDD.n7164 VDD.n7163 23.1255
R28178 VDD.n1886 VDD.n1882 23.1255
R28179 VDD.n7160 VDD.n1882 23.1255
R28180 VDD.n7154 VDD.n1893 23.1255
R28181 VDD.n7154 VDD.n7153 23.1255
R28182 VDD.n1898 VDD.n1894 23.1255
R28183 VDD.n7150 VDD.n1894 23.1255
R28184 VDD.n1912 VDD.n1911 23.1255
R28185 VDD.n1915 VDD.n1912 23.1255
R28186 VDD.n1917 VDD.n1907 23.1255
R28187 VDD.n1916 VDD.n1907 23.1255
R28188 VDD.n1918 VDD.n1908 23.1255
R28189 VDD.n7134 VDD.n1908 23.1255
R28190 VDD.n7132 VDD.n7131 23.1255
R28191 VDD.n7133 VDD.n7132 23.1255
R28192 VDD.n7129 VDD.n7128 23.1255
R28193 VDD.n7128 VDD.n7127 23.1255
R28194 VDD.n1928 VDD.n1924 23.1255
R28195 VDD.n7126 VDD.n1924 23.1255
R28196 VDD.n7120 VDD.n1935 23.1255
R28197 VDD.n7120 VDD.n7119 23.1255
R28198 VDD.n1940 VDD.n1936 23.1255
R28199 VDD.n7116 VDD.n1936 23.1255
R28200 VDD.n7110 VDD.n1948 23.1255
R28201 VDD.n7110 VDD.n7109 23.1255
R28202 VDD.n1953 VDD.n1949 23.1255
R28203 VDD.n7106 VDD.n1949 23.1255
R28204 VDD.n7100 VDD.n1959 23.1255
R28205 VDD.n7100 VDD.n7099 23.1255
R28206 VDD.n1964 VDD.n1960 23.1255
R28207 VDD.n7096 VDD.n1960 23.1255
R28208 VDD.n7090 VDD.n1969 23.1255
R28209 VDD.n7090 VDD.n7089 23.1255
R28210 VDD.n1974 VDD.n1970 23.1255
R28211 VDD.n7086 VDD.n1970 23.1255
R28212 VDD.n7080 VDD.n7076 23.1255
R28213 VDD.n7080 VDD.n7079 23.1255
R28214 VDD.n1846 VDD.n1842 23.1255
R28215 VDD.n7193 VDD.n7192 23.1255
R28216 VDD.n7192 VDD.n7191 23.1255
R28217 VDD.n7189 VDD.n7188 23.1255
R28218 VDD.n7190 VDD.n7189 23.1255
R28219 VDD.n7182 VDD.n7181 23.1255
R28220 VDD.n7183 VDD.n7182 23.1255
R28221 VDD.n7179 VDD.n7178 23.1255
R28222 VDD.n7180 VDD.n7179 23.1255
R28223 VDD.n7172 VDD.n7171 23.1255
R28224 VDD.n7173 VDD.n7172 23.1255
R28225 VDD.n7169 VDD.n7168 23.1255
R28226 VDD.n7170 VDD.n7169 23.1255
R28227 VDD.n7162 VDD.n7161 23.1255
R28228 VDD.n7163 VDD.n7162 23.1255
R28229 VDD.n7159 VDD.n7158 23.1255
R28230 VDD.n7160 VDD.n7159 23.1255
R28231 VDD.n7152 VDD.n7151 23.1255
R28232 VDD.n7153 VDD.n7152 23.1255
R28233 VDD.n7137 VDD.n7135 23.1255
R28234 VDD.n7135 VDD.n1916 23.1255
R28235 VDD.n7138 VDD.n7136 23.1255
R28236 VDD.n7136 VDD.n7134 23.1255
R28237 VDD.n7125 VDD.n7124 23.1255
R28238 VDD.n7126 VDD.n7125 23.1255
R28239 VDD.n7118 VDD.n7117 23.1255
R28240 VDD.n7119 VDD.n7118 23.1255
R28241 VDD.n7115 VDD.n7114 23.1255
R28242 VDD.n7116 VDD.n7115 23.1255
R28243 VDD.n7108 VDD.n7107 23.1255
R28244 VDD.n7109 VDD.n7108 23.1255
R28245 VDD.n7105 VDD.n7104 23.1255
R28246 VDD.n7106 VDD.n7105 23.1255
R28247 VDD.n7098 VDD.n7097 23.1255
R28248 VDD.n7099 VDD.n7098 23.1255
R28249 VDD.n7095 VDD.n7094 23.1255
R28250 VDD.n7096 VDD.n7095 23.1255
R28251 VDD.n7088 VDD.n7087 23.1255
R28252 VDD.n7089 VDD.n7088 23.1255
R28253 VDD.n7085 VDD.n7084 23.1255
R28254 VDD.n7086 VDD.n7085 23.1255
R28255 VDD.n7078 VDD.n7077 23.1255
R28256 VDD.n7079 VDD.n7078 23.1255
R28257 VDD.n1914 VDD.n1913 23.1255
R28258 VDD.n1915 VDD.n1914 23.1255
R28259 VDD.n7149 VDD.n7148 23.1255
R28260 VDD.n7150 VDD.n7149 23.1255
R28261 VDD.n6941 VDD.n6940 23.1255
R28262 VDD.n6942 VDD.n6941 23.1255
R28263 VDD.n6938 VDD.n6937 23.1255
R28264 VDD.n6945 VDD.n6944 23.1255
R28265 VDD.n6944 VDD.n6943 23.1255
R28266 VDD.n6930 VDD.n6926 23.1255
R28267 VDD.n6962 VDD.n6961 23.1255
R28268 VDD.n6963 VDD.n6962 23.1255
R28269 VDD.n6959 VDD.n6958 23.1255
R28270 VDD.n6958 VDD.n6957 23.1255
R28271 VDD.n6955 VDD.n6954 23.1255
R28272 VDD.n6956 VDD.n6955 23.1255
R28273 VDD.n6952 VDD.n6951 23.1255
R28274 VDD.n6966 VDD.n6965 23.1255
R28275 VDD.n6965 VDD.n6964 23.1255
R28276 VDD.n6914 VDD.n6910 23.1255
R28277 VDD.n6976 VDD.n6975 23.1255
R28278 VDD.n6977 VDD.n6976 23.1255
R28279 VDD.n6973 VDD.n6972 23.1255
R28280 VDD.n6980 VDD.n6979 23.1255
R28281 VDD.n6979 VDD.n6978 23.1255
R28282 VDD.n6905 VDD.n6901 23.1255
R28283 VDD.n6997 VDD.n6996 23.1255
R28284 VDD.n6998 VDD.n6997 23.1255
R28285 VDD.n6994 VDD.n6993 23.1255
R28286 VDD.n6993 VDD.n6992 23.1255
R28287 VDD.n6990 VDD.n6989 23.1255
R28288 VDD.n6991 VDD.n6990 23.1255
R28289 VDD.n6987 VDD.n6986 23.1255
R28290 VDD.n7001 VDD.n7000 23.1255
R28291 VDD.n7000 VDD.n6999 23.1255
R28292 VDD.n6889 VDD.n6885 23.1255
R28293 VDD.n7011 VDD.n7010 23.1255
R28294 VDD.n7012 VDD.n7011 23.1255
R28295 VDD.n7008 VDD.n7007 23.1255
R28296 VDD.n7015 VDD.n7014 23.1255
R28297 VDD.n7014 VDD.n7013 23.1255
R28298 VDD.n6880 VDD.n6876 23.1255
R28299 VDD.n7032 VDD.n7031 23.1255
R28300 VDD.n7033 VDD.n7032 23.1255
R28301 VDD.n7029 VDD.n7028 23.1255
R28302 VDD.n7028 VDD.n7027 23.1255
R28303 VDD.n7025 VDD.n7024 23.1255
R28304 VDD.n7026 VDD.n7025 23.1255
R28305 VDD.n7022 VDD.n7021 23.1255
R28306 VDD.n7036 VDD.n7035 23.1255
R28307 VDD.n7035 VDD.n7034 23.1255
R28308 VDD.n6864 VDD.n6860 23.1255
R28309 VDD.n7046 VDD.n7045 23.1255
R28310 VDD.n7047 VDD.n7046 23.1255
R28311 VDD.n7043 VDD.n7042 23.1255
R28312 VDD.n7050 VDD.n7049 23.1255
R28313 VDD.n7049 VDD.n7048 23.1255
R28314 VDD.n6855 VDD.n6851 23.1255
R28315 VDD.n6833 VDD.n6831 23.1255
R28316 VDD.n6846 VDD.n6833 23.1255
R28317 VDD.n6834 VDD.n6832 23.1255
R28318 VDD.n7062 VDD.n6834 23.1255
R28319 VDD.n7060 VDD.n7059 23.1255
R28320 VDD.n7061 VDD.n7060 23.1255
R28321 VDD.n7057 VDD.n7056 23.1255
R28322 VDD.n6844 VDD.n6843 23.1255
R28323 VDD.n6845 VDD.n6844 23.1255
R28324 VDD.n6841 VDD.n6840 23.1255
R28325 VDD.n5839 VDD.n5836 23.1255
R28326 VDD.n5838 VDD.n5836 23.1255
R28327 VDD.n5840 VDD.n5837 23.1255
R28328 VDD.n6079 VDD.n5837 23.1255
R28329 VDD.n5847 VDD.n5843 23.1255
R28330 VDD.n6078 VDD.n5843 23.1255
R28331 VDD.n6072 VDD.n5852 23.1255
R28332 VDD.n6072 VDD.n6071 23.1255
R28333 VDD.n5857 VDD.n5853 23.1255
R28334 VDD.n6068 VDD.n5853 23.1255
R28335 VDD.n6062 VDD.n5862 23.1255
R28336 VDD.n6062 VDD.n6061 23.1255
R28337 VDD.n5867 VDD.n5863 23.1255
R28338 VDD.n6058 VDD.n5863 23.1255
R28339 VDD.n6052 VDD.n5873 23.1255
R28340 VDD.n6052 VDD.n6051 23.1255
R28341 VDD.n5878 VDD.n5874 23.1255
R28342 VDD.n6048 VDD.n5874 23.1255
R28343 VDD.n6042 VDD.n5886 23.1255
R28344 VDD.n6042 VDD.n6041 23.1255
R28345 VDD.n6037 VDD.n6036 23.1255
R28346 VDD.n6038 VDD.n6037 23.1255
R28347 VDD.n6034 VDD.n6033 23.1255
R28348 VDD.n6033 VDD.n6032 23.1255
R28349 VDD.n5894 VDD.n5890 23.1255
R28350 VDD.n6031 VDD.n5890 23.1255
R28351 VDD.n6025 VDD.n5901 23.1255
R28352 VDD.n6025 VDD.n6024 23.1255
R28353 VDD.n5906 VDD.n5902 23.1255
R28354 VDD.n6021 VDD.n5902 23.1255
R28355 VDD.n6015 VDD.n5914 23.1255
R28356 VDD.n6015 VDD.n6014 23.1255
R28357 VDD.n5919 VDD.n5915 23.1255
R28358 VDD.n6011 VDD.n5915 23.1255
R28359 VDD.n6005 VDD.n5924 23.1255
R28360 VDD.n6005 VDD.n6004 23.1255
R28361 VDD.n5929 VDD.n5925 23.1255
R28362 VDD.n6001 VDD.n5925 23.1255
R28363 VDD.n5995 VDD.n5935 23.1255
R28364 VDD.n5995 VDD.n5994 23.1255
R28365 VDD.n5940 VDD.n5936 23.1255
R28366 VDD.n5991 VDD.n5936 23.1255
R28367 VDD.n5985 VDD.n5948 23.1255
R28368 VDD.n5985 VDD.n5984 23.1255
R28369 VDD.n5953 VDD.n5949 23.1255
R28370 VDD.n5981 VDD.n5949 23.1255
R28371 VDD.n5975 VDD.n5958 23.1255
R28372 VDD.n5975 VDD.n5974 23.1255
R28373 VDD.n6077 VDD.n6076 23.1255
R28374 VDD.n6078 VDD.n6077 23.1255
R28375 VDD.n6070 VDD.n6069 23.1255
R28376 VDD.n6071 VDD.n6070 23.1255
R28377 VDD.n6067 VDD.n6066 23.1255
R28378 VDD.n6068 VDD.n6067 23.1255
R28379 VDD.n6060 VDD.n6059 23.1255
R28380 VDD.n6061 VDD.n6060 23.1255
R28381 VDD.n6057 VDD.n6056 23.1255
R28382 VDD.n6058 VDD.n6057 23.1255
R28383 VDD.n6050 VDD.n6049 23.1255
R28384 VDD.n6051 VDD.n6050 23.1255
R28385 VDD.n6047 VDD.n6046 23.1255
R28386 VDD.n6048 VDD.n6047 23.1255
R28387 VDD.n6040 VDD.n6039 23.1255
R28388 VDD.n6041 VDD.n6040 23.1255
R28389 VDD.n6030 VDD.n6029 23.1255
R28390 VDD.n6031 VDD.n6030 23.1255
R28391 VDD.n6023 VDD.n6022 23.1255
R28392 VDD.n6024 VDD.n6023 23.1255
R28393 VDD.n6020 VDD.n6019 23.1255
R28394 VDD.n6021 VDD.n6020 23.1255
R28395 VDD.n6013 VDD.n6012 23.1255
R28396 VDD.n6014 VDD.n6013 23.1255
R28397 VDD.n6010 VDD.n6009 23.1255
R28398 VDD.n6011 VDD.n6010 23.1255
R28399 VDD.n6003 VDD.n6002 23.1255
R28400 VDD.n6004 VDD.n6003 23.1255
R28401 VDD.n6000 VDD.n5999 23.1255
R28402 VDD.n6001 VDD.n6000 23.1255
R28403 VDD.n5993 VDD.n5992 23.1255
R28404 VDD.n5994 VDD.n5993 23.1255
R28405 VDD.n5990 VDD.n5989 23.1255
R28406 VDD.n5991 VDD.n5990 23.1255
R28407 VDD.n5983 VDD.n5982 23.1255
R28408 VDD.n5984 VDD.n5983 23.1255
R28409 VDD.n5980 VDD.n5979 23.1255
R28410 VDD.n5981 VDD.n5980 23.1255
R28411 VDD.n5973 VDD.n5972 23.1255
R28412 VDD.n5974 VDD.n5973 23.1255
R28413 VDD.n5970 VDD.n5969 23.1255
R28414 VDD.n5971 VDD.n5970 23.1255
R28415 VDD.n5964 VDD.n5963 23.1255
R28416 VDD.n6083 VDD.n6081 23.1255
R28417 VDD.n6081 VDD.n6079 23.1255
R28418 VDD.n6082 VDD.n6080 23.1255
R28419 VDD.n6080 VDD.n5838 23.1255
R28420 VDD.n5703 VDD.n5700 23.1255
R28421 VDD.n5702 VDD.n5700 23.1255
R28422 VDD.n5704 VDD.n5701 23.1255
R28423 VDD.n6202 VDD.n5701 23.1255
R28424 VDD.n5711 VDD.n5707 23.1255
R28425 VDD.n6201 VDD.n5707 23.1255
R28426 VDD.n6195 VDD.n5716 23.1255
R28427 VDD.n6195 VDD.n6194 23.1255
R28428 VDD.n5721 VDD.n5717 23.1255
R28429 VDD.n6191 VDD.n5717 23.1255
R28430 VDD.n6185 VDD.n5726 23.1255
R28431 VDD.n6185 VDD.n6184 23.1255
R28432 VDD.n5731 VDD.n5727 23.1255
R28433 VDD.n6181 VDD.n5727 23.1255
R28434 VDD.n6175 VDD.n5737 23.1255
R28435 VDD.n6175 VDD.n6174 23.1255
R28436 VDD.n5742 VDD.n5738 23.1255
R28437 VDD.n6171 VDD.n5738 23.1255
R28438 VDD.n6165 VDD.n5750 23.1255
R28439 VDD.n6165 VDD.n6164 23.1255
R28440 VDD.n6160 VDD.n6159 23.1255
R28441 VDD.n6161 VDD.n6160 23.1255
R28442 VDD.n6157 VDD.n6156 23.1255
R28443 VDD.n6156 VDD.n6155 23.1255
R28444 VDD.n5758 VDD.n5754 23.1255
R28445 VDD.n6154 VDD.n5754 23.1255
R28446 VDD.n6148 VDD.n5765 23.1255
R28447 VDD.n6148 VDD.n6147 23.1255
R28448 VDD.n5770 VDD.n5766 23.1255
R28449 VDD.n6144 VDD.n5766 23.1255
R28450 VDD.n6138 VDD.n5778 23.1255
R28451 VDD.n6138 VDD.n6137 23.1255
R28452 VDD.n5783 VDD.n5779 23.1255
R28453 VDD.n6134 VDD.n5779 23.1255
R28454 VDD.n6128 VDD.n5788 23.1255
R28455 VDD.n6128 VDD.n6127 23.1255
R28456 VDD.n5793 VDD.n5789 23.1255
R28457 VDD.n6124 VDD.n5789 23.1255
R28458 VDD.n6118 VDD.n5799 23.1255
R28459 VDD.n6118 VDD.n6117 23.1255
R28460 VDD.n5804 VDD.n5800 23.1255
R28461 VDD.n6114 VDD.n5800 23.1255
R28462 VDD.n6108 VDD.n5812 23.1255
R28463 VDD.n6108 VDD.n6107 23.1255
R28464 VDD.n5817 VDD.n5813 23.1255
R28465 VDD.n6104 VDD.n5813 23.1255
R28466 VDD.n6098 VDD.n5822 23.1255
R28467 VDD.n6098 VDD.n6097 23.1255
R28468 VDD.n6200 VDD.n6199 23.1255
R28469 VDD.n6201 VDD.n6200 23.1255
R28470 VDD.n6193 VDD.n6192 23.1255
R28471 VDD.n6194 VDD.n6193 23.1255
R28472 VDD.n6190 VDD.n6189 23.1255
R28473 VDD.n6191 VDD.n6190 23.1255
R28474 VDD.n6183 VDD.n6182 23.1255
R28475 VDD.n6184 VDD.n6183 23.1255
R28476 VDD.n6180 VDD.n6179 23.1255
R28477 VDD.n6181 VDD.n6180 23.1255
R28478 VDD.n6173 VDD.n6172 23.1255
R28479 VDD.n6174 VDD.n6173 23.1255
R28480 VDD.n6170 VDD.n6169 23.1255
R28481 VDD.n6171 VDD.n6170 23.1255
R28482 VDD.n6163 VDD.n6162 23.1255
R28483 VDD.n6164 VDD.n6163 23.1255
R28484 VDD.n6153 VDD.n6152 23.1255
R28485 VDD.n6154 VDD.n6153 23.1255
R28486 VDD.n6146 VDD.n6145 23.1255
R28487 VDD.n6147 VDD.n6146 23.1255
R28488 VDD.n6143 VDD.n6142 23.1255
R28489 VDD.n6144 VDD.n6143 23.1255
R28490 VDD.n6136 VDD.n6135 23.1255
R28491 VDD.n6137 VDD.n6136 23.1255
R28492 VDD.n6133 VDD.n6132 23.1255
R28493 VDD.n6134 VDD.n6133 23.1255
R28494 VDD.n6126 VDD.n6125 23.1255
R28495 VDD.n6127 VDD.n6126 23.1255
R28496 VDD.n6123 VDD.n6122 23.1255
R28497 VDD.n6124 VDD.n6123 23.1255
R28498 VDD.n6116 VDD.n6115 23.1255
R28499 VDD.n6117 VDD.n6116 23.1255
R28500 VDD.n6113 VDD.n6112 23.1255
R28501 VDD.n6114 VDD.n6113 23.1255
R28502 VDD.n6106 VDD.n6105 23.1255
R28503 VDD.n6107 VDD.n6106 23.1255
R28504 VDD.n6103 VDD.n6102 23.1255
R28505 VDD.n6104 VDD.n6103 23.1255
R28506 VDD.n6096 VDD.n6095 23.1255
R28507 VDD.n6097 VDD.n6096 23.1255
R28508 VDD.n6093 VDD.n6092 23.1255
R28509 VDD.n6094 VDD.n6093 23.1255
R28510 VDD.n5828 VDD.n5827 23.1255
R28511 VDD.n6206 VDD.n6204 23.1255
R28512 VDD.n6204 VDD.n6202 23.1255
R28513 VDD.n6205 VDD.n6203 23.1255
R28514 VDD.n6203 VDD.n5702 23.1255
R28515 VDD.n5567 VDD.n5564 23.1255
R28516 VDD.n5566 VDD.n5564 23.1255
R28517 VDD.n5568 VDD.n5565 23.1255
R28518 VDD.n6325 VDD.n5565 23.1255
R28519 VDD.n5575 VDD.n5571 23.1255
R28520 VDD.n6324 VDD.n5571 23.1255
R28521 VDD.n6318 VDD.n5580 23.1255
R28522 VDD.n6318 VDD.n6317 23.1255
R28523 VDD.n5585 VDD.n5581 23.1255
R28524 VDD.n6314 VDD.n5581 23.1255
R28525 VDD.n6308 VDD.n5590 23.1255
R28526 VDD.n6308 VDD.n6307 23.1255
R28527 VDD.n5595 VDD.n5591 23.1255
R28528 VDD.n6304 VDD.n5591 23.1255
R28529 VDD.n6298 VDD.n5601 23.1255
R28530 VDD.n6298 VDD.n6297 23.1255
R28531 VDD.n5606 VDD.n5602 23.1255
R28532 VDD.n6294 VDD.n5602 23.1255
R28533 VDD.n6288 VDD.n5614 23.1255
R28534 VDD.n6288 VDD.n6287 23.1255
R28535 VDD.n6283 VDD.n6282 23.1255
R28536 VDD.n6284 VDD.n6283 23.1255
R28537 VDD.n6280 VDD.n6279 23.1255
R28538 VDD.n6279 VDD.n6278 23.1255
R28539 VDD.n5622 VDD.n5618 23.1255
R28540 VDD.n6277 VDD.n5618 23.1255
R28541 VDD.n6271 VDD.n5629 23.1255
R28542 VDD.n6271 VDD.n6270 23.1255
R28543 VDD.n5634 VDD.n5630 23.1255
R28544 VDD.n6267 VDD.n5630 23.1255
R28545 VDD.n6261 VDD.n5642 23.1255
R28546 VDD.n6261 VDD.n6260 23.1255
R28547 VDD.n5647 VDD.n5643 23.1255
R28548 VDD.n6257 VDD.n5643 23.1255
R28549 VDD.n6251 VDD.n5652 23.1255
R28550 VDD.n6251 VDD.n6250 23.1255
R28551 VDD.n5657 VDD.n5653 23.1255
R28552 VDD.n6247 VDD.n5653 23.1255
R28553 VDD.n6241 VDD.n5663 23.1255
R28554 VDD.n6241 VDD.n6240 23.1255
R28555 VDD.n5668 VDD.n5664 23.1255
R28556 VDD.n6237 VDD.n5664 23.1255
R28557 VDD.n6231 VDD.n5676 23.1255
R28558 VDD.n6231 VDD.n6230 23.1255
R28559 VDD.n5681 VDD.n5677 23.1255
R28560 VDD.n6227 VDD.n5677 23.1255
R28561 VDD.n6221 VDD.n5686 23.1255
R28562 VDD.n6221 VDD.n6220 23.1255
R28563 VDD.n6323 VDD.n6322 23.1255
R28564 VDD.n6324 VDD.n6323 23.1255
R28565 VDD.n6316 VDD.n6315 23.1255
R28566 VDD.n6317 VDD.n6316 23.1255
R28567 VDD.n6313 VDD.n6312 23.1255
R28568 VDD.n6314 VDD.n6313 23.1255
R28569 VDD.n6306 VDD.n6305 23.1255
R28570 VDD.n6307 VDD.n6306 23.1255
R28571 VDD.n6303 VDD.n6302 23.1255
R28572 VDD.n6304 VDD.n6303 23.1255
R28573 VDD.n6296 VDD.n6295 23.1255
R28574 VDD.n6297 VDD.n6296 23.1255
R28575 VDD.n6293 VDD.n6292 23.1255
R28576 VDD.n6294 VDD.n6293 23.1255
R28577 VDD.n6286 VDD.n6285 23.1255
R28578 VDD.n6287 VDD.n6286 23.1255
R28579 VDD.n6276 VDD.n6275 23.1255
R28580 VDD.n6277 VDD.n6276 23.1255
R28581 VDD.n6269 VDD.n6268 23.1255
R28582 VDD.n6270 VDD.n6269 23.1255
R28583 VDD.n6266 VDD.n6265 23.1255
R28584 VDD.n6267 VDD.n6266 23.1255
R28585 VDD.n6259 VDD.n6258 23.1255
R28586 VDD.n6260 VDD.n6259 23.1255
R28587 VDD.n6256 VDD.n6255 23.1255
R28588 VDD.n6257 VDD.n6256 23.1255
R28589 VDD.n6249 VDD.n6248 23.1255
R28590 VDD.n6250 VDD.n6249 23.1255
R28591 VDD.n6246 VDD.n6245 23.1255
R28592 VDD.n6247 VDD.n6246 23.1255
R28593 VDD.n6239 VDD.n6238 23.1255
R28594 VDD.n6240 VDD.n6239 23.1255
R28595 VDD.n6236 VDD.n6235 23.1255
R28596 VDD.n6237 VDD.n6236 23.1255
R28597 VDD.n6229 VDD.n6228 23.1255
R28598 VDD.n6230 VDD.n6229 23.1255
R28599 VDD.n6226 VDD.n6225 23.1255
R28600 VDD.n6227 VDD.n6226 23.1255
R28601 VDD.n6219 VDD.n6218 23.1255
R28602 VDD.n6220 VDD.n6219 23.1255
R28603 VDD.n6216 VDD.n6215 23.1255
R28604 VDD.n6217 VDD.n6216 23.1255
R28605 VDD.n5692 VDD.n5691 23.1255
R28606 VDD.n6329 VDD.n6327 23.1255
R28607 VDD.n6327 VDD.n6325 23.1255
R28608 VDD.n6328 VDD.n6326 23.1255
R28609 VDD.n6326 VDD.n5566 23.1255
R28610 VDD.n5431 VDD.n5428 23.1255
R28611 VDD.n5430 VDD.n5428 23.1255
R28612 VDD.n5432 VDD.n5429 23.1255
R28613 VDD.n6448 VDD.n5429 23.1255
R28614 VDD.n5439 VDD.n5435 23.1255
R28615 VDD.n6447 VDD.n5435 23.1255
R28616 VDD.n6441 VDD.n5444 23.1255
R28617 VDD.n6441 VDD.n6440 23.1255
R28618 VDD.n5449 VDD.n5445 23.1255
R28619 VDD.n6437 VDD.n5445 23.1255
R28620 VDD.n6431 VDD.n5454 23.1255
R28621 VDD.n6431 VDD.n6430 23.1255
R28622 VDD.n5459 VDD.n5455 23.1255
R28623 VDD.n6427 VDD.n5455 23.1255
R28624 VDD.n6421 VDD.n5465 23.1255
R28625 VDD.n6421 VDD.n6420 23.1255
R28626 VDD.n5470 VDD.n5466 23.1255
R28627 VDD.n6417 VDD.n5466 23.1255
R28628 VDD.n6411 VDD.n5478 23.1255
R28629 VDD.n6411 VDD.n6410 23.1255
R28630 VDD.n6406 VDD.n6405 23.1255
R28631 VDD.n6407 VDD.n6406 23.1255
R28632 VDD.n6403 VDD.n6402 23.1255
R28633 VDD.n6402 VDD.n6401 23.1255
R28634 VDD.n5486 VDD.n5482 23.1255
R28635 VDD.n6400 VDD.n5482 23.1255
R28636 VDD.n6394 VDD.n5493 23.1255
R28637 VDD.n6394 VDD.n6393 23.1255
R28638 VDD.n5498 VDD.n5494 23.1255
R28639 VDD.n6390 VDD.n5494 23.1255
R28640 VDD.n6384 VDD.n5506 23.1255
R28641 VDD.n6384 VDD.n6383 23.1255
R28642 VDD.n5511 VDD.n5507 23.1255
R28643 VDD.n6380 VDD.n5507 23.1255
R28644 VDD.n6374 VDD.n5516 23.1255
R28645 VDD.n6374 VDD.n6373 23.1255
R28646 VDD.n5521 VDD.n5517 23.1255
R28647 VDD.n6370 VDD.n5517 23.1255
R28648 VDD.n6364 VDD.n5527 23.1255
R28649 VDD.n6364 VDD.n6363 23.1255
R28650 VDD.n5532 VDD.n5528 23.1255
R28651 VDD.n6360 VDD.n5528 23.1255
R28652 VDD.n6354 VDD.n5540 23.1255
R28653 VDD.n6354 VDD.n6353 23.1255
R28654 VDD.n5545 VDD.n5541 23.1255
R28655 VDD.n6350 VDD.n5541 23.1255
R28656 VDD.n6344 VDD.n5550 23.1255
R28657 VDD.n6344 VDD.n6343 23.1255
R28658 VDD.n6446 VDD.n6445 23.1255
R28659 VDD.n6447 VDD.n6446 23.1255
R28660 VDD.n6439 VDD.n6438 23.1255
R28661 VDD.n6440 VDD.n6439 23.1255
R28662 VDD.n6436 VDD.n6435 23.1255
R28663 VDD.n6437 VDD.n6436 23.1255
R28664 VDD.n6429 VDD.n6428 23.1255
R28665 VDD.n6430 VDD.n6429 23.1255
R28666 VDD.n6426 VDD.n6425 23.1255
R28667 VDD.n6427 VDD.n6426 23.1255
R28668 VDD.n6419 VDD.n6418 23.1255
R28669 VDD.n6420 VDD.n6419 23.1255
R28670 VDD.n6416 VDD.n6415 23.1255
R28671 VDD.n6417 VDD.n6416 23.1255
R28672 VDD.n6409 VDD.n6408 23.1255
R28673 VDD.n6410 VDD.n6409 23.1255
R28674 VDD.n6399 VDD.n6398 23.1255
R28675 VDD.n6400 VDD.n6399 23.1255
R28676 VDD.n6392 VDD.n6391 23.1255
R28677 VDD.n6393 VDD.n6392 23.1255
R28678 VDD.n6389 VDD.n6388 23.1255
R28679 VDD.n6390 VDD.n6389 23.1255
R28680 VDD.n6382 VDD.n6381 23.1255
R28681 VDD.n6383 VDD.n6382 23.1255
R28682 VDD.n6379 VDD.n6378 23.1255
R28683 VDD.n6380 VDD.n6379 23.1255
R28684 VDD.n6372 VDD.n6371 23.1255
R28685 VDD.n6373 VDD.n6372 23.1255
R28686 VDD.n6369 VDD.n6368 23.1255
R28687 VDD.n6370 VDD.n6369 23.1255
R28688 VDD.n6362 VDD.n6361 23.1255
R28689 VDD.n6363 VDD.n6362 23.1255
R28690 VDD.n6359 VDD.n6358 23.1255
R28691 VDD.n6360 VDD.n6359 23.1255
R28692 VDD.n6352 VDD.n6351 23.1255
R28693 VDD.n6353 VDD.n6352 23.1255
R28694 VDD.n6349 VDD.n6348 23.1255
R28695 VDD.n6350 VDD.n6349 23.1255
R28696 VDD.n6342 VDD.n6341 23.1255
R28697 VDD.n6343 VDD.n6342 23.1255
R28698 VDD.n6339 VDD.n6338 23.1255
R28699 VDD.n6340 VDD.n6339 23.1255
R28700 VDD.n5556 VDD.n5555 23.1255
R28701 VDD.n6452 VDD.n6450 23.1255
R28702 VDD.n6450 VDD.n6448 23.1255
R28703 VDD.n6451 VDD.n6449 23.1255
R28704 VDD.n6449 VDD.n5430 23.1255
R28705 VDD.n5295 VDD.n5292 23.1255
R28706 VDD.n5294 VDD.n5292 23.1255
R28707 VDD.n5296 VDD.n5293 23.1255
R28708 VDD.n6571 VDD.n5293 23.1255
R28709 VDD.n5303 VDD.n5299 23.1255
R28710 VDD.n6570 VDD.n5299 23.1255
R28711 VDD.n6564 VDD.n5308 23.1255
R28712 VDD.n6564 VDD.n6563 23.1255
R28713 VDD.n5313 VDD.n5309 23.1255
R28714 VDD.n6560 VDD.n5309 23.1255
R28715 VDD.n6554 VDD.n5318 23.1255
R28716 VDD.n6554 VDD.n6553 23.1255
R28717 VDD.n5323 VDD.n5319 23.1255
R28718 VDD.n6550 VDD.n5319 23.1255
R28719 VDD.n6544 VDD.n5329 23.1255
R28720 VDD.n6544 VDD.n6543 23.1255
R28721 VDD.n5334 VDD.n5330 23.1255
R28722 VDD.n6540 VDD.n5330 23.1255
R28723 VDD.n6534 VDD.n5342 23.1255
R28724 VDD.n6534 VDD.n6533 23.1255
R28725 VDD.n6529 VDD.n6528 23.1255
R28726 VDD.n6530 VDD.n6529 23.1255
R28727 VDD.n6526 VDD.n6525 23.1255
R28728 VDD.n6525 VDD.n6524 23.1255
R28729 VDD.n5350 VDD.n5346 23.1255
R28730 VDD.n6523 VDD.n5346 23.1255
R28731 VDD.n6517 VDD.n5357 23.1255
R28732 VDD.n6517 VDD.n6516 23.1255
R28733 VDD.n5362 VDD.n5358 23.1255
R28734 VDD.n6513 VDD.n5358 23.1255
R28735 VDD.n6507 VDD.n5370 23.1255
R28736 VDD.n6507 VDD.n6506 23.1255
R28737 VDD.n5375 VDD.n5371 23.1255
R28738 VDD.n6503 VDD.n5371 23.1255
R28739 VDD.n6497 VDD.n5380 23.1255
R28740 VDD.n6497 VDD.n6496 23.1255
R28741 VDD.n5385 VDD.n5381 23.1255
R28742 VDD.n6493 VDD.n5381 23.1255
R28743 VDD.n6487 VDD.n5391 23.1255
R28744 VDD.n6487 VDD.n6486 23.1255
R28745 VDD.n5396 VDD.n5392 23.1255
R28746 VDD.n6483 VDD.n5392 23.1255
R28747 VDD.n6477 VDD.n5404 23.1255
R28748 VDD.n6477 VDD.n6476 23.1255
R28749 VDD.n5409 VDD.n5405 23.1255
R28750 VDD.n6473 VDD.n5405 23.1255
R28751 VDD.n6467 VDD.n5414 23.1255
R28752 VDD.n6467 VDD.n6466 23.1255
R28753 VDD.n6569 VDD.n6568 23.1255
R28754 VDD.n6570 VDD.n6569 23.1255
R28755 VDD.n6562 VDD.n6561 23.1255
R28756 VDD.n6563 VDD.n6562 23.1255
R28757 VDD.n6559 VDD.n6558 23.1255
R28758 VDD.n6560 VDD.n6559 23.1255
R28759 VDD.n6552 VDD.n6551 23.1255
R28760 VDD.n6553 VDD.n6552 23.1255
R28761 VDD.n6549 VDD.n6548 23.1255
R28762 VDD.n6550 VDD.n6549 23.1255
R28763 VDD.n6542 VDD.n6541 23.1255
R28764 VDD.n6543 VDD.n6542 23.1255
R28765 VDD.n6539 VDD.n6538 23.1255
R28766 VDD.n6540 VDD.n6539 23.1255
R28767 VDD.n6532 VDD.n6531 23.1255
R28768 VDD.n6533 VDD.n6532 23.1255
R28769 VDD.n6522 VDD.n6521 23.1255
R28770 VDD.n6523 VDD.n6522 23.1255
R28771 VDD.n6515 VDD.n6514 23.1255
R28772 VDD.n6516 VDD.n6515 23.1255
R28773 VDD.n6512 VDD.n6511 23.1255
R28774 VDD.n6513 VDD.n6512 23.1255
R28775 VDD.n6505 VDD.n6504 23.1255
R28776 VDD.n6506 VDD.n6505 23.1255
R28777 VDD.n6502 VDD.n6501 23.1255
R28778 VDD.n6503 VDD.n6502 23.1255
R28779 VDD.n6495 VDD.n6494 23.1255
R28780 VDD.n6496 VDD.n6495 23.1255
R28781 VDD.n6492 VDD.n6491 23.1255
R28782 VDD.n6493 VDD.n6492 23.1255
R28783 VDD.n6485 VDD.n6484 23.1255
R28784 VDD.n6486 VDD.n6485 23.1255
R28785 VDD.n6482 VDD.n6481 23.1255
R28786 VDD.n6483 VDD.n6482 23.1255
R28787 VDD.n6475 VDD.n6474 23.1255
R28788 VDD.n6476 VDD.n6475 23.1255
R28789 VDD.n6472 VDD.n6471 23.1255
R28790 VDD.n6473 VDD.n6472 23.1255
R28791 VDD.n6465 VDD.n6464 23.1255
R28792 VDD.n6466 VDD.n6465 23.1255
R28793 VDD.n6462 VDD.n6461 23.1255
R28794 VDD.n6463 VDD.n6462 23.1255
R28795 VDD.n5420 VDD.n5419 23.1255
R28796 VDD.n6575 VDD.n6573 23.1255
R28797 VDD.n6573 VDD.n6571 23.1255
R28798 VDD.n6574 VDD.n6572 23.1255
R28799 VDD.n6572 VDD.n5294 23.1255
R28800 VDD.n5159 VDD.n5156 23.1255
R28801 VDD.n5158 VDD.n5156 23.1255
R28802 VDD.n5160 VDD.n5157 23.1255
R28803 VDD.n6694 VDD.n5157 23.1255
R28804 VDD.n5167 VDD.n5163 23.1255
R28805 VDD.n6693 VDD.n5163 23.1255
R28806 VDD.n6687 VDD.n5172 23.1255
R28807 VDD.n6687 VDD.n6686 23.1255
R28808 VDD.n5177 VDD.n5173 23.1255
R28809 VDD.n6683 VDD.n5173 23.1255
R28810 VDD.n6677 VDD.n5182 23.1255
R28811 VDD.n6677 VDD.n6676 23.1255
R28812 VDD.n5187 VDD.n5183 23.1255
R28813 VDD.n6673 VDD.n5183 23.1255
R28814 VDD.n6667 VDD.n5193 23.1255
R28815 VDD.n6667 VDD.n6666 23.1255
R28816 VDD.n5198 VDD.n5194 23.1255
R28817 VDD.n6663 VDD.n5194 23.1255
R28818 VDD.n6657 VDD.n5206 23.1255
R28819 VDD.n6657 VDD.n6656 23.1255
R28820 VDD.n6652 VDD.n6651 23.1255
R28821 VDD.n6653 VDD.n6652 23.1255
R28822 VDD.n6649 VDD.n6648 23.1255
R28823 VDD.n6648 VDD.n6647 23.1255
R28824 VDD.n5214 VDD.n5210 23.1255
R28825 VDD.n6646 VDD.n5210 23.1255
R28826 VDD.n6640 VDD.n5221 23.1255
R28827 VDD.n6640 VDD.n6639 23.1255
R28828 VDD.n5226 VDD.n5222 23.1255
R28829 VDD.n6636 VDD.n5222 23.1255
R28830 VDD.n6630 VDD.n5234 23.1255
R28831 VDD.n6630 VDD.n6629 23.1255
R28832 VDD.n5239 VDD.n5235 23.1255
R28833 VDD.n6626 VDD.n5235 23.1255
R28834 VDD.n6620 VDD.n5244 23.1255
R28835 VDD.n6620 VDD.n6619 23.1255
R28836 VDD.n5249 VDD.n5245 23.1255
R28837 VDD.n6616 VDD.n5245 23.1255
R28838 VDD.n6610 VDD.n5255 23.1255
R28839 VDD.n6610 VDD.n6609 23.1255
R28840 VDD.n5260 VDD.n5256 23.1255
R28841 VDD.n6606 VDD.n5256 23.1255
R28842 VDD.n6600 VDD.n5268 23.1255
R28843 VDD.n6600 VDD.n6599 23.1255
R28844 VDD.n5273 VDD.n5269 23.1255
R28845 VDD.n6596 VDD.n5269 23.1255
R28846 VDD.n6590 VDD.n5278 23.1255
R28847 VDD.n6590 VDD.n6589 23.1255
R28848 VDD.n6692 VDD.n6691 23.1255
R28849 VDD.n6693 VDD.n6692 23.1255
R28850 VDD.n6685 VDD.n6684 23.1255
R28851 VDD.n6686 VDD.n6685 23.1255
R28852 VDD.n6682 VDD.n6681 23.1255
R28853 VDD.n6683 VDD.n6682 23.1255
R28854 VDD.n6675 VDD.n6674 23.1255
R28855 VDD.n6676 VDD.n6675 23.1255
R28856 VDD.n6672 VDD.n6671 23.1255
R28857 VDD.n6673 VDD.n6672 23.1255
R28858 VDD.n6665 VDD.n6664 23.1255
R28859 VDD.n6666 VDD.n6665 23.1255
R28860 VDD.n6662 VDD.n6661 23.1255
R28861 VDD.n6663 VDD.n6662 23.1255
R28862 VDD.n6655 VDD.n6654 23.1255
R28863 VDD.n6656 VDD.n6655 23.1255
R28864 VDD.n6645 VDD.n6644 23.1255
R28865 VDD.n6646 VDD.n6645 23.1255
R28866 VDD.n6638 VDD.n6637 23.1255
R28867 VDD.n6639 VDD.n6638 23.1255
R28868 VDD.n6635 VDD.n6634 23.1255
R28869 VDD.n6636 VDD.n6635 23.1255
R28870 VDD.n6628 VDD.n6627 23.1255
R28871 VDD.n6629 VDD.n6628 23.1255
R28872 VDD.n6625 VDD.n6624 23.1255
R28873 VDD.n6626 VDD.n6625 23.1255
R28874 VDD.n6618 VDD.n6617 23.1255
R28875 VDD.n6619 VDD.n6618 23.1255
R28876 VDD.n6615 VDD.n6614 23.1255
R28877 VDD.n6616 VDD.n6615 23.1255
R28878 VDD.n6608 VDD.n6607 23.1255
R28879 VDD.n6609 VDD.n6608 23.1255
R28880 VDD.n6605 VDD.n6604 23.1255
R28881 VDD.n6606 VDD.n6605 23.1255
R28882 VDD.n6598 VDD.n6597 23.1255
R28883 VDD.n6599 VDD.n6598 23.1255
R28884 VDD.n6595 VDD.n6594 23.1255
R28885 VDD.n6596 VDD.n6595 23.1255
R28886 VDD.n6588 VDD.n6587 23.1255
R28887 VDD.n6589 VDD.n6588 23.1255
R28888 VDD.n6585 VDD.n6584 23.1255
R28889 VDD.n6586 VDD.n6585 23.1255
R28890 VDD.n5284 VDD.n5283 23.1255
R28891 VDD.n6698 VDD.n6696 23.1255
R28892 VDD.n6696 VDD.n6694 23.1255
R28893 VDD.n6697 VDD.n6695 23.1255
R28894 VDD.n6695 VDD.n5158 23.1255
R28895 VDD.n5023 VDD.n5020 23.1255
R28896 VDD.n5022 VDD.n5020 23.1255
R28897 VDD.n5024 VDD.n5021 23.1255
R28898 VDD.n6817 VDD.n5021 23.1255
R28899 VDD.n5031 VDD.n5027 23.1255
R28900 VDD.n6816 VDD.n5027 23.1255
R28901 VDD.n6810 VDD.n5036 23.1255
R28902 VDD.n6810 VDD.n6809 23.1255
R28903 VDD.n5041 VDD.n5037 23.1255
R28904 VDD.n6806 VDD.n5037 23.1255
R28905 VDD.n6800 VDD.n5046 23.1255
R28906 VDD.n6800 VDD.n6799 23.1255
R28907 VDD.n5051 VDD.n5047 23.1255
R28908 VDD.n6796 VDD.n5047 23.1255
R28909 VDD.n6790 VDD.n5057 23.1255
R28910 VDD.n6790 VDD.n6789 23.1255
R28911 VDD.n5062 VDD.n5058 23.1255
R28912 VDD.n6786 VDD.n5058 23.1255
R28913 VDD.n6780 VDD.n5070 23.1255
R28914 VDD.n6780 VDD.n6779 23.1255
R28915 VDD.n6775 VDD.n6774 23.1255
R28916 VDD.n6776 VDD.n6775 23.1255
R28917 VDD.n6772 VDD.n6771 23.1255
R28918 VDD.n6771 VDD.n6770 23.1255
R28919 VDD.n5078 VDD.n5074 23.1255
R28920 VDD.n6769 VDD.n5074 23.1255
R28921 VDD.n6763 VDD.n5085 23.1255
R28922 VDD.n6763 VDD.n6762 23.1255
R28923 VDD.n5090 VDD.n5086 23.1255
R28924 VDD.n6759 VDD.n5086 23.1255
R28925 VDD.n6753 VDD.n5098 23.1255
R28926 VDD.n6753 VDD.n6752 23.1255
R28927 VDD.n5103 VDD.n5099 23.1255
R28928 VDD.n6749 VDD.n5099 23.1255
R28929 VDD.n6743 VDD.n5108 23.1255
R28930 VDD.n6743 VDD.n6742 23.1255
R28931 VDD.n5113 VDD.n5109 23.1255
R28932 VDD.n6739 VDD.n5109 23.1255
R28933 VDD.n6733 VDD.n5119 23.1255
R28934 VDD.n6733 VDD.n6732 23.1255
R28935 VDD.n5124 VDD.n5120 23.1255
R28936 VDD.n6729 VDD.n5120 23.1255
R28937 VDD.n6723 VDD.n5132 23.1255
R28938 VDD.n6723 VDD.n6722 23.1255
R28939 VDD.n5137 VDD.n5133 23.1255
R28940 VDD.n6719 VDD.n5133 23.1255
R28941 VDD.n6713 VDD.n5142 23.1255
R28942 VDD.n6713 VDD.n6712 23.1255
R28943 VDD.n6815 VDD.n6814 23.1255
R28944 VDD.n6816 VDD.n6815 23.1255
R28945 VDD.n6808 VDD.n6807 23.1255
R28946 VDD.n6809 VDD.n6808 23.1255
R28947 VDD.n6805 VDD.n6804 23.1255
R28948 VDD.n6806 VDD.n6805 23.1255
R28949 VDD.n6798 VDD.n6797 23.1255
R28950 VDD.n6799 VDD.n6798 23.1255
R28951 VDD.n6795 VDD.n6794 23.1255
R28952 VDD.n6796 VDD.n6795 23.1255
R28953 VDD.n6788 VDD.n6787 23.1255
R28954 VDD.n6789 VDD.n6788 23.1255
R28955 VDD.n6785 VDD.n6784 23.1255
R28956 VDD.n6786 VDD.n6785 23.1255
R28957 VDD.n6778 VDD.n6777 23.1255
R28958 VDD.n6779 VDD.n6778 23.1255
R28959 VDD.n6768 VDD.n6767 23.1255
R28960 VDD.n6769 VDD.n6768 23.1255
R28961 VDD.n6761 VDD.n6760 23.1255
R28962 VDD.n6762 VDD.n6761 23.1255
R28963 VDD.n6758 VDD.n6757 23.1255
R28964 VDD.n6759 VDD.n6758 23.1255
R28965 VDD.n6751 VDD.n6750 23.1255
R28966 VDD.n6752 VDD.n6751 23.1255
R28967 VDD.n6748 VDD.n6747 23.1255
R28968 VDD.n6749 VDD.n6748 23.1255
R28969 VDD.n6741 VDD.n6740 23.1255
R28970 VDD.n6742 VDD.n6741 23.1255
R28971 VDD.n6738 VDD.n6737 23.1255
R28972 VDD.n6739 VDD.n6738 23.1255
R28973 VDD.n6731 VDD.n6730 23.1255
R28974 VDD.n6732 VDD.n6731 23.1255
R28975 VDD.n6728 VDD.n6727 23.1255
R28976 VDD.n6729 VDD.n6728 23.1255
R28977 VDD.n6721 VDD.n6720 23.1255
R28978 VDD.n6722 VDD.n6721 23.1255
R28979 VDD.n6718 VDD.n6717 23.1255
R28980 VDD.n6719 VDD.n6718 23.1255
R28981 VDD.n6711 VDD.n6710 23.1255
R28982 VDD.n6712 VDD.n6711 23.1255
R28983 VDD.n6708 VDD.n6707 23.1255
R28984 VDD.n6709 VDD.n6708 23.1255
R28985 VDD.n5148 VDD.n5147 23.1255
R28986 VDD.n6821 VDD.n6819 23.1255
R28987 VDD.n6819 VDD.n6817 23.1255
R28988 VDD.n6820 VDD.n6818 23.1255
R28989 VDD.n6818 VDD.n5022 23.1255
R28990 VDD.n4889 VDD.n4885 23.1255
R28991 VDD.n4889 VDD.n4888 23.1255
R28992 VDD.n4881 VDD.n4877 23.1255
R28993 VDD.n4898 VDD.n4877 23.1255
R28994 VDD.n4902 VDD.n4876 23.1255
R28995 VDD.n4902 VDD.n4901 23.1255
R28996 VDD.n4871 VDD.n4867 23.1255
R28997 VDD.n4908 VDD.n4867 23.1255
R28998 VDD.n4912 VDD.n4866 23.1255
R28999 VDD.n4912 VDD.n4911 23.1255
R29000 VDD.n4860 VDD.n4856 23.1255
R29001 VDD.n4918 VDD.n4856 23.1255
R29002 VDD.n4922 VDD.n4855 23.1255
R29003 VDD.n4922 VDD.n4921 23.1255
R29004 VDD.n4847 VDD.n4843 23.1255
R29005 VDD.n4928 VDD.n4843 23.1255
R29006 VDD.n4932 VDD.n4842 23.1255
R29007 VDD.n4932 VDD.n4931 23.1255
R29008 VDD.n4835 VDD.n4831 23.1255
R29009 VDD.n4938 VDD.n4831 23.1255
R29010 VDD.n4941 VDD.n4940 23.1255
R29011 VDD.n4940 VDD.n4939 23.1255
R29012 VDD.n4944 VDD.n4943 23.1255
R29013 VDD.n4945 VDD.n4944 23.1255
R29014 VDD.n4949 VDD.n4827 23.1255
R29015 VDD.n4949 VDD.n4948 23.1255
R29016 VDD.n4819 VDD.n4815 23.1255
R29017 VDD.n4955 VDD.n4815 23.1255
R29018 VDD.n4959 VDD.n4814 23.1255
R29019 VDD.n4959 VDD.n4958 23.1255
R29020 VDD.n4809 VDD.n4805 23.1255
R29021 VDD.n4965 VDD.n4805 23.1255
R29022 VDD.n4969 VDD.n4804 23.1255
R29023 VDD.n4969 VDD.n4968 23.1255
R29024 VDD.n4798 VDD.n4794 23.1255
R29025 VDD.n4975 VDD.n4794 23.1255
R29026 VDD.n4979 VDD.n4793 23.1255
R29027 VDD.n4979 VDD.n4978 23.1255
R29028 VDD.n4785 VDD.n4781 23.1255
R29029 VDD.n4985 VDD.n4781 23.1255
R29030 VDD.n4989 VDD.n4780 23.1255
R29031 VDD.n4989 VDD.n4988 23.1255
R29032 VDD.n4775 VDD.n4771 23.1255
R29033 VDD.n4995 VDD.n4771 23.1255
R29034 VDD.n4999 VDD.n4770 23.1255
R29035 VDD.n4999 VDD.n4998 23.1255
R29036 VDD.n4764 VDD.n4760 23.1255
R29037 VDD.n5005 VDD.n4760 23.1255
R29038 VDD.n4900 VDD.n4899 23.1255
R29039 VDD.n4901 VDD.n4900 23.1255
R29040 VDD.n4907 VDD.n4906 23.1255
R29041 VDD.n4908 VDD.n4907 23.1255
R29042 VDD.n4910 VDD.n4909 23.1255
R29043 VDD.n4911 VDD.n4910 23.1255
R29044 VDD.n4917 VDD.n4916 23.1255
R29045 VDD.n4918 VDD.n4917 23.1255
R29046 VDD.n4920 VDD.n4919 23.1255
R29047 VDD.n4921 VDD.n4920 23.1255
R29048 VDD.n4927 VDD.n4926 23.1255
R29049 VDD.n4928 VDD.n4927 23.1255
R29050 VDD.n4930 VDD.n4929 23.1255
R29051 VDD.n4931 VDD.n4930 23.1255
R29052 VDD.n4937 VDD.n4936 23.1255
R29053 VDD.n4938 VDD.n4937 23.1255
R29054 VDD.n4947 VDD.n4946 23.1255
R29055 VDD.n4948 VDD.n4947 23.1255
R29056 VDD.n4954 VDD.n4953 23.1255
R29057 VDD.n4955 VDD.n4954 23.1255
R29058 VDD.n4957 VDD.n4956 23.1255
R29059 VDD.n4958 VDD.n4957 23.1255
R29060 VDD.n4964 VDD.n4963 23.1255
R29061 VDD.n4965 VDD.n4964 23.1255
R29062 VDD.n4967 VDD.n4966 23.1255
R29063 VDD.n4968 VDD.n4967 23.1255
R29064 VDD.n4974 VDD.n4973 23.1255
R29065 VDD.n4975 VDD.n4974 23.1255
R29066 VDD.n4977 VDD.n4976 23.1255
R29067 VDD.n4978 VDD.n4977 23.1255
R29068 VDD.n4984 VDD.n4983 23.1255
R29069 VDD.n4985 VDD.n4984 23.1255
R29070 VDD.n4987 VDD.n4986 23.1255
R29071 VDD.n4988 VDD.n4987 23.1255
R29072 VDD.n4994 VDD.n4993 23.1255
R29073 VDD.n4995 VDD.n4994 23.1255
R29074 VDD.n4997 VDD.n4996 23.1255
R29075 VDD.n4998 VDD.n4997 23.1255
R29076 VDD.n5004 VDD.n5003 23.1255
R29077 VDD.n5005 VDD.n5004 23.1255
R29078 VDD.n5006 VDD.n4756 23.1255
R29079 VDD.n5007 VDD.n5006 23.1255
R29080 VDD.n5010 VDD.n5009 23.1255
R29081 VDD.n4897 VDD.n4896 23.1255
R29082 VDD.n4898 VDD.n4897 23.1255
R29083 VDD.n4887 VDD.n4886 23.1255
R29084 VDD.n4888 VDD.n4887 23.1255
R29085 VDD.n1988 VDD.n1984 23.1255
R29086 VDD.n4749 VDD.n1984 23.1255
R29087 VDD.n4743 VDD.n1994 23.1255
R29088 VDD.n4743 VDD.n4742 23.1255
R29089 VDD.n1999 VDD.n1995 23.1255
R29090 VDD.n4739 VDD.n1995 23.1255
R29091 VDD.n4733 VDD.n2004 23.1255
R29092 VDD.n4733 VDD.n4732 23.1255
R29093 VDD.n2009 VDD.n2005 23.1255
R29094 VDD.n4729 VDD.n2005 23.1255
R29095 VDD.n4723 VDD.n2017 23.1255
R29096 VDD.n4723 VDD.n4722 23.1255
R29097 VDD.n2022 VDD.n2018 23.1255
R29098 VDD.n4719 VDD.n2018 23.1255
R29099 VDD.n4713 VDD.n2029 23.1255
R29100 VDD.n4713 VDD.n4712 23.1255
R29101 VDD.n2034 VDD.n2030 23.1255
R29102 VDD.n4709 VDD.n2030 23.1255
R29103 VDD.n2048 VDD.n2047 23.1255
R29104 VDD.n2051 VDD.n2048 23.1255
R29105 VDD.n2053 VDD.n2043 23.1255
R29106 VDD.n2052 VDD.n2043 23.1255
R29107 VDD.n2054 VDD.n2044 23.1255
R29108 VDD.n4693 VDD.n2044 23.1255
R29109 VDD.n4691 VDD.n4690 23.1255
R29110 VDD.n4692 VDD.n4691 23.1255
R29111 VDD.n4688 VDD.n4687 23.1255
R29112 VDD.n4687 VDD.n4686 23.1255
R29113 VDD.n2064 VDD.n2060 23.1255
R29114 VDD.n4685 VDD.n2060 23.1255
R29115 VDD.n4679 VDD.n2071 23.1255
R29116 VDD.n4679 VDD.n4678 23.1255
R29117 VDD.n2076 VDD.n2072 23.1255
R29118 VDD.n4675 VDD.n2072 23.1255
R29119 VDD.n4669 VDD.n2084 23.1255
R29120 VDD.n4669 VDD.n4668 23.1255
R29121 VDD.n2089 VDD.n2085 23.1255
R29122 VDD.n4665 VDD.n2085 23.1255
R29123 VDD.n4659 VDD.n2095 23.1255
R29124 VDD.n4659 VDD.n4658 23.1255
R29125 VDD.n2100 VDD.n2096 23.1255
R29126 VDD.n4655 VDD.n2096 23.1255
R29127 VDD.n4649 VDD.n2105 23.1255
R29128 VDD.n4649 VDD.n4648 23.1255
R29129 VDD.n2110 VDD.n2106 23.1255
R29130 VDD.n4645 VDD.n2106 23.1255
R29131 VDD.n4639 VDD.n4635 23.1255
R29132 VDD.n4639 VDD.n4638 23.1255
R29133 VDD.n1982 VDD.n1978 23.1255
R29134 VDD.n4752 VDD.n4751 23.1255
R29135 VDD.n4751 VDD.n4750 23.1255
R29136 VDD.n4748 VDD.n4747 23.1255
R29137 VDD.n4749 VDD.n4748 23.1255
R29138 VDD.n4741 VDD.n4740 23.1255
R29139 VDD.n4742 VDD.n4741 23.1255
R29140 VDD.n4738 VDD.n4737 23.1255
R29141 VDD.n4739 VDD.n4738 23.1255
R29142 VDD.n4731 VDD.n4730 23.1255
R29143 VDD.n4732 VDD.n4731 23.1255
R29144 VDD.n4728 VDD.n4727 23.1255
R29145 VDD.n4729 VDD.n4728 23.1255
R29146 VDD.n4721 VDD.n4720 23.1255
R29147 VDD.n4722 VDD.n4721 23.1255
R29148 VDD.n4718 VDD.n4717 23.1255
R29149 VDD.n4719 VDD.n4718 23.1255
R29150 VDD.n4711 VDD.n4710 23.1255
R29151 VDD.n4712 VDD.n4711 23.1255
R29152 VDD.n4696 VDD.n4694 23.1255
R29153 VDD.n4694 VDD.n2052 23.1255
R29154 VDD.n4697 VDD.n4695 23.1255
R29155 VDD.n4695 VDD.n4693 23.1255
R29156 VDD.n4684 VDD.n4683 23.1255
R29157 VDD.n4685 VDD.n4684 23.1255
R29158 VDD.n4677 VDD.n4676 23.1255
R29159 VDD.n4678 VDD.n4677 23.1255
R29160 VDD.n4674 VDD.n4673 23.1255
R29161 VDD.n4675 VDD.n4674 23.1255
R29162 VDD.n4667 VDD.n4666 23.1255
R29163 VDD.n4668 VDD.n4667 23.1255
R29164 VDD.n4664 VDD.n4663 23.1255
R29165 VDD.n4665 VDD.n4664 23.1255
R29166 VDD.n4657 VDD.n4656 23.1255
R29167 VDD.n4658 VDD.n4657 23.1255
R29168 VDD.n4654 VDD.n4653 23.1255
R29169 VDD.n4655 VDD.n4654 23.1255
R29170 VDD.n4647 VDD.n4646 23.1255
R29171 VDD.n4648 VDD.n4647 23.1255
R29172 VDD.n4644 VDD.n4643 23.1255
R29173 VDD.n4645 VDD.n4644 23.1255
R29174 VDD.n4637 VDD.n4636 23.1255
R29175 VDD.n4638 VDD.n4637 23.1255
R29176 VDD.n2050 VDD.n2049 23.1255
R29177 VDD.n2051 VDD.n2050 23.1255
R29178 VDD.n4708 VDD.n4707 23.1255
R29179 VDD.n4709 VDD.n4708 23.1255
R29180 VDD.n2124 VDD.n2120 23.1255
R29181 VDD.n4624 VDD.n2120 23.1255
R29182 VDD.n4618 VDD.n2130 23.1255
R29183 VDD.n4618 VDD.n4617 23.1255
R29184 VDD.n2135 VDD.n2131 23.1255
R29185 VDD.n4614 VDD.n2131 23.1255
R29186 VDD.n4608 VDD.n2140 23.1255
R29187 VDD.n4608 VDD.n4607 23.1255
R29188 VDD.n2145 VDD.n2141 23.1255
R29189 VDD.n4604 VDD.n2141 23.1255
R29190 VDD.n4598 VDD.n2153 23.1255
R29191 VDD.n4598 VDD.n4597 23.1255
R29192 VDD.n2158 VDD.n2154 23.1255
R29193 VDD.n4594 VDD.n2154 23.1255
R29194 VDD.n4588 VDD.n2165 23.1255
R29195 VDD.n4588 VDD.n4587 23.1255
R29196 VDD.n2170 VDD.n2166 23.1255
R29197 VDD.n4584 VDD.n2166 23.1255
R29198 VDD.n2184 VDD.n2183 23.1255
R29199 VDD.n2187 VDD.n2184 23.1255
R29200 VDD.n2189 VDD.n2179 23.1255
R29201 VDD.n2188 VDD.n2179 23.1255
R29202 VDD.n2190 VDD.n2180 23.1255
R29203 VDD.n4568 VDD.n2180 23.1255
R29204 VDD.n4566 VDD.n4565 23.1255
R29205 VDD.n4567 VDD.n4566 23.1255
R29206 VDD.n4563 VDD.n4562 23.1255
R29207 VDD.n4562 VDD.n4561 23.1255
R29208 VDD.n2200 VDD.n2196 23.1255
R29209 VDD.n4560 VDD.n2196 23.1255
R29210 VDD.n4554 VDD.n2207 23.1255
R29211 VDD.n4554 VDD.n4553 23.1255
R29212 VDD.n2212 VDD.n2208 23.1255
R29213 VDD.n4550 VDD.n2208 23.1255
R29214 VDD.n4544 VDD.n2220 23.1255
R29215 VDD.n4544 VDD.n4543 23.1255
R29216 VDD.n2225 VDD.n2221 23.1255
R29217 VDD.n4540 VDD.n2221 23.1255
R29218 VDD.n4534 VDD.n2231 23.1255
R29219 VDD.n4534 VDD.n4533 23.1255
R29220 VDD.n2236 VDD.n2232 23.1255
R29221 VDD.n4530 VDD.n2232 23.1255
R29222 VDD.n4524 VDD.n2241 23.1255
R29223 VDD.n4524 VDD.n4523 23.1255
R29224 VDD.n2246 VDD.n2242 23.1255
R29225 VDD.n4520 VDD.n2242 23.1255
R29226 VDD.n4514 VDD.n4510 23.1255
R29227 VDD.n4514 VDD.n4513 23.1255
R29228 VDD.n2118 VDD.n2114 23.1255
R29229 VDD.n4627 VDD.n4626 23.1255
R29230 VDD.n4626 VDD.n4625 23.1255
R29231 VDD.n4623 VDD.n4622 23.1255
R29232 VDD.n4624 VDD.n4623 23.1255
R29233 VDD.n4616 VDD.n4615 23.1255
R29234 VDD.n4617 VDD.n4616 23.1255
R29235 VDD.n4613 VDD.n4612 23.1255
R29236 VDD.n4614 VDD.n4613 23.1255
R29237 VDD.n4606 VDD.n4605 23.1255
R29238 VDD.n4607 VDD.n4606 23.1255
R29239 VDD.n4603 VDD.n4602 23.1255
R29240 VDD.n4604 VDD.n4603 23.1255
R29241 VDD.n4596 VDD.n4595 23.1255
R29242 VDD.n4597 VDD.n4596 23.1255
R29243 VDD.n4593 VDD.n4592 23.1255
R29244 VDD.n4594 VDD.n4593 23.1255
R29245 VDD.n4586 VDD.n4585 23.1255
R29246 VDD.n4587 VDD.n4586 23.1255
R29247 VDD.n4571 VDD.n4569 23.1255
R29248 VDD.n4569 VDD.n2188 23.1255
R29249 VDD.n4572 VDD.n4570 23.1255
R29250 VDD.n4570 VDD.n4568 23.1255
R29251 VDD.n4559 VDD.n4558 23.1255
R29252 VDD.n4560 VDD.n4559 23.1255
R29253 VDD.n4552 VDD.n4551 23.1255
R29254 VDD.n4553 VDD.n4552 23.1255
R29255 VDD.n4549 VDD.n4548 23.1255
R29256 VDD.n4550 VDD.n4549 23.1255
R29257 VDD.n4542 VDD.n4541 23.1255
R29258 VDD.n4543 VDD.n4542 23.1255
R29259 VDD.n4539 VDD.n4538 23.1255
R29260 VDD.n4540 VDD.n4539 23.1255
R29261 VDD.n4532 VDD.n4531 23.1255
R29262 VDD.n4533 VDD.n4532 23.1255
R29263 VDD.n4529 VDD.n4528 23.1255
R29264 VDD.n4530 VDD.n4529 23.1255
R29265 VDD.n4522 VDD.n4521 23.1255
R29266 VDD.n4523 VDD.n4522 23.1255
R29267 VDD.n4519 VDD.n4518 23.1255
R29268 VDD.n4520 VDD.n4519 23.1255
R29269 VDD.n4512 VDD.n4511 23.1255
R29270 VDD.n4513 VDD.n4512 23.1255
R29271 VDD.n2186 VDD.n2185 23.1255
R29272 VDD.n2187 VDD.n2186 23.1255
R29273 VDD.n4583 VDD.n4582 23.1255
R29274 VDD.n4584 VDD.n4583 23.1255
R29275 VDD.n2260 VDD.n2256 23.1255
R29276 VDD.n4499 VDD.n2256 23.1255
R29277 VDD.n4493 VDD.n2266 23.1255
R29278 VDD.n4493 VDD.n4492 23.1255
R29279 VDD.n2271 VDD.n2267 23.1255
R29280 VDD.n4489 VDD.n2267 23.1255
R29281 VDD.n4483 VDD.n2276 23.1255
R29282 VDD.n4483 VDD.n4482 23.1255
R29283 VDD.n2281 VDD.n2277 23.1255
R29284 VDD.n4479 VDD.n2277 23.1255
R29285 VDD.n4473 VDD.n2289 23.1255
R29286 VDD.n4473 VDD.n4472 23.1255
R29287 VDD.n2294 VDD.n2290 23.1255
R29288 VDD.n4469 VDD.n2290 23.1255
R29289 VDD.n4463 VDD.n2301 23.1255
R29290 VDD.n4463 VDD.n4462 23.1255
R29291 VDD.n2306 VDD.n2302 23.1255
R29292 VDD.n4459 VDD.n2302 23.1255
R29293 VDD.n2320 VDD.n2319 23.1255
R29294 VDD.n2323 VDD.n2320 23.1255
R29295 VDD.n2325 VDD.n2315 23.1255
R29296 VDD.n2324 VDD.n2315 23.1255
R29297 VDD.n2326 VDD.n2316 23.1255
R29298 VDD.n4443 VDD.n2316 23.1255
R29299 VDD.n4441 VDD.n4440 23.1255
R29300 VDD.n4442 VDD.n4441 23.1255
R29301 VDD.n4438 VDD.n4437 23.1255
R29302 VDD.n4437 VDD.n4436 23.1255
R29303 VDD.n2336 VDD.n2332 23.1255
R29304 VDD.n4435 VDD.n2332 23.1255
R29305 VDD.n4429 VDD.n2343 23.1255
R29306 VDD.n4429 VDD.n4428 23.1255
R29307 VDD.n2348 VDD.n2344 23.1255
R29308 VDD.n4425 VDD.n2344 23.1255
R29309 VDD.n4419 VDD.n2356 23.1255
R29310 VDD.n4419 VDD.n4418 23.1255
R29311 VDD.n2361 VDD.n2357 23.1255
R29312 VDD.n4415 VDD.n2357 23.1255
R29313 VDD.n4409 VDD.n2367 23.1255
R29314 VDD.n4409 VDD.n4408 23.1255
R29315 VDD.n2372 VDD.n2368 23.1255
R29316 VDD.n4405 VDD.n2368 23.1255
R29317 VDD.n4399 VDD.n2377 23.1255
R29318 VDD.n4399 VDD.n4398 23.1255
R29319 VDD.n2382 VDD.n2378 23.1255
R29320 VDD.n4395 VDD.n2378 23.1255
R29321 VDD.n4389 VDD.n4385 23.1255
R29322 VDD.n4389 VDD.n4388 23.1255
R29323 VDD.n2254 VDD.n2250 23.1255
R29324 VDD.n4502 VDD.n4501 23.1255
R29325 VDD.n4501 VDD.n4500 23.1255
R29326 VDD.n4498 VDD.n4497 23.1255
R29327 VDD.n4499 VDD.n4498 23.1255
R29328 VDD.n4491 VDD.n4490 23.1255
R29329 VDD.n4492 VDD.n4491 23.1255
R29330 VDD.n4488 VDD.n4487 23.1255
R29331 VDD.n4489 VDD.n4488 23.1255
R29332 VDD.n4481 VDD.n4480 23.1255
R29333 VDD.n4482 VDD.n4481 23.1255
R29334 VDD.n4478 VDD.n4477 23.1255
R29335 VDD.n4479 VDD.n4478 23.1255
R29336 VDD.n4471 VDD.n4470 23.1255
R29337 VDD.n4472 VDD.n4471 23.1255
R29338 VDD.n4468 VDD.n4467 23.1255
R29339 VDD.n4469 VDD.n4468 23.1255
R29340 VDD.n4461 VDD.n4460 23.1255
R29341 VDD.n4462 VDD.n4461 23.1255
R29342 VDD.n4446 VDD.n4444 23.1255
R29343 VDD.n4444 VDD.n2324 23.1255
R29344 VDD.n4447 VDD.n4445 23.1255
R29345 VDD.n4445 VDD.n4443 23.1255
R29346 VDD.n4434 VDD.n4433 23.1255
R29347 VDD.n4435 VDD.n4434 23.1255
R29348 VDD.n4427 VDD.n4426 23.1255
R29349 VDD.n4428 VDD.n4427 23.1255
R29350 VDD.n4424 VDD.n4423 23.1255
R29351 VDD.n4425 VDD.n4424 23.1255
R29352 VDD.n4417 VDD.n4416 23.1255
R29353 VDD.n4418 VDD.n4417 23.1255
R29354 VDD.n4414 VDD.n4413 23.1255
R29355 VDD.n4415 VDD.n4414 23.1255
R29356 VDD.n4407 VDD.n4406 23.1255
R29357 VDD.n4408 VDD.n4407 23.1255
R29358 VDD.n4404 VDD.n4403 23.1255
R29359 VDD.n4405 VDD.n4404 23.1255
R29360 VDD.n4397 VDD.n4396 23.1255
R29361 VDD.n4398 VDD.n4397 23.1255
R29362 VDD.n4394 VDD.n4393 23.1255
R29363 VDD.n4395 VDD.n4394 23.1255
R29364 VDD.n4387 VDD.n4386 23.1255
R29365 VDD.n4388 VDD.n4387 23.1255
R29366 VDD.n2322 VDD.n2321 23.1255
R29367 VDD.n2323 VDD.n2322 23.1255
R29368 VDD.n4458 VDD.n4457 23.1255
R29369 VDD.n4459 VDD.n4458 23.1255
R29370 VDD.n2396 VDD.n2392 23.1255
R29371 VDD.n4374 VDD.n2392 23.1255
R29372 VDD.n4368 VDD.n2402 23.1255
R29373 VDD.n4368 VDD.n4367 23.1255
R29374 VDD.n2407 VDD.n2403 23.1255
R29375 VDD.n4364 VDD.n2403 23.1255
R29376 VDD.n4358 VDD.n2412 23.1255
R29377 VDD.n4358 VDD.n4357 23.1255
R29378 VDD.n2417 VDD.n2413 23.1255
R29379 VDD.n4354 VDD.n2413 23.1255
R29380 VDD.n4348 VDD.n2425 23.1255
R29381 VDD.n4348 VDD.n4347 23.1255
R29382 VDD.n2430 VDD.n2426 23.1255
R29383 VDD.n4344 VDD.n2426 23.1255
R29384 VDD.n4338 VDD.n2437 23.1255
R29385 VDD.n4338 VDD.n4337 23.1255
R29386 VDD.n2442 VDD.n2438 23.1255
R29387 VDD.n4334 VDD.n2438 23.1255
R29388 VDD.n2456 VDD.n2455 23.1255
R29389 VDD.n2459 VDD.n2456 23.1255
R29390 VDD.n2461 VDD.n2451 23.1255
R29391 VDD.n2460 VDD.n2451 23.1255
R29392 VDD.n2462 VDD.n2452 23.1255
R29393 VDD.n4318 VDD.n2452 23.1255
R29394 VDD.n4316 VDD.n4315 23.1255
R29395 VDD.n4317 VDD.n4316 23.1255
R29396 VDD.n4313 VDD.n4312 23.1255
R29397 VDD.n4312 VDD.n4311 23.1255
R29398 VDD.n2472 VDD.n2468 23.1255
R29399 VDD.n4310 VDD.n2468 23.1255
R29400 VDD.n4304 VDD.n2479 23.1255
R29401 VDD.n4304 VDD.n4303 23.1255
R29402 VDD.n2484 VDD.n2480 23.1255
R29403 VDD.n4300 VDD.n2480 23.1255
R29404 VDD.n4294 VDD.n2492 23.1255
R29405 VDD.n4294 VDD.n4293 23.1255
R29406 VDD.n2497 VDD.n2493 23.1255
R29407 VDD.n4290 VDD.n2493 23.1255
R29408 VDD.n4284 VDD.n2503 23.1255
R29409 VDD.n4284 VDD.n4283 23.1255
R29410 VDD.n2508 VDD.n2504 23.1255
R29411 VDD.n4280 VDD.n2504 23.1255
R29412 VDD.n4274 VDD.n2513 23.1255
R29413 VDD.n4274 VDD.n4273 23.1255
R29414 VDD.n2518 VDD.n2514 23.1255
R29415 VDD.n4270 VDD.n2514 23.1255
R29416 VDD.n4264 VDD.n4260 23.1255
R29417 VDD.n4264 VDD.n4263 23.1255
R29418 VDD.n2390 VDD.n2386 23.1255
R29419 VDD.n4377 VDD.n4376 23.1255
R29420 VDD.n4376 VDD.n4375 23.1255
R29421 VDD.n4373 VDD.n4372 23.1255
R29422 VDD.n4374 VDD.n4373 23.1255
R29423 VDD.n4366 VDD.n4365 23.1255
R29424 VDD.n4367 VDD.n4366 23.1255
R29425 VDD.n4363 VDD.n4362 23.1255
R29426 VDD.n4364 VDD.n4363 23.1255
R29427 VDD.n4356 VDD.n4355 23.1255
R29428 VDD.n4357 VDD.n4356 23.1255
R29429 VDD.n4353 VDD.n4352 23.1255
R29430 VDD.n4354 VDD.n4353 23.1255
R29431 VDD.n4346 VDD.n4345 23.1255
R29432 VDD.n4347 VDD.n4346 23.1255
R29433 VDD.n4343 VDD.n4342 23.1255
R29434 VDD.n4344 VDD.n4343 23.1255
R29435 VDD.n4336 VDD.n4335 23.1255
R29436 VDD.n4337 VDD.n4336 23.1255
R29437 VDD.n4321 VDD.n4319 23.1255
R29438 VDD.n4319 VDD.n2460 23.1255
R29439 VDD.n4322 VDD.n4320 23.1255
R29440 VDD.n4320 VDD.n4318 23.1255
R29441 VDD.n4309 VDD.n4308 23.1255
R29442 VDD.n4310 VDD.n4309 23.1255
R29443 VDD.n4302 VDD.n4301 23.1255
R29444 VDD.n4303 VDD.n4302 23.1255
R29445 VDD.n4299 VDD.n4298 23.1255
R29446 VDD.n4300 VDD.n4299 23.1255
R29447 VDD.n4292 VDD.n4291 23.1255
R29448 VDD.n4293 VDD.n4292 23.1255
R29449 VDD.n4289 VDD.n4288 23.1255
R29450 VDD.n4290 VDD.n4289 23.1255
R29451 VDD.n4282 VDD.n4281 23.1255
R29452 VDD.n4283 VDD.n4282 23.1255
R29453 VDD.n4279 VDD.n4278 23.1255
R29454 VDD.n4280 VDD.n4279 23.1255
R29455 VDD.n4272 VDD.n4271 23.1255
R29456 VDD.n4273 VDD.n4272 23.1255
R29457 VDD.n4269 VDD.n4268 23.1255
R29458 VDD.n4270 VDD.n4269 23.1255
R29459 VDD.n4262 VDD.n4261 23.1255
R29460 VDD.n4263 VDD.n4262 23.1255
R29461 VDD.n2458 VDD.n2457 23.1255
R29462 VDD.n2459 VDD.n2458 23.1255
R29463 VDD.n4333 VDD.n4332 23.1255
R29464 VDD.n4334 VDD.n4333 23.1255
R29465 VDD.n2532 VDD.n2528 23.1255
R29466 VDD.n4249 VDD.n2528 23.1255
R29467 VDD.n4243 VDD.n2538 23.1255
R29468 VDD.n4243 VDD.n4242 23.1255
R29469 VDD.n2543 VDD.n2539 23.1255
R29470 VDD.n4239 VDD.n2539 23.1255
R29471 VDD.n4233 VDD.n2548 23.1255
R29472 VDD.n4233 VDD.n4232 23.1255
R29473 VDD.n2553 VDD.n2549 23.1255
R29474 VDD.n4229 VDD.n2549 23.1255
R29475 VDD.n4223 VDD.n2561 23.1255
R29476 VDD.n4223 VDD.n4222 23.1255
R29477 VDD.n2566 VDD.n2562 23.1255
R29478 VDD.n4219 VDD.n2562 23.1255
R29479 VDD.n4213 VDD.n2573 23.1255
R29480 VDD.n4213 VDD.n4212 23.1255
R29481 VDD.n2578 VDD.n2574 23.1255
R29482 VDD.n4209 VDD.n2574 23.1255
R29483 VDD.n2592 VDD.n2591 23.1255
R29484 VDD.n2595 VDD.n2592 23.1255
R29485 VDD.n2597 VDD.n2587 23.1255
R29486 VDD.n2596 VDD.n2587 23.1255
R29487 VDD.n2598 VDD.n2588 23.1255
R29488 VDD.n4193 VDD.n2588 23.1255
R29489 VDD.n4191 VDD.n4190 23.1255
R29490 VDD.n4192 VDD.n4191 23.1255
R29491 VDD.n4188 VDD.n4187 23.1255
R29492 VDD.n4187 VDD.n4186 23.1255
R29493 VDD.n2608 VDD.n2604 23.1255
R29494 VDD.n4185 VDD.n2604 23.1255
R29495 VDD.n4179 VDD.n2615 23.1255
R29496 VDD.n4179 VDD.n4178 23.1255
R29497 VDD.n2620 VDD.n2616 23.1255
R29498 VDD.n4175 VDD.n2616 23.1255
R29499 VDD.n4169 VDD.n2628 23.1255
R29500 VDD.n4169 VDD.n4168 23.1255
R29501 VDD.n2633 VDD.n2629 23.1255
R29502 VDD.n4165 VDD.n2629 23.1255
R29503 VDD.n4159 VDD.n2639 23.1255
R29504 VDD.n4159 VDD.n4158 23.1255
R29505 VDD.n2644 VDD.n2640 23.1255
R29506 VDD.n4155 VDD.n2640 23.1255
R29507 VDD.n4149 VDD.n2649 23.1255
R29508 VDD.n4149 VDD.n4148 23.1255
R29509 VDD.n2654 VDD.n2650 23.1255
R29510 VDD.n4145 VDD.n2650 23.1255
R29511 VDD.n4139 VDD.n4135 23.1255
R29512 VDD.n4139 VDD.n4138 23.1255
R29513 VDD.n2526 VDD.n2522 23.1255
R29514 VDD.n4252 VDD.n4251 23.1255
R29515 VDD.n4251 VDD.n4250 23.1255
R29516 VDD.n4248 VDD.n4247 23.1255
R29517 VDD.n4249 VDD.n4248 23.1255
R29518 VDD.n4241 VDD.n4240 23.1255
R29519 VDD.n4242 VDD.n4241 23.1255
R29520 VDD.n4238 VDD.n4237 23.1255
R29521 VDD.n4239 VDD.n4238 23.1255
R29522 VDD.n4231 VDD.n4230 23.1255
R29523 VDD.n4232 VDD.n4231 23.1255
R29524 VDD.n4228 VDD.n4227 23.1255
R29525 VDD.n4229 VDD.n4228 23.1255
R29526 VDD.n4221 VDD.n4220 23.1255
R29527 VDD.n4222 VDD.n4221 23.1255
R29528 VDD.n4218 VDD.n4217 23.1255
R29529 VDD.n4219 VDD.n4218 23.1255
R29530 VDD.n4211 VDD.n4210 23.1255
R29531 VDD.n4212 VDD.n4211 23.1255
R29532 VDD.n4196 VDD.n4194 23.1255
R29533 VDD.n4194 VDD.n2596 23.1255
R29534 VDD.n4197 VDD.n4195 23.1255
R29535 VDD.n4195 VDD.n4193 23.1255
R29536 VDD.n4184 VDD.n4183 23.1255
R29537 VDD.n4185 VDD.n4184 23.1255
R29538 VDD.n4177 VDD.n4176 23.1255
R29539 VDD.n4178 VDD.n4177 23.1255
R29540 VDD.n4174 VDD.n4173 23.1255
R29541 VDD.n4175 VDD.n4174 23.1255
R29542 VDD.n4167 VDD.n4166 23.1255
R29543 VDD.n4168 VDD.n4167 23.1255
R29544 VDD.n4164 VDD.n4163 23.1255
R29545 VDD.n4165 VDD.n4164 23.1255
R29546 VDD.n4157 VDD.n4156 23.1255
R29547 VDD.n4158 VDD.n4157 23.1255
R29548 VDD.n4154 VDD.n4153 23.1255
R29549 VDD.n4155 VDD.n4154 23.1255
R29550 VDD.n4147 VDD.n4146 23.1255
R29551 VDD.n4148 VDD.n4147 23.1255
R29552 VDD.n4144 VDD.n4143 23.1255
R29553 VDD.n4145 VDD.n4144 23.1255
R29554 VDD.n4137 VDD.n4136 23.1255
R29555 VDD.n4138 VDD.n4137 23.1255
R29556 VDD.n2594 VDD.n2593 23.1255
R29557 VDD.n2595 VDD.n2594 23.1255
R29558 VDD.n4208 VDD.n4207 23.1255
R29559 VDD.n4209 VDD.n4208 23.1255
R29560 VDD.n2668 VDD.n2664 23.1255
R29561 VDD.n4124 VDD.n2664 23.1255
R29562 VDD.n4118 VDD.n2674 23.1255
R29563 VDD.n4118 VDD.n4117 23.1255
R29564 VDD.n2679 VDD.n2675 23.1255
R29565 VDD.n4114 VDD.n2675 23.1255
R29566 VDD.n4108 VDD.n2684 23.1255
R29567 VDD.n4108 VDD.n4107 23.1255
R29568 VDD.n2689 VDD.n2685 23.1255
R29569 VDD.n4104 VDD.n2685 23.1255
R29570 VDD.n4098 VDD.n2697 23.1255
R29571 VDD.n4098 VDD.n4097 23.1255
R29572 VDD.n2702 VDD.n2698 23.1255
R29573 VDD.n4094 VDD.n2698 23.1255
R29574 VDD.n4088 VDD.n2709 23.1255
R29575 VDD.n4088 VDD.n4087 23.1255
R29576 VDD.n2714 VDD.n2710 23.1255
R29577 VDD.n4084 VDD.n2710 23.1255
R29578 VDD.n2728 VDD.n2727 23.1255
R29579 VDD.n2731 VDD.n2728 23.1255
R29580 VDD.n2733 VDD.n2723 23.1255
R29581 VDD.n2732 VDD.n2723 23.1255
R29582 VDD.n2734 VDD.n2724 23.1255
R29583 VDD.n4068 VDD.n2724 23.1255
R29584 VDD.n4066 VDD.n4065 23.1255
R29585 VDD.n4067 VDD.n4066 23.1255
R29586 VDD.n4063 VDD.n4062 23.1255
R29587 VDD.n4062 VDD.n4061 23.1255
R29588 VDD.n2744 VDD.n2740 23.1255
R29589 VDD.n4060 VDD.n2740 23.1255
R29590 VDD.n4054 VDD.n2751 23.1255
R29591 VDD.n4054 VDD.n4053 23.1255
R29592 VDD.n2756 VDD.n2752 23.1255
R29593 VDD.n4050 VDD.n2752 23.1255
R29594 VDD.n4044 VDD.n2764 23.1255
R29595 VDD.n4044 VDD.n4043 23.1255
R29596 VDD.n2769 VDD.n2765 23.1255
R29597 VDD.n4040 VDD.n2765 23.1255
R29598 VDD.n4034 VDD.n2775 23.1255
R29599 VDD.n4034 VDD.n4033 23.1255
R29600 VDD.n2780 VDD.n2776 23.1255
R29601 VDD.n4030 VDD.n2776 23.1255
R29602 VDD.n4024 VDD.n2785 23.1255
R29603 VDD.n4024 VDD.n4023 23.1255
R29604 VDD.n2790 VDD.n2786 23.1255
R29605 VDD.n4020 VDD.n2786 23.1255
R29606 VDD.n4014 VDD.n4010 23.1255
R29607 VDD.n4014 VDD.n4013 23.1255
R29608 VDD.n2662 VDD.n2658 23.1255
R29609 VDD.n4127 VDD.n4126 23.1255
R29610 VDD.n4126 VDD.n4125 23.1255
R29611 VDD.n4123 VDD.n4122 23.1255
R29612 VDD.n4124 VDD.n4123 23.1255
R29613 VDD.n4116 VDD.n4115 23.1255
R29614 VDD.n4117 VDD.n4116 23.1255
R29615 VDD.n4113 VDD.n4112 23.1255
R29616 VDD.n4114 VDD.n4113 23.1255
R29617 VDD.n4106 VDD.n4105 23.1255
R29618 VDD.n4107 VDD.n4106 23.1255
R29619 VDD.n4103 VDD.n4102 23.1255
R29620 VDD.n4104 VDD.n4103 23.1255
R29621 VDD.n4096 VDD.n4095 23.1255
R29622 VDD.n4097 VDD.n4096 23.1255
R29623 VDD.n4093 VDD.n4092 23.1255
R29624 VDD.n4094 VDD.n4093 23.1255
R29625 VDD.n4086 VDD.n4085 23.1255
R29626 VDD.n4087 VDD.n4086 23.1255
R29627 VDD.n4071 VDD.n4069 23.1255
R29628 VDD.n4069 VDD.n2732 23.1255
R29629 VDD.n4072 VDD.n4070 23.1255
R29630 VDD.n4070 VDD.n4068 23.1255
R29631 VDD.n4059 VDD.n4058 23.1255
R29632 VDD.n4060 VDD.n4059 23.1255
R29633 VDD.n4052 VDD.n4051 23.1255
R29634 VDD.n4053 VDD.n4052 23.1255
R29635 VDD.n4049 VDD.n4048 23.1255
R29636 VDD.n4050 VDD.n4049 23.1255
R29637 VDD.n4042 VDD.n4041 23.1255
R29638 VDD.n4043 VDD.n4042 23.1255
R29639 VDD.n4039 VDD.n4038 23.1255
R29640 VDD.n4040 VDD.n4039 23.1255
R29641 VDD.n4032 VDD.n4031 23.1255
R29642 VDD.n4033 VDD.n4032 23.1255
R29643 VDD.n4029 VDD.n4028 23.1255
R29644 VDD.n4030 VDD.n4029 23.1255
R29645 VDD.n4022 VDD.n4021 23.1255
R29646 VDD.n4023 VDD.n4022 23.1255
R29647 VDD.n4019 VDD.n4018 23.1255
R29648 VDD.n4020 VDD.n4019 23.1255
R29649 VDD.n4012 VDD.n4011 23.1255
R29650 VDD.n4013 VDD.n4012 23.1255
R29651 VDD.n2730 VDD.n2729 23.1255
R29652 VDD.n2731 VDD.n2730 23.1255
R29653 VDD.n4083 VDD.n4082 23.1255
R29654 VDD.n4084 VDD.n4083 23.1255
R29655 VDD.n2804 VDD.n2800 23.1255
R29656 VDD.n3999 VDD.n2800 23.1255
R29657 VDD.n3993 VDD.n2810 23.1255
R29658 VDD.n3993 VDD.n3992 23.1255
R29659 VDD.n2815 VDD.n2811 23.1255
R29660 VDD.n3989 VDD.n2811 23.1255
R29661 VDD.n3983 VDD.n2820 23.1255
R29662 VDD.n3983 VDD.n3982 23.1255
R29663 VDD.n2825 VDD.n2821 23.1255
R29664 VDD.n3979 VDD.n2821 23.1255
R29665 VDD.n3973 VDD.n2833 23.1255
R29666 VDD.n3973 VDD.n3972 23.1255
R29667 VDD.n2838 VDD.n2834 23.1255
R29668 VDD.n3969 VDD.n2834 23.1255
R29669 VDD.n3963 VDD.n2845 23.1255
R29670 VDD.n3963 VDD.n3962 23.1255
R29671 VDD.n2850 VDD.n2846 23.1255
R29672 VDD.n3959 VDD.n2846 23.1255
R29673 VDD.n2864 VDD.n2863 23.1255
R29674 VDD.n2867 VDD.n2864 23.1255
R29675 VDD.n2869 VDD.n2859 23.1255
R29676 VDD.n2868 VDD.n2859 23.1255
R29677 VDD.n2870 VDD.n2860 23.1255
R29678 VDD.n3943 VDD.n2860 23.1255
R29679 VDD.n3941 VDD.n3940 23.1255
R29680 VDD.n3942 VDD.n3941 23.1255
R29681 VDD.n3938 VDD.n3937 23.1255
R29682 VDD.n3937 VDD.n3936 23.1255
R29683 VDD.n2880 VDD.n2876 23.1255
R29684 VDD.n3935 VDD.n2876 23.1255
R29685 VDD.n3929 VDD.n2887 23.1255
R29686 VDD.n3929 VDD.n3928 23.1255
R29687 VDD.n2892 VDD.n2888 23.1255
R29688 VDD.n3925 VDD.n2888 23.1255
R29689 VDD.n3919 VDD.n2900 23.1255
R29690 VDD.n3919 VDD.n3918 23.1255
R29691 VDD.n2905 VDD.n2901 23.1255
R29692 VDD.n3915 VDD.n2901 23.1255
R29693 VDD.n3909 VDD.n2911 23.1255
R29694 VDD.n3909 VDD.n3908 23.1255
R29695 VDD.n2916 VDD.n2912 23.1255
R29696 VDD.n3905 VDD.n2912 23.1255
R29697 VDD.n3899 VDD.n2921 23.1255
R29698 VDD.n3899 VDD.n3898 23.1255
R29699 VDD.n2926 VDD.n2922 23.1255
R29700 VDD.n3895 VDD.n2922 23.1255
R29701 VDD.n3889 VDD.n3885 23.1255
R29702 VDD.n3889 VDD.n3888 23.1255
R29703 VDD.n2798 VDD.n2794 23.1255
R29704 VDD.n4002 VDD.n4001 23.1255
R29705 VDD.n4001 VDD.n4000 23.1255
R29706 VDD.n3998 VDD.n3997 23.1255
R29707 VDD.n3999 VDD.n3998 23.1255
R29708 VDD.n3991 VDD.n3990 23.1255
R29709 VDD.n3992 VDD.n3991 23.1255
R29710 VDD.n3988 VDD.n3987 23.1255
R29711 VDD.n3989 VDD.n3988 23.1255
R29712 VDD.n3981 VDD.n3980 23.1255
R29713 VDD.n3982 VDD.n3981 23.1255
R29714 VDD.n3978 VDD.n3977 23.1255
R29715 VDD.n3979 VDD.n3978 23.1255
R29716 VDD.n3971 VDD.n3970 23.1255
R29717 VDD.n3972 VDD.n3971 23.1255
R29718 VDD.n3968 VDD.n3967 23.1255
R29719 VDD.n3969 VDD.n3968 23.1255
R29720 VDD.n3961 VDD.n3960 23.1255
R29721 VDD.n3962 VDD.n3961 23.1255
R29722 VDD.n3946 VDD.n3944 23.1255
R29723 VDD.n3944 VDD.n2868 23.1255
R29724 VDD.n3947 VDD.n3945 23.1255
R29725 VDD.n3945 VDD.n3943 23.1255
R29726 VDD.n3934 VDD.n3933 23.1255
R29727 VDD.n3935 VDD.n3934 23.1255
R29728 VDD.n3927 VDD.n3926 23.1255
R29729 VDD.n3928 VDD.n3927 23.1255
R29730 VDD.n3924 VDD.n3923 23.1255
R29731 VDD.n3925 VDD.n3924 23.1255
R29732 VDD.n3917 VDD.n3916 23.1255
R29733 VDD.n3918 VDD.n3917 23.1255
R29734 VDD.n3914 VDD.n3913 23.1255
R29735 VDD.n3915 VDD.n3914 23.1255
R29736 VDD.n3907 VDD.n3906 23.1255
R29737 VDD.n3908 VDD.n3907 23.1255
R29738 VDD.n3904 VDD.n3903 23.1255
R29739 VDD.n3905 VDD.n3904 23.1255
R29740 VDD.n3897 VDD.n3896 23.1255
R29741 VDD.n3898 VDD.n3897 23.1255
R29742 VDD.n3894 VDD.n3893 23.1255
R29743 VDD.n3895 VDD.n3894 23.1255
R29744 VDD.n3887 VDD.n3886 23.1255
R29745 VDD.n3888 VDD.n3887 23.1255
R29746 VDD.n2866 VDD.n2865 23.1255
R29747 VDD.n2867 VDD.n2866 23.1255
R29748 VDD.n3958 VDD.n3957 23.1255
R29749 VDD.n3959 VDD.n3958 23.1255
R29750 VDD.n3212 VDD.n3209 23.1255
R29751 VDD.n3211 VDD.n3209 23.1255
R29752 VDD.n3213 VDD.n3210 23.1255
R29753 VDD.n3548 VDD.n3210 23.1255
R29754 VDD.n3220 VDD.n3216 23.1255
R29755 VDD.n3547 VDD.n3216 23.1255
R29756 VDD.n3541 VDD.n3225 23.1255
R29757 VDD.n3541 VDD.n3540 23.1255
R29758 VDD.n3230 VDD.n3226 23.1255
R29759 VDD.n3537 VDD.n3226 23.1255
R29760 VDD.n3238 VDD.n3234 23.1255
R29761 VDD.n3238 VDD.n3237 23.1255
R29762 VDD.n3551 VDD.n3549 23.1255
R29763 VDD.n3549 VDD.n3211 23.1255
R29764 VDD.n3552 VDD.n3550 23.1255
R29765 VDD.n3550 VDD.n3548 23.1255
R29766 VDD.n3546 VDD.n3545 23.1255
R29767 VDD.n3547 VDD.n3546 23.1255
R29768 VDD.n3539 VDD.n3538 23.1255
R29769 VDD.n3540 VDD.n3539 23.1255
R29770 VDD.n3236 VDD.n3235 23.1255
R29771 VDD.n3237 VDD.n3236 23.1255
R29772 VDD.n3536 VDD.n3535 23.1255
R29773 VDD.n3537 VDD.n3536 23.1255
R29774 VDD.n3369 VDD.n3290 23.1255
R29775 VDD.n3370 VDD.n3369 23.1255
R29776 VDD.n3381 VDD.n3380 23.1255
R29777 VDD.n3382 VDD.n3381 23.1255
R29778 VDD.n3383 VDD.n3283 23.1255
R29779 VDD.n3384 VDD.n3383 23.1255
R29780 VDD.n3387 VDD.n3386 23.1255
R29781 VDD.n3373 VDD.n3372 23.1255
R29782 VDD.n3372 VDD.n3371 23.1255
R29783 VDD.n3367 VDD.n3363 23.1255
R29784 VDD.n3407 VDD.n3399 23.1255
R29785 VDD.n3408 VDD.n3407 23.1255
R29786 VDD.n3418 VDD.n3417 23.1255
R29787 VDD.n3419 VDD.n3418 23.1255
R29788 VDD.n3420 VDD.n3392 23.1255
R29789 VDD.n3421 VDD.n3420 23.1255
R29790 VDD.n3424 VDD.n3423 23.1255
R29791 VDD.n3411 VDD.n3410 23.1255
R29792 VDD.n3410 VDD.n3409 23.1255
R29793 VDD.n3405 VDD.n3401 23.1255
R29794 VDD.n3447 VDD.n3446 23.1255
R29795 VDD.n3448 VDD.n3447 23.1255
R29796 VDD.n3270 VDD.n3265 23.1255
R29797 VDD.n3271 VDD.n3270 23.1255
R29798 VDD.n3272 VDD.n3266 23.1255
R29799 VDD.n3273 VDD.n3272 23.1255
R29800 VDD.n3276 VDD.n3275 23.1255
R29801 VDD.n3451 VDD.n3450 23.1255
R29802 VDD.n3450 VDD.n3449 23.1255
R29803 VDD.n3260 VDD.n3256 23.1255
R29804 VDD.n3464 VDD.n3253 23.1255
R29805 VDD.n3465 VDD.n3464 23.1255
R29806 VDD.n3476 VDD.n3475 23.1255
R29807 VDD.n3477 VDD.n3476 23.1255
R29808 VDD.n3478 VDD.n3246 23.1255
R29809 VDD.n3479 VDD.n3478 23.1255
R29810 VDD.n3482 VDD.n3481 23.1255
R29811 VDD.n3468 VDD.n3467 23.1255
R29812 VDD.n3467 VDD.n3466 23.1255
R29813 VDD.n3462 VDD.n3458 23.1255
R29814 VDD.n3501 VDD.n3493 23.1255
R29815 VDD.n3502 VDD.n3501 23.1255
R29816 VDD.n3512 VDD.n3511 23.1255
R29817 VDD.n3513 VDD.n3512 23.1255
R29818 VDD.n3514 VDD.n3486 23.1255
R29819 VDD.n3515 VDD.n3514 23.1255
R29820 VDD.n3518 VDD.n3517 23.1255
R29821 VDD.n3505 VDD.n3504 23.1255
R29822 VDD.n3504 VDD.n3503 23.1255
R29823 VDD.n3499 VDD.n3495 23.1255
R29824 VDD.n3352 VDD.n3351 23.1255
R29825 VDD.n3353 VDD.n3352 23.1255
R29826 VDD.n3326 VDD.n3321 23.1255
R29827 VDD.n3327 VDD.n3326 23.1255
R29828 VDD.n3328 VDD.n3322 23.1255
R29829 VDD.n3329 VDD.n3328 23.1255
R29830 VDD.n3332 VDD.n3331 23.1255
R29831 VDD.n3356 VDD.n3355 23.1255
R29832 VDD.n3355 VDD.n3354 23.1255
R29833 VDD.n3316 VDD.n3312 23.1255
R29834 VDD.n2940 VDD.n2936 23.1255
R29835 VDD.n3874 VDD.n2936 23.1255
R29836 VDD.n3868 VDD.n2946 23.1255
R29837 VDD.n3868 VDD.n3867 23.1255
R29838 VDD.n2951 VDD.n2947 23.1255
R29839 VDD.n3864 VDD.n2947 23.1255
R29840 VDD.n3858 VDD.n2956 23.1255
R29841 VDD.n3858 VDD.n3857 23.1255
R29842 VDD.n2961 VDD.n2957 23.1255
R29843 VDD.n3854 VDD.n2957 23.1255
R29844 VDD.n3848 VDD.n2969 23.1255
R29845 VDD.n3848 VDD.n3847 23.1255
R29846 VDD.n2974 VDD.n2970 23.1255
R29847 VDD.n3844 VDD.n2970 23.1255
R29848 VDD.n3838 VDD.n3671 23.1255
R29849 VDD.n3838 VDD.n3837 23.1255
R29850 VDD.n3676 VDD.n3672 23.1255
R29851 VDD.n3834 VDD.n3672 23.1255
R29852 VDD.n3690 VDD.n3689 23.1255
R29853 VDD.n3693 VDD.n3690 23.1255
R29854 VDD.n3695 VDD.n3685 23.1255
R29855 VDD.n3694 VDD.n3685 23.1255
R29856 VDD.n3696 VDD.n3686 23.1255
R29857 VDD.n3818 VDD.n3686 23.1255
R29858 VDD.n3816 VDD.n3815 23.1255
R29859 VDD.n3817 VDD.n3816 23.1255
R29860 VDD.n3813 VDD.n3812 23.1255
R29861 VDD.n3812 VDD.n3811 23.1255
R29862 VDD.n3706 VDD.n3702 23.1255
R29863 VDD.n3810 VDD.n3702 23.1255
R29864 VDD.n3804 VDD.n3713 23.1255
R29865 VDD.n3804 VDD.n3803 23.1255
R29866 VDD.n3718 VDD.n3714 23.1255
R29867 VDD.n3800 VDD.n3714 23.1255
R29868 VDD.n3794 VDD.n3726 23.1255
R29869 VDD.n3794 VDD.n3793 23.1255
R29870 VDD.n3731 VDD.n3727 23.1255
R29871 VDD.n3790 VDD.n3727 23.1255
R29872 VDD.n3784 VDD.n3737 23.1255
R29873 VDD.n3784 VDD.n3783 23.1255
R29874 VDD.n3742 VDD.n3738 23.1255
R29875 VDD.n3780 VDD.n3738 23.1255
R29876 VDD.n3774 VDD.n3747 23.1255
R29877 VDD.n3774 VDD.n3773 23.1255
R29878 VDD.n3752 VDD.n3748 23.1255
R29879 VDD.n3770 VDD.n3748 23.1255
R29880 VDD.n3764 VDD.n3760 23.1255
R29881 VDD.n3764 VDD.n3763 23.1255
R29882 VDD.n2934 VDD.n2930 23.1255
R29883 VDD.n3877 VDD.n3876 23.1255
R29884 VDD.n3876 VDD.n3875 23.1255
R29885 VDD.n3873 VDD.n3872 23.1255
R29886 VDD.n3874 VDD.n3873 23.1255
R29887 VDD.n3866 VDD.n3865 23.1255
R29888 VDD.n3867 VDD.n3866 23.1255
R29889 VDD.n3863 VDD.n3862 23.1255
R29890 VDD.n3864 VDD.n3863 23.1255
R29891 VDD.n3856 VDD.n3855 23.1255
R29892 VDD.n3857 VDD.n3856 23.1255
R29893 VDD.n3853 VDD.n3852 23.1255
R29894 VDD.n3854 VDD.n3853 23.1255
R29895 VDD.n3846 VDD.n3845 23.1255
R29896 VDD.n3847 VDD.n3846 23.1255
R29897 VDD.n3843 VDD.n3842 23.1255
R29898 VDD.n3844 VDD.n3843 23.1255
R29899 VDD.n3836 VDD.n3835 23.1255
R29900 VDD.n3837 VDD.n3836 23.1255
R29901 VDD.n3821 VDD.n3819 23.1255
R29902 VDD.n3819 VDD.n3694 23.1255
R29903 VDD.n3822 VDD.n3820 23.1255
R29904 VDD.n3820 VDD.n3818 23.1255
R29905 VDD.n3809 VDD.n3808 23.1255
R29906 VDD.n3810 VDD.n3809 23.1255
R29907 VDD.n3802 VDD.n3801 23.1255
R29908 VDD.n3803 VDD.n3802 23.1255
R29909 VDD.n3799 VDD.n3798 23.1255
R29910 VDD.n3800 VDD.n3799 23.1255
R29911 VDD.n3792 VDD.n3791 23.1255
R29912 VDD.n3793 VDD.n3792 23.1255
R29913 VDD.n3789 VDD.n3788 23.1255
R29914 VDD.n3790 VDD.n3789 23.1255
R29915 VDD.n3782 VDD.n3781 23.1255
R29916 VDD.n3783 VDD.n3782 23.1255
R29917 VDD.n3779 VDD.n3778 23.1255
R29918 VDD.n3780 VDD.n3779 23.1255
R29919 VDD.n3772 VDD.n3771 23.1255
R29920 VDD.n3773 VDD.n3772 23.1255
R29921 VDD.n3769 VDD.n3768 23.1255
R29922 VDD.n3770 VDD.n3769 23.1255
R29923 VDD.n3762 VDD.n3761 23.1255
R29924 VDD.n3763 VDD.n3762 23.1255
R29925 VDD.n3692 VDD.n3691 23.1255
R29926 VDD.n3693 VDD.n3692 23.1255
R29927 VDD.n3833 VDD.n3832 23.1255
R29928 VDD.n3834 VDD.n3833 23.1255
R29929 VDD.n265 VDD.n246 21.3068
R29930 VDD.n265 VDD.n264 21.3068
R29931 VDD.n267 VDD.t463 20.9643
R29932 VDD.n272 VDD.n271 20.7726
R29933 VDD.n275 VDD.n274 20.7726
R29934 VDD VDD.n3245 19.2885
R29935 VDD.n3134 VDD 18.5394
R29936 VDD.n241 VDD.t702 18.427
R29937 VDD.n241 VDD.t700 18.427
R29938 VDD.n3109 VDD.n3108 15.5222
R29939 VDD.n3173 VDD.n3172 15.5222
R29940 VDD.n3197 VDD.n3196 15.5222
R29941 VDD.n3574 VDD.n3573 15.5222
R29942 VDD.n3031 VDD.n3030 15.5222
R29943 VDD.n3618 VDD.n3617 15.5222
R29944 VDD.n3641 VDD.n3640 15.5222
R29945 VDD.n3128 VDD.n3127 15.5222
R29946 VDD.n3662 VDD.n3661 15.5222
R29947 VDD.n3485 VDD 14.6853
R29948 VDD.n281 VDD.n280 11.8208
R29949 VDD.n7071 VDD.n7070 10.9545
R29950 VDD VDD.n3240 9.59289
R29951 VDD.n3390 VDD 9.58202
R29952 VDD VDD.n3391 9.58202
R29953 VDD.n3485 VDD 9.58202
R29954 VDD.n1841 VDD.n1840 9.00833
R29955 VDD.n1581 VDD.n1580 9.00833
R29956 VDD.n1321 VDD.n1320 9.00833
R29957 VDD.n1061 VDD.n1060 9.00833
R29958 VDD.n801 VDD.n800 9.00833
R29959 VDD.n541 VDD.n540 9.00833
R29960 VDD.n7457 VDD.n7456 9.00833
R29961 VDD.n7459 VDD.n7458 9.00833
R29962 VDD.n3362 VDD.n3361 8.94311
R29963 VDD.n3400 VDD.n3254 8.94311
R29964 VDD.n3455 VDD.n3454 8.94311
R29965 VDD.n3457 VDD.n3456 8.94311
R29966 VDD.n3494 VDD.n3204 8.94311
R29967 VDD.n3360 VDD.n3359 8.94311
R29968 VDD.n3559 VDD.n3558 8.94311
R29969 VDD.n3094 VDD.n3081 8.48148
R29970 VDD.n3158 VDD.n3145 8.48148
R29971 VDD.n3055 VDD.n3042 8.48148
R29972 VDD.n3309 VDD.n3296 8.48148
R29973 VDD.n3016 VDD.n3003 8.48148
R29974 VDD.n3603 VDD.n3590 8.48148
R29975 VDD.n2996 VDD.n2983 8.48148
R29976 VDD.n3074 VDD.n3061 8.48148
R29977 VDD VDD.n3282 8.38365
R29978 VDD.n2995 VDD.n2988 8.26552
R29979 VDD.n7070 VDD.n7069 7.9105
R29980 VDD.n3341 VDD.n3281 7.9105
R29981 VDD.n3428 VDD.n3427 7.9105
R29982 VDD.n3442 VDD.n3441 7.9105
R29983 VDD.n3436 VDD.n3244 7.9105
R29984 VDD.n3522 VDD.n3521 7.9105
R29985 VDD.n3347 VDD.n3346 7.9105
R29986 VDD.n3531 VDD.n3530 7.9105
R29987 VDD.n3667 VDD.n3666 7.9105
R29988 VDD.n3645 VDD.n2841 7.9105
R29989 VDD.n3622 VDD.n2705 7.9105
R29990 VDD.n3035 VDD.n2569 7.9105
R29991 VDD.n3578 VDD.n2433 7.9105
R29992 VDD.n3201 VDD.n2297 7.9105
R29993 VDD.n3177 VDD.n2161 7.9105
R29994 VDD.n3113 VDD.n2025 7.9105
R29995 VDD.n3132 VDD.n1889 7.9105
R29996 VDD.n3093 VDD 7.85707
R29997 VDD.n3109 VDD 7.85707
R29998 VDD.n3157 VDD 7.85707
R29999 VDD.n3173 VDD 7.85707
R30000 VDD.n3054 VDD 7.85707
R30001 VDD.n3197 VDD 7.85707
R30002 VDD.n3308 VDD 7.85707
R30003 VDD.n3574 VDD 7.85707
R30004 VDD.n3015 VDD 7.85707
R30005 VDD.n3031 VDD 7.85707
R30006 VDD.n3602 VDD 7.85707
R30007 VDD.n3618 VDD 7.85707
R30008 VDD.n3641 VDD 7.85707
R30009 VDD.n3073 VDD 7.85707
R30010 VDD.n3128 VDD 7.85707
R30011 VDD.n3662 VDD 7.85707
R30012 VDD.n7606 VDD.n7605 7.39606
R30013 VDD.n7605 VDD.n7596 7.39606
R30014 VDD.n7616 VDD.n7615 7.39606
R30015 VDD.n7615 VDD.n7583 7.39606
R30016 VDD.n7626 VDD.n7625 7.39606
R30017 VDD.n7625 VDD.n7573 7.39606
R30018 VDD.n7636 VDD.n7635 7.39606
R30019 VDD.n7635 VDD.n7562 7.39606
R30020 VDD.n7646 VDD.n7645 7.39606
R30021 VDD.n7645 VDD.n7549 7.39606
R30022 VDD.n7663 VDD.n7662 7.39606
R30023 VDD.n7662 VDD.n7534 7.39606
R30024 VDD.n7673 VDD.n7672 7.39606
R30025 VDD.n7672 VDD.n7521 7.39606
R30026 VDD.n7683 VDD.n7682 7.39606
R30027 VDD.n7682 VDD.n7511 7.39606
R30028 VDD.n7693 VDD.n7692 7.39606
R30029 VDD.n7692 VDD.n7500 7.39606
R30030 VDD.n7703 VDD.n7702 7.39606
R30031 VDD.n7702 VDD.n7487 7.39606
R30032 VDD.n7715 VDD.n7462 7.39606
R30033 VDD.n7715 VDD.n7464 7.39606
R30034 VDD.n1724 VDD.n1723 7.39606
R30035 VDD.n1723 VDD.n1714 7.39606
R30036 VDD.n1734 VDD.n1733 7.39606
R30037 VDD.n1733 VDD.n1701 7.39606
R30038 VDD.n1744 VDD.n1743 7.39606
R30039 VDD.n1743 VDD.n1691 7.39606
R30040 VDD.n1754 VDD.n1753 7.39606
R30041 VDD.n1753 VDD.n1680 7.39606
R30042 VDD.n1764 VDD.n1763 7.39606
R30043 VDD.n1763 VDD.n1667 7.39606
R30044 VDD.n1781 VDD.n1780 7.39606
R30045 VDD.n1780 VDD.n1652 7.39606
R30046 VDD.n1791 VDD.n1790 7.39606
R30047 VDD.n1790 VDD.n1639 7.39606
R30048 VDD.n1801 VDD.n1800 7.39606
R30049 VDD.n1800 VDD.n1629 7.39606
R30050 VDD.n1811 VDD.n1810 7.39606
R30051 VDD.n1810 VDD.n1618 7.39606
R30052 VDD.n1821 VDD.n1820 7.39606
R30053 VDD.n1820 VDD.n1605 7.39606
R30054 VDD.n1831 VDD.n1830 7.39606
R30055 VDD.n1830 VDD.n1595 7.39606
R30056 VDD.n1464 VDD.n1463 7.39606
R30057 VDD.n1463 VDD.n1454 7.39606
R30058 VDD.n1474 VDD.n1473 7.39606
R30059 VDD.n1473 VDD.n1441 7.39606
R30060 VDD.n1484 VDD.n1483 7.39606
R30061 VDD.n1483 VDD.n1431 7.39606
R30062 VDD.n1494 VDD.n1493 7.39606
R30063 VDD.n1493 VDD.n1420 7.39606
R30064 VDD.n1504 VDD.n1503 7.39606
R30065 VDD.n1503 VDD.n1407 7.39606
R30066 VDD.n1521 VDD.n1520 7.39606
R30067 VDD.n1520 VDD.n1392 7.39606
R30068 VDD.n1531 VDD.n1530 7.39606
R30069 VDD.n1530 VDD.n1379 7.39606
R30070 VDD.n1541 VDD.n1540 7.39606
R30071 VDD.n1540 VDD.n1369 7.39606
R30072 VDD.n1551 VDD.n1550 7.39606
R30073 VDD.n1550 VDD.n1358 7.39606
R30074 VDD.n1561 VDD.n1560 7.39606
R30075 VDD.n1560 VDD.n1345 7.39606
R30076 VDD.n1571 VDD.n1570 7.39606
R30077 VDD.n1570 VDD.n1335 7.39606
R30078 VDD.n1204 VDD.n1203 7.39606
R30079 VDD.n1203 VDD.n1194 7.39606
R30080 VDD.n1214 VDD.n1213 7.39606
R30081 VDD.n1213 VDD.n1181 7.39606
R30082 VDD.n1224 VDD.n1223 7.39606
R30083 VDD.n1223 VDD.n1171 7.39606
R30084 VDD.n1234 VDD.n1233 7.39606
R30085 VDD.n1233 VDD.n1160 7.39606
R30086 VDD.n1244 VDD.n1243 7.39606
R30087 VDD.n1243 VDD.n1147 7.39606
R30088 VDD.n1261 VDD.n1260 7.39606
R30089 VDD.n1260 VDD.n1132 7.39606
R30090 VDD.n1271 VDD.n1270 7.39606
R30091 VDD.n1270 VDD.n1119 7.39606
R30092 VDD.n1281 VDD.n1280 7.39606
R30093 VDD.n1280 VDD.n1109 7.39606
R30094 VDD.n1291 VDD.n1290 7.39606
R30095 VDD.n1290 VDD.n1098 7.39606
R30096 VDD.n1301 VDD.n1300 7.39606
R30097 VDD.n1300 VDD.n1085 7.39606
R30098 VDD.n1311 VDD.n1310 7.39606
R30099 VDD.n1310 VDD.n1075 7.39606
R30100 VDD.n944 VDD.n943 7.39606
R30101 VDD.n943 VDD.n934 7.39606
R30102 VDD.n954 VDD.n953 7.39606
R30103 VDD.n953 VDD.n921 7.39606
R30104 VDD.n964 VDD.n963 7.39606
R30105 VDD.n963 VDD.n911 7.39606
R30106 VDD.n974 VDD.n973 7.39606
R30107 VDD.n973 VDD.n900 7.39606
R30108 VDD.n984 VDD.n983 7.39606
R30109 VDD.n983 VDD.n887 7.39606
R30110 VDD.n1001 VDD.n1000 7.39606
R30111 VDD.n1000 VDD.n872 7.39606
R30112 VDD.n1011 VDD.n1010 7.39606
R30113 VDD.n1010 VDD.n859 7.39606
R30114 VDD.n1021 VDD.n1020 7.39606
R30115 VDD.n1020 VDD.n849 7.39606
R30116 VDD.n1031 VDD.n1030 7.39606
R30117 VDD.n1030 VDD.n838 7.39606
R30118 VDD.n1041 VDD.n1040 7.39606
R30119 VDD.n1040 VDD.n825 7.39606
R30120 VDD.n1051 VDD.n1050 7.39606
R30121 VDD.n1050 VDD.n815 7.39606
R30122 VDD.n684 VDD.n683 7.39606
R30123 VDD.n683 VDD.n674 7.39606
R30124 VDD.n694 VDD.n693 7.39606
R30125 VDD.n693 VDD.n661 7.39606
R30126 VDD.n704 VDD.n703 7.39606
R30127 VDD.n703 VDD.n651 7.39606
R30128 VDD.n714 VDD.n713 7.39606
R30129 VDD.n713 VDD.n640 7.39606
R30130 VDD.n724 VDD.n723 7.39606
R30131 VDD.n723 VDD.n627 7.39606
R30132 VDD.n741 VDD.n740 7.39606
R30133 VDD.n740 VDD.n612 7.39606
R30134 VDD.n751 VDD.n750 7.39606
R30135 VDD.n750 VDD.n599 7.39606
R30136 VDD.n761 VDD.n760 7.39606
R30137 VDD.n760 VDD.n589 7.39606
R30138 VDD.n771 VDD.n770 7.39606
R30139 VDD.n770 VDD.n578 7.39606
R30140 VDD.n781 VDD.n780 7.39606
R30141 VDD.n780 VDD.n565 7.39606
R30142 VDD.n791 VDD.n790 7.39606
R30143 VDD.n790 VDD.n555 7.39606
R30144 VDD.n424 VDD.n423 7.39606
R30145 VDD.n423 VDD.n414 7.39606
R30146 VDD.n434 VDD.n433 7.39606
R30147 VDD.n433 VDD.n401 7.39606
R30148 VDD.n444 VDD.n443 7.39606
R30149 VDD.n443 VDD.n391 7.39606
R30150 VDD.n454 VDD.n453 7.39606
R30151 VDD.n453 VDD.n380 7.39606
R30152 VDD.n464 VDD.n463 7.39606
R30153 VDD.n463 VDD.n367 7.39606
R30154 VDD.n481 VDD.n480 7.39606
R30155 VDD.n480 VDD.n352 7.39606
R30156 VDD.n491 VDD.n490 7.39606
R30157 VDD.n490 VDD.n339 7.39606
R30158 VDD.n501 VDD.n500 7.39606
R30159 VDD.n500 VDD.n329 7.39606
R30160 VDD.n511 VDD.n510 7.39606
R30161 VDD.n510 VDD.n318 7.39606
R30162 VDD.n521 VDD.n520 7.39606
R30163 VDD.n520 VDD.n305 7.39606
R30164 VDD.n531 VDD.n530 7.39606
R30165 VDD.n530 VDD.n295 7.39606
R30166 VDD.n7340 VDD.n7339 7.39606
R30167 VDD.n7339 VDD.n7330 7.39606
R30168 VDD.n7350 VDD.n7349 7.39606
R30169 VDD.n7349 VDD.n7317 7.39606
R30170 VDD.n7360 VDD.n7359 7.39606
R30171 VDD.n7359 VDD.n7307 7.39606
R30172 VDD.n7370 VDD.n7369 7.39606
R30173 VDD.n7369 VDD.n7296 7.39606
R30174 VDD.n7380 VDD.n7379 7.39606
R30175 VDD.n7379 VDD.n7283 7.39606
R30176 VDD.n7397 VDD.n7396 7.39606
R30177 VDD.n7396 VDD.n7268 7.39606
R30178 VDD.n7407 VDD.n7406 7.39606
R30179 VDD.n7406 VDD.n7255 7.39606
R30180 VDD.n7417 VDD.n7416 7.39606
R30181 VDD.n7416 VDD.n7245 7.39606
R30182 VDD.n7427 VDD.n7426 7.39606
R30183 VDD.n7426 VDD.n7234 7.39606
R30184 VDD.n7437 VDD.n7436 7.39606
R30185 VDD.n7436 VDD.n7221 7.39606
R30186 VDD.n7447 VDD.n7446 7.39606
R30187 VDD.n7446 VDD.n7211 7.39606
R30188 VDD.n7083 VDD.n7082 7.39606
R30189 VDD.n7082 VDD.n7073 7.39606
R30190 VDD.n7093 VDD.n7092 7.39606
R30191 VDD.n7092 VDD.n1966 7.39606
R30192 VDD.n7103 VDD.n7102 7.39606
R30193 VDD.n7102 VDD.n1956 7.39606
R30194 VDD.n7113 VDD.n7112 7.39606
R30195 VDD.n7112 VDD.n1945 7.39606
R30196 VDD.n7123 VDD.n7122 7.39606
R30197 VDD.n7122 VDD.n1932 7.39606
R30198 VDD.n7142 VDD.n1904 7.39606
R30199 VDD.n7142 VDD.n1906 7.39606
R30200 VDD.n7157 VDD.n7156 7.39606
R30201 VDD.n7156 VDD.n1890 7.39606
R30202 VDD.n7167 VDD.n7166 7.39606
R30203 VDD.n7166 VDD.n1878 7.39606
R30204 VDD.n7177 VDD.n7176 7.39606
R30205 VDD.n7176 VDD.n1865 7.39606
R30206 VDD.n7187 VDD.n7186 7.39606
R30207 VDD.n7186 VDD.n1855 7.39606
R30208 VDD.n7147 VDD.n7146 7.39606
R30209 VDD.n7146 VDD.n1899 7.39606
R30210 VDD.n5978 VDD.n5977 7.39606
R30211 VDD.n5977 VDD.n5955 7.39606
R30212 VDD.n5988 VDD.n5987 7.39606
R30213 VDD.n5987 VDD.n5945 7.39606
R30214 VDD.n5998 VDD.n5997 7.39606
R30215 VDD.n5997 VDD.n5932 7.39606
R30216 VDD.n6008 VDD.n6007 7.39606
R30217 VDD.n6007 VDD.n5921 7.39606
R30218 VDD.n6018 VDD.n6017 7.39606
R30219 VDD.n6017 VDD.n5911 7.39606
R30220 VDD.n6028 VDD.n6027 7.39606
R30221 VDD.n6027 VDD.n5898 7.39606
R30222 VDD.n6045 VDD.n6044 7.39606
R30223 VDD.n6044 VDD.n5883 7.39606
R30224 VDD.n6055 VDD.n6054 7.39606
R30225 VDD.n6054 VDD.n5870 7.39606
R30226 VDD.n6065 VDD.n6064 7.39606
R30227 VDD.n6064 VDD.n5859 7.39606
R30228 VDD.n6075 VDD.n6074 7.39606
R30229 VDD.n6074 VDD.n5849 7.39606
R30230 VDD.n6087 VDD.n5833 7.39606
R30231 VDD.n6087 VDD.n5835 7.39606
R30232 VDD.n6101 VDD.n6100 7.39606
R30233 VDD.n6100 VDD.n5819 7.39606
R30234 VDD.n6111 VDD.n6110 7.39606
R30235 VDD.n6110 VDD.n5809 7.39606
R30236 VDD.n6121 VDD.n6120 7.39606
R30237 VDD.n6120 VDD.n5796 7.39606
R30238 VDD.n6131 VDD.n6130 7.39606
R30239 VDD.n6130 VDD.n5785 7.39606
R30240 VDD.n6141 VDD.n6140 7.39606
R30241 VDD.n6140 VDD.n5775 7.39606
R30242 VDD.n6151 VDD.n6150 7.39606
R30243 VDD.n6150 VDD.n5762 7.39606
R30244 VDD.n6168 VDD.n6167 7.39606
R30245 VDD.n6167 VDD.n5747 7.39606
R30246 VDD.n6178 VDD.n6177 7.39606
R30247 VDD.n6177 VDD.n5734 7.39606
R30248 VDD.n6188 VDD.n6187 7.39606
R30249 VDD.n6187 VDD.n5723 7.39606
R30250 VDD.n6198 VDD.n6197 7.39606
R30251 VDD.n6197 VDD.n5713 7.39606
R30252 VDD.n6210 VDD.n5697 7.39606
R30253 VDD.n6210 VDD.n5699 7.39606
R30254 VDD.n6224 VDD.n6223 7.39606
R30255 VDD.n6223 VDD.n5683 7.39606
R30256 VDD.n6234 VDD.n6233 7.39606
R30257 VDD.n6233 VDD.n5673 7.39606
R30258 VDD.n6244 VDD.n6243 7.39606
R30259 VDD.n6243 VDD.n5660 7.39606
R30260 VDD.n6254 VDD.n6253 7.39606
R30261 VDD.n6253 VDD.n5649 7.39606
R30262 VDD.n6264 VDD.n6263 7.39606
R30263 VDD.n6263 VDD.n5639 7.39606
R30264 VDD.n6274 VDD.n6273 7.39606
R30265 VDD.n6273 VDD.n5626 7.39606
R30266 VDD.n6291 VDD.n6290 7.39606
R30267 VDD.n6290 VDD.n5611 7.39606
R30268 VDD.n6301 VDD.n6300 7.39606
R30269 VDD.n6300 VDD.n5598 7.39606
R30270 VDD.n6311 VDD.n6310 7.39606
R30271 VDD.n6310 VDD.n5587 7.39606
R30272 VDD.n6321 VDD.n6320 7.39606
R30273 VDD.n6320 VDD.n5577 7.39606
R30274 VDD.n6333 VDD.n5561 7.39606
R30275 VDD.n6333 VDD.n5563 7.39606
R30276 VDD.n6347 VDD.n6346 7.39606
R30277 VDD.n6346 VDD.n5547 7.39606
R30278 VDD.n6357 VDD.n6356 7.39606
R30279 VDD.n6356 VDD.n5537 7.39606
R30280 VDD.n6367 VDD.n6366 7.39606
R30281 VDD.n6366 VDD.n5524 7.39606
R30282 VDD.n6377 VDD.n6376 7.39606
R30283 VDD.n6376 VDD.n5513 7.39606
R30284 VDD.n6387 VDD.n6386 7.39606
R30285 VDD.n6386 VDD.n5503 7.39606
R30286 VDD.n6397 VDD.n6396 7.39606
R30287 VDD.n6396 VDD.n5490 7.39606
R30288 VDD.n6414 VDD.n6413 7.39606
R30289 VDD.n6413 VDD.n5475 7.39606
R30290 VDD.n6424 VDD.n6423 7.39606
R30291 VDD.n6423 VDD.n5462 7.39606
R30292 VDD.n6434 VDD.n6433 7.39606
R30293 VDD.n6433 VDD.n5451 7.39606
R30294 VDD.n6444 VDD.n6443 7.39606
R30295 VDD.n6443 VDD.n5441 7.39606
R30296 VDD.n6456 VDD.n5425 7.39606
R30297 VDD.n6456 VDD.n5427 7.39606
R30298 VDD.n6470 VDD.n6469 7.39606
R30299 VDD.n6469 VDD.n5411 7.39606
R30300 VDD.n6480 VDD.n6479 7.39606
R30301 VDD.n6479 VDD.n5401 7.39606
R30302 VDD.n6490 VDD.n6489 7.39606
R30303 VDD.n6489 VDD.n5388 7.39606
R30304 VDD.n6500 VDD.n6499 7.39606
R30305 VDD.n6499 VDD.n5377 7.39606
R30306 VDD.n6510 VDD.n6509 7.39606
R30307 VDD.n6509 VDD.n5367 7.39606
R30308 VDD.n6520 VDD.n6519 7.39606
R30309 VDD.n6519 VDD.n5354 7.39606
R30310 VDD.n6537 VDD.n6536 7.39606
R30311 VDD.n6536 VDD.n5339 7.39606
R30312 VDD.n6547 VDD.n6546 7.39606
R30313 VDD.n6546 VDD.n5326 7.39606
R30314 VDD.n6557 VDD.n6556 7.39606
R30315 VDD.n6556 VDD.n5315 7.39606
R30316 VDD.n6567 VDD.n6566 7.39606
R30317 VDD.n6566 VDD.n5305 7.39606
R30318 VDD.n6579 VDD.n5289 7.39606
R30319 VDD.n6579 VDD.n5291 7.39606
R30320 VDD.n6593 VDD.n6592 7.39606
R30321 VDD.n6592 VDD.n5275 7.39606
R30322 VDD.n6603 VDD.n6602 7.39606
R30323 VDD.n6602 VDD.n5265 7.39606
R30324 VDD.n6613 VDD.n6612 7.39606
R30325 VDD.n6612 VDD.n5252 7.39606
R30326 VDD.n6623 VDD.n6622 7.39606
R30327 VDD.n6622 VDD.n5241 7.39606
R30328 VDD.n6633 VDD.n6632 7.39606
R30329 VDD.n6632 VDD.n5231 7.39606
R30330 VDD.n6643 VDD.n6642 7.39606
R30331 VDD.n6642 VDD.n5218 7.39606
R30332 VDD.n6660 VDD.n6659 7.39606
R30333 VDD.n6659 VDD.n5203 7.39606
R30334 VDD.n6670 VDD.n6669 7.39606
R30335 VDD.n6669 VDD.n5190 7.39606
R30336 VDD.n6680 VDD.n6679 7.39606
R30337 VDD.n6679 VDD.n5179 7.39606
R30338 VDD.n6690 VDD.n6689 7.39606
R30339 VDD.n6689 VDD.n5169 7.39606
R30340 VDD.n6702 VDD.n5153 7.39606
R30341 VDD.n6702 VDD.n5155 7.39606
R30342 VDD.n6716 VDD.n6715 7.39606
R30343 VDD.n6715 VDD.n5139 7.39606
R30344 VDD.n6726 VDD.n6725 7.39606
R30345 VDD.n6725 VDD.n5129 7.39606
R30346 VDD.n6736 VDD.n6735 7.39606
R30347 VDD.n6735 VDD.n5116 7.39606
R30348 VDD.n6746 VDD.n6745 7.39606
R30349 VDD.n6745 VDD.n5105 7.39606
R30350 VDD.n6756 VDD.n6755 7.39606
R30351 VDD.n6755 VDD.n5095 7.39606
R30352 VDD.n6766 VDD.n6765 7.39606
R30353 VDD.n6765 VDD.n5082 7.39606
R30354 VDD.n6783 VDD.n6782 7.39606
R30355 VDD.n6782 VDD.n5067 7.39606
R30356 VDD.n6793 VDD.n6792 7.39606
R30357 VDD.n6792 VDD.n5054 7.39606
R30358 VDD.n6803 VDD.n6802 7.39606
R30359 VDD.n6802 VDD.n5043 7.39606
R30360 VDD.n6813 VDD.n6812 7.39606
R30361 VDD.n6812 VDD.n5033 7.39606
R30362 VDD.n6825 VDD.n5017 7.39606
R30363 VDD.n6825 VDD.n5019 7.39606
R30364 VDD.n5001 VDD.n4765 7.39606
R30365 VDD.n5002 VDD.n5001 7.39606
R30366 VDD.n4991 VDD.n4776 7.39606
R30367 VDD.n4992 VDD.n4991 7.39606
R30368 VDD.n4981 VDD.n4786 7.39606
R30369 VDD.n4982 VDD.n4981 7.39606
R30370 VDD.n4971 VDD.n4799 7.39606
R30371 VDD.n4972 VDD.n4971 7.39606
R30372 VDD.n4961 VDD.n4810 7.39606
R30373 VDD.n4962 VDD.n4961 7.39606
R30374 VDD.n4951 VDD.n4820 7.39606
R30375 VDD.n4952 VDD.n4951 7.39606
R30376 VDD.n4934 VDD.n4836 7.39606
R30377 VDD.n4935 VDD.n4934 7.39606
R30378 VDD.n4924 VDD.n4848 7.39606
R30379 VDD.n4925 VDD.n4924 7.39606
R30380 VDD.n4914 VDD.n4861 7.39606
R30381 VDD.n4915 VDD.n4914 7.39606
R30382 VDD.n4904 VDD.n4872 7.39606
R30383 VDD.n4905 VDD.n4904 7.39606
R30384 VDD.n4894 VDD.n4882 7.39606
R30385 VDD.n4895 VDD.n4894 7.39606
R30386 VDD.n4642 VDD.n4641 7.39606
R30387 VDD.n4641 VDD.n4632 7.39606
R30388 VDD.n4652 VDD.n4651 7.39606
R30389 VDD.n4651 VDD.n2102 7.39606
R30390 VDD.n4662 VDD.n4661 7.39606
R30391 VDD.n4661 VDD.n2092 7.39606
R30392 VDD.n4672 VDD.n4671 7.39606
R30393 VDD.n4671 VDD.n2081 7.39606
R30394 VDD.n4682 VDD.n4681 7.39606
R30395 VDD.n4681 VDD.n2068 7.39606
R30396 VDD.n4701 VDD.n2040 7.39606
R30397 VDD.n4701 VDD.n2042 7.39606
R30398 VDD.n4716 VDD.n4715 7.39606
R30399 VDD.n4715 VDD.n2026 7.39606
R30400 VDD.n4726 VDD.n4725 7.39606
R30401 VDD.n4725 VDD.n2014 7.39606
R30402 VDD.n4736 VDD.n4735 7.39606
R30403 VDD.n4735 VDD.n2001 7.39606
R30404 VDD.n4746 VDD.n4745 7.39606
R30405 VDD.n4745 VDD.n1991 7.39606
R30406 VDD.n4706 VDD.n4705 7.39606
R30407 VDD.n4705 VDD.n2035 7.39606
R30408 VDD.n4517 VDD.n4516 7.39606
R30409 VDD.n4516 VDD.n4507 7.39606
R30410 VDD.n4527 VDD.n4526 7.39606
R30411 VDD.n4526 VDD.n2238 7.39606
R30412 VDD.n4537 VDD.n4536 7.39606
R30413 VDD.n4536 VDD.n2228 7.39606
R30414 VDD.n4547 VDD.n4546 7.39606
R30415 VDD.n4546 VDD.n2217 7.39606
R30416 VDD.n4557 VDD.n4556 7.39606
R30417 VDD.n4556 VDD.n2204 7.39606
R30418 VDD.n4576 VDD.n2176 7.39606
R30419 VDD.n4576 VDD.n2178 7.39606
R30420 VDD.n4591 VDD.n4590 7.39606
R30421 VDD.n4590 VDD.n2162 7.39606
R30422 VDD.n4601 VDD.n4600 7.39606
R30423 VDD.n4600 VDD.n2150 7.39606
R30424 VDD.n4611 VDD.n4610 7.39606
R30425 VDD.n4610 VDD.n2137 7.39606
R30426 VDD.n4621 VDD.n4620 7.39606
R30427 VDD.n4620 VDD.n2127 7.39606
R30428 VDD.n4581 VDD.n4580 7.39606
R30429 VDD.n4580 VDD.n2171 7.39606
R30430 VDD.n4392 VDD.n4391 7.39606
R30431 VDD.n4391 VDD.n4382 7.39606
R30432 VDD.n4402 VDD.n4401 7.39606
R30433 VDD.n4401 VDD.n2374 7.39606
R30434 VDD.n4412 VDD.n4411 7.39606
R30435 VDD.n4411 VDD.n2364 7.39606
R30436 VDD.n4422 VDD.n4421 7.39606
R30437 VDD.n4421 VDD.n2353 7.39606
R30438 VDD.n4432 VDD.n4431 7.39606
R30439 VDD.n4431 VDD.n2340 7.39606
R30440 VDD.n4451 VDD.n2312 7.39606
R30441 VDD.n4451 VDD.n2314 7.39606
R30442 VDD.n4466 VDD.n4465 7.39606
R30443 VDD.n4465 VDD.n2298 7.39606
R30444 VDD.n4476 VDD.n4475 7.39606
R30445 VDD.n4475 VDD.n2286 7.39606
R30446 VDD.n4486 VDD.n4485 7.39606
R30447 VDD.n4485 VDD.n2273 7.39606
R30448 VDD.n4496 VDD.n4495 7.39606
R30449 VDD.n4495 VDD.n2263 7.39606
R30450 VDD.n4456 VDD.n4455 7.39606
R30451 VDD.n4455 VDD.n2307 7.39606
R30452 VDD.n4267 VDD.n4266 7.39606
R30453 VDD.n4266 VDD.n4257 7.39606
R30454 VDD.n4277 VDD.n4276 7.39606
R30455 VDD.n4276 VDD.n2510 7.39606
R30456 VDD.n4287 VDD.n4286 7.39606
R30457 VDD.n4286 VDD.n2500 7.39606
R30458 VDD.n4297 VDD.n4296 7.39606
R30459 VDD.n4296 VDD.n2489 7.39606
R30460 VDD.n4307 VDD.n4306 7.39606
R30461 VDD.n4306 VDD.n2476 7.39606
R30462 VDD.n4326 VDD.n2448 7.39606
R30463 VDD.n4326 VDD.n2450 7.39606
R30464 VDD.n4341 VDD.n4340 7.39606
R30465 VDD.n4340 VDD.n2434 7.39606
R30466 VDD.n4351 VDD.n4350 7.39606
R30467 VDD.n4350 VDD.n2422 7.39606
R30468 VDD.n4361 VDD.n4360 7.39606
R30469 VDD.n4360 VDD.n2409 7.39606
R30470 VDD.n4371 VDD.n4370 7.39606
R30471 VDD.n4370 VDD.n2399 7.39606
R30472 VDD.n4331 VDD.n4330 7.39606
R30473 VDD.n4330 VDD.n2443 7.39606
R30474 VDD.n4142 VDD.n4141 7.39606
R30475 VDD.n4141 VDD.n4132 7.39606
R30476 VDD.n4152 VDD.n4151 7.39606
R30477 VDD.n4151 VDD.n2646 7.39606
R30478 VDD.n4162 VDD.n4161 7.39606
R30479 VDD.n4161 VDD.n2636 7.39606
R30480 VDD.n4172 VDD.n4171 7.39606
R30481 VDD.n4171 VDD.n2625 7.39606
R30482 VDD.n4182 VDD.n4181 7.39606
R30483 VDD.n4181 VDD.n2612 7.39606
R30484 VDD.n4201 VDD.n2584 7.39606
R30485 VDD.n4201 VDD.n2586 7.39606
R30486 VDD.n4216 VDD.n4215 7.39606
R30487 VDD.n4215 VDD.n2570 7.39606
R30488 VDD.n4226 VDD.n4225 7.39606
R30489 VDD.n4225 VDD.n2558 7.39606
R30490 VDD.n4236 VDD.n4235 7.39606
R30491 VDD.n4235 VDD.n2545 7.39606
R30492 VDD.n4246 VDD.n4245 7.39606
R30493 VDD.n4245 VDD.n2535 7.39606
R30494 VDD.n4206 VDD.n4205 7.39606
R30495 VDD.n4205 VDD.n2579 7.39606
R30496 VDD.n4017 VDD.n4016 7.39606
R30497 VDD.n4016 VDD.n4007 7.39606
R30498 VDD.n4027 VDD.n4026 7.39606
R30499 VDD.n4026 VDD.n2782 7.39606
R30500 VDD.n4037 VDD.n4036 7.39606
R30501 VDD.n4036 VDD.n2772 7.39606
R30502 VDD.n4047 VDD.n4046 7.39606
R30503 VDD.n4046 VDD.n2761 7.39606
R30504 VDD.n4057 VDD.n4056 7.39606
R30505 VDD.n4056 VDD.n2748 7.39606
R30506 VDD.n4076 VDD.n2720 7.39606
R30507 VDD.n4076 VDD.n2722 7.39606
R30508 VDD.n4091 VDD.n4090 7.39606
R30509 VDD.n4090 VDD.n2706 7.39606
R30510 VDD.n4101 VDD.n4100 7.39606
R30511 VDD.n4100 VDD.n2694 7.39606
R30512 VDD.n4111 VDD.n4110 7.39606
R30513 VDD.n4110 VDD.n2681 7.39606
R30514 VDD.n4121 VDD.n4120 7.39606
R30515 VDD.n4120 VDD.n2671 7.39606
R30516 VDD.n4081 VDD.n4080 7.39606
R30517 VDD.n4080 VDD.n2715 7.39606
R30518 VDD.n3892 VDD.n3891 7.39606
R30519 VDD.n3891 VDD.n3882 7.39606
R30520 VDD.n3902 VDD.n3901 7.39606
R30521 VDD.n3901 VDD.n2918 7.39606
R30522 VDD.n3912 VDD.n3911 7.39606
R30523 VDD.n3911 VDD.n2908 7.39606
R30524 VDD.n3922 VDD.n3921 7.39606
R30525 VDD.n3921 VDD.n2897 7.39606
R30526 VDD.n3932 VDD.n3931 7.39606
R30527 VDD.n3931 VDD.n2884 7.39606
R30528 VDD.n3951 VDD.n2856 7.39606
R30529 VDD.n3951 VDD.n2858 7.39606
R30530 VDD.n3966 VDD.n3965 7.39606
R30531 VDD.n3965 VDD.n2842 7.39606
R30532 VDD.n3976 VDD.n3975 7.39606
R30533 VDD.n3975 VDD.n2830 7.39606
R30534 VDD.n3986 VDD.n3985 7.39606
R30535 VDD.n3985 VDD.n2817 7.39606
R30536 VDD.n3996 VDD.n3995 7.39606
R30537 VDD.n3995 VDD.n2807 7.39606
R30538 VDD.n3956 VDD.n3955 7.39606
R30539 VDD.n3955 VDD.n2851 7.39606
R30540 VDD.n3544 VDD.n3543 7.39606
R30541 VDD.n3543 VDD.n3222 7.39606
R30542 VDD.n3556 VDD.n3206 7.39606
R30543 VDD.n3556 VDD.n3208 7.39606
R30544 VDD.n3534 VDD.n3533 7.39606
R30545 VDD.n3533 VDD.n3231 7.39606
R30546 VDD.n3767 VDD.n3766 7.39606
R30547 VDD.n3766 VDD.n3757 7.39606
R30548 VDD.n3777 VDD.n3776 7.39606
R30549 VDD.n3776 VDD.n3744 7.39606
R30550 VDD.n3787 VDD.n3786 7.39606
R30551 VDD.n3786 VDD.n3734 7.39606
R30552 VDD.n3797 VDD.n3796 7.39606
R30553 VDD.n3796 VDD.n3723 7.39606
R30554 VDD.n3807 VDD.n3806 7.39606
R30555 VDD.n3806 VDD.n3710 7.39606
R30556 VDD.n3826 VDD.n3682 7.39606
R30557 VDD.n3826 VDD.n3684 7.39606
R30558 VDD.n3841 VDD.n3840 7.39606
R30559 VDD.n3840 VDD.n3668 7.39606
R30560 VDD.n3851 VDD.n3850 7.39606
R30561 VDD.n3850 VDD.n2966 7.39606
R30562 VDD.n3861 VDD.n3860 7.39606
R30563 VDD.n3860 VDD.n2953 7.39606
R30564 VDD.n3871 VDD.n3870 7.39606
R30565 VDD.n3870 VDD.n2943 7.39606
R30566 VDD.n3831 VDD.n3830 7.39606
R30567 VDD.n3830 VDD.n3677 7.39606
R30568 VDD.n102 VDD.t197 7.31106
R30569 VDD.t379 VDD.n97 7.31106
R30570 VDD.n116 VDD.t250 7.31106
R30571 VDD.t859 VDD.n81 7.31106
R30572 VDD.n137 VDD.t827 7.31106
R30573 VDD.t993 VDD.n72 7.31106
R30574 VDD.n151 VDD.t7 7.31106
R30575 VDD.t326 VDD.n56 7.31106
R30576 VDD.n172 VDD.t153 7.31106
R30577 VDD.t568 VDD.n47 7.31106
R30578 VDD.n186 VDD.t821 7.31106
R30579 VDD.t637 VDD.n31 7.31106
R30580 VDD.n207 VDD.t201 7.31106
R30581 VDD.t910 VDD.n22 7.31106
R30582 VDD.n221 VDD.t539 7.31106
R30583 VDD.t834 VDD.n6 7.31106
R30584 VDD.n6936 VDD.t694 7.31106
R30585 VDD.t329 VDD.n6931 7.31106
R30586 VDD.n6950 VDD.t1036 7.31106
R30587 VDD.t324 VDD.n6915 7.31106
R30588 VDD.n6971 VDD.t878 7.31106
R30589 VDD.t357 VDD.n6906 7.31106
R30590 VDD.n6985 VDD.t1012 7.31106
R30591 VDD.t576 VDD.n6890 7.31106
R30592 VDD.n7006 VDD.t905 7.31106
R30593 VDD.t582 VDD.n6881 7.31106
R30594 VDD.n7020 VDD.t1040 7.31106
R30595 VDD.t600 VDD.n6865 7.31106
R30596 VDD.n7041 VDD.t870 7.31106
R30597 VDD.t367 VDD.n6856 7.31106
R30598 VDD.n7055 VDD.t1008 7.31106
R30599 VDD.n6839 VDD.t589 7.31106
R30600 VDD.t384 VDD.n3368 7.31106
R30601 VDD.n3385 VDD.t307 7.31106
R30602 VDD.t990 VDD.n3406 7.31106
R30603 VDD.n3422 VDD.t618 7.31106
R30604 VDD.t464 VDD.n3261 7.31106
R30605 VDD.n3274 VDD.t381 7.31106
R30606 VDD.t405 VDD.n3463 7.31106
R30607 VDD.n3480 VDD.t867 7.31106
R30608 VDD.t640 VDD.n3500 7.31106
R30609 VDD.n3516 VDD.t966 7.31106
R30610 VDD.t211 VDD.n3317 7.31106
R30611 VDD.n3330 VDD.t533 7.31106
R30612 VDD VDD.n6703 7.20159
R30613 VDD VDD.n6580 7.20159
R30614 VDD VDD.n6457 7.20159
R30615 VDD VDD.n6334 7.20159
R30616 VDD VDD.n6211 7.20159
R30617 VDD VDD.n6088 7.20159
R30618 VDD.n3094 VDD.n3093 6.96517
R30619 VDD.n3158 VDD.n3157 6.96517
R30620 VDD.n3055 VDD.n3054 6.96517
R30621 VDD.n3309 VDD.n3308 6.96517
R30622 VDD.n3016 VDD.n3015 6.96517
R30623 VDD.n3603 VDD.n3602 6.96517
R30624 VDD.n2996 VDD.n2995 6.96517
R30625 VDD.n3074 VDD.n3073 6.96517
R30626 VDD VDD.n3880 6.79126
R30627 VDD VDD.n4005 6.79126
R30628 VDD VDD.n4130 6.79126
R30629 VDD VDD.n4255 6.79126
R30630 VDD VDD.n4380 6.79126
R30631 VDD VDD.n4505 6.79126
R30632 VDD VDD.n4630 6.79126
R30633 VDD.n3456 VDD.n3455 5.59193
R30634 VDD.n3626 VDD.n2996 5.50827
R30635 VDD.n3240 VDD 4.96789
R30636 VDD.n6827 VDD.n6826 4.92985
R30637 VDD.n266 VDD.n244 4.65539
R30638 VDD.n7071 VDD.n4755 4.51952
R30639 VDD.n3093 VDD.n3092 4.5005
R30640 VDD.n3110 VDD.n3109 4.5005
R30641 VDD.n3157 VDD.n3156 4.5005
R30642 VDD.n3174 VDD.n3173 4.5005
R30643 VDD.n3054 VDD.n3053 4.5005
R30644 VDD.n3198 VDD.n3197 4.5005
R30645 VDD.n3308 VDD.n3307 4.5005
R30646 VDD.n3575 VDD.n3574 4.5005
R30647 VDD.n3015 VDD.n3014 4.5005
R30648 VDD.n3032 VDD.n3031 4.5005
R30649 VDD.n3602 VDD.n3601 4.5005
R30650 VDD.n3619 VDD.n3618 4.5005
R30651 VDD.n2995 VDD.n2994 4.5005
R30652 VDD.n3642 VDD.n3641 4.5005
R30653 VDD.n3073 VDD.n3072 4.5005
R30654 VDD.n3129 VDD.n3128 4.5005
R30655 VDD.n3663 VDD.n3662 4.5005
R30656 VDD.n1581 VDD.n1321 4.44435
R30657 VDD.n3441 VDD.n3440 4.44122
R30658 VDD.n2976 VDD 4.43528
R30659 VDD.n2840 VDD 4.43528
R30660 VDD.n2704 VDD 4.43528
R30661 VDD.n2568 VDD 4.43528
R30662 VDD.n2432 VDD 4.43528
R30663 VDD.n2296 VDD 4.43528
R30664 VDD.n2160 VDD 4.43528
R30665 VDD.n2024 VDD 4.43528
R30666 VDD.n1888 VDD 4.43528
R30667 VDD.n7470 VDD.t943 4.27344
R30668 VDD.t939 VDD.n1587 4.27344
R30669 VDD.t852 VDD.n1327 4.27344
R30670 VDD.t976 VDD.n1067 4.27344
R30671 VDD.t941 VDD.n807 4.27344
R30672 VDD.t848 VDD.n547 4.27344
R30673 VDD.t978 VDD.n287 4.27344
R30674 VDD.t850 VDD.n7203 4.27344
R30675 VDD.t913 VDD.n1847 4.27344
R30676 VDD.n5962 VDD.t345 4.27344
R30677 VDD.n5826 VDD.t946 4.27344
R30678 VDD.n5690 VDD.t209 4.27344
R30679 VDD.n5554 VDD.t829 4.27344
R30680 VDD.n5418 VDD.t837 4.27344
R30681 VDD.n5282 VDD.t155 4.27344
R30682 VDD.n5146 VDD.t566 4.27344
R30683 VDD.n5008 VDD.t203 4.27344
R30684 VDD.t2 VDD.n1983 4.27344
R30685 VDD.t920 VDD.n2119 4.27344
R30686 VDD.t291 VDD.n2255 4.27344
R30687 VDD.t903 VDD.n2391 4.27344
R30688 VDD.t571 VDD.n2527 4.27344
R30689 VDD.t876 VDD.n2663 4.27344
R30690 VDD.t1102 VDD.n2799 4.27344
R30691 VDD.t696 VDD.n2935 4.27344
R30692 VDD.n3138 VDD.n3094 4.23927
R30693 VDD.n3179 VDD.n3158 4.23927
R30694 VDD.n3182 VDD.n3055 4.23927
R30695 VDD.n3310 VDD.n3309 4.23927
R30696 VDD.n3583 VDD.n3016 4.23927
R30697 VDD.n3624 VDD.n3603 4.23927
R30698 VDD.n3075 VDD.n3074 4.23927
R30699 VDD.n3362 VDD 3.73292
R30700 VDD.n3400 VDD 3.73292
R30701 VDD.n3454 VDD 3.73292
R30702 VDD.n3457 VDD 3.73292
R30703 VDD.n3494 VDD 3.73292
R30704 VDD.n3359 VDD 3.73292
R30705 VDD.n3558 VDD 3.73292
R30706 VDD.n3360 VDD.n3310 3.53255
R30707 VDD.n3134 VDD.n3133 3.473
R30708 VDD.n3625 VDD.n3624 3.4105
R30709 VDD.n3584 VDD.n3583 3.4105
R30710 VDD.n3310 VDD.n2997 3.4105
R30711 VDD.n3182 VDD.n3181 3.4105
R30712 VDD.n3180 VDD.n3179 3.4105
R30713 VDD.n3139 VDD.n3138 3.4105
R30714 VDD.n3137 VDD.n3136 3.4105
R30715 VDD.n3178 VDD.n3036 3.4105
R30716 VDD.n3203 VDD.n3202 3.4105
R30717 VDD.n3580 VDD.n3579 3.4105
R30718 VDD.n3582 VDD.n3581 3.4105
R30719 VDD.n3623 VDD.n2977 3.4105
R30720 VDD.n3647 VDD.n3646 3.4105
R30721 VDD.n267 VDD.n266 3.29941
R30722 VDD.n4894 VDD.n4893 3.15974
R30723 VDD.n3579 VDD.n3559 3.08605
R30724 VDD.n3679 VDD 3.063
R30725 VDD.n2853 VDD 3.063
R30726 VDD.n2717 VDD 3.063
R30727 VDD.n2581 VDD 3.063
R30728 VDD.n2445 VDD 3.063
R30729 VDD.n2309 VDD 3.063
R30730 VDD.n2173 VDD 3.063
R30731 VDD.n2037 VDD 3.063
R30732 VDD.n1901 VDD 3.063
R30733 VDD.n3559 VDD.n3204 2.797
R30734 VDD.n3456 VDD.n3204 2.79387
R30735 VDD.n3455 VDD.n3254 2.79387
R30736 VDD.n3361 VDD.n3254 2.79387
R30737 VDD.n801 VDD.n541 2.7876
R30738 VDD.n1061 VDD.n801 2.7876
R30739 VDD.n1321 VDD.n1061 2.7876
R30740 VDD.n1841 VDD.n1581 2.7876
R30741 VDD.n7458 VDD.n1841 2.7876
R30742 VDD.n7458 VDD.n7457 2.7876
R30743 VDD.n6838 VDD.n6837 2.73583
R30744 VDD.n7068 VDD 2.60011
R30745 VDD.n242 VDD.t703 2.59419
R30746 VDD.n3361 VDD.n3360 2.44842
R30747 VDD.n1839 VDD.n1838 2.3255
R30748 VDD.n1830 VDD.n1594 2.3255
R30749 VDD.n1820 VDD.n1604 2.3255
R30750 VDD.n1810 VDD.n1617 2.3255
R30751 VDD.n1800 VDD.n1628 2.3255
R30752 VDD.n1790 VDD.n1638 2.3255
R30753 VDD.n1780 VDD.n1651 2.3255
R30754 VDD.n1665 VDD.n1658 2.3255
R30755 VDD.n1763 VDD.n1666 2.3255
R30756 VDD.n1753 VDD.n1679 2.3255
R30757 VDD.n1743 VDD.n1690 2.3255
R30758 VDD.n1733 VDD.n1700 2.3255
R30759 VDD.n1723 VDD.n1713 2.3255
R30760 VDD.n1579 VDD.n1578 2.3255
R30761 VDD.n1570 VDD.n1334 2.3255
R30762 VDD.n1560 VDD.n1344 2.3255
R30763 VDD.n1550 VDD.n1357 2.3255
R30764 VDD.n1540 VDD.n1368 2.3255
R30765 VDD.n1530 VDD.n1378 2.3255
R30766 VDD.n1520 VDD.n1391 2.3255
R30767 VDD.n1405 VDD.n1398 2.3255
R30768 VDD.n1503 VDD.n1406 2.3255
R30769 VDD.n1493 VDD.n1419 2.3255
R30770 VDD.n1483 VDD.n1430 2.3255
R30771 VDD.n1473 VDD.n1440 2.3255
R30772 VDD.n1463 VDD.n1453 2.3255
R30773 VDD.n1319 VDD.n1318 2.3255
R30774 VDD.n1310 VDD.n1074 2.3255
R30775 VDD.n1300 VDD.n1084 2.3255
R30776 VDD.n1290 VDD.n1097 2.3255
R30777 VDD.n1280 VDD.n1108 2.3255
R30778 VDD.n1270 VDD.n1118 2.3255
R30779 VDD.n1260 VDD.n1131 2.3255
R30780 VDD.n1145 VDD.n1138 2.3255
R30781 VDD.n1243 VDD.n1146 2.3255
R30782 VDD.n1233 VDD.n1159 2.3255
R30783 VDD.n1223 VDD.n1170 2.3255
R30784 VDD.n1213 VDD.n1180 2.3255
R30785 VDD.n1203 VDD.n1193 2.3255
R30786 VDD.n1059 VDD.n1058 2.3255
R30787 VDD.n1050 VDD.n814 2.3255
R30788 VDD.n1040 VDD.n824 2.3255
R30789 VDD.n1030 VDD.n837 2.3255
R30790 VDD.n1020 VDD.n848 2.3255
R30791 VDD.n1010 VDD.n858 2.3255
R30792 VDD.n1000 VDD.n871 2.3255
R30793 VDD.n885 VDD.n878 2.3255
R30794 VDD.n983 VDD.n886 2.3255
R30795 VDD.n973 VDD.n899 2.3255
R30796 VDD.n963 VDD.n910 2.3255
R30797 VDD.n953 VDD.n920 2.3255
R30798 VDD.n943 VDD.n933 2.3255
R30799 VDD.n799 VDD.n798 2.3255
R30800 VDD.n790 VDD.n554 2.3255
R30801 VDD.n780 VDD.n564 2.3255
R30802 VDD.n770 VDD.n577 2.3255
R30803 VDD.n760 VDD.n588 2.3255
R30804 VDD.n750 VDD.n598 2.3255
R30805 VDD.n740 VDD.n611 2.3255
R30806 VDD.n625 VDD.n618 2.3255
R30807 VDD.n723 VDD.n626 2.3255
R30808 VDD.n713 VDD.n639 2.3255
R30809 VDD.n703 VDD.n650 2.3255
R30810 VDD.n693 VDD.n660 2.3255
R30811 VDD.n683 VDD.n673 2.3255
R30812 VDD.n539 VDD.n538 2.3255
R30813 VDD.n530 VDD.n294 2.3255
R30814 VDD.n520 VDD.n304 2.3255
R30815 VDD.n510 VDD.n317 2.3255
R30816 VDD.n500 VDD.n328 2.3255
R30817 VDD.n490 VDD.n338 2.3255
R30818 VDD.n480 VDD.n351 2.3255
R30819 VDD.n365 VDD.n358 2.3255
R30820 VDD.n463 VDD.n366 2.3255
R30821 VDD.n453 VDD.n379 2.3255
R30822 VDD.n443 VDD.n390 2.3255
R30823 VDD.n433 VDD.n400 2.3255
R30824 VDD.n423 VDD.n413 2.3255
R30825 VDD.n239 VDD.n238 2.3255
R30826 VDD.n13 VDD.n9 2.3255
R30827 VDD.n220 VDD.n219 2.3255
R30828 VDD.n218 VDD.n217 2.3255
R30829 VDD.n206 VDD.n205 2.3255
R30830 VDD.n204 VDD.n203 2.3255
R30831 VDD.n38 VDD.n34 2.3255
R30832 VDD.n185 VDD.n184 2.3255
R30833 VDD.n183 VDD.n182 2.3255
R30834 VDD.n171 VDD.n170 2.3255
R30835 VDD.n169 VDD.n168 2.3255
R30836 VDD.n63 VDD.n59 2.3255
R30837 VDD.n150 VDD.n149 2.3255
R30838 VDD.n148 VDD.n147 2.3255
R30839 VDD.n136 VDD.n135 2.3255
R30840 VDD.n134 VDD.n133 2.3255
R30841 VDD.n88 VDD.n84 2.3255
R30842 VDD.n115 VDD.n114 2.3255
R30843 VDD.n113 VDD.n112 2.3255
R30844 VDD.n101 VDD.n100 2.3255
R30845 VDD.n7455 VDD.n7454 2.3255
R30846 VDD.n7446 VDD.n7210 2.3255
R30847 VDD.n7436 VDD.n7220 2.3255
R30848 VDD.n7426 VDD.n7233 2.3255
R30849 VDD.n7416 VDD.n7244 2.3255
R30850 VDD.n7406 VDD.n7254 2.3255
R30851 VDD.n7396 VDD.n7267 2.3255
R30852 VDD.n7281 VDD.n7274 2.3255
R30853 VDD.n7379 VDD.n7282 2.3255
R30854 VDD.n7369 VDD.n7295 2.3255
R30855 VDD.n7359 VDD.n7306 2.3255
R30856 VDD.n7349 VDD.n7316 2.3255
R30857 VDD.n7339 VDD.n7329 2.3255
R30858 VDD.n7054 VDD.n7053 2.3255
R30859 VDD.n7052 VDD.n7051 2.3255
R30860 VDD.n7040 VDD.n7039 2.3255
R30861 VDD.n7038 VDD.n7037 2.3255
R30862 VDD.n6872 VDD.n6868 2.3255
R30863 VDD.n7019 VDD.n7018 2.3255
R30864 VDD.n7017 VDD.n7016 2.3255
R30865 VDD.n7005 VDD.n7004 2.3255
R30866 VDD.n7003 VDD.n7002 2.3255
R30867 VDD.n6897 VDD.n6893 2.3255
R30868 VDD.n6984 VDD.n6983 2.3255
R30869 VDD.n6982 VDD.n6981 2.3255
R30870 VDD.n6970 VDD.n6969 2.3255
R30871 VDD.n6968 VDD.n6967 2.3255
R30872 VDD.n6922 VDD.n6918 2.3255
R30873 VDD.n6949 VDD.n6948 2.3255
R30874 VDD.n6947 VDD.n6946 2.3255
R30875 VDD.n6935 VDD.n6934 2.3255
R30876 VDD.n7067 VDD.n7066 2.3255
R30877 VDD.n6826 VDD.n6825 2.3255
R30878 VDD.n6812 VDD.n5032 2.3255
R30879 VDD.n6802 VDD.n5042 2.3255
R30880 VDD.n6792 VDD.n5053 2.3255
R30881 VDD.n6782 VDD.n5066 2.3255
R30882 VDD.n5079 VDD.n5073 2.3255
R30883 VDD.n6765 VDD.n5081 2.3255
R30884 VDD.n6755 VDD.n5094 2.3255
R30885 VDD.n6745 VDD.n5104 2.3255
R30886 VDD.n6735 VDD.n5115 2.3255
R30887 VDD.n6725 VDD.n5128 2.3255
R30888 VDD.n6715 VDD.n5138 2.3255
R30889 VDD.n6706 VDD.n6705 2.3255
R30890 VDD.n6703 VDD.n6702 2.3255
R30891 VDD.n6689 VDD.n5168 2.3255
R30892 VDD.n6679 VDD.n5178 2.3255
R30893 VDD.n6669 VDD.n5189 2.3255
R30894 VDD.n6659 VDD.n5202 2.3255
R30895 VDD.n5215 VDD.n5209 2.3255
R30896 VDD.n6642 VDD.n5217 2.3255
R30897 VDD.n6632 VDD.n5230 2.3255
R30898 VDD.n6622 VDD.n5240 2.3255
R30899 VDD.n6612 VDD.n5251 2.3255
R30900 VDD.n6602 VDD.n5264 2.3255
R30901 VDD.n6592 VDD.n5274 2.3255
R30902 VDD.n6583 VDD.n6582 2.3255
R30903 VDD.n6580 VDD.n6579 2.3255
R30904 VDD.n6566 VDD.n5304 2.3255
R30905 VDD.n6556 VDD.n5314 2.3255
R30906 VDD.n6546 VDD.n5325 2.3255
R30907 VDD.n6536 VDD.n5338 2.3255
R30908 VDD.n5351 VDD.n5345 2.3255
R30909 VDD.n6519 VDD.n5353 2.3255
R30910 VDD.n6509 VDD.n5366 2.3255
R30911 VDD.n6499 VDD.n5376 2.3255
R30912 VDD.n6489 VDD.n5387 2.3255
R30913 VDD.n6479 VDD.n5400 2.3255
R30914 VDD.n6469 VDD.n5410 2.3255
R30915 VDD.n6460 VDD.n6459 2.3255
R30916 VDD.n6457 VDD.n6456 2.3255
R30917 VDD.n6443 VDD.n5440 2.3255
R30918 VDD.n6433 VDD.n5450 2.3255
R30919 VDD.n6423 VDD.n5461 2.3255
R30920 VDD.n6413 VDD.n5474 2.3255
R30921 VDD.n5487 VDD.n5481 2.3255
R30922 VDD.n6396 VDD.n5489 2.3255
R30923 VDD.n6386 VDD.n5502 2.3255
R30924 VDD.n6376 VDD.n5512 2.3255
R30925 VDD.n6366 VDD.n5523 2.3255
R30926 VDD.n6356 VDD.n5536 2.3255
R30927 VDD.n6346 VDD.n5546 2.3255
R30928 VDD.n6337 VDD.n6336 2.3255
R30929 VDD.n6334 VDD.n6333 2.3255
R30930 VDD.n6320 VDD.n5576 2.3255
R30931 VDD.n6310 VDD.n5586 2.3255
R30932 VDD.n6300 VDD.n5597 2.3255
R30933 VDD.n6290 VDD.n5610 2.3255
R30934 VDD.n5623 VDD.n5617 2.3255
R30935 VDD.n6273 VDD.n5625 2.3255
R30936 VDD.n6263 VDD.n5638 2.3255
R30937 VDD.n6253 VDD.n5648 2.3255
R30938 VDD.n6243 VDD.n5659 2.3255
R30939 VDD.n6233 VDD.n5672 2.3255
R30940 VDD.n6223 VDD.n5682 2.3255
R30941 VDD.n6214 VDD.n6213 2.3255
R30942 VDD.n6211 VDD.n6210 2.3255
R30943 VDD.n6197 VDD.n5712 2.3255
R30944 VDD.n6187 VDD.n5722 2.3255
R30945 VDD.n6177 VDD.n5733 2.3255
R30946 VDD.n6167 VDD.n5746 2.3255
R30947 VDD.n5759 VDD.n5753 2.3255
R30948 VDD.n6150 VDD.n5761 2.3255
R30949 VDD.n6140 VDD.n5774 2.3255
R30950 VDD.n6130 VDD.n5784 2.3255
R30951 VDD.n6120 VDD.n5795 2.3255
R30952 VDD.n6110 VDD.n5808 2.3255
R30953 VDD.n6100 VDD.n5818 2.3255
R30954 VDD.n6091 VDD.n6090 2.3255
R30955 VDD.n6088 VDD.n6087 2.3255
R30956 VDD.n6074 VDD.n5848 2.3255
R30957 VDD.n6064 VDD.n5858 2.3255
R30958 VDD.n6054 VDD.n5869 2.3255
R30959 VDD.n6044 VDD.n5882 2.3255
R30960 VDD.n5895 VDD.n5889 2.3255
R30961 VDD.n6027 VDD.n5897 2.3255
R30962 VDD.n6017 VDD.n5910 2.3255
R30963 VDD.n6007 VDD.n5920 2.3255
R30964 VDD.n5997 VDD.n5931 2.3255
R30965 VDD.n5987 VDD.n5944 2.3255
R30966 VDD.n5977 VDD.n5954 2.3255
R30967 VDD.n5968 VDD.n5967 2.3255
R30968 VDD.n4904 VDD.n4873 2.3255
R30969 VDD.n4914 VDD.n4863 2.3255
R30970 VDD.n4924 VDD.n4852 2.3255
R30971 VDD.n4934 VDD.n4839 2.3255
R30972 VDD.n4838 VDD.n4830 2.3255
R30973 VDD.n4951 VDD.n4824 2.3255
R30974 VDD.n4961 VDD.n4811 2.3255
R30975 VDD.n4971 VDD.n4801 2.3255
R30976 VDD.n4981 VDD.n4790 2.3255
R30977 VDD.n4991 VDD.n4777 2.3255
R30978 VDD.n5001 VDD.n4767 2.3255
R30979 VDD.n5012 VDD.n5011 2.3255
R30980 VDD.n3375 VDD.n3374 2.3255
R30981 VDD.n3379 VDD.n3378 2.3255
R30982 VDD.n3413 VDD.n3412 2.3255
R30983 VDD.n3416 VDD.n3415 2.3255
R30984 VDD.n3453 VDD.n3452 2.3255
R30985 VDD.n3445 VDD.n3444 2.3255
R30986 VDD.n3470 VDD.n3469 2.3255
R30987 VDD.n3474 VDD.n3473 2.3255
R30988 VDD.n3507 VDD.n3506 2.3255
R30989 VDD.n3510 VDD.n3509 2.3255
R30990 VDD.n3358 VDD.n3357 2.3255
R30991 VDD.n3350 VDD.n3349 2.3255
R30992 VDD.n3334 VDD.n3333 2.3255
R30993 VDD.n3389 VDD.n3388 2.3255
R30994 VDD.n3426 VDD.n3425 2.3255
R30995 VDD.n3278 VDD.n3277 2.3255
R30996 VDD.n3484 VDD.n3483 2.3255
R30997 VDD.n3520 VDD.n3519 2.3255
R30998 VDD.n3533 VDD.n3532 2.3255
R30999 VDD.n3557 VDD.n3556 2.3255
R31000 VDD.n3543 VDD.n3221 2.3255
R31001 VDD.n3830 VDD.n3829 2.3255
R31002 VDD.n3827 VDD.n3826 2.3255
R31003 VDD.n3708 VDD.n3701 2.3255
R31004 VDD.n3806 VDD.n3709 2.3255
R31005 VDD.n3796 VDD.n3722 2.3255
R31006 VDD.n3786 VDD.n3733 2.3255
R31007 VDD.n3776 VDD.n3743 2.3255
R31008 VDD.n3766 VDD.n3756 2.3255
R31009 VDD.n3840 VDD.n3667 2.3255
R31010 VDD.n3955 VDD.n3954 2.3255
R31011 VDD.n3952 VDD.n3951 2.3255
R31012 VDD.n2882 VDD.n2875 2.3255
R31013 VDD.n3931 VDD.n2883 2.3255
R31014 VDD.n3921 VDD.n2896 2.3255
R31015 VDD.n3911 VDD.n2907 2.3255
R31016 VDD.n3901 VDD.n2917 2.3255
R31017 VDD.n3891 VDD.n3881 2.3255
R31018 VDD.n3879 VDD.n3878 2.3255
R31019 VDD.n3870 VDD.n2942 2.3255
R31020 VDD.n3860 VDD.n2952 2.3255
R31021 VDD.n3850 VDD.n2965 2.3255
R31022 VDD.n3965 VDD.n2841 2.3255
R31023 VDD.n4080 VDD.n4079 2.3255
R31024 VDD.n4077 VDD.n4076 2.3255
R31025 VDD.n2746 VDD.n2739 2.3255
R31026 VDD.n4056 VDD.n2747 2.3255
R31027 VDD.n4046 VDD.n2760 2.3255
R31028 VDD.n4036 VDD.n2771 2.3255
R31029 VDD.n4026 VDD.n2781 2.3255
R31030 VDD.n4016 VDD.n4006 2.3255
R31031 VDD.n4004 VDD.n4003 2.3255
R31032 VDD.n3995 VDD.n2806 2.3255
R31033 VDD.n3985 VDD.n2816 2.3255
R31034 VDD.n3975 VDD.n2829 2.3255
R31035 VDD.n4090 VDD.n2705 2.3255
R31036 VDD.n4205 VDD.n4204 2.3255
R31037 VDD.n4202 VDD.n4201 2.3255
R31038 VDD.n2610 VDD.n2603 2.3255
R31039 VDD.n4181 VDD.n2611 2.3255
R31040 VDD.n4171 VDD.n2624 2.3255
R31041 VDD.n4161 VDD.n2635 2.3255
R31042 VDD.n4151 VDD.n2645 2.3255
R31043 VDD.n4141 VDD.n4131 2.3255
R31044 VDD.n4129 VDD.n4128 2.3255
R31045 VDD.n4120 VDD.n2670 2.3255
R31046 VDD.n4110 VDD.n2680 2.3255
R31047 VDD.n4100 VDD.n2693 2.3255
R31048 VDD.n4215 VDD.n2569 2.3255
R31049 VDD.n4330 VDD.n4329 2.3255
R31050 VDD.n4327 VDD.n4326 2.3255
R31051 VDD.n2474 VDD.n2467 2.3255
R31052 VDD.n4306 VDD.n2475 2.3255
R31053 VDD.n4296 VDD.n2488 2.3255
R31054 VDD.n4286 VDD.n2499 2.3255
R31055 VDD.n4276 VDD.n2509 2.3255
R31056 VDD.n4266 VDD.n4256 2.3255
R31057 VDD.n4254 VDD.n4253 2.3255
R31058 VDD.n4245 VDD.n2534 2.3255
R31059 VDD.n4235 VDD.n2544 2.3255
R31060 VDD.n4225 VDD.n2557 2.3255
R31061 VDD.n4340 VDD.n2433 2.3255
R31062 VDD.n4455 VDD.n4454 2.3255
R31063 VDD.n4452 VDD.n4451 2.3255
R31064 VDD.n2338 VDD.n2331 2.3255
R31065 VDD.n4431 VDD.n2339 2.3255
R31066 VDD.n4421 VDD.n2352 2.3255
R31067 VDD.n4411 VDD.n2363 2.3255
R31068 VDD.n4401 VDD.n2373 2.3255
R31069 VDD.n4391 VDD.n4381 2.3255
R31070 VDD.n4379 VDD.n4378 2.3255
R31071 VDD.n4370 VDD.n2398 2.3255
R31072 VDD.n4360 VDD.n2408 2.3255
R31073 VDD.n4350 VDD.n2421 2.3255
R31074 VDD.n4465 VDD.n2297 2.3255
R31075 VDD.n4580 VDD.n4579 2.3255
R31076 VDD.n4577 VDD.n4576 2.3255
R31077 VDD.n2202 VDD.n2195 2.3255
R31078 VDD.n4556 VDD.n2203 2.3255
R31079 VDD.n4546 VDD.n2216 2.3255
R31080 VDD.n4536 VDD.n2227 2.3255
R31081 VDD.n4526 VDD.n2237 2.3255
R31082 VDD.n4516 VDD.n4506 2.3255
R31083 VDD.n4504 VDD.n4503 2.3255
R31084 VDD.n4495 VDD.n2262 2.3255
R31085 VDD.n4485 VDD.n2272 2.3255
R31086 VDD.n4475 VDD.n2285 2.3255
R31087 VDD.n4590 VDD.n2161 2.3255
R31088 VDD.n4705 VDD.n4704 2.3255
R31089 VDD.n4702 VDD.n4701 2.3255
R31090 VDD.n2066 VDD.n2059 2.3255
R31091 VDD.n4681 VDD.n2067 2.3255
R31092 VDD.n4671 VDD.n2080 2.3255
R31093 VDD.n4661 VDD.n2091 2.3255
R31094 VDD.n4651 VDD.n2101 2.3255
R31095 VDD.n4641 VDD.n4631 2.3255
R31096 VDD.n4629 VDD.n4628 2.3255
R31097 VDD.n4620 VDD.n2126 2.3255
R31098 VDD.n4610 VDD.n2136 2.3255
R31099 VDD.n4600 VDD.n2149 2.3255
R31100 VDD.n4715 VDD.n2025 2.3255
R31101 VDD.n4754 VDD.n4753 2.3255
R31102 VDD.n4745 VDD.n1990 2.3255
R31103 VDD.n4735 VDD.n2000 2.3255
R31104 VDD.n4725 VDD.n2013 2.3255
R31105 VDD.n7146 VDD.n7145 2.3255
R31106 VDD.n7143 VDD.n7142 2.3255
R31107 VDD.n1930 VDD.n1923 2.3255
R31108 VDD.n7122 VDD.n1931 2.3255
R31109 VDD.n7112 VDD.n1944 2.3255
R31110 VDD.n7102 VDD.n1955 2.3255
R31111 VDD.n7092 VDD.n1965 2.3255
R31112 VDD.n7082 VDD.n7072 2.3255
R31113 VDD.n7156 VDD.n1889 2.3255
R31114 VDD.n7195 VDD.n7194 2.3255
R31115 VDD.n7186 VDD.n1854 2.3255
R31116 VDD.n7176 VDD.n1864 2.3255
R31117 VDD.n7166 VDD.n1877 2.3255
R31118 VDD.n7473 VDD.n7460 2.3255
R31119 VDD.n7716 VDD.n7715 2.3255
R31120 VDD.n7702 VDD.n7461 2.3255
R31121 VDD.n7692 VDD.n7499 2.3255
R31122 VDD.n7682 VDD.n7510 2.3255
R31123 VDD.n7672 VDD.n7520 2.3255
R31124 VDD.n7662 VDD.n7533 2.3255
R31125 VDD.n7547 VDD.n7540 2.3255
R31126 VDD.n7645 VDD.n7548 2.3255
R31127 VDD.n7635 VDD.n7561 2.3255
R31128 VDD.n7625 VDD.n7572 2.3255
R31129 VDD.n7615 VDD.n7582 2.3255
R31130 VDD.n7605 VDD.n7595 2.3255
R31131 VDD.n6827 VDD 2.22333
R31132 VDD VDD.n7071 2.22333
R31133 VDD.n541 VDD.n281 1.71757
R31134 VDD.n1604 VDD.n1594 1.66898
R31135 VDD.n1638 VDD.n1628 1.66898
R31136 VDD.n1700 VDD.n1690 1.66898
R31137 VDD.n1344 VDD.n1334 1.66898
R31138 VDD.n1378 VDD.n1368 1.66898
R31139 VDD.n1440 VDD.n1430 1.66898
R31140 VDD.n1084 VDD.n1074 1.66898
R31141 VDD.n1118 VDD.n1108 1.66898
R31142 VDD.n1180 VDD.n1170 1.66898
R31143 VDD.n824 VDD.n814 1.66898
R31144 VDD.n858 VDD.n848 1.66898
R31145 VDD.n920 VDD.n910 1.66898
R31146 VDD.n564 VDD.n554 1.66898
R31147 VDD.n598 VDD.n588 1.66898
R31148 VDD.n660 VDD.n650 1.66898
R31149 VDD.n304 VDD.n294 1.66898
R31150 VDD.n338 VDD.n328 1.66898
R31151 VDD.n400 VDD.n390 1.66898
R31152 VDD.n7220 VDD.n7210 1.66898
R31153 VDD.n7254 VDD.n7244 1.66898
R31154 VDD.n7316 VDD.n7306 1.66898
R31155 VDD.n5042 VDD.n5032 1.66898
R31156 VDD.n5104 VDD.n5094 1.66898
R31157 VDD.n5138 VDD.n5128 1.66898
R31158 VDD.n5178 VDD.n5168 1.66898
R31159 VDD.n5240 VDD.n5230 1.66898
R31160 VDD.n5274 VDD.n5264 1.66898
R31161 VDD.n5314 VDD.n5304 1.66898
R31162 VDD.n5376 VDD.n5366 1.66898
R31163 VDD.n5410 VDD.n5400 1.66898
R31164 VDD.n5450 VDD.n5440 1.66898
R31165 VDD.n5512 VDD.n5502 1.66898
R31166 VDD.n5546 VDD.n5536 1.66898
R31167 VDD.n5586 VDD.n5576 1.66898
R31168 VDD.n5648 VDD.n5638 1.66898
R31169 VDD.n5682 VDD.n5672 1.66898
R31170 VDD.n5722 VDD.n5712 1.66898
R31171 VDD.n5784 VDD.n5774 1.66898
R31172 VDD.n5818 VDD.n5808 1.66898
R31173 VDD.n5858 VDD.n5848 1.66898
R31174 VDD.n5920 VDD.n5910 1.66898
R31175 VDD.n5954 VDD.n5944 1.66898
R31176 VDD.n4873 VDD.n4863 1.66898
R31177 VDD.n4811 VDD.n4801 1.66898
R31178 VDD.n4777 VDD.n4767 1.66898
R31179 VDD.n3743 VDD.n3733 1.66898
R31180 VDD.n2917 VDD.n2907 1.66898
R31181 VDD.n2952 VDD.n2942 1.66898
R31182 VDD.n2781 VDD.n2771 1.66898
R31183 VDD.n2816 VDD.n2806 1.66898
R31184 VDD.n2645 VDD.n2635 1.66898
R31185 VDD.n2680 VDD.n2670 1.66898
R31186 VDD.n2509 VDD.n2499 1.66898
R31187 VDD.n2544 VDD.n2534 1.66898
R31188 VDD.n2373 VDD.n2363 1.66898
R31189 VDD.n2408 VDD.n2398 1.66898
R31190 VDD.n2237 VDD.n2227 1.66898
R31191 VDD.n2272 VDD.n2262 1.66898
R31192 VDD.n2101 VDD.n2091 1.66898
R31193 VDD.n2136 VDD.n2126 1.66898
R31194 VDD.n2000 VDD.n1990 1.66898
R31195 VDD.n1965 VDD.n1955 1.66898
R31196 VDD.n1864 VDD.n1854 1.66898
R31197 VDD.n7716 VDD.n7461 1.66898
R31198 VDD.n7520 VDD.n7510 1.66898
R31199 VDD.n7582 VDD.n7572 1.66898
R31200 VDD.n3523 VDD.n3522 1.64628
R31201 VDD.n3436 VDD.n3435 1.64315
R31202 VDD.n3429 VDD.n3428 1.64315
R31203 VDD.n3341 VDD.n3340 1.64315
R31204 VDD.n3829 VDD.n3679 1.58202
R31205 VDD.n3954 VDD.n2853 1.58202
R31206 VDD.n4079 VDD.n2717 1.58202
R31207 VDD.n4204 VDD.n2581 1.58202
R31208 VDD.n4329 VDD.n2445 1.58202
R31209 VDD.n4454 VDD.n2309 1.58202
R31210 VDD.n4579 VDD.n2173 1.58202
R31211 VDD.n4704 VDD.n2037 1.58202
R31212 VDD.n7145 VDD.n1901 1.58202
R31213 VDD.n3377 VDD 1.53854
R31214 VDD.n3280 VDD 1.53854
R31215 VDD.n3443 VDD 1.53854
R31216 VDD.n3472 VDD 1.53854
R31217 VDD.n3243 VDD 1.53854
R31218 VDD.n3348 VDD 1.53854
R31219 VDD.n3241 VDD 1.53854
R31220 VDD.n242 VDD 1.50356
R31221 VDD.n3137 VDD.n3113 1.46377
R31222 VDD.n3178 VDD.n3177 1.46377
R31223 VDD.n3202 VDD.n3201 1.46377
R31224 VDD.n3579 VDD.n3578 1.46377
R31225 VDD.n3582 VDD.n3035 1.46377
R31226 VDD.n3623 VDD.n3622 1.46377
R31227 VDD.n3646 VDD.n3645 1.46377
R31228 VDD.n3133 VDD.n3132 1.46377
R31229 VDD.n240 VDD 1.33448
R31230 VDD.n7197 VDD 1.33448
R31231 VDD.n3346 VDD.n3345 1.2977
R31232 VDD.n3378 VDD.n3376 1.26409
R31233 VDD.n3415 VDD.n3414 1.26409
R31234 VDD.n3444 VDD.n3255 1.26409
R31235 VDD.n3473 VDD.n3471 1.26409
R31236 VDD.n3509 VDD.n3508 1.26409
R31237 VDD.n3349 VDD.n3311 1.26409
R31238 VDD.n3221 VDD.n3205 1.26409
R31239 VDD.n251 VDD.n245 1.22567
R31240 VDD.n251 VDD.n250 1.22567
R31241 VDD.n249 VDD.n247 1.22567
R31242 VDD.n254 VDD.n253 1.22567
R31243 VDD.n3083 VDD.n3082 1.19615
R31244 VDD.n3099 VDD.n3098 1.19615
R31245 VDD.n3147 VDD.n3146 1.19615
R31246 VDD.n3163 VDD.n3162 1.19615
R31247 VDD.n3044 VDD.n3043 1.19615
R31248 VDD.n3187 VDD.n3186 1.19615
R31249 VDD.n3298 VDD.n3297 1.19615
R31250 VDD.n3564 VDD.n3563 1.19615
R31251 VDD.n3005 VDD.n3004 1.19615
R31252 VDD.n3021 VDD.n3020 1.19615
R31253 VDD.n3592 VDD.n3591 1.19615
R31254 VDD.n3608 VDD.n3607 1.19615
R31255 VDD.n2986 VDD.n2985 1.19615
R31256 VDD.n3631 VDD.n3630 1.19615
R31257 VDD.n3063 VDD.n3062 1.19615
R31258 VDD.n3118 VDD.n3117 1.19615
R31259 VDD.n3652 VDD.n3651 1.19615
R31260 VDD.n278 VDD.n277 1.163
R31261 VDD.n3378 VDD.n3377 1.1418
R31262 VDD.n3415 VDD.n3280 1.1418
R31263 VDD.n3444 VDD.n3443 1.1418
R31264 VDD.n3473 VDD.n3472 1.1418
R31265 VDD.n3509 VDD.n3243 1.1418
R31266 VDD.n3349 VDD.n3348 1.1418
R31267 VDD.n3241 VDD.n3221 1.1418
R31268 VDD.n3088 VDD 1.09561
R31269 VDD.n3077 VDD 1.09561
R31270 VDD.n3104 VDD 1.09561
R31271 VDD.n3111 VDD 1.09561
R31272 VDD.n3152 VDD 1.09561
R31273 VDD.n3141 VDD 1.09561
R31274 VDD.n3168 VDD 1.09561
R31275 VDD.n3175 VDD 1.09561
R31276 VDD.n3049 VDD 1.09561
R31277 VDD.n3038 VDD 1.09561
R31278 VDD.n3192 VDD 1.09561
R31279 VDD.n3199 VDD 1.09561
R31280 VDD.n3303 VDD 1.09561
R31281 VDD.n3292 VDD 1.09561
R31282 VDD.n3569 VDD 1.09561
R31283 VDD.n3576 VDD 1.09561
R31284 VDD.n3010 VDD 1.09561
R31285 VDD.n2999 VDD 1.09561
R31286 VDD.n3026 VDD 1.09561
R31287 VDD.n3033 VDD 1.09561
R31288 VDD.n3597 VDD 1.09561
R31289 VDD.n3586 VDD 1.09561
R31290 VDD.n3613 VDD 1.09561
R31291 VDD.n3620 VDD 1.09561
R31292 VDD.n3636 VDD 1.09561
R31293 VDD.n3643 VDD 1.09561
R31294 VDD.n3068 VDD 1.09561
R31295 VDD.n3057 VDD 1.09561
R31296 VDD.n3123 VDD 1.09561
R31297 VDD.n3130 VDD 1.09561
R31298 VDD.n3657 VDD 1.09561
R31299 VDD.n3664 VDD 1.09561
R31300 VDD.n244 VDD 1.04639
R31301 VDD.n276 VDD.n275 1.02828
R31302 VDD.n272 VDD.n268 1.02828
R31303 VDD.n1839 VDD 1.01137
R31304 VDD VDD.n1617 1.01137
R31305 VDD VDD.n1651 1.01137
R31306 VDD VDD.n1665 1.01137
R31307 VDD.n1666 VDD 1.01137
R31308 VDD VDD.n1679 1.01137
R31309 VDD.n1713 VDD 1.01137
R31310 VDD.n1579 VDD 1.01137
R31311 VDD VDD.n1357 1.01137
R31312 VDD VDD.n1391 1.01137
R31313 VDD VDD.n1405 1.01137
R31314 VDD.n1406 VDD 1.01137
R31315 VDD VDD.n1419 1.01137
R31316 VDD.n1453 VDD 1.01137
R31317 VDD.n1319 VDD 1.01137
R31318 VDD VDD.n1097 1.01137
R31319 VDD VDD.n1131 1.01137
R31320 VDD VDD.n1145 1.01137
R31321 VDD.n1146 VDD 1.01137
R31322 VDD VDD.n1159 1.01137
R31323 VDD.n1193 VDD 1.01137
R31324 VDD.n1059 VDD 1.01137
R31325 VDD VDD.n837 1.01137
R31326 VDD VDD.n871 1.01137
R31327 VDD VDD.n885 1.01137
R31328 VDD.n886 VDD 1.01137
R31329 VDD VDD.n899 1.01137
R31330 VDD.n933 VDD 1.01137
R31331 VDD.n799 VDD 1.01137
R31332 VDD VDD.n577 1.01137
R31333 VDD VDD.n611 1.01137
R31334 VDD VDD.n625 1.01137
R31335 VDD.n626 VDD 1.01137
R31336 VDD VDD.n639 1.01137
R31337 VDD.n673 VDD 1.01137
R31338 VDD.n539 VDD 1.01137
R31339 VDD VDD.n317 1.01137
R31340 VDD VDD.n351 1.01137
R31341 VDD VDD.n365 1.01137
R31342 VDD.n366 VDD 1.01137
R31343 VDD VDD.n379 1.01137
R31344 VDD.n413 VDD 1.01137
R31345 VDD.n13 VDD 1.01137
R31346 VDD.n219 VDD 1.01137
R31347 VDD.n205 VDD 1.01137
R31348 VDD.n38 VDD 1.01137
R31349 VDD.n184 VDD 1.01137
R31350 VDD.n170 VDD 1.01137
R31351 VDD.n63 VDD 1.01137
R31352 VDD.n149 VDD 1.01137
R31353 VDD.n135 VDD 1.01137
R31354 VDD.n88 VDD 1.01137
R31355 VDD.n114 VDD 1.01137
R31356 VDD.n100 VDD 1.01137
R31357 VDD.n7455 VDD 1.01137
R31358 VDD VDD.n7233 1.01137
R31359 VDD VDD.n7267 1.01137
R31360 VDD VDD.n7281 1.01137
R31361 VDD.n7282 VDD 1.01137
R31362 VDD VDD.n7295 1.01137
R31363 VDD.n7329 VDD 1.01137
R31364 VDD.n7053 VDD 1.01137
R31365 VDD.n7039 VDD 1.01137
R31366 VDD.n6872 VDD 1.01137
R31367 VDD.n7018 VDD 1.01137
R31368 VDD.n7004 VDD 1.01137
R31369 VDD.n6897 VDD 1.01137
R31370 VDD.n6983 VDD 1.01137
R31371 VDD.n6969 VDD 1.01137
R31372 VDD.n6922 VDD 1.01137
R31373 VDD.n6948 VDD 1.01137
R31374 VDD.n6934 VDD 1.01137
R31375 VDD.n5053 VDD 1.01137
R31376 VDD VDD.n5066 1.01137
R31377 VDD.n5079 VDD 1.01137
R31378 VDD.n5081 VDD 1.01137
R31379 VDD.n5115 VDD 1.01137
R31380 VDD.n6705 VDD 1.01137
R31381 VDD.n5189 VDD 1.01137
R31382 VDD VDD.n5202 1.01137
R31383 VDD.n5215 VDD 1.01137
R31384 VDD.n5217 VDD 1.01137
R31385 VDD.n5251 VDD 1.01137
R31386 VDD.n6582 VDD 1.01137
R31387 VDD.n5325 VDD 1.01137
R31388 VDD VDD.n5338 1.01137
R31389 VDD.n5351 VDD 1.01137
R31390 VDD.n5353 VDD 1.01137
R31391 VDD.n5387 VDD 1.01137
R31392 VDD.n6459 VDD 1.01137
R31393 VDD.n5461 VDD 1.01137
R31394 VDD VDD.n5474 1.01137
R31395 VDD.n5487 VDD 1.01137
R31396 VDD.n5489 VDD 1.01137
R31397 VDD.n5523 VDD 1.01137
R31398 VDD.n6336 VDD 1.01137
R31399 VDD.n5597 VDD 1.01137
R31400 VDD VDD.n5610 1.01137
R31401 VDD.n5623 VDD 1.01137
R31402 VDD.n5625 VDD 1.01137
R31403 VDD.n5659 VDD 1.01137
R31404 VDD.n6213 VDD 1.01137
R31405 VDD.n5733 VDD 1.01137
R31406 VDD VDD.n5746 1.01137
R31407 VDD.n5759 VDD 1.01137
R31408 VDD.n5761 VDD 1.01137
R31409 VDD.n5795 VDD 1.01137
R31410 VDD.n6090 VDD 1.01137
R31411 VDD.n5869 VDD 1.01137
R31412 VDD VDD.n5882 1.01137
R31413 VDD.n5895 VDD 1.01137
R31414 VDD.n5897 VDD 1.01137
R31415 VDD.n5931 VDD 1.01137
R31416 VDD.n5967 VDD 1.01137
R31417 VDD VDD.n4852 1.01137
R31418 VDD.n4839 VDD 1.01137
R31419 VDD VDD.n4838 1.01137
R31420 VDD VDD.n4824 1.01137
R31421 VDD VDD.n4790 1.01137
R31422 VDD.n5012 VDD 1.01137
R31423 VDD.n3827 VDD 1.01137
R31424 VDD VDD.n3708 1.01137
R31425 VDD.n3709 VDD 1.01137
R31426 VDD VDD.n3722 1.01137
R31427 VDD.n3756 VDD 1.01137
R31428 VDD.n3952 VDD 1.01137
R31429 VDD VDD.n2882 1.01137
R31430 VDD.n2883 VDD 1.01137
R31431 VDD VDD.n2896 1.01137
R31432 VDD.n3881 VDD 1.01137
R31433 VDD.n3879 VDD 1.01137
R31434 VDD VDD.n2965 1.01137
R31435 VDD.n4077 VDD 1.01137
R31436 VDD VDD.n2746 1.01137
R31437 VDD.n2747 VDD 1.01137
R31438 VDD VDD.n2760 1.01137
R31439 VDD.n4006 VDD 1.01137
R31440 VDD.n4004 VDD 1.01137
R31441 VDD VDD.n2829 1.01137
R31442 VDD.n4202 VDD 1.01137
R31443 VDD VDD.n2610 1.01137
R31444 VDD.n2611 VDD 1.01137
R31445 VDD VDD.n2624 1.01137
R31446 VDD.n4131 VDD 1.01137
R31447 VDD.n4129 VDD 1.01137
R31448 VDD VDD.n2693 1.01137
R31449 VDD.n4327 VDD 1.01137
R31450 VDD VDD.n2474 1.01137
R31451 VDD.n2475 VDD 1.01137
R31452 VDD VDD.n2488 1.01137
R31453 VDD.n4256 VDD 1.01137
R31454 VDD.n4254 VDD 1.01137
R31455 VDD VDD.n2557 1.01137
R31456 VDD.n4452 VDD 1.01137
R31457 VDD VDD.n2338 1.01137
R31458 VDD.n2339 VDD 1.01137
R31459 VDD VDD.n2352 1.01137
R31460 VDD.n4381 VDD 1.01137
R31461 VDD.n4379 VDD 1.01137
R31462 VDD VDD.n2421 1.01137
R31463 VDD.n4577 VDD 1.01137
R31464 VDD VDD.n2202 1.01137
R31465 VDD.n2203 VDD 1.01137
R31466 VDD VDD.n2216 1.01137
R31467 VDD.n4506 VDD 1.01137
R31468 VDD.n4504 VDD 1.01137
R31469 VDD VDD.n2285 1.01137
R31470 VDD.n4702 VDD 1.01137
R31471 VDD VDD.n2066 1.01137
R31472 VDD.n2067 VDD 1.01137
R31473 VDD VDD.n2080 1.01137
R31474 VDD.n4631 VDD 1.01137
R31475 VDD.n4629 VDD 1.01137
R31476 VDD VDD.n2149 1.01137
R31477 VDD.n4754 VDD 1.01137
R31478 VDD VDD.n2013 1.01137
R31479 VDD.n7143 VDD 1.01137
R31480 VDD VDD.n1930 1.01137
R31481 VDD.n1931 VDD 1.01137
R31482 VDD VDD.n1944 1.01137
R31483 VDD.n7072 VDD 1.01137
R31484 VDD.n7195 VDD 1.01137
R31485 VDD VDD.n1877 1.01137
R31486 VDD VDD.n7460 1.01137
R31487 VDD VDD.n7499 1.01137
R31488 VDD VDD.n7533 1.01137
R31489 VDD VDD.n7547 1.01137
R31490 VDD.n7548 VDD 1.01137
R31491 VDD VDD.n7561 1.01137
R31492 VDD.n7595 VDD 1.01137
R31493 VDD.n3389 VDD 0.980969
R31494 VDD.n3426 VDD 0.980969
R31495 VDD.n3278 VDD 0.980969
R31496 VDD.n3484 VDD 0.980969
R31497 VDD.n3334 VDD 0.980969
R31498 VDD.n3532 VDD 0.980969
R31499 VDD.n3520 VDD 0.965885
R31500 VDD.n7068 VDD.n7067 0.938
R31501 VDD.n240 VDD.n239 0.845609
R31502 VDD.n3375 VDD.n3362 0.845609
R31503 VDD.n3413 VDD.n3400 0.845609
R31504 VDD.n3454 VDD.n3453 0.845609
R31505 VDD.n3470 VDD.n3457 0.845609
R31506 VDD.n3507 VDD.n3494 0.845609
R31507 VDD.n3359 VDD.n3358 0.845609
R31508 VDD.n3558 VDD.n3557 0.845609
R31509 VDD.n1616 VDD.n1604 0.834739
R31510 VDD.n1617 VDD.n1616 0.834739
R31511 VDD.n1650 VDD.n1638 0.834739
R31512 VDD.n1651 VDD.n1650 0.834739
R31513 VDD.n1678 VDD.n1666 0.834739
R31514 VDD.n1679 VDD.n1678 0.834739
R31515 VDD.n1712 VDD.n1700 0.834739
R31516 VDD.n1713 VDD.n1712 0.834739
R31517 VDD.n1356 VDD.n1344 0.834739
R31518 VDD.n1357 VDD.n1356 0.834739
R31519 VDD.n1390 VDD.n1378 0.834739
R31520 VDD.n1391 VDD.n1390 0.834739
R31521 VDD.n1418 VDD.n1406 0.834739
R31522 VDD.n1419 VDD.n1418 0.834739
R31523 VDD.n1452 VDD.n1440 0.834739
R31524 VDD.n1453 VDD.n1452 0.834739
R31525 VDD.n1096 VDD.n1084 0.834739
R31526 VDD.n1097 VDD.n1096 0.834739
R31527 VDD.n1130 VDD.n1118 0.834739
R31528 VDD.n1131 VDD.n1130 0.834739
R31529 VDD.n1158 VDD.n1146 0.834739
R31530 VDD.n1159 VDD.n1158 0.834739
R31531 VDD.n1192 VDD.n1180 0.834739
R31532 VDD.n1193 VDD.n1192 0.834739
R31533 VDD.n836 VDD.n824 0.834739
R31534 VDD.n837 VDD.n836 0.834739
R31535 VDD.n870 VDD.n858 0.834739
R31536 VDD.n871 VDD.n870 0.834739
R31537 VDD.n898 VDD.n886 0.834739
R31538 VDD.n899 VDD.n898 0.834739
R31539 VDD.n932 VDD.n920 0.834739
R31540 VDD.n933 VDD.n932 0.834739
R31541 VDD.n576 VDD.n564 0.834739
R31542 VDD.n577 VDD.n576 0.834739
R31543 VDD.n610 VDD.n598 0.834739
R31544 VDD.n611 VDD.n610 0.834739
R31545 VDD.n638 VDD.n626 0.834739
R31546 VDD.n639 VDD.n638 0.834739
R31547 VDD.n672 VDD.n660 0.834739
R31548 VDD.n673 VDD.n672 0.834739
R31549 VDD.n316 VDD.n304 0.834739
R31550 VDD.n317 VDD.n316 0.834739
R31551 VDD.n350 VDD.n338 0.834739
R31552 VDD.n351 VDD.n350 0.834739
R31553 VDD.n378 VDD.n366 0.834739
R31554 VDD.n379 VDD.n378 0.834739
R31555 VDD.n412 VDD.n400 0.834739
R31556 VDD.n413 VDD.n412 0.834739
R31557 VDD.n14 VDD.n13 0.834739
R31558 VDD.n219 VDD.n14 0.834739
R31559 VDD.n218 VDD.n16 0.834739
R31560 VDD.n205 VDD.n16 0.834739
R31561 VDD.n39 VDD.n38 0.834739
R31562 VDD.n184 VDD.n39 0.834739
R31563 VDD.n183 VDD.n41 0.834739
R31564 VDD.n170 VDD.n41 0.834739
R31565 VDD.n64 VDD.n63 0.834739
R31566 VDD.n149 VDD.n64 0.834739
R31567 VDD.n148 VDD.n66 0.834739
R31568 VDD.n135 VDD.n66 0.834739
R31569 VDD.n89 VDD.n88 0.834739
R31570 VDD.n114 VDD.n89 0.834739
R31571 VDD.n113 VDD.n91 0.834739
R31572 VDD.n100 VDD.n91 0.834739
R31573 VDD.n7232 VDD.n7220 0.834739
R31574 VDD.n7233 VDD.n7232 0.834739
R31575 VDD.n7266 VDD.n7254 0.834739
R31576 VDD.n7267 VDD.n7266 0.834739
R31577 VDD.n7294 VDD.n7282 0.834739
R31578 VDD.n7295 VDD.n7294 0.834739
R31579 VDD.n7328 VDD.n7316 0.834739
R31580 VDD.n7329 VDD.n7328 0.834739
R31581 VDD.n7067 VDD.n6830 0.834739
R31582 VDD.n7053 VDD.n6830 0.834739
R31583 VDD.n7052 VDD.n6850 0.834739
R31584 VDD.n7039 VDD.n6850 0.834739
R31585 VDD.n6873 VDD.n6872 0.834739
R31586 VDD.n7018 VDD.n6873 0.834739
R31587 VDD.n7017 VDD.n6875 0.834739
R31588 VDD.n7004 VDD.n6875 0.834739
R31589 VDD.n6898 VDD.n6897 0.834739
R31590 VDD.n6983 VDD.n6898 0.834739
R31591 VDD.n6982 VDD.n6900 0.834739
R31592 VDD.n6969 VDD.n6900 0.834739
R31593 VDD.n6923 VDD.n6922 0.834739
R31594 VDD.n6948 VDD.n6923 0.834739
R31595 VDD.n6947 VDD.n6925 0.834739
R31596 VDD.n6934 VDD.n6925 0.834739
R31597 VDD.n6826 VDD.n5016 0.834739
R31598 VDD.n5032 VDD.n5016 0.834739
R31599 VDD.n5065 VDD.n5053 0.834739
R31600 VDD.n5066 VDD.n5065 0.834739
R31601 VDD.n5093 VDD.n5081 0.834739
R31602 VDD.n5094 VDD.n5093 0.834739
R31603 VDD.n5127 VDD.n5115 0.834739
R31604 VDD.n5128 VDD.n5127 0.834739
R31605 VDD.n6703 VDD.n5152 0.834739
R31606 VDD.n5168 VDD.n5152 0.834739
R31607 VDD.n5201 VDD.n5189 0.834739
R31608 VDD.n5202 VDD.n5201 0.834739
R31609 VDD.n5229 VDD.n5217 0.834739
R31610 VDD.n5230 VDD.n5229 0.834739
R31611 VDD.n5263 VDD.n5251 0.834739
R31612 VDD.n5264 VDD.n5263 0.834739
R31613 VDD.n6580 VDD.n5288 0.834739
R31614 VDD.n5304 VDD.n5288 0.834739
R31615 VDD.n5337 VDD.n5325 0.834739
R31616 VDD.n5338 VDD.n5337 0.834739
R31617 VDD.n5365 VDD.n5353 0.834739
R31618 VDD.n5366 VDD.n5365 0.834739
R31619 VDD.n5399 VDD.n5387 0.834739
R31620 VDD.n5400 VDD.n5399 0.834739
R31621 VDD.n6457 VDD.n5424 0.834739
R31622 VDD.n5440 VDD.n5424 0.834739
R31623 VDD.n5473 VDD.n5461 0.834739
R31624 VDD.n5474 VDD.n5473 0.834739
R31625 VDD.n5501 VDD.n5489 0.834739
R31626 VDD.n5502 VDD.n5501 0.834739
R31627 VDD.n5535 VDD.n5523 0.834739
R31628 VDD.n5536 VDD.n5535 0.834739
R31629 VDD.n6334 VDD.n5560 0.834739
R31630 VDD.n5576 VDD.n5560 0.834739
R31631 VDD.n5609 VDD.n5597 0.834739
R31632 VDD.n5610 VDD.n5609 0.834739
R31633 VDD.n5637 VDD.n5625 0.834739
R31634 VDD.n5638 VDD.n5637 0.834739
R31635 VDD.n5671 VDD.n5659 0.834739
R31636 VDD.n5672 VDD.n5671 0.834739
R31637 VDD.n6211 VDD.n5696 0.834739
R31638 VDD.n5712 VDD.n5696 0.834739
R31639 VDD.n5745 VDD.n5733 0.834739
R31640 VDD.n5746 VDD.n5745 0.834739
R31641 VDD.n5773 VDD.n5761 0.834739
R31642 VDD.n5774 VDD.n5773 0.834739
R31643 VDD.n5807 VDD.n5795 0.834739
R31644 VDD.n5808 VDD.n5807 0.834739
R31645 VDD.n6088 VDD.n5832 0.834739
R31646 VDD.n5848 VDD.n5832 0.834739
R31647 VDD.n5881 VDD.n5869 0.834739
R31648 VDD.n5882 VDD.n5881 0.834739
R31649 VDD.n5909 VDD.n5897 0.834739
R31650 VDD.n5910 VDD.n5909 0.834739
R31651 VDD.n5943 VDD.n5931 0.834739
R31652 VDD.n5944 VDD.n5943 0.834739
R31653 VDD.n4893 VDD.n4873 0.834739
R31654 VDD.n4852 VDD.n4851 0.834739
R31655 VDD.n4851 VDD.n4839 0.834739
R31656 VDD.n4824 VDD.n4823 0.834739
R31657 VDD.n4823 VDD.n4811 0.834739
R31658 VDD.n4790 VDD.n4789 0.834739
R31659 VDD.n4789 VDD.n4777 0.834739
R31660 VDD.n3829 VDD.n3828 0.834739
R31661 VDD.n3828 VDD.n3827 0.834739
R31662 VDD.n3721 VDD.n3709 0.834739
R31663 VDD.n3722 VDD.n3721 0.834739
R31664 VDD.n3755 VDD.n3743 0.834739
R31665 VDD.n3756 VDD.n3755 0.834739
R31666 VDD.n3954 VDD.n3953 0.834739
R31667 VDD.n3953 VDD.n3952 0.834739
R31668 VDD.n2895 VDD.n2883 0.834739
R31669 VDD.n2896 VDD.n2895 0.834739
R31670 VDD.n2929 VDD.n2917 0.834739
R31671 VDD.n3881 VDD.n2929 0.834739
R31672 VDD.n2964 VDD.n2952 0.834739
R31673 VDD.n2965 VDD.n2964 0.834739
R31674 VDD.n4079 VDD.n4078 0.834739
R31675 VDD.n4078 VDD.n4077 0.834739
R31676 VDD.n2759 VDD.n2747 0.834739
R31677 VDD.n2760 VDD.n2759 0.834739
R31678 VDD.n2793 VDD.n2781 0.834739
R31679 VDD.n4006 VDD.n2793 0.834739
R31680 VDD.n2828 VDD.n2816 0.834739
R31681 VDD.n2829 VDD.n2828 0.834739
R31682 VDD.n4204 VDD.n4203 0.834739
R31683 VDD.n4203 VDD.n4202 0.834739
R31684 VDD.n2623 VDD.n2611 0.834739
R31685 VDD.n2624 VDD.n2623 0.834739
R31686 VDD.n2657 VDD.n2645 0.834739
R31687 VDD.n4131 VDD.n2657 0.834739
R31688 VDD.n2692 VDD.n2680 0.834739
R31689 VDD.n2693 VDD.n2692 0.834739
R31690 VDD.n4329 VDD.n4328 0.834739
R31691 VDD.n4328 VDD.n4327 0.834739
R31692 VDD.n2487 VDD.n2475 0.834739
R31693 VDD.n2488 VDD.n2487 0.834739
R31694 VDD.n2521 VDD.n2509 0.834739
R31695 VDD.n4256 VDD.n2521 0.834739
R31696 VDD.n2556 VDD.n2544 0.834739
R31697 VDD.n2557 VDD.n2556 0.834739
R31698 VDD.n4454 VDD.n4453 0.834739
R31699 VDD.n4453 VDD.n4452 0.834739
R31700 VDD.n2351 VDD.n2339 0.834739
R31701 VDD.n2352 VDD.n2351 0.834739
R31702 VDD.n2385 VDD.n2373 0.834739
R31703 VDD.n4381 VDD.n2385 0.834739
R31704 VDD.n2420 VDD.n2408 0.834739
R31705 VDD.n2421 VDD.n2420 0.834739
R31706 VDD.n4579 VDD.n4578 0.834739
R31707 VDD.n4578 VDD.n4577 0.834739
R31708 VDD.n2215 VDD.n2203 0.834739
R31709 VDD.n2216 VDD.n2215 0.834739
R31710 VDD.n2249 VDD.n2237 0.834739
R31711 VDD.n4506 VDD.n2249 0.834739
R31712 VDD.n2284 VDD.n2272 0.834739
R31713 VDD.n2285 VDD.n2284 0.834739
R31714 VDD.n4704 VDD.n4703 0.834739
R31715 VDD.n4703 VDD.n4702 0.834739
R31716 VDD.n2079 VDD.n2067 0.834739
R31717 VDD.n2080 VDD.n2079 0.834739
R31718 VDD.n2113 VDD.n2101 0.834739
R31719 VDD.n4631 VDD.n2113 0.834739
R31720 VDD.n2148 VDD.n2136 0.834739
R31721 VDD.n2149 VDD.n2148 0.834739
R31722 VDD.n2012 VDD.n2000 0.834739
R31723 VDD.n2013 VDD.n2012 0.834739
R31724 VDD.n7145 VDD.n7144 0.834739
R31725 VDD.n7144 VDD.n7143 0.834739
R31726 VDD.n1943 VDD.n1931 0.834739
R31727 VDD.n1944 VDD.n1943 0.834739
R31728 VDD.n1977 VDD.n1965 0.834739
R31729 VDD.n7072 VDD.n1977 0.834739
R31730 VDD.n1876 VDD.n1864 0.834739
R31731 VDD.n1877 VDD.n1876 0.834739
R31732 VDD.n7498 VDD.n7461 0.834739
R31733 VDD.n7499 VDD.n7498 0.834739
R31734 VDD.n7532 VDD.n7520 0.834739
R31735 VDD.n7533 VDD.n7532 0.834739
R31736 VDD.n7560 VDD.n7548 0.834739
R31737 VDD.n7561 VDD.n7560 0.834739
R31738 VDD.n7594 VDD.n7582 0.834739
R31739 VDD.n7595 VDD.n7594 0.834739
R31740 VDD.n1616 VDD.n1614 0.807565
R31741 VDD.n1616 VDD.n1615 0.807565
R31742 VDD.n1650 VDD.n1648 0.807565
R31743 VDD.n1650 VDD.n1649 0.807565
R31744 VDD.n1678 VDD.n1676 0.807565
R31745 VDD.n1678 VDD.n1677 0.807565
R31746 VDD.n1712 VDD.n1710 0.807565
R31747 VDD.n1712 VDD.n1711 0.807565
R31748 VDD.n1356 VDD.n1354 0.807565
R31749 VDD.n1356 VDD.n1355 0.807565
R31750 VDD.n1390 VDD.n1388 0.807565
R31751 VDD.n1390 VDD.n1389 0.807565
R31752 VDD.n1418 VDD.n1416 0.807565
R31753 VDD.n1418 VDD.n1417 0.807565
R31754 VDD.n1452 VDD.n1450 0.807565
R31755 VDD.n1452 VDD.n1451 0.807565
R31756 VDD.n1096 VDD.n1094 0.807565
R31757 VDD.n1096 VDD.n1095 0.807565
R31758 VDD.n1130 VDD.n1128 0.807565
R31759 VDD.n1130 VDD.n1129 0.807565
R31760 VDD.n1158 VDD.n1156 0.807565
R31761 VDD.n1158 VDD.n1157 0.807565
R31762 VDD.n1192 VDD.n1190 0.807565
R31763 VDD.n1192 VDD.n1191 0.807565
R31764 VDD.n836 VDD.n834 0.807565
R31765 VDD.n836 VDD.n835 0.807565
R31766 VDD.n870 VDD.n868 0.807565
R31767 VDD.n870 VDD.n869 0.807565
R31768 VDD.n898 VDD.n896 0.807565
R31769 VDD.n898 VDD.n897 0.807565
R31770 VDD.n932 VDD.n930 0.807565
R31771 VDD.n932 VDD.n931 0.807565
R31772 VDD.n576 VDD.n574 0.807565
R31773 VDD.n576 VDD.n575 0.807565
R31774 VDD.n610 VDD.n608 0.807565
R31775 VDD.n610 VDD.n609 0.807565
R31776 VDD.n638 VDD.n636 0.807565
R31777 VDD.n638 VDD.n637 0.807565
R31778 VDD.n672 VDD.n670 0.807565
R31779 VDD.n672 VDD.n671 0.807565
R31780 VDD.n316 VDD.n314 0.807565
R31781 VDD.n316 VDD.n315 0.807565
R31782 VDD.n350 VDD.n348 0.807565
R31783 VDD.n350 VDD.n349 0.807565
R31784 VDD.n378 VDD.n376 0.807565
R31785 VDD.n378 VDD.n377 0.807565
R31786 VDD.n412 VDD.n410 0.807565
R31787 VDD.n412 VDD.n411 0.807565
R31788 VDD.n266 VDD.n241 0.807565
R31789 VDD.n279 VDD.n278 0.807565
R31790 VDD.n91 VDD.n90 0.807565
R31791 VDD.n89 VDD.n87 0.807565
R31792 VDD.n66 VDD.n65 0.807565
R31793 VDD.n64 VDD.n62 0.807565
R31794 VDD.n41 VDD.n40 0.807565
R31795 VDD.n39 VDD.n37 0.807565
R31796 VDD.n16 VDD.n15 0.807565
R31797 VDD.n14 VDD.n12 0.807565
R31798 VDD.n7232 VDD.n7230 0.807565
R31799 VDD.n7232 VDD.n7231 0.807565
R31800 VDD.n7266 VDD.n7264 0.807565
R31801 VDD.n7266 VDD.n7265 0.807565
R31802 VDD.n7294 VDD.n7292 0.807565
R31803 VDD.n7294 VDD.n7293 0.807565
R31804 VDD.n7328 VDD.n7326 0.807565
R31805 VDD.n7328 VDD.n7327 0.807565
R31806 VDD.n6925 VDD.n6924 0.807565
R31807 VDD.n6923 VDD.n6921 0.807565
R31808 VDD.n6900 VDD.n6899 0.807565
R31809 VDD.n6898 VDD.n6896 0.807565
R31810 VDD.n6875 VDD.n6874 0.807565
R31811 VDD.n6873 VDD.n6871 0.807565
R31812 VDD.n6850 VDD.n6849 0.807565
R31813 VDD.n6830 VDD.n6829 0.807565
R31814 VDD.n5016 VDD.n5014 0.807565
R31815 VDD.n5016 VDD.n5015 0.807565
R31816 VDD.n5065 VDD.n5063 0.807565
R31817 VDD.n5065 VDD.n5064 0.807565
R31818 VDD.n5093 VDD.n5091 0.807565
R31819 VDD.n5093 VDD.n5092 0.807565
R31820 VDD.n5127 VDD.n5125 0.807565
R31821 VDD.n5127 VDD.n5126 0.807565
R31822 VDD.n5152 VDD.n5150 0.807565
R31823 VDD.n5152 VDD.n5151 0.807565
R31824 VDD.n5201 VDD.n5199 0.807565
R31825 VDD.n5201 VDD.n5200 0.807565
R31826 VDD.n5229 VDD.n5227 0.807565
R31827 VDD.n5229 VDD.n5228 0.807565
R31828 VDD.n5263 VDD.n5261 0.807565
R31829 VDD.n5263 VDD.n5262 0.807565
R31830 VDD.n5288 VDD.n5286 0.807565
R31831 VDD.n5288 VDD.n5287 0.807565
R31832 VDD.n5337 VDD.n5335 0.807565
R31833 VDD.n5337 VDD.n5336 0.807565
R31834 VDD.n5365 VDD.n5363 0.807565
R31835 VDD.n5365 VDD.n5364 0.807565
R31836 VDD.n5399 VDD.n5397 0.807565
R31837 VDD.n5399 VDD.n5398 0.807565
R31838 VDD.n5424 VDD.n5422 0.807565
R31839 VDD.n5424 VDD.n5423 0.807565
R31840 VDD.n5473 VDD.n5471 0.807565
R31841 VDD.n5473 VDD.n5472 0.807565
R31842 VDD.n5501 VDD.n5499 0.807565
R31843 VDD.n5501 VDD.n5500 0.807565
R31844 VDD.n5535 VDD.n5533 0.807565
R31845 VDD.n5535 VDD.n5534 0.807565
R31846 VDD.n5560 VDD.n5558 0.807565
R31847 VDD.n5560 VDD.n5559 0.807565
R31848 VDD.n5609 VDD.n5607 0.807565
R31849 VDD.n5609 VDD.n5608 0.807565
R31850 VDD.n5637 VDD.n5635 0.807565
R31851 VDD.n5637 VDD.n5636 0.807565
R31852 VDD.n5671 VDD.n5669 0.807565
R31853 VDD.n5671 VDD.n5670 0.807565
R31854 VDD.n5696 VDD.n5694 0.807565
R31855 VDD.n5696 VDD.n5695 0.807565
R31856 VDD.n5745 VDD.n5743 0.807565
R31857 VDD.n5745 VDD.n5744 0.807565
R31858 VDD.n5773 VDD.n5771 0.807565
R31859 VDD.n5773 VDD.n5772 0.807565
R31860 VDD.n5807 VDD.n5805 0.807565
R31861 VDD.n5807 VDD.n5806 0.807565
R31862 VDD.n5832 VDD.n5830 0.807565
R31863 VDD.n5832 VDD.n5831 0.807565
R31864 VDD.n5881 VDD.n5879 0.807565
R31865 VDD.n5881 VDD.n5880 0.807565
R31866 VDD.n5909 VDD.n5907 0.807565
R31867 VDD.n5909 VDD.n5908 0.807565
R31868 VDD.n5943 VDD.n5941 0.807565
R31869 VDD.n5943 VDD.n5942 0.807565
R31870 VDD.n4893 VDD.n4891 0.807565
R31871 VDD.n4893 VDD.n4892 0.807565
R31872 VDD.n4851 VDD.n4849 0.807565
R31873 VDD.n4851 VDD.n4850 0.807565
R31874 VDD.n4823 VDD.n4821 0.807565
R31875 VDD.n4823 VDD.n4822 0.807565
R31876 VDD.n4789 VDD.n4787 0.807565
R31877 VDD.n4789 VDD.n4788 0.807565
R31878 VDD.n3828 VDD.n3680 0.807565
R31879 VDD.n3828 VDD.n3681 0.807565
R31880 VDD.n3721 VDD.n3719 0.807565
R31881 VDD.n3721 VDD.n3720 0.807565
R31882 VDD.n3755 VDD.n3753 0.807565
R31883 VDD.n3755 VDD.n3754 0.807565
R31884 VDD.n3953 VDD.n2854 0.807565
R31885 VDD.n3953 VDD.n2855 0.807565
R31886 VDD.n2895 VDD.n2893 0.807565
R31887 VDD.n2895 VDD.n2894 0.807565
R31888 VDD.n2929 VDD.n2927 0.807565
R31889 VDD.n2929 VDD.n2928 0.807565
R31890 VDD.n2964 VDD.n2962 0.807565
R31891 VDD.n2964 VDD.n2963 0.807565
R31892 VDD.n4078 VDD.n2718 0.807565
R31893 VDD.n4078 VDD.n2719 0.807565
R31894 VDD.n2759 VDD.n2757 0.807565
R31895 VDD.n2759 VDD.n2758 0.807565
R31896 VDD.n2793 VDD.n2791 0.807565
R31897 VDD.n2793 VDD.n2792 0.807565
R31898 VDD.n2828 VDD.n2826 0.807565
R31899 VDD.n2828 VDD.n2827 0.807565
R31900 VDD.n4203 VDD.n2582 0.807565
R31901 VDD.n4203 VDD.n2583 0.807565
R31902 VDD.n2623 VDD.n2621 0.807565
R31903 VDD.n2623 VDD.n2622 0.807565
R31904 VDD.n2657 VDD.n2655 0.807565
R31905 VDD.n2657 VDD.n2656 0.807565
R31906 VDD.n2692 VDD.n2690 0.807565
R31907 VDD.n2692 VDD.n2691 0.807565
R31908 VDD.n4328 VDD.n2446 0.807565
R31909 VDD.n4328 VDD.n2447 0.807565
R31910 VDD.n2487 VDD.n2485 0.807565
R31911 VDD.n2487 VDD.n2486 0.807565
R31912 VDD.n2521 VDD.n2519 0.807565
R31913 VDD.n2521 VDD.n2520 0.807565
R31914 VDD.n2556 VDD.n2554 0.807565
R31915 VDD.n2556 VDD.n2555 0.807565
R31916 VDD.n4453 VDD.n2310 0.807565
R31917 VDD.n4453 VDD.n2311 0.807565
R31918 VDD.n2351 VDD.n2349 0.807565
R31919 VDD.n2351 VDD.n2350 0.807565
R31920 VDD.n2385 VDD.n2383 0.807565
R31921 VDD.n2385 VDD.n2384 0.807565
R31922 VDD.n2420 VDD.n2418 0.807565
R31923 VDD.n2420 VDD.n2419 0.807565
R31924 VDD.n4578 VDD.n2174 0.807565
R31925 VDD.n4578 VDD.n2175 0.807565
R31926 VDD.n2215 VDD.n2213 0.807565
R31927 VDD.n2215 VDD.n2214 0.807565
R31928 VDD.n2249 VDD.n2247 0.807565
R31929 VDD.n2249 VDD.n2248 0.807565
R31930 VDD.n2284 VDD.n2282 0.807565
R31931 VDD.n2284 VDD.n2283 0.807565
R31932 VDD.n4703 VDD.n2038 0.807565
R31933 VDD.n4703 VDD.n2039 0.807565
R31934 VDD.n2079 VDD.n2077 0.807565
R31935 VDD.n2079 VDD.n2078 0.807565
R31936 VDD.n2113 VDD.n2111 0.807565
R31937 VDD.n2113 VDD.n2112 0.807565
R31938 VDD.n2148 VDD.n2146 0.807565
R31939 VDD.n2148 VDD.n2147 0.807565
R31940 VDD.n2012 VDD.n2010 0.807565
R31941 VDD.n2012 VDD.n2011 0.807565
R31942 VDD.n7144 VDD.n1902 0.807565
R31943 VDD.n7144 VDD.n1903 0.807565
R31944 VDD.n1943 VDD.n1941 0.807565
R31945 VDD.n1943 VDD.n1942 0.807565
R31946 VDD.n1977 VDD.n1975 0.807565
R31947 VDD.n1977 VDD.n1976 0.807565
R31948 VDD.n1876 VDD.n1874 0.807565
R31949 VDD.n1876 VDD.n1875 0.807565
R31950 VDD.n7498 VDD.n7496 0.807565
R31951 VDD.n7498 VDD.n7497 0.807565
R31952 VDD.n7532 VDD.n7530 0.807565
R31953 VDD.n7532 VDD.n7531 0.807565
R31954 VDD.n7560 VDD.n7558 0.807565
R31955 VDD.n7560 VDD.n7559 0.807565
R31956 VDD.n7594 VDD.n7592 0.807565
R31957 VDD.n7594 VDD.n7593 0.807565
R31958 VDD.n3091 VDD.n3090 0.796696
R31959 VDD.n3080 VDD.n3079 0.796696
R31960 VDD.n3107 VDD.n3106 0.796696
R31961 VDD.n3097 VDD.n3096 0.796696
R31962 VDD.n3155 VDD.n3154 0.796696
R31963 VDD.n3144 VDD.n3143 0.796696
R31964 VDD.n3171 VDD.n3170 0.796696
R31965 VDD.n3161 VDD.n3160 0.796696
R31966 VDD.n3052 VDD.n3051 0.796696
R31967 VDD.n3041 VDD.n3040 0.796696
R31968 VDD.n3195 VDD.n3194 0.796696
R31969 VDD.n3185 VDD.n3184 0.796696
R31970 VDD.n3306 VDD.n3305 0.796696
R31971 VDD.n3295 VDD.n3294 0.796696
R31972 VDD.n3572 VDD.n3571 0.796696
R31973 VDD.n3562 VDD.n3561 0.796696
R31974 VDD.n3013 VDD.n3012 0.796696
R31975 VDD.n3002 VDD.n3001 0.796696
R31976 VDD.n3029 VDD.n3028 0.796696
R31977 VDD.n3019 VDD.n3018 0.796696
R31978 VDD.n3600 VDD.n3599 0.796696
R31979 VDD.n3589 VDD.n3588 0.796696
R31980 VDD.n3616 VDD.n3615 0.796696
R31981 VDD.n3606 VDD.n3605 0.796696
R31982 VDD.n2990 VDD.n2989 0.796696
R31983 VDD.n2979 VDD.n2978 0.796696
R31984 VDD.n3639 VDD.n3638 0.796696
R31985 VDD.n3629 VDD.n3628 0.796696
R31986 VDD.n3071 VDD.n3070 0.796696
R31987 VDD.n3060 VDD.n3059 0.796696
R31988 VDD.n3126 VDD.n3125 0.796696
R31989 VDD.n3116 VDD.n3115 0.796696
R31990 VDD.n3660 VDD.n3659 0.796696
R31991 VDD.n3650 VDD.n3649 0.796696
R31992 VDD.n3086 VDD.n3085 0.783833
R31993 VDD.n3102 VDD.n3101 0.783833
R31994 VDD.n3150 VDD.n3149 0.783833
R31995 VDD.n3166 VDD.n3165 0.783833
R31996 VDD.n3047 VDD.n3046 0.783833
R31997 VDD.n3190 VDD.n3189 0.783833
R31998 VDD.n3301 VDD.n3300 0.783833
R31999 VDD.n3567 VDD.n3566 0.783833
R32000 VDD.n3008 VDD.n3007 0.783833
R32001 VDD.n3024 VDD.n3023 0.783833
R32002 VDD.n3595 VDD.n3594 0.783833
R32003 VDD.n3611 VDD.n3610 0.783833
R32004 VDD.n2988 VDD.n2987 0.783833
R32005 VDD.n3634 VDD.n3633 0.783833
R32006 VDD.n3066 VDD.n3065 0.783833
R32007 VDD.n3121 VDD.n3120 0.783833
R32008 VDD.n3655 VDD.n3654 0.783833
R32009 VDD.n3085 VDD 0.716182
R32010 VDD.n3101 VDD 0.716182
R32011 VDD.n3149 VDD 0.716182
R32012 VDD.n3165 VDD 0.716182
R32013 VDD.n3046 VDD 0.716182
R32014 VDD.n3189 VDD 0.716182
R32015 VDD.n3300 VDD 0.716182
R32016 VDD.n3566 VDD 0.716182
R32017 VDD.n3007 VDD 0.716182
R32018 VDD.n3023 VDD 0.716182
R32019 VDD.n3594 VDD 0.716182
R32020 VDD.n3610 VDD 0.716182
R32021 VDD.n2988 VDD 0.716182
R32022 VDD.n3633 VDD 0.716182
R32023 VDD.n3065 VDD 0.716182
R32024 VDD.n3120 VDD 0.716182
R32025 VDD.n3654 VDD 0.716182
R32026 VDD.n243 VDD 0.685334
R32027 VDD.n3091 VDD 0.662609
R32028 VDD.n3080 VDD 0.662609
R32029 VDD.n3107 VDD 0.662609
R32030 VDD.n3097 VDD 0.662609
R32031 VDD.n3155 VDD 0.662609
R32032 VDD.n3144 VDD 0.662609
R32033 VDD.n3171 VDD 0.662609
R32034 VDD.n3161 VDD 0.662609
R32035 VDD.n3052 VDD 0.662609
R32036 VDD.n3041 VDD 0.662609
R32037 VDD.n3195 VDD 0.662609
R32038 VDD.n3185 VDD 0.662609
R32039 VDD.n3306 VDD 0.662609
R32040 VDD.n3295 VDD 0.662609
R32041 VDD.n3572 VDD 0.662609
R32042 VDD.n3562 VDD 0.662609
R32043 VDD.n3013 VDD 0.662609
R32044 VDD.n3002 VDD 0.662609
R32045 VDD.n3029 VDD 0.662609
R32046 VDD.n3019 VDD 0.662609
R32047 VDD.n3600 VDD 0.662609
R32048 VDD.n3589 VDD 0.662609
R32049 VDD.n3616 VDD 0.662609
R32050 VDD.n3606 VDD 0.662609
R32051 VDD.n3639 VDD 0.662609
R32052 VDD.n3629 VDD 0.662609
R32053 VDD.n3071 VDD 0.662609
R32054 VDD.n3060 VDD 0.662609
R32055 VDD.n3126 VDD 0.662609
R32056 VDD.n3116 VDD 0.662609
R32057 VDD.n3660 VDD 0.662609
R32058 VDD.n3650 VDD 0.662609
R32059 VDD.n3336 VDD.n3335 0.648317
R32060 VDD.n3528 VDD.n3527 0.648317
R32061 VDD.n3525 VDD.n3524 0.648317
R32062 VDD.n3434 VDD.n3433 0.648317
R32063 VDD.n3439 VDD.n3438 0.648317
R32064 VDD.n3431 VDD.n3430 0.648317
R32065 VDD.n3339 VDD.n3338 0.648317
R32066 VDD.n3344 VDD.n3343 0.648317
R32067 VDD.n266 VDD.n265 0.6205
R32068 VDD.n1593 VDD 0.601043
R32069 VDD.n1627 VDD 0.601043
R32070 VDD.n1664 VDD 0.601043
R32071 VDD.n1689 VDD 0.601043
R32072 VDD.n1333 VDD 0.601043
R32073 VDD.n1367 VDD 0.601043
R32074 VDD.n1404 VDD 0.601043
R32075 VDD.n1429 VDD 0.601043
R32076 VDD.n1073 VDD 0.601043
R32077 VDD.n1107 VDD 0.601043
R32078 VDD.n1144 VDD 0.601043
R32079 VDD.n1169 VDD 0.601043
R32080 VDD.n813 VDD 0.601043
R32081 VDD.n847 VDD 0.601043
R32082 VDD.n884 VDD 0.601043
R32083 VDD.n909 VDD 0.601043
R32084 VDD.n553 VDD 0.601043
R32085 VDD.n587 VDD 0.601043
R32086 VDD.n624 VDD 0.601043
R32087 VDD.n649 VDD 0.601043
R32088 VDD.n293 VDD 0.601043
R32089 VDD.n327 VDD 0.601043
R32090 VDD.n364 VDD 0.601043
R32091 VDD.n389 VDD 0.601043
R32092 VDD VDD.n0 0.601043
R32093 VDD VDD.n25 0.601043
R32094 VDD VDD.n50 0.601043
R32095 VDD VDD.n75 0.601043
R32096 VDD.n7209 VDD 0.601043
R32097 VDD.n7243 VDD 0.601043
R32098 VDD.n7280 VDD 0.601043
R32099 VDD.n7305 VDD 0.601043
R32100 VDD VDD.n6859 0.601043
R32101 VDD VDD.n6884 0.601043
R32102 VDD VDD.n6909 0.601043
R32103 VDD VDD.n5052 0.601043
R32104 VDD VDD.n5080 0.601043
R32105 VDD VDD.n5114 0.601043
R32106 VDD VDD.n5149 0.601043
R32107 VDD.n6704 VDD 0.601043
R32108 VDD VDD.n5188 0.601043
R32109 VDD VDD.n5216 0.601043
R32110 VDD VDD.n5250 0.601043
R32111 VDD VDD.n5285 0.601043
R32112 VDD.n6581 VDD 0.601043
R32113 VDD VDD.n5324 0.601043
R32114 VDD VDD.n5352 0.601043
R32115 VDD VDD.n5386 0.601043
R32116 VDD VDD.n5421 0.601043
R32117 VDD.n6458 VDD 0.601043
R32118 VDD VDD.n5460 0.601043
R32119 VDD VDD.n5488 0.601043
R32120 VDD VDD.n5522 0.601043
R32121 VDD VDD.n5557 0.601043
R32122 VDD.n6335 VDD 0.601043
R32123 VDD VDD.n5596 0.601043
R32124 VDD VDD.n5624 0.601043
R32125 VDD VDD.n5658 0.601043
R32126 VDD VDD.n5693 0.601043
R32127 VDD.n6212 VDD 0.601043
R32128 VDD VDD.n5732 0.601043
R32129 VDD VDD.n5760 0.601043
R32130 VDD VDD.n5794 0.601043
R32131 VDD VDD.n5829 0.601043
R32132 VDD.n6089 VDD 0.601043
R32133 VDD VDD.n5868 0.601043
R32134 VDD VDD.n5896 0.601043
R32135 VDD VDD.n5930 0.601043
R32136 VDD VDD.n5965 0.601043
R32137 VDD.n5966 VDD 0.601043
R32138 VDD.n4862 VDD 0.601043
R32139 VDD.n4837 VDD 0.601043
R32140 VDD.n4800 VDD 0.601043
R32141 VDD.n4766 VDD 0.601043
R32142 VDD VDD.n5013 0.601043
R32143 VDD.n3707 VDD 0.601043
R32144 VDD.n3732 VDD 0.601043
R32145 VDD.n2881 VDD 0.601043
R32146 VDD.n2906 VDD 0.601043
R32147 VDD.n2941 VDD 0.601043
R32148 VDD.n2975 VDD 0.601043
R32149 VDD.n2745 VDD 0.601043
R32150 VDD.n2770 VDD 0.601043
R32151 VDD.n2805 VDD 0.601043
R32152 VDD.n2839 VDD 0.601043
R32153 VDD.n2609 VDD 0.601043
R32154 VDD.n2634 VDD 0.601043
R32155 VDD.n2669 VDD 0.601043
R32156 VDD.n2703 VDD 0.601043
R32157 VDD.n2473 VDD 0.601043
R32158 VDD.n2498 VDD 0.601043
R32159 VDD.n2533 VDD 0.601043
R32160 VDD.n2567 VDD 0.601043
R32161 VDD.n2337 VDD 0.601043
R32162 VDD.n2362 VDD 0.601043
R32163 VDD.n2397 VDD 0.601043
R32164 VDD.n2431 VDD 0.601043
R32165 VDD.n2201 VDD 0.601043
R32166 VDD.n2226 VDD 0.601043
R32167 VDD.n2261 VDD 0.601043
R32168 VDD.n2295 VDD 0.601043
R32169 VDD.n2065 VDD 0.601043
R32170 VDD.n2090 VDD 0.601043
R32171 VDD.n2125 VDD 0.601043
R32172 VDD.n2159 VDD 0.601043
R32173 VDD.n1989 VDD 0.601043
R32174 VDD.n2023 VDD 0.601043
R32175 VDD.n1929 VDD 0.601043
R32176 VDD.n1954 VDD 0.601043
R32177 VDD.n1853 VDD 0.601043
R32178 VDD.n1887 VDD 0.601043
R32179 VDD VDD.n7717 0.601043
R32180 VDD.n7509 VDD 0.601043
R32181 VDD.n7546 VDD 0.601043
R32182 VDD.n7571 VDD 0.601043
R32183 VDD.n3335 VDD 0.592985
R32184 VDD.n3528 VDD 0.592985
R32185 VDD.n3524 VDD 0.592985
R32186 VDD.n3434 VDD 0.592985
R32187 VDD.n3439 VDD 0.592985
R32188 VDD.n3430 VDD 0.592985
R32189 VDD.n3339 VDD 0.592985
R32190 VDD.n3344 VDD 0.592985
R32191 VDD.n2990 VDD 0.524957
R32192 VDD.n2979 VDD 0.524957
R32193 VDD.n6837 VDD.n6828 0.5005
R32194 VDD.n278 VDD.n267 0.486913
R32195 VDD.n3087 VDD 0.447191
R32196 VDD.n3076 VDD 0.447191
R32197 VDD.n3103 VDD 0.447191
R32198 VDD.n3112 VDD 0.447191
R32199 VDD.n3151 VDD 0.447191
R32200 VDD.n3140 VDD 0.447191
R32201 VDD.n3167 VDD 0.447191
R32202 VDD.n3176 VDD 0.447191
R32203 VDD.n3048 VDD 0.447191
R32204 VDD.n3037 VDD 0.447191
R32205 VDD.n3191 VDD 0.447191
R32206 VDD.n3200 VDD 0.447191
R32207 VDD.n3302 VDD 0.447191
R32208 VDD.n3291 VDD 0.447191
R32209 VDD.n3568 VDD 0.447191
R32210 VDD.n3577 VDD 0.447191
R32211 VDD.n3009 VDD 0.447191
R32212 VDD.n2998 VDD 0.447191
R32213 VDD.n3025 VDD 0.447191
R32214 VDD.n3034 VDD 0.447191
R32215 VDD.n3596 VDD 0.447191
R32216 VDD.n3585 VDD 0.447191
R32217 VDD.n3612 VDD 0.447191
R32218 VDD.n3621 VDD 0.447191
R32219 VDD.n2986 VDD 0.447191
R32220 VDD.n3635 VDD 0.447191
R32221 VDD.n3644 VDD 0.447191
R32222 VDD.n3067 VDD 0.447191
R32223 VDD.n3056 VDD 0.447191
R32224 VDD.n3122 VDD 0.447191
R32225 VDD.n3131 VDD 0.447191
R32226 VDD.n3656 VDD 0.447191
R32227 VDD.n3665 VDD 0.447191
R32228 VDD.n3346 VDD.n3337 0.447
R32229 VDD.n3530 VDD.n3529 0.447
R32230 VDD.n3530 VDD.n3526 0.447
R32231 VDD.n3437 VDD.n3436 0.447
R32232 VDD.n3441 VDD.n3432 0.447
R32233 VDD.n3428 VDD.n3279 0.447
R32234 VDD.n3342 VDD.n3341 0.447
R32235 VDD.n3522 VDD.n3242 0.446929
R32236 VDD.n7197 VDD.n7196 0.435283
R32237 VDD.n1840 VDD.n1839 0.410826
R32238 VDD.n1594 VDD.n1593 0.410826
R32239 VDD.n1628 VDD.n1627 0.410826
R32240 VDD.n1665 VDD.n1664 0.410826
R32241 VDD.n1690 VDD.n1689 0.410826
R32242 VDD.n1580 VDD.n1579 0.410826
R32243 VDD.n1334 VDD.n1333 0.410826
R32244 VDD.n1368 VDD.n1367 0.410826
R32245 VDD.n1405 VDD.n1404 0.410826
R32246 VDD.n1430 VDD.n1429 0.410826
R32247 VDD.n1320 VDD.n1319 0.410826
R32248 VDD.n1074 VDD.n1073 0.410826
R32249 VDD.n1108 VDD.n1107 0.410826
R32250 VDD.n1145 VDD.n1144 0.410826
R32251 VDD.n1170 VDD.n1169 0.410826
R32252 VDD.n1060 VDD.n1059 0.410826
R32253 VDD.n814 VDD.n813 0.410826
R32254 VDD.n848 VDD.n847 0.410826
R32255 VDD.n885 VDD.n884 0.410826
R32256 VDD.n910 VDD.n909 0.410826
R32257 VDD.n800 VDD.n799 0.410826
R32258 VDD.n554 VDD.n553 0.410826
R32259 VDD.n588 VDD.n587 0.410826
R32260 VDD.n625 VDD.n624 0.410826
R32261 VDD.n650 VDD.n649 0.410826
R32262 VDD.n540 VDD.n539 0.410826
R32263 VDD.n294 VDD.n293 0.410826
R32264 VDD.n328 VDD.n327 0.410826
R32265 VDD.n365 VDD.n364 0.410826
R32266 VDD.n390 VDD.n389 0.410826
R32267 VDD.n239 VDD.n0 0.410826
R32268 VDD.n204 VDD.n25 0.410826
R32269 VDD.n169 VDD.n50 0.410826
R32270 VDD.n134 VDD.n75 0.410826
R32271 VDD.n7456 VDD.n7455 0.410826
R32272 VDD.n7210 VDD.n7209 0.410826
R32273 VDD.n7244 VDD.n7243 0.410826
R32274 VDD.n7281 VDD.n7280 0.410826
R32275 VDD.n7306 VDD.n7305 0.410826
R32276 VDD.n7038 VDD.n6859 0.410826
R32277 VDD.n7003 VDD.n6884 0.410826
R32278 VDD.n6968 VDD.n6909 0.410826
R32279 VDD.n5052 VDD.n5042 0.410826
R32280 VDD.n5080 VDD.n5079 0.410826
R32281 VDD.n5114 VDD.n5104 0.410826
R32282 VDD.n5149 VDD.n5138 0.410826
R32283 VDD.n6705 VDD.n6704 0.410826
R32284 VDD.n5188 VDD.n5178 0.410826
R32285 VDD.n5216 VDD.n5215 0.410826
R32286 VDD.n5250 VDD.n5240 0.410826
R32287 VDD.n5285 VDD.n5274 0.410826
R32288 VDD.n6582 VDD.n6581 0.410826
R32289 VDD.n5324 VDD.n5314 0.410826
R32290 VDD.n5352 VDD.n5351 0.410826
R32291 VDD.n5386 VDD.n5376 0.410826
R32292 VDD.n5421 VDD.n5410 0.410826
R32293 VDD.n6459 VDD.n6458 0.410826
R32294 VDD.n5460 VDD.n5450 0.410826
R32295 VDD.n5488 VDD.n5487 0.410826
R32296 VDD.n5522 VDD.n5512 0.410826
R32297 VDD.n5557 VDD.n5546 0.410826
R32298 VDD.n6336 VDD.n6335 0.410826
R32299 VDD.n5596 VDD.n5586 0.410826
R32300 VDD.n5624 VDD.n5623 0.410826
R32301 VDD.n5658 VDD.n5648 0.410826
R32302 VDD.n5693 VDD.n5682 0.410826
R32303 VDD.n6213 VDD.n6212 0.410826
R32304 VDD.n5732 VDD.n5722 0.410826
R32305 VDD.n5760 VDD.n5759 0.410826
R32306 VDD.n5794 VDD.n5784 0.410826
R32307 VDD.n5829 VDD.n5818 0.410826
R32308 VDD.n6090 VDD.n6089 0.410826
R32309 VDD.n5868 VDD.n5858 0.410826
R32310 VDD.n5896 VDD.n5895 0.410826
R32311 VDD.n5930 VDD.n5920 0.410826
R32312 VDD.n5965 VDD.n5954 0.410826
R32313 VDD.n5967 VDD.n5966 0.410826
R32314 VDD.n4863 VDD.n4862 0.410826
R32315 VDD.n4838 VDD.n4837 0.410826
R32316 VDD.n4801 VDD.n4800 0.410826
R32317 VDD.n4767 VDD.n4766 0.410826
R32318 VDD.n5013 VDD.n5012 0.410826
R32319 VDD.n3708 VDD.n3707 0.410826
R32320 VDD.n3733 VDD.n3732 0.410826
R32321 VDD.n2882 VDD.n2881 0.410826
R32322 VDD.n2907 VDD.n2906 0.410826
R32323 VDD.n3880 VDD.n3879 0.410826
R32324 VDD.n2942 VDD.n2941 0.410826
R32325 VDD.n2746 VDD.n2745 0.410826
R32326 VDD.n2771 VDD.n2770 0.410826
R32327 VDD.n4005 VDD.n4004 0.410826
R32328 VDD.n2806 VDD.n2805 0.410826
R32329 VDD.n2610 VDD.n2609 0.410826
R32330 VDD.n2635 VDD.n2634 0.410826
R32331 VDD.n4130 VDD.n4129 0.410826
R32332 VDD.n2670 VDD.n2669 0.410826
R32333 VDD.n2474 VDD.n2473 0.410826
R32334 VDD.n2499 VDD.n2498 0.410826
R32335 VDD.n4255 VDD.n4254 0.410826
R32336 VDD.n2534 VDD.n2533 0.410826
R32337 VDD.n2338 VDD.n2337 0.410826
R32338 VDD.n2363 VDD.n2362 0.410826
R32339 VDD.n4380 VDD.n4379 0.410826
R32340 VDD.n2398 VDD.n2397 0.410826
R32341 VDD.n2202 VDD.n2201 0.410826
R32342 VDD.n2227 VDD.n2226 0.410826
R32343 VDD.n4505 VDD.n4504 0.410826
R32344 VDD.n2262 VDD.n2261 0.410826
R32345 VDD.n2066 VDD.n2065 0.410826
R32346 VDD.n2091 VDD.n2090 0.410826
R32347 VDD.n4630 VDD.n4629 0.410826
R32348 VDD.n2126 VDD.n2125 0.410826
R32349 VDD.n4755 VDD.n4754 0.410826
R32350 VDD.n1990 VDD.n1989 0.410826
R32351 VDD.n1930 VDD.n1929 0.410826
R32352 VDD.n1955 VDD.n1954 0.410826
R32353 VDD.n7196 VDD.n7195 0.410826
R32354 VDD.n1854 VDD.n1853 0.410826
R32355 VDD.n7460 VDD.n7459 0.410826
R32356 VDD.n7717 VDD.n7716 0.410826
R32357 VDD.n7510 VDD.n7509 0.410826
R32358 VDD.n7547 VDD.n7546 0.410826
R32359 VDD.n7572 VDD.n7571 0.410826
R32360 VDD.n3376 VDD.n3375 0.405391
R32361 VDD.n3414 VDD.n3413 0.405391
R32362 VDD.n3453 VDD.n3255 0.405391
R32363 VDD.n3471 VDD.n3470 0.405391
R32364 VDD.n3508 VDD.n3507 0.405391
R32365 VDD.n3358 VDD.n3311 0.405391
R32366 VDD.n3557 VDD.n3205 0.405391
R32367 VDD.n2976 VDD.n2975 0.32387
R32368 VDD.n2840 VDD.n2839 0.32387
R32369 VDD.n2704 VDD.n2703 0.32387
R32370 VDD.n2568 VDD.n2567 0.32387
R32371 VDD.n2432 VDD.n2431 0.32387
R32372 VDD.n2296 VDD.n2295 0.32387
R32373 VDD.n2160 VDD.n2159 0.32387
R32374 VDD.n2024 VDD.n2023 0.32387
R32375 VDD.n1888 VDD.n1887 0.32387
R32376 VDD.n2993 VDD 0.252453
R32377 VDD.n2982 VDD 0.252453
R32378 VDD.n3088 VDD.n3087 0.226043
R32379 VDD.n3077 VDD.n3076 0.226043
R32380 VDD.n3104 VDD.n3103 0.226043
R32381 VDD.n3112 VDD.n3111 0.226043
R32382 VDD.n3152 VDD.n3151 0.226043
R32383 VDD.n3141 VDD.n3140 0.226043
R32384 VDD.n3168 VDD.n3167 0.226043
R32385 VDD.n3176 VDD.n3175 0.226043
R32386 VDD.n3049 VDD.n3048 0.226043
R32387 VDD.n3038 VDD.n3037 0.226043
R32388 VDD.n3192 VDD.n3191 0.226043
R32389 VDD.n3200 VDD.n3199 0.226043
R32390 VDD.n3303 VDD.n3302 0.226043
R32391 VDD.n3292 VDD.n3291 0.226043
R32392 VDD.n3569 VDD.n3568 0.226043
R32393 VDD.n3577 VDD.n3576 0.226043
R32394 VDD.n3010 VDD.n3009 0.226043
R32395 VDD.n2999 VDD.n2998 0.226043
R32396 VDD.n3026 VDD.n3025 0.226043
R32397 VDD.n3034 VDD.n3033 0.226043
R32398 VDD.n3597 VDD.n3596 0.226043
R32399 VDD.n3586 VDD.n3585 0.226043
R32400 VDD.n3613 VDD.n3612 0.226043
R32401 VDD.n3621 VDD.n3620 0.226043
R32402 VDD.n2993 VDD.n2992 0.226043
R32403 VDD.n2982 VDD.n2981 0.226043
R32404 VDD.n3636 VDD.n3635 0.226043
R32405 VDD.n3644 VDD.n3643 0.226043
R32406 VDD.n3068 VDD.n3067 0.226043
R32407 VDD.n3057 VDD.n3056 0.226043
R32408 VDD.n3123 VDD.n3122 0.226043
R32409 VDD.n3131 VDD.n3130 0.226043
R32410 VDD.n3657 VDD.n3656 0.226043
R32411 VDD.n3665 VDD.n3664 0.226043
R32412 VDD.n3082 VDD 0.217464
R32413 VDD.n3098 VDD 0.217464
R32414 VDD.n3146 VDD 0.217464
R32415 VDD.n3162 VDD 0.217464
R32416 VDD.n3043 VDD 0.217464
R32417 VDD.n3186 VDD 0.217464
R32418 VDD.n3297 VDD 0.217464
R32419 VDD.n3563 VDD 0.217464
R32420 VDD.n3004 VDD 0.217464
R32421 VDD.n3020 VDD 0.217464
R32422 VDD.n3591 VDD 0.217464
R32423 VDD.n3607 VDD 0.217464
R32424 VDD.n2989 VDD 0.217464
R32425 VDD.n2978 VDD 0.217464
R32426 VDD.n3630 VDD 0.217464
R32427 VDD.n3062 VDD 0.217464
R32428 VDD.n3117 VDD 0.217464
R32429 VDD.n3651 VDD 0.217464
R32430 VDD.n279 VDD 0.166261
R32431 VDD.n3090 VDD 0.1255
R32432 VDD.n3083 VDD 0.1255
R32433 VDD.n3079 VDD 0.1255
R32434 VDD.n3106 VDD 0.1255
R32435 VDD.n3099 VDD 0.1255
R32436 VDD.n3096 VDD 0.1255
R32437 VDD.n3154 VDD 0.1255
R32438 VDD.n3147 VDD 0.1255
R32439 VDD.n3143 VDD 0.1255
R32440 VDD.n3170 VDD 0.1255
R32441 VDD.n3163 VDD 0.1255
R32442 VDD.n3160 VDD 0.1255
R32443 VDD.n3051 VDD 0.1255
R32444 VDD.n3044 VDD 0.1255
R32445 VDD.n3040 VDD 0.1255
R32446 VDD.n3194 VDD 0.1255
R32447 VDD.n3187 VDD 0.1255
R32448 VDD.n3184 VDD 0.1255
R32449 VDD.n3305 VDD 0.1255
R32450 VDD.n3298 VDD 0.1255
R32451 VDD.n3294 VDD 0.1255
R32452 VDD.n3571 VDD 0.1255
R32453 VDD.n3564 VDD 0.1255
R32454 VDD.n3561 VDD 0.1255
R32455 VDD.n3012 VDD 0.1255
R32456 VDD.n3005 VDD 0.1255
R32457 VDD.n3001 VDD 0.1255
R32458 VDD.n3028 VDD 0.1255
R32459 VDD.n3021 VDD 0.1255
R32460 VDD.n3018 VDD 0.1255
R32461 VDD.n3599 VDD 0.1255
R32462 VDD.n3592 VDD 0.1255
R32463 VDD.n3588 VDD 0.1255
R32464 VDD.n3615 VDD 0.1255
R32465 VDD.n3608 VDD 0.1255
R32466 VDD.n3605 VDD 0.1255
R32467 VDD.n2992 VDD 0.1255
R32468 VDD.n2985 VDD 0.1255
R32469 VDD.n2981 VDD 0.1255
R32470 VDD.n3638 VDD 0.1255
R32471 VDD.n3631 VDD 0.1255
R32472 VDD.n3628 VDD 0.1255
R32473 VDD.n3070 VDD 0.1255
R32474 VDD.n3063 VDD 0.1255
R32475 VDD.n3059 VDD 0.1255
R32476 VDD.n3125 VDD 0.1255
R32477 VDD.n3118 VDD 0.1255
R32478 VDD.n3115 VDD 0.1255
R32479 VDD.n3659 VDD 0.1255
R32480 VDD.n3652 VDD 0.1255
R32481 VDD.n3649 VDD 0.1255
R32482 VDD.n243 VDD.n242 0.112862
R32483 VDD.n6828 VDD 0.101043
R32484 VDD.t701 VDD.n262 0.086419
R32485 VDD.t699 VDD.n256 0.086419
R32486 VDD.n280 VDD.n279 0.063
R32487 VDD.n7069 VDD.n6828 0.063
R32488 VDD.n3092 VDD.n3088 0.063
R32489 VDD.n3092 VDD.n3091 0.063
R32490 VDD.n3081 VDD.n3077 0.063
R32491 VDD.n3081 VDD.n3080 0.063
R32492 VDD.n3108 VDD.n3104 0.063
R32493 VDD.n3108 VDD.n3107 0.063
R32494 VDD.n3111 VDD.n3110 0.063
R32495 VDD.n3110 VDD.n3097 0.063
R32496 VDD.n3156 VDD.n3152 0.063
R32497 VDD.n3156 VDD.n3155 0.063
R32498 VDD.n3145 VDD.n3141 0.063
R32499 VDD.n3145 VDD.n3144 0.063
R32500 VDD.n3172 VDD.n3168 0.063
R32501 VDD.n3172 VDD.n3171 0.063
R32502 VDD.n3175 VDD.n3174 0.063
R32503 VDD.n3174 VDD.n3161 0.063
R32504 VDD.n3053 VDD.n3049 0.063
R32505 VDD.n3053 VDD.n3052 0.063
R32506 VDD.n3042 VDD.n3038 0.063
R32507 VDD.n3042 VDD.n3041 0.063
R32508 VDD.n3196 VDD.n3192 0.063
R32509 VDD.n3196 VDD.n3195 0.063
R32510 VDD.n3199 VDD.n3198 0.063
R32511 VDD.n3198 VDD.n3185 0.063
R32512 VDD.n3307 VDD.n3303 0.063
R32513 VDD.n3307 VDD.n3306 0.063
R32514 VDD.n3296 VDD.n3292 0.063
R32515 VDD.n3296 VDD.n3295 0.063
R32516 VDD.n3377 VDD.n3281 0.063
R32517 VDD.n3389 VDD.n3281 0.063
R32518 VDD.n3427 VDD.n3280 0.063
R32519 VDD.n3427 VDD.n3426 0.063
R32520 VDD.n3443 VDD.n3442 0.063
R32521 VDD.n3442 VDD.n3278 0.063
R32522 VDD.n3472 VDD.n3244 0.063
R32523 VDD.n3484 VDD.n3244 0.063
R32524 VDD.n3348 VDD.n3347 0.063
R32525 VDD.n3347 VDD.n3334 0.063
R32526 VDD.n3531 VDD.n3241 0.063
R32527 VDD.n3532 VDD.n3531 0.063
R32528 VDD.n3573 VDD.n3569 0.063
R32529 VDD.n3573 VDD.n3572 0.063
R32530 VDD.n3576 VDD.n3575 0.063
R32531 VDD.n3575 VDD.n3562 0.063
R32532 VDD.n3014 VDD.n3010 0.063
R32533 VDD.n3014 VDD.n3013 0.063
R32534 VDD.n3003 VDD.n2999 0.063
R32535 VDD.n3003 VDD.n3002 0.063
R32536 VDD.n3030 VDD.n3026 0.063
R32537 VDD.n3030 VDD.n3029 0.063
R32538 VDD.n3033 VDD.n3032 0.063
R32539 VDD.n3032 VDD.n3019 0.063
R32540 VDD.n3601 VDD.n3597 0.063
R32541 VDD.n3601 VDD.n3600 0.063
R32542 VDD.n3590 VDD.n3586 0.063
R32543 VDD.n3590 VDD.n3589 0.063
R32544 VDD.n3617 VDD.n3613 0.063
R32545 VDD.n3617 VDD.n3616 0.063
R32546 VDD.n3620 VDD.n3619 0.063
R32547 VDD.n3619 VDD.n3606 0.063
R32548 VDD.n2994 VDD.n2990 0.063
R32549 VDD.n2994 VDD.n2993 0.063
R32550 VDD.n2983 VDD.n2979 0.063
R32551 VDD.n2983 VDD.n2982 0.063
R32552 VDD.n3640 VDD.n3636 0.063
R32553 VDD.n3640 VDD.n3639 0.063
R32554 VDD.n3643 VDD.n3642 0.063
R32555 VDD.n3642 VDD.n3629 0.063
R32556 VDD.n3072 VDD.n3068 0.063
R32557 VDD.n3072 VDD.n3071 0.063
R32558 VDD.n3061 VDD.n3057 0.063
R32559 VDD.n3061 VDD.n3060 0.063
R32560 VDD.n3127 VDD.n3123 0.063
R32561 VDD.n3127 VDD.n3126 0.063
R32562 VDD.n3130 VDD.n3129 0.063
R32563 VDD.n3129 VDD.n3116 0.063
R32564 VDD.n3661 VDD.n3657 0.063
R32565 VDD.n3661 VDD.n3660 0.063
R32566 VDD.n3664 VDD.n3663 0.063
R32567 VDD.n3663 VDD.n3650 0.063
R32568 VDD.n3667 VDD.n2976 0.063
R32569 VDD.n3679 VDD.n3667 0.063
R32570 VDD.n2841 VDD.n2840 0.063
R32571 VDD.n2853 VDD.n2841 0.063
R32572 VDD.n2705 VDD.n2704 0.063
R32573 VDD.n2717 VDD.n2705 0.063
R32574 VDD.n2569 VDD.n2568 0.063
R32575 VDD.n2581 VDD.n2569 0.063
R32576 VDD.n2433 VDD.n2432 0.063
R32577 VDD.n2445 VDD.n2433 0.063
R32578 VDD.n2297 VDD.n2296 0.063
R32579 VDD.n2309 VDD.n2297 0.063
R32580 VDD.n2161 VDD.n2160 0.063
R32581 VDD.n2173 VDD.n2161 0.063
R32582 VDD.n2025 VDD.n2024 0.063
R32583 VDD.n2037 VDD.n2025 0.063
R32584 VDD.n1889 VDD.n1888 0.063
R32585 VDD.n1901 VDD.n1889 0.063
R32586 VDD.n3521 VDD.n3243 0.0620385
R32587 VDD.n3521 VDD.n3520 0.0620385
R32588 VDD.n274 VDD.t462 0.0617545
R32589 VDD.n271 VDD.t462 0.0617545
R32590 VDD.n280 VDD 0.0571406
R32591 VDD VDD.n7068 0.0532344
R32592 VDD.n3136 VDD 0.0477973
R32593 VDD.n3135 VDD 0.0249565
R32594 VDD.n3529 VDD.n3528 0.024
R32595 VDD.n3524 VDD.n3523 0.024
R32596 VDD.n3435 VDD.n3434 0.024
R32597 VDD.n3440 VDD.n3439 0.024
R32598 VDD.n3430 VDD.n3429 0.024
R32599 VDD.n3340 VDD.n3339 0.024
R32600 VDD.n3345 VDD.n3344 0.024
R32601 VDD.n3084 VDD.n3083 0.0216397
R32602 VDD.n3084 VDD 0.0216397
R32603 VDD.n3100 VDD.n3099 0.0216397
R32604 VDD.n3100 VDD 0.0216397
R32605 VDD.n3148 VDD.n3147 0.0216397
R32606 VDD.n3148 VDD 0.0216397
R32607 VDD.n3164 VDD.n3163 0.0216397
R32608 VDD.n3164 VDD 0.0216397
R32609 VDD.n3045 VDD.n3044 0.0216397
R32610 VDD.n3045 VDD 0.0216397
R32611 VDD.n3188 VDD.n3187 0.0216397
R32612 VDD.n3188 VDD 0.0216397
R32613 VDD.n3299 VDD.n3298 0.0216397
R32614 VDD.n3299 VDD 0.0216397
R32615 VDD.n3565 VDD.n3564 0.0216397
R32616 VDD.n3565 VDD 0.0216397
R32617 VDD.n3006 VDD.n3005 0.0216397
R32618 VDD.n3006 VDD 0.0216397
R32619 VDD.n3022 VDD.n3021 0.0216397
R32620 VDD.n3022 VDD 0.0216397
R32621 VDD.n3593 VDD.n3592 0.0216397
R32622 VDD.n3593 VDD 0.0216397
R32623 VDD.n3609 VDD.n3608 0.0216397
R32624 VDD.n3609 VDD 0.0216397
R32625 VDD.n2992 VDD.n2991 0.0216397
R32626 VDD.n2991 VDD 0.0216397
R32627 VDD.n2981 VDD.n2980 0.0216397
R32628 VDD.n2980 VDD 0.0216397
R32629 VDD.n3632 VDD.n3631 0.0216397
R32630 VDD.n3632 VDD 0.0216397
R32631 VDD.n3064 VDD.n3063 0.0216397
R32632 VDD.n3064 VDD 0.0216397
R32633 VDD.n3119 VDD.n3118 0.0216397
R32634 VDD.n3119 VDD 0.0216397
R32635 VDD.n3653 VDD.n3652 0.0216397
R32636 VDD.n3653 VDD 0.0216397
R32637 VDD.n3337 VDD 0.0204394
R32638 VDD.n3526 VDD 0.0204394
R32639 VDD VDD.n3242 0.0204394
R32640 VDD VDD.n3437 0.0204394
R32641 VDD.n3432 VDD 0.0204394
R32642 VDD VDD.n3279 0.0204394
R32643 VDD VDD.n3342 0.0204394
R32644 VDD VDD.n3135 0.0157027
R32645 VDD.n3090 VDD.n3089 0.0107679
R32646 VDD.n3089 VDD 0.0107679
R32647 VDD.n3079 VDD.n3078 0.0107679
R32648 VDD.n3078 VDD 0.0107679
R32649 VDD.n3106 VDD.n3105 0.0107679
R32650 VDD.n3105 VDD 0.0107679
R32651 VDD.n3096 VDD.n3095 0.0107679
R32652 VDD.n3095 VDD 0.0107679
R32653 VDD.n3154 VDD.n3153 0.0107679
R32654 VDD.n3153 VDD 0.0107679
R32655 VDD.n3143 VDD.n3142 0.0107679
R32656 VDD.n3142 VDD 0.0107679
R32657 VDD.n3170 VDD.n3169 0.0107679
R32658 VDD.n3169 VDD 0.0107679
R32659 VDD.n3160 VDD.n3159 0.0107679
R32660 VDD.n3159 VDD 0.0107679
R32661 VDD.n3051 VDD.n3050 0.0107679
R32662 VDD.n3050 VDD 0.0107679
R32663 VDD.n3040 VDD.n3039 0.0107679
R32664 VDD.n3039 VDD 0.0107679
R32665 VDD.n3194 VDD.n3193 0.0107679
R32666 VDD.n3193 VDD 0.0107679
R32667 VDD.n3184 VDD.n3183 0.0107679
R32668 VDD.n3183 VDD 0.0107679
R32669 VDD.n3305 VDD.n3304 0.0107679
R32670 VDD.n3304 VDD 0.0107679
R32671 VDD.n3294 VDD.n3293 0.0107679
R32672 VDD.n3293 VDD 0.0107679
R32673 VDD.n3571 VDD.n3570 0.0107679
R32674 VDD.n3570 VDD 0.0107679
R32675 VDD.n3561 VDD.n3560 0.0107679
R32676 VDD.n3560 VDD 0.0107679
R32677 VDD.n3012 VDD.n3011 0.0107679
R32678 VDD.n3011 VDD 0.0107679
R32679 VDD.n3001 VDD.n3000 0.0107679
R32680 VDD.n3000 VDD 0.0107679
R32681 VDD.n3028 VDD.n3027 0.0107679
R32682 VDD.n3027 VDD 0.0107679
R32683 VDD.n3018 VDD.n3017 0.0107679
R32684 VDD.n3017 VDD 0.0107679
R32685 VDD.n3599 VDD.n3598 0.0107679
R32686 VDD.n3598 VDD 0.0107679
R32687 VDD.n3588 VDD.n3587 0.0107679
R32688 VDD.n3587 VDD 0.0107679
R32689 VDD.n3615 VDD.n3614 0.0107679
R32690 VDD.n3614 VDD 0.0107679
R32691 VDD.n3605 VDD.n3604 0.0107679
R32692 VDD.n3604 VDD 0.0107679
R32693 VDD.n2985 VDD.n2984 0.0107679
R32694 VDD.n2984 VDD 0.0107679
R32695 VDD.n3638 VDD.n3637 0.0107679
R32696 VDD.n3637 VDD 0.0107679
R32697 VDD.n3628 VDD.n3627 0.0107679
R32698 VDD.n3627 VDD 0.0107679
R32699 VDD.n3070 VDD.n3069 0.0107679
R32700 VDD.n3069 VDD 0.0107679
R32701 VDD.n3059 VDD.n3058 0.0107679
R32702 VDD.n3058 VDD 0.0107679
R32703 VDD.n3125 VDD.n3124 0.0107679
R32704 VDD.n3124 VDD 0.0107679
R32705 VDD.n3115 VDD.n3114 0.0107679
R32706 VDD.n3114 VDD 0.0107679
R32707 VDD.n3659 VDD.n3658 0.0107679
R32708 VDD.n3658 VDD 0.0107679
R32709 VDD.n3649 VDD.n3648 0.0107679
R32710 VDD.n3648 VDD 0.0107679
R32711 VDD.n7069 VDD 0.0102656
R32712 VDD.n3334 VDD 0.00534007
R32713 VDD.n3389 VDD.n3282 0.00534007
R32714 VDD VDD.n3389 0.00534007
R32715 VDD.n3426 VDD.n3390 0.00534007
R32716 VDD.n3426 VDD 0.00534007
R32717 VDD.n3391 VDD.n3278 0.00534007
R32718 VDD.n3278 VDD 0.00534007
R32719 VDD.n3484 VDD.n3245 0.00534007
R32720 VDD VDD.n3484 0.00534007
R32721 VDD.n3520 VDD.n3485 0.00534007
R32722 VDD.n3520 VDD 0.00534007
R32723 VDD.n3532 VDD.n3240 0.00534007
R32724 VDD.n3532 VDD 0.00534007
R32725 VDD.n3086 VDD 0.00441667
R32726 VDD.n3102 VDD 0.00441667
R32727 VDD.n3150 VDD 0.00441667
R32728 VDD.n3166 VDD 0.00441667
R32729 VDD.n3047 VDD 0.00441667
R32730 VDD.n3190 VDD 0.00441667
R32731 VDD.n3301 VDD 0.00441667
R32732 VDD.n3336 VDD 0.00441667
R32733 VDD.n3527 VDD 0.00441667
R32734 VDD.n3525 VDD 0.00441667
R32735 VDD.n3433 VDD 0.00441667
R32736 VDD.n3438 VDD 0.00441667
R32737 VDD.n3431 VDD 0.00441667
R32738 VDD.n3338 VDD 0.00441667
R32739 VDD.n3343 VDD 0.00441667
R32740 VDD.n3567 VDD 0.00441667
R32741 VDD.n3008 VDD 0.00441667
R32742 VDD.n3024 VDD 0.00441667
R32743 VDD.n3595 VDD 0.00441667
R32744 VDD.n3611 VDD 0.00441667
R32745 VDD.n2987 VDD 0.00441667
R32746 VDD.n3634 VDD 0.00441667
R32747 VDD.n3066 VDD 0.00441667
R32748 VDD.n3121 VDD 0.00441667
R32749 VDD.n3655 VDD 0.00441667
R32750 VDD VDD.n3086 0.00406061
R32751 VDD VDD.n3102 0.00406061
R32752 VDD VDD.n3150 0.00406061
R32753 VDD VDD.n3166 0.00406061
R32754 VDD VDD.n3047 0.00406061
R32755 VDD VDD.n3190 0.00406061
R32756 VDD VDD.n3301 0.00406061
R32757 VDD VDD.n3336 0.00406061
R32758 VDD.n3527 VDD 0.00406061
R32759 VDD VDD.n3525 0.00406061
R32760 VDD.n3433 VDD 0.00406061
R32761 VDD.n3438 VDD 0.00406061
R32762 VDD VDD.n3431 0.00406061
R32763 VDD.n3338 VDD 0.00406061
R32764 VDD.n3343 VDD 0.00406061
R32765 VDD VDD.n3567 0.00406061
R32766 VDD VDD.n3008 0.00406061
R32767 VDD VDD.n3024 0.00406061
R32768 VDD VDD.n3595 0.00406061
R32769 VDD VDD.n3611 0.00406061
R32770 VDD.n2987 VDD 0.00406061
R32771 VDD VDD.n3634 0.00406061
R32772 VDD VDD.n3066 0.00406061
R32773 VDD VDD.n3121 0.00406061
R32774 VDD VDD.n3655 0.00406061
R32775 VDD.n244 VDD.n243 0.00170773
R32776 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C.t1 169.46
R32777 D_FlipFlop_6.3-input-nand_2.C.n4 D_FlipFlop_6.3-input-nand_2.C.t2 167.809
R32778 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C.t3 167.809
R32779 D_FlipFlop_6.3-input-nand_2.C.n3 D_FlipFlop_6.3-input-nand_2.C.t5 167.226
R32780 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.t7 150.273
R32781 D_FlipFlop_6.3-input-nand_2.C.t5 D_FlipFlop_6.3-input-nand_2.C.n2 150.273
R32782 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C.t6 73.6406
R32783 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C.t4 73.6304
R32784 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.t0 60.4568
R32785 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.n11 12.3891
R32786 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C.n4 11.4489
R32787 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C 1.68257
R32788 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C.n13 1.38365
R32789 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C.n0 1.19615
R32790 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C.n9 1.1717
R32791 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C 1.08448
R32792 D_FlipFlop_6.3-input-nand_2.C.n10 D_FlipFlop_6.3-input-nand_2.C 0.932141
R32793 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C 0.720633
R32794 D_FlipFlop_6.3-input-nand_2.C.n5 D_FlipFlop_6.3-input-nand_2.C.n3 0.280391
R32795 D_FlipFlop_6.3-input-nand_2.C.n0 D_FlipFlop_6.3-input-nand_2.C 0.217464
R32796 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C 0.1255
R32797 D_FlipFlop_6.3-input-nand_2.C.n1 D_FlipFlop_6.3-input-nand_2.C 0.1255
R32798 D_FlipFlop_6.3-input-nand_2.C.n14 D_FlipFlop_6.3-input-nand_2.C 0.1255
R32799 D_FlipFlop_6.3-input-nand_2.C.n7 D_FlipFlop_6.3-input-nand_2.C.n6 0.0874565
R32800 D_FlipFlop_6.3-input-nand_2.C.n11 D_FlipFlop_6.3-input-nand_2.C.n10 0.063
R32801 D_FlipFlop_6.3-input-nand_2.C.n12 D_FlipFlop_6.3-input-nand_2.C.n7 0.063
R32802 D_FlipFlop_6.3-input-nand_2.C.n13 D_FlipFlop_6.3-input-nand_2.C.n12 0.063
R32803 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.C.n14 0.063
R32804 D_FlipFlop_6.3-input-nand_2.C.n6 D_FlipFlop_6.3-input-nand_2.C.n5 0.0435206
R32805 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C.n1 0.0216397
R32806 D_FlipFlop_6.3-input-nand_2.C.n2 D_FlipFlop_6.3-input-nand_2.C 0.0216397
R32807 D_FlipFlop_6.3-input-nand_2.C.n9 D_FlipFlop_6.3-input-nand_2.C.n8 0.0107679
R32808 D_FlipFlop_6.3-input-nand_2.C.n8 D_FlipFlop_6.3-input-nand_2.C 0.0107679
R32809 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 169.46
R32810 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 167.809
R32811 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 167.809
R32812 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 167.226
R32813 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 150.273
R32814 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 150.273
R32815 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 73.6406
R32816 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 73.6304
R32817 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 60.3943
R32818 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 12.3891
R32819 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 11.4489
R32820 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 1.68257
R32821 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 1.38365
R32822 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 1.19615
R32823 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 1.1717
R32824 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 1.08448
R32825 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.932141
R32826 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.720633
R32827 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 0.280391
R32828 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.217464
R32829 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R32830 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R32831 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.1255
R32832 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 0.0874565
R32833 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 0.063
R32834 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 0.063
R32835 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 0.063
R32836 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 0.063
R32837 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 0.0435206
R32838 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 0.0216397
R32839 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.0216397
R32840 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 0.0107679
R32841 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.0107679
R32842 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 169.46
R32843 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 168.089
R32844 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 167.809
R32845 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 150.293
R32846 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 73.6304
R32847 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 60.4568
R32848 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 12.0358
R32849 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 11.4489
R32850 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.981478
R32851 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 0.788543
R32852 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.769522
R32853 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 0.720633
R32854 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 0.682565
R32855 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.580578
R32856 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 0.55213
R32857 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 0.470609
R32858 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.447191
R32859 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.428234
R32860 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.1255
R32861 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.1255
R32862 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 0.063
R32863 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 0.063
R32864 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.063
R32865 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 0.063
R32866 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 0.063
R32867 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 0.0435206
R32868 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 0.0107679
R32869 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.0107679
R32870 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z.t0 168.635
R32871 CDAC8_0.switch_8.Z CDAC8_0.switch_8.Z.t1 168.571
R32872 CDAC8_0.switch_8.Z.n0 CDAC8_0.switch_8.Z.t2 60.321
R32873 CDAC8_0.switch_8.Z.n0 CDAC8_0.switch_8.Z.t3 60.321
R32874 CDAC8_0.switch_8.Z.n20 CDAC8_0.switch_8.Z.n19 11.3205
R32875 CDAC8_0.switch_8.Z.n15 CDAC8_0.switch_8.Z.n14 5.49497
R32876 CDAC8_0.switch_8.Z.n19 CDAC8_0.switch_8.Z.n3 2.98587
R32877 CDAC8_0.switch_8.Z.n19 CDAC8_0.switch_8.Z.n18 2.5049
R32878 CDAC8_0.switch_8.Z.n2 CDAC8_0.switch_8.Z 1.36463
R32879 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z.n21 1.04126
R32880 CDAC8_0.switch_8.Z.n21 CDAC8_0.switch_8.Z 0.838391
R32881 CDAC8_0.switch_8.Z.n4 CDAC8_0.switch_8.Z.t4 0.77316
R32882 CDAC8_0.switch_8.Z.n10 CDAC8_0.switch_8.Z.t12 0.77316
R32883 CDAC8_0.switch_8.Z.n3 CDAC8_0.switch_8.Z.t14 0.658247
R32884 CDAC8_0.switch_8.Z.n18 CDAC8_0.switch_8.Z.t6 0.658247
R32885 CDAC8_0.switch_8.Z.n8 CDAC8_0.switch_8.Z.t13 0.611304
R32886 CDAC8_0.switch_8.Z.n9 CDAC8_0.switch_8.Z.t18 0.611304
R32887 CDAC8_0.switch_8.Z.n17 CDAC8_0.switch_8.Z.t5 0.611304
R32888 CDAC8_0.switch_8.Z.n16 CDAC8_0.switch_8.Z.t11 0.611304
R32889 CDAC8_0.switch_8.Z.n7 CDAC8_0.switch_8.Z.t9 0.611304
R32890 CDAC8_0.switch_8.Z.n6 CDAC8_0.switch_8.Z.t15 0.611304
R32891 CDAC8_0.switch_8.Z.n5 CDAC8_0.switch_8.Z.t19 0.611304
R32892 CDAC8_0.switch_8.Z.n4 CDAC8_0.switch_8.Z.t17 0.611304
R32893 CDAC8_0.switch_8.Z.n13 CDAC8_0.switch_8.Z.t16 0.611304
R32894 CDAC8_0.switch_8.Z.n12 CDAC8_0.switch_8.Z.t7 0.611304
R32895 CDAC8_0.switch_8.Z.n11 CDAC8_0.switch_8.Z.t10 0.611304
R32896 CDAC8_0.switch_8.Z.n10 CDAC8_0.switch_8.Z.t8 0.611304
R32897 CDAC8_0.switch_8.Z.n2 CDAC8_0.switch_8.Z.n1 0.405391
R32898 CDAC8_0.switch_8.Z.n1 CDAC8_0.switch_8.Z 0.259656
R32899 CDAC8_0.switch_8.Z.n17 CDAC8_0.switch_8.Z.n16 0.162356
R32900 CDAC8_0.switch_8.Z.n7 CDAC8_0.switch_8.Z.n6 0.162356
R32901 CDAC8_0.switch_8.Z.n6 CDAC8_0.switch_8.Z.n5 0.162356
R32902 CDAC8_0.switch_8.Z.n5 CDAC8_0.switch_8.Z.n4 0.162356
R32903 CDAC8_0.switch_8.Z.n9 CDAC8_0.switch_8.Z.n8 0.162356
R32904 CDAC8_0.switch_8.Z.n13 CDAC8_0.switch_8.Z.n12 0.162356
R32905 CDAC8_0.switch_8.Z.n12 CDAC8_0.switch_8.Z.n11 0.162356
R32906 CDAC8_0.switch_8.Z.n11 CDAC8_0.switch_8.Z.n10 0.162356
R32907 CDAC8_0.switch_8.Z.n22 CDAC8_0.switch_8.Z 0.1255
R32908 CDAC8_0.switch_8.Z.n18 CDAC8_0.switch_8.Z.n17 0.115412
R32909 CDAC8_0.switch_8.Z.n8 CDAC8_0.switch_8.Z.n3 0.115412
R32910 CDAC8_0.switch_8.Z.n15 CDAC8_0.switch_8.Z.n7 0.0845094
R32911 CDAC8_0.switch_8.Z.n14 CDAC8_0.switch_8.Z.n13 0.0845094
R32912 CDAC8_0.switch_8.Z.n21 CDAC8_0.switch_8.Z.n20 0.0805781
R32913 CDAC8_0.switch_8.Z.n16 CDAC8_0.switch_8.Z.n15 0.0783469
R32914 CDAC8_0.switch_8.Z.n14 CDAC8_0.switch_8.Z.n9 0.0783469
R32915 CDAC8_0.switch_8.Z.n20 CDAC8_0.switch_8.Z.n2 0.063
R32916 CDAC8_0.switch_8.Z CDAC8_0.switch_8.Z.n22 0.063
R32917 CDAC8_0.switch_8.Z.n1 CDAC8_0.switch_8.Z.n0 0.0188121
R32918 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 179.256
R32919 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 168.089
R32920 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 150.293
R32921 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 73.6304
R32922 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 60.4568
R32923 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 12.0358
R32924 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.981478
R32925 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 0.788543
R32926 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.769522
R32927 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 0.720633
R32928 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 0.682565
R32929 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.580578
R32930 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 0.55213
R32931 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 0.470609
R32932 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.447191
R32933 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.428234
R32934 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1255
R32935 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1255
R32936 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 0.063
R32937 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 0.063
R32938 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.063
R32939 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 0.063
R32940 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 0.063
R32941 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 0.0435206
R32942 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 0.0107679
R32943 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.0107679
R32944 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.t3 168.548
R32945 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.t0 168.548
R32946 CDAC8_0.switch_6.Z.n0 CDAC8_0.switch_6.Z.t1 60.321
R32947 CDAC8_0.switch_6.Z.n0 CDAC8_0.switch_6.Z.t2 60.321
R32948 CDAC8_0.switch_6.Z.n102 CDAC8_0.switch_6.Z.n101 22.979
R32949 CDAC8_0.switch_6.Z.n124 CDAC8_0.switch_6.Z.n123 11.3711
R32950 CDAC8_0.switch_6.Z.n123 CDAC8_0.switch_6.Z.n3 11.3479
R32951 CDAC8_0.switch_6.Z.n123 CDAC8_0.switch_6.Z.n122 10.8669
R32952 CDAC8_0.switch_6.Z.n54 CDAC8_0.switch_6.Z.n53 4.99363
R32953 CDAC8_0.switch_6.Z.n57 CDAC8_0.switch_6.Z.n56 4.99363
R32954 CDAC8_0.switch_6.Z.n65 CDAC8_0.switch_6.Z.n64 4.99363
R32955 CDAC8_0.switch_6.Z.n70 CDAC8_0.switch_6.Z.n69 4.99363
R32956 CDAC8_0.switch_6.Z.n73 CDAC8_0.switch_6.Z.n72 4.99363
R32957 CDAC8_0.switch_6.Z.n76 CDAC8_0.switch_6.Z.n75 4.99363
R32958 CDAC8_0.switch_6.Z.n79 CDAC8_0.switch_6.Z.n78 4.99363
R32959 CDAC8_0.switch_6.Z.n83 CDAC8_0.switch_6.Z.n82 4.99363
R32960 CDAC8_0.switch_6.Z.n85 CDAC8_0.switch_6.Z.n43 4.99363
R32961 CDAC8_0.switch_6.Z.n9 CDAC8_0.switch_6.Z.n8 4.99363
R32962 CDAC8_0.switch_6.Z.n12 CDAC8_0.switch_6.Z.n11 4.99363
R32963 CDAC8_0.switch_6.Z.n15 CDAC8_0.switch_6.Z.n14 4.99363
R32964 CDAC8_0.switch_6.Z.n19 CDAC8_0.switch_6.Z.n18 4.99363
R32965 CDAC8_0.switch_6.Z.n119 CDAC8_0.switch_6.Z.n118 4.99363
R32966 CDAC8_0.switch_6.Z.n116 CDAC8_0.switch_6.Z.n115 4.99363
R32967 CDAC8_0.switch_6.Z.n113 CDAC8_0.switch_6.Z.n112 4.99363
R32968 CDAC8_0.switch_6.Z.n110 CDAC8_0.switch_6.Z.n109 4.99363
R32969 CDAC8_0.switch_6.Z.n107 CDAC8_0.switch_6.Z.n106 4.99363
R32970 CDAC8_0.switch_6.Z.n104 CDAC8_0.switch_6.Z.n103 4.99363
R32971 CDAC8_0.switch_6.Z.n41 CDAC8_0.switch_6.Z.n40 4.99363
R32972 CDAC8_0.switch_6.Z.n38 CDAC8_0.switch_6.Z.n37 4.99363
R32973 CDAC8_0.switch_6.Z.n35 CDAC8_0.switch_6.Z.n34 4.99363
R32974 CDAC8_0.switch_6.Z.n32 CDAC8_0.switch_6.Z.n31 4.99363
R32975 CDAC8_0.switch_6.Z.n99 CDAC8_0.switch_6.Z.n98 4.99363
R32976 CDAC8_0.switch_6.Z.n96 CDAC8_0.switch_6.Z.n95 4.99363
R32977 CDAC8_0.switch_6.Z.n93 CDAC8_0.switch_6.Z.n92 4.99363
R32978 CDAC8_0.switch_6.Z.n90 CDAC8_0.switch_6.Z.n89 4.99363
R32979 CDAC8_0.switch_6.Z.n122 CDAC8_0.switch_6.Z.n4 4.61363
R32980 CDAC8_0.switch_6.Z.n62 CDAC8_0.switch_6.Z.n3 4.61363
R32981 CDAC8_0.switch_6.Z.n60 CDAC8_0.switch_6.Z.n59 3.9471
R32982 CDAC8_0.switch_6.Z.n2 CDAC8_0.switch_6.Z.n1 1.58202
R32983 CDAC8_0.switch_6.Z.n32 CDAC8_0.switch_6.Z.t5 0.726216
R32984 CDAC8_0.switch_6.Z.n31 CDAC8_0.switch_6.Z.t37 0.726216
R32985 CDAC8_0.switch_6.Z.n89 CDAC8_0.switch_6.Z.t50 0.726216
R32986 CDAC8_0.switch_6.Z.n90 CDAC8_0.switch_6.Z.t36 0.726216
R32987 CDAC8_0.switch_6.Z.n54 CDAC8_0.switch_6.Z.t31 0.658247
R32988 CDAC8_0.switch_6.Z.n53 CDAC8_0.switch_6.Z.t47 0.658247
R32989 CDAC8_0.switch_6.Z.n8 CDAC8_0.switch_6.Z.t32 0.658247
R32990 CDAC8_0.switch_6.Z.n9 CDAC8_0.switch_6.Z.t63 0.658247
R32991 CDAC8_0.switch_6.Z.n55 CDAC8_0.switch_6.Z.t28 0.611304
R32992 CDAC8_0.switch_6.Z.n51 CDAC8_0.switch_6.Z.t44 0.611304
R32993 CDAC8_0.switch_6.Z.n61 CDAC8_0.switch_6.Z.t40 0.611304
R32994 CDAC8_0.switch_6.Z.n63 CDAC8_0.switch_6.Z.t66 0.611304
R32995 CDAC8_0.switch_6.Z.n49 CDAC8_0.switch_6.Z.t11 0.611304
R32996 CDAC8_0.switch_6.Z.n71 CDAC8_0.switch_6.Z.t8 0.611304
R32997 CDAC8_0.switch_6.Z.n47 CDAC8_0.switch_6.Z.t19 0.611304
R32998 CDAC8_0.switch_6.Z.n77 CDAC8_0.switch_6.Z.t16 0.611304
R32999 CDAC8_0.switch_6.Z.n45 CDAC8_0.switch_6.Z.t48 0.611304
R33000 CDAC8_0.switch_6.Z.n84 CDAC8_0.switch_6.Z.t57 0.611304
R33001 CDAC8_0.switch_6.Z.n86 CDAC8_0.switch_6.Z.t55 0.611304
R33002 CDAC8_0.switch_6.Z.n97 CDAC8_0.switch_6.Z.t64 0.611304
R33003 CDAC8_0.switch_6.Z.n87 CDAC8_0.switch_6.Z.t26 0.611304
R33004 CDAC8_0.switch_6.Z.n91 CDAC8_0.switch_6.Z.t24 0.611304
R33005 CDAC8_0.switch_6.Z.n52 CDAC8_0.switch_6.Z.t43 0.611304
R33006 CDAC8_0.switch_6.Z.n58 CDAC8_0.switch_6.Z.t54 0.611304
R33007 CDAC8_0.switch_6.Z.n50 CDAC8_0.switch_6.Z.t52 0.611304
R33008 CDAC8_0.switch_6.Z.n66 CDAC8_0.switch_6.Z.t14 0.611304
R33009 CDAC8_0.switch_6.Z.n68 CDAC8_0.switch_6.Z.t21 0.611304
R33010 CDAC8_0.switch_6.Z.n48 CDAC8_0.switch_6.Z.t18 0.611304
R33011 CDAC8_0.switch_6.Z.n74 CDAC8_0.switch_6.Z.t35 0.611304
R33012 CDAC8_0.switch_6.Z.n46 CDAC8_0.switch_6.Z.t30 0.611304
R33013 CDAC8_0.switch_6.Z.n80 CDAC8_0.switch_6.Z.t60 0.611304
R33014 CDAC8_0.switch_6.Z.n81 CDAC8_0.switch_6.Z.t6 0.611304
R33015 CDAC8_0.switch_6.Z.n7 CDAC8_0.switch_6.Z.t29 0.611304
R33016 CDAC8_0.switch_6.Z.n13 CDAC8_0.switch_6.Z.t45 0.611304
R33017 CDAC8_0.switch_6.Z.n5 CDAC8_0.switch_6.Z.t41 0.611304
R33018 CDAC8_0.switch_6.Z.n20 CDAC8_0.switch_6.Z.t67 0.611304
R33019 CDAC8_0.switch_6.Z.n120 CDAC8_0.switch_6.Z.t12 0.611304
R33020 CDAC8_0.switch_6.Z.n21 CDAC8_0.switch_6.Z.t9 0.611304
R33021 CDAC8_0.switch_6.Z.n114 CDAC8_0.switch_6.Z.t20 0.611304
R33022 CDAC8_0.switch_6.Z.n24 CDAC8_0.switch_6.Z.t17 0.611304
R33023 CDAC8_0.switch_6.Z.n108 CDAC8_0.switch_6.Z.t49 0.611304
R33024 CDAC8_0.switch_6.Z.n26 CDAC8_0.switch_6.Z.t58 0.611304
R33025 CDAC8_0.switch_6.Z.n42 CDAC8_0.switch_6.Z.t56 0.611304
R33026 CDAC8_0.switch_6.Z.n28 CDAC8_0.switch_6.Z.t65 0.611304
R33027 CDAC8_0.switch_6.Z.n36 CDAC8_0.switch_6.Z.t27 0.611304
R33028 CDAC8_0.switch_6.Z.n30 CDAC8_0.switch_6.Z.t25 0.611304
R33029 CDAC8_0.switch_6.Z.n10 CDAC8_0.switch_6.Z.t62 0.611304
R33030 CDAC8_0.switch_6.Z.n6 CDAC8_0.switch_6.Z.t10 0.611304
R33031 CDAC8_0.switch_6.Z.n16 CDAC8_0.switch_6.Z.t7 0.611304
R33032 CDAC8_0.switch_6.Z.n17 CDAC8_0.switch_6.Z.t34 0.611304
R33033 CDAC8_0.switch_6.Z.n22 CDAC8_0.switch_6.Z.t46 0.611304
R33034 CDAC8_0.switch_6.Z.n117 CDAC8_0.switch_6.Z.t42 0.611304
R33035 CDAC8_0.switch_6.Z.n23 CDAC8_0.switch_6.Z.t53 0.611304
R33036 CDAC8_0.switch_6.Z.n111 CDAC8_0.switch_6.Z.t51 0.611304
R33037 CDAC8_0.switch_6.Z.n25 CDAC8_0.switch_6.Z.t15 0.611304
R33038 CDAC8_0.switch_6.Z.n105 CDAC8_0.switch_6.Z.t23 0.611304
R33039 CDAC8_0.switch_6.Z.n27 CDAC8_0.switch_6.Z.t22 0.611304
R33040 CDAC8_0.switch_6.Z.n39 CDAC8_0.switch_6.Z.t33 0.611304
R33041 CDAC8_0.switch_6.Z.n29 CDAC8_0.switch_6.Z.t61 0.611304
R33042 CDAC8_0.switch_6.Z.n33 CDAC8_0.switch_6.Z.t59 0.611304
R33043 CDAC8_0.switch_6.Z.n100 CDAC8_0.switch_6.Z.t4 0.611304
R33044 CDAC8_0.switch_6.Z.n44 CDAC8_0.switch_6.Z.t13 0.611304
R33045 CDAC8_0.switch_6.Z.n94 CDAC8_0.switch_6.Z.t39 0.611304
R33046 CDAC8_0.switch_6.Z.n88 CDAC8_0.switch_6.Z.t38 0.611304
R33047 CDAC8_0.switch_6.Z.n122 CDAC8_0.switch_6.Z.n121 0.3805
R33048 CDAC8_0.switch_6.Z.n67 CDAC8_0.switch_6.Z.n3 0.3805
R33049 CDAC8_0.switch_6.Z.n1 CDAC8_0.switch_6.Z 0.259656
R33050 CDAC8_0.switch_6.Z.n2 CDAC8_0.switch_6.Z 0.188
R33051 CDAC8_0.switch_6.Z.n10 CDAC8_0.switch_6.Z.n9 0.115412
R33052 CDAC8_0.switch_6.Z.n11 CDAC8_0.switch_6.Z.n6 0.115412
R33053 CDAC8_0.switch_6.Z.n16 CDAC8_0.switch_6.Z.n15 0.115412
R33054 CDAC8_0.switch_6.Z.n18 CDAC8_0.switch_6.Z.n17 0.115412
R33055 CDAC8_0.switch_6.Z.n22 CDAC8_0.switch_6.Z.n4 0.115412
R33056 CDAC8_0.switch_6.Z.n118 CDAC8_0.switch_6.Z.n117 0.115412
R33057 CDAC8_0.switch_6.Z.n116 CDAC8_0.switch_6.Z.n23 0.115412
R33058 CDAC8_0.switch_6.Z.n112 CDAC8_0.switch_6.Z.n111 0.115412
R33059 CDAC8_0.switch_6.Z.n110 CDAC8_0.switch_6.Z.n25 0.115412
R33060 CDAC8_0.switch_6.Z.n106 CDAC8_0.switch_6.Z.n105 0.115412
R33061 CDAC8_0.switch_6.Z.n104 CDAC8_0.switch_6.Z.n27 0.115412
R33062 CDAC8_0.switch_6.Z.n40 CDAC8_0.switch_6.Z.n39 0.115412
R33063 CDAC8_0.switch_6.Z.n38 CDAC8_0.switch_6.Z.n29 0.115412
R33064 CDAC8_0.switch_6.Z.n34 CDAC8_0.switch_6.Z.n33 0.115412
R33065 CDAC8_0.switch_6.Z.n8 CDAC8_0.switch_6.Z.n7 0.115412
R33066 CDAC8_0.switch_6.Z.n13 CDAC8_0.switch_6.Z.n12 0.115412
R33067 CDAC8_0.switch_6.Z.n14 CDAC8_0.switch_6.Z.n5 0.115412
R33068 CDAC8_0.switch_6.Z.n20 CDAC8_0.switch_6.Z.n19 0.115412
R33069 CDAC8_0.switch_6.Z.n121 CDAC8_0.switch_6.Z.n120 0.115412
R33070 CDAC8_0.switch_6.Z.n119 CDAC8_0.switch_6.Z.n21 0.115412
R33071 CDAC8_0.switch_6.Z.n115 CDAC8_0.switch_6.Z.n114 0.115412
R33072 CDAC8_0.switch_6.Z.n113 CDAC8_0.switch_6.Z.n24 0.115412
R33073 CDAC8_0.switch_6.Z.n109 CDAC8_0.switch_6.Z.n108 0.115412
R33074 CDAC8_0.switch_6.Z.n107 CDAC8_0.switch_6.Z.n26 0.115412
R33075 CDAC8_0.switch_6.Z.n41 CDAC8_0.switch_6.Z.n28 0.115412
R33076 CDAC8_0.switch_6.Z.n37 CDAC8_0.switch_6.Z.n36 0.115412
R33077 CDAC8_0.switch_6.Z.n35 CDAC8_0.switch_6.Z.n30 0.115412
R33078 CDAC8_0.switch_6.Z.n53 CDAC8_0.switch_6.Z.n52 0.115412
R33079 CDAC8_0.switch_6.Z.n58 CDAC8_0.switch_6.Z.n57 0.115412
R33080 CDAC8_0.switch_6.Z.n59 CDAC8_0.switch_6.Z.n50 0.115412
R33081 CDAC8_0.switch_6.Z.n66 CDAC8_0.switch_6.Z.n65 0.115412
R33082 CDAC8_0.switch_6.Z.n68 CDAC8_0.switch_6.Z.n67 0.115412
R33083 CDAC8_0.switch_6.Z.n69 CDAC8_0.switch_6.Z.n48 0.115412
R33084 CDAC8_0.switch_6.Z.n74 CDAC8_0.switch_6.Z.n73 0.115412
R33085 CDAC8_0.switch_6.Z.n75 CDAC8_0.switch_6.Z.n46 0.115412
R33086 CDAC8_0.switch_6.Z.n80 CDAC8_0.switch_6.Z.n79 0.115412
R33087 CDAC8_0.switch_6.Z.n82 CDAC8_0.switch_6.Z.n81 0.115412
R33088 CDAC8_0.switch_6.Z.n99 CDAC8_0.switch_6.Z.n44 0.115412
R33089 CDAC8_0.switch_6.Z.n95 CDAC8_0.switch_6.Z.n94 0.115412
R33090 CDAC8_0.switch_6.Z.n93 CDAC8_0.switch_6.Z.n88 0.115412
R33091 CDAC8_0.switch_6.Z.n55 CDAC8_0.switch_6.Z.n54 0.115412
R33092 CDAC8_0.switch_6.Z.n56 CDAC8_0.switch_6.Z.n51 0.115412
R33093 CDAC8_0.switch_6.Z.n61 CDAC8_0.switch_6.Z.n60 0.115412
R33094 CDAC8_0.switch_6.Z.n64 CDAC8_0.switch_6.Z.n63 0.115412
R33095 CDAC8_0.switch_6.Z.n62 CDAC8_0.switch_6.Z.n49 0.115412
R33096 CDAC8_0.switch_6.Z.n71 CDAC8_0.switch_6.Z.n70 0.115412
R33097 CDAC8_0.switch_6.Z.n72 CDAC8_0.switch_6.Z.n47 0.115412
R33098 CDAC8_0.switch_6.Z.n77 CDAC8_0.switch_6.Z.n76 0.115412
R33099 CDAC8_0.switch_6.Z.n78 CDAC8_0.switch_6.Z.n45 0.115412
R33100 CDAC8_0.switch_6.Z.n84 CDAC8_0.switch_6.Z.n83 0.115412
R33101 CDAC8_0.switch_6.Z.n86 CDAC8_0.switch_6.Z.n85 0.115412
R33102 CDAC8_0.switch_6.Z.n98 CDAC8_0.switch_6.Z.n97 0.115412
R33103 CDAC8_0.switch_6.Z.n96 CDAC8_0.switch_6.Z.n87 0.115412
R33104 CDAC8_0.switch_6.Z.n92 CDAC8_0.switch_6.Z.n91 0.115412
R33105 CDAC8_0.switch_6.Z.n102 CDAC8_0.switch_6.Z.n42 0.0845094
R33106 CDAC8_0.switch_6.Z.n101 CDAC8_0.switch_6.Z.n100 0.0845094
R33107 CDAC8_0.switch_6.Z.n124 CDAC8_0.switch_6.Z.n2 0.063
R33108 CDAC8_0.switch_6.Z.n11 CDAC8_0.switch_6.Z.n10 0.0474438
R33109 CDAC8_0.switch_6.Z.n15 CDAC8_0.switch_6.Z.n6 0.0474438
R33110 CDAC8_0.switch_6.Z.n18 CDAC8_0.switch_6.Z.n16 0.0474438
R33111 CDAC8_0.switch_6.Z.n17 CDAC8_0.switch_6.Z.n4 0.0474438
R33112 CDAC8_0.switch_6.Z.n118 CDAC8_0.switch_6.Z.n22 0.0474438
R33113 CDAC8_0.switch_6.Z.n117 CDAC8_0.switch_6.Z.n116 0.0474438
R33114 CDAC8_0.switch_6.Z.n112 CDAC8_0.switch_6.Z.n23 0.0474438
R33115 CDAC8_0.switch_6.Z.n111 CDAC8_0.switch_6.Z.n110 0.0474438
R33116 CDAC8_0.switch_6.Z.n106 CDAC8_0.switch_6.Z.n25 0.0474438
R33117 CDAC8_0.switch_6.Z.n105 CDAC8_0.switch_6.Z.n104 0.0474438
R33118 CDAC8_0.switch_6.Z.n40 CDAC8_0.switch_6.Z.n27 0.0474438
R33119 CDAC8_0.switch_6.Z.n39 CDAC8_0.switch_6.Z.n38 0.0474438
R33120 CDAC8_0.switch_6.Z.n34 CDAC8_0.switch_6.Z.n29 0.0474438
R33121 CDAC8_0.switch_6.Z.n33 CDAC8_0.switch_6.Z.n32 0.0474438
R33122 CDAC8_0.switch_6.Z.n12 CDAC8_0.switch_6.Z.n7 0.0474438
R33123 CDAC8_0.switch_6.Z.n14 CDAC8_0.switch_6.Z.n13 0.0474438
R33124 CDAC8_0.switch_6.Z.n19 CDAC8_0.switch_6.Z.n5 0.0474438
R33125 CDAC8_0.switch_6.Z.n121 CDAC8_0.switch_6.Z.n20 0.0474438
R33126 CDAC8_0.switch_6.Z.n120 CDAC8_0.switch_6.Z.n119 0.0474438
R33127 CDAC8_0.switch_6.Z.n115 CDAC8_0.switch_6.Z.n21 0.0474438
R33128 CDAC8_0.switch_6.Z.n114 CDAC8_0.switch_6.Z.n113 0.0474438
R33129 CDAC8_0.switch_6.Z.n109 CDAC8_0.switch_6.Z.n24 0.0474438
R33130 CDAC8_0.switch_6.Z.n108 CDAC8_0.switch_6.Z.n107 0.0474438
R33131 CDAC8_0.switch_6.Z.n103 CDAC8_0.switch_6.Z.n26 0.0474438
R33132 CDAC8_0.switch_6.Z.n42 CDAC8_0.switch_6.Z.n41 0.0474438
R33133 CDAC8_0.switch_6.Z.n37 CDAC8_0.switch_6.Z.n28 0.0474438
R33134 CDAC8_0.switch_6.Z.n36 CDAC8_0.switch_6.Z.n35 0.0474438
R33135 CDAC8_0.switch_6.Z.n31 CDAC8_0.switch_6.Z.n30 0.0474438
R33136 CDAC8_0.switch_6.Z.n57 CDAC8_0.switch_6.Z.n52 0.0474438
R33137 CDAC8_0.switch_6.Z.n59 CDAC8_0.switch_6.Z.n58 0.0474438
R33138 CDAC8_0.switch_6.Z.n65 CDAC8_0.switch_6.Z.n50 0.0474438
R33139 CDAC8_0.switch_6.Z.n67 CDAC8_0.switch_6.Z.n66 0.0474438
R33140 CDAC8_0.switch_6.Z.n69 CDAC8_0.switch_6.Z.n68 0.0474438
R33141 CDAC8_0.switch_6.Z.n73 CDAC8_0.switch_6.Z.n48 0.0474438
R33142 CDAC8_0.switch_6.Z.n75 CDAC8_0.switch_6.Z.n74 0.0474438
R33143 CDAC8_0.switch_6.Z.n79 CDAC8_0.switch_6.Z.n46 0.0474438
R33144 CDAC8_0.switch_6.Z.n82 CDAC8_0.switch_6.Z.n80 0.0474438
R33145 CDAC8_0.switch_6.Z.n81 CDAC8_0.switch_6.Z.n43 0.0474438
R33146 CDAC8_0.switch_6.Z.n100 CDAC8_0.switch_6.Z.n99 0.0474438
R33147 CDAC8_0.switch_6.Z.n95 CDAC8_0.switch_6.Z.n44 0.0474438
R33148 CDAC8_0.switch_6.Z.n94 CDAC8_0.switch_6.Z.n93 0.0474438
R33149 CDAC8_0.switch_6.Z.n89 CDAC8_0.switch_6.Z.n88 0.0474438
R33150 CDAC8_0.switch_6.Z.n56 CDAC8_0.switch_6.Z.n55 0.0474438
R33151 CDAC8_0.switch_6.Z.n60 CDAC8_0.switch_6.Z.n51 0.0474438
R33152 CDAC8_0.switch_6.Z.n64 CDAC8_0.switch_6.Z.n61 0.0474438
R33153 CDAC8_0.switch_6.Z.n63 CDAC8_0.switch_6.Z.n62 0.0474438
R33154 CDAC8_0.switch_6.Z.n70 CDAC8_0.switch_6.Z.n49 0.0474438
R33155 CDAC8_0.switch_6.Z.n72 CDAC8_0.switch_6.Z.n71 0.0474438
R33156 CDAC8_0.switch_6.Z.n76 CDAC8_0.switch_6.Z.n47 0.0474438
R33157 CDAC8_0.switch_6.Z.n78 CDAC8_0.switch_6.Z.n77 0.0474438
R33158 CDAC8_0.switch_6.Z.n83 CDAC8_0.switch_6.Z.n45 0.0474438
R33159 CDAC8_0.switch_6.Z.n85 CDAC8_0.switch_6.Z.n84 0.0474438
R33160 CDAC8_0.switch_6.Z.n98 CDAC8_0.switch_6.Z.n86 0.0474438
R33161 CDAC8_0.switch_6.Z.n97 CDAC8_0.switch_6.Z.n96 0.0474438
R33162 CDAC8_0.switch_6.Z.n92 CDAC8_0.switch_6.Z.n87 0.0474438
R33163 CDAC8_0.switch_6.Z.n91 CDAC8_0.switch_6.Z.n90 0.0474438
R33164 CDAC8_0.switch_6.Z CDAC8_0.switch_6.Z.n125 0.0454219
R33165 CDAC8_0.switch_6.Z.n103 CDAC8_0.switch_6.Z.n102 0.0314031
R33166 CDAC8_0.switch_6.Z.n101 CDAC8_0.switch_6.Z.n43 0.0314031
R33167 CDAC8_0.switch_6.Z.n125 CDAC8_0.switch_6.Z.n124 0.0278438
R33168 CDAC8_0.switch_6.Z.n1 CDAC8_0.switch_6.Z.n0 0.0188121
R33169 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout.t3 169.46
R33170 D_FlipFlop_1.3-input-nand_2.Vout.n4 D_FlipFlop_1.3-input-nand_2.Vout.t2 167.809
R33171 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout.t1 167.809
R33172 D_FlipFlop_1.3-input-nand_2.Vout.n3 D_FlipFlop_1.3-input-nand_2.Vout.t4 167.227
R33173 D_FlipFlop_1.3-input-nand_2.Vout.t4 D_FlipFlop_1.3-input-nand_2.Vout.n2 150.293
R33174 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.t7 150.273
R33175 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout.t5 73.6406
R33176 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout.t6 73.6304
R33177 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.t0 60.3809
R33178 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout.n9 12.3891
R33179 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.n4 11.4489
R33180 D_FlipFlop_1.3-input-nand_2.Vout.n12 D_FlipFlop_1.3-input-nand_2.Vout.n11 1.38365
R33181 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout.n1 1.19615
R33182 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout.n8 1.1717
R33183 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.Vout.n12 0.848156
R33184 D_FlipFlop_1.3-input-nand_2.Vout.n2 D_FlipFlop_1.3-input-nand_2.Vout 0.447191
R33185 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R33186 D_FlipFlop_1.3-input-nand_2.Vout.n5 D_FlipFlop_1.3-input-nand_2.Vout.n3 0.280391
R33187 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout.n5 0.262643
R33188 D_FlipFlop_1.3-input-nand_2.Vout.n8 D_FlipFlop_1.3-input-nand_2.Vout 0.217464
R33189 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R33190 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R33191 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R33192 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R33193 D_FlipFlop_1.3-input-nand_2.Vout.n7 D_FlipFlop_1.3-input-nand_2.Vout.n6 0.0874565
R33194 D_FlipFlop_1.3-input-nand_2.Vout.n6 D_FlipFlop_1.3-input-nand_2.Vout 0.063
R33195 D_FlipFlop_1.3-input-nand_2.Vout.n11 D_FlipFlop_1.3-input-nand_2.Vout.n10 0.063
R33196 D_FlipFlop_1.3-input-nand_2.Vout.n10 D_FlipFlop_1.3-input-nand_2.Vout.n7 0.063
R33197 D_FlipFlop_1.3-input-nand_2.Vout.n9 D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R33198 D_FlipFlop_1.3-input-nand_2.Vout.n1 D_FlipFlop_1.3-input-nand_2.Vout.n0 0.0107679
R33199 D_FlipFlop_1.3-input-nand_2.Vout.n0 D_FlipFlop_1.3-input-nand_2.Vout 0.0107679
R33200 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t0 169.46
R33201 D_FlipFlop_1.3-input-nand_2.C.n11 D_FlipFlop_1.3-input-nand_2.C.t1 167.809
R33202 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.t3 167.809
R33203 D_FlipFlop_1.3-input-nand_2.C.t7 D_FlipFlop_1.3-input-nand_2.C.n13 167.226
R33204 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C.t4 150.273
R33205 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.t7 150.273
R33206 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C.t6 73.6406
R33207 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C.t5 73.6304
R33208 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C.t2 60.4568
R33209 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C.n7 12.3891
R33210 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.n11 11.4489
R33211 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C 1.68257
R33212 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C.n2 1.38365
R33213 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C.n0 1.19615
R33214 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C.n5 1.1717
R33215 D_FlipFlop_1.3-input-nand_2.C.n3 D_FlipFlop_1.3-input-nand_2.C 1.08448
R33216 D_FlipFlop_1.3-input-nand_2.C.n6 D_FlipFlop_1.3-input-nand_2.C 0.932141
R33217 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C 0.720633
R33218 D_FlipFlop_1.3-input-nand_2.C.n13 D_FlipFlop_1.3-input-nand_2.C.n12 0.280391
R33219 D_FlipFlop_1.3-input-nand_2.C.n0 D_FlipFlop_1.3-input-nand_2.C 0.217464
R33220 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C 0.1255
R33221 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C 0.1255
R33222 D_FlipFlop_1.3-input-nand_2.C.n1 D_FlipFlop_1.3-input-nand_2.C 0.1255
R33223 D_FlipFlop_1.3-input-nand_2.C.n10 D_FlipFlop_1.3-input-nand_2.C.n9 0.0874565
R33224 D_FlipFlop_1.3-input-nand_2.C.n7 D_FlipFlop_1.3-input-nand_2.C.n6 0.063
R33225 D_FlipFlop_1.3-input-nand_2.C.n2 D_FlipFlop_1.3-input-nand_2.C 0.063
R33226 D_FlipFlop_1.3-input-nand_2.C.n9 D_FlipFlop_1.3-input-nand_2.C.n8 0.063
R33227 D_FlipFlop_1.3-input-nand_2.C.n8 D_FlipFlop_1.3-input-nand_2.C.n3 0.063
R33228 D_FlipFlop_1.3-input-nand_2.C.n12 D_FlipFlop_1.3-input-nand_2.C.n10 0.0435206
R33229 D_FlipFlop_1.3-input-nand_2.C.n14 D_FlipFlop_1.3-input-nand_2.C.n1 0.0216397
R33230 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.C.n14 0.0216397
R33231 D_FlipFlop_1.3-input-nand_2.C.n5 D_FlipFlop_1.3-input-nand_2.C.n4 0.0107679
R33232 D_FlipFlop_1.3-input-nand_2.C.n4 D_FlipFlop_1.3-input-nand_2.C 0.0107679
R33233 D_FlipFlop_0.D.n104 D_FlipFlop_0.D.t16 150.273
R33234 D_FlipFlop_0.D.n110 D_FlipFlop_0.D.t7 150.273
R33235 D_FlipFlop_0.D.n7 D_FlipFlop_0.D.t30 150.273
R33236 D_FlipFlop_0.D.n13 D_FlipFlop_0.D.t23 150.273
R33237 D_FlipFlop_0.D.n20 D_FlipFlop_0.D.t11 150.273
R33238 D_FlipFlop_0.D.n26 D_FlipFlop_0.D.t32 150.273
R33239 D_FlipFlop_0.D.n34 D_FlipFlop_0.D.t17 150.273
R33240 D_FlipFlop_0.D.n40 D_FlipFlop_0.D.t8 150.273
R33241 D_FlipFlop_0.D.n48 D_FlipFlop_0.D.t29 150.273
R33242 D_FlipFlop_0.D.n54 D_FlipFlop_0.D.t22 150.273
R33243 D_FlipFlop_0.D.n62 D_FlipFlop_0.D.t13 150.273
R33244 D_FlipFlop_0.D.n68 D_FlipFlop_0.D.t3 150.273
R33245 D_FlipFlop_0.D.n89 D_FlipFlop_0.D.t18 150.273
R33246 D_FlipFlop_0.D.n95 D_FlipFlop_0.D.t9 150.273
R33247 D_FlipFlop_0.D.n76 D_FlipFlop_0.D.t12 150.273
R33248 D_FlipFlop_0.D.n82 D_FlipFlop_0.D.t34 150.273
R33249 D_FlipFlop_0.D.n102 D_FlipFlop_0.D.t5 73.6406
R33250 D_FlipFlop_0.D.n108 D_FlipFlop_0.D.t10 73.6406
R33251 D_FlipFlop_0.D.n5 D_FlipFlop_0.D.t20 73.6406
R33252 D_FlipFlop_0.D.n11 D_FlipFlop_0.D.t27 73.6406
R33253 D_FlipFlop_0.D.n18 D_FlipFlop_0.D.t31 73.6406
R33254 D_FlipFlop_0.D.n24 D_FlipFlop_0.D.t4 73.6406
R33255 D_FlipFlop_0.D.n32 D_FlipFlop_0.D.t14 73.6406
R33256 D_FlipFlop_0.D.n38 D_FlipFlop_0.D.t24 73.6406
R33257 D_FlipFlop_0.D.n46 D_FlipFlop_0.D.t19 73.6406
R33258 D_FlipFlop_0.D.n52 D_FlipFlop_0.D.t26 73.6406
R33259 D_FlipFlop_0.D.n60 D_FlipFlop_0.D.t21 73.6406
R33260 D_FlipFlop_0.D.n66 D_FlipFlop_0.D.t28 73.6406
R33261 D_FlipFlop_0.D.n87 D_FlipFlop_0.D.t15 73.6406
R33262 D_FlipFlop_0.D.n93 D_FlipFlop_0.D.t25 73.6406
R33263 D_FlipFlop_0.D.n74 D_FlipFlop_0.D.t33 73.6406
R33264 D_FlipFlop_0.D.n80 D_FlipFlop_0.D.t6 73.6406
R33265 D_FlipFlop_0.D.n1 D_FlipFlop_0.D.t2 33.6184
R33266 D_FlipFlop_0.D.n1 D_FlipFlop_0.D.t1 28.6263
R33267 D_FlipFlop_0.D.n114 D_FlipFlop_0.D.n113 8.12822
R33268 D_FlipFlop_0.D.n17 D_FlipFlop_0.D.n16 8.12822
R33269 D_FlipFlop_0.D.n30 D_FlipFlop_0.D.n29 8.12822
R33270 D_FlipFlop_0.D.n44 D_FlipFlop_0.D.n43 8.12822
R33271 D_FlipFlop_0.D.n58 D_FlipFlop_0.D.n57 8.12822
R33272 D_FlipFlop_0.D.n72 D_FlipFlop_0.D.n71 8.12822
R33273 D_FlipFlop_0.D.n99 D_FlipFlop_0.D.n98 8.12822
R33274 D_FlipFlop_0.D.n86 D_FlipFlop_0.D.n85 8.12822
R33275 D_FlipFlop_0.D.n31 D_FlipFlop_0.D.n17 7.52349
R33276 D_FlipFlop_0.D.n100 D_FlipFlop_0.D.n86 7.52349
R33277 D_FlipFlop_0.D.n31 D_FlipFlop_0.D.n30 7.2005
R33278 D_FlipFlop_0.D.n45 D_FlipFlop_0.D.n44 7.2005
R33279 D_FlipFlop_0.D.n59 D_FlipFlop_0.D.n58 7.2005
R33280 D_FlipFlop_0.D.n73 D_FlipFlop_0.D.n72 7.2005
R33281 D_FlipFlop_0.D.n100 D_FlipFlop_0.D.n99 7.2005
R33282 D_FlipFlop_0.D.n115 D_FlipFlop_0.D.n114 6.8205
R33283 D_FlipFlop_0.D.n114 D_FlipFlop_0.D.n107 4.5005
R33284 D_FlipFlop_0.D.n17 D_FlipFlop_0.D.n10 4.5005
R33285 D_FlipFlop_0.D.n30 D_FlipFlop_0.D.n23 4.5005
R33286 D_FlipFlop_0.D.n44 D_FlipFlop_0.D.n37 4.5005
R33287 D_FlipFlop_0.D.n58 D_FlipFlop_0.D.n51 4.5005
R33288 D_FlipFlop_0.D.n72 D_FlipFlop_0.D.n65 4.5005
R33289 D_FlipFlop_0.D.n99 D_FlipFlop_0.D.n92 4.5005
R33290 D_FlipFlop_0.D.n86 D_FlipFlop_0.D.n79 4.5005
R33291 D_FlipFlop_0.D.n4 D_FlipFlop_0.D.n1 3.8456
R33292 D_FlipFlop_0.D.n116 D_FlipFlop_0.D.n115 2.08738
R33293 D_FlipFlop_0.D.n0 D_FlipFlop_0.D.t35 1.13717
R33294 D_FlipFlop_0.D.n3 D_FlipFlop_0.D.n2 0.855396
R33295 D_FlipFlop_0.D.n103 D_FlipFlop_5.Inverter_0.Vin 0.851043
R33296 D_FlipFlop_0.D.n109 D_FlipFlop_5.3-input-nand_0.B 0.851043
R33297 D_FlipFlop_0.D.n6 D_FlipFlop_0.Inverter_0.Vin 0.851043
R33298 D_FlipFlop_0.D.n12 D_FlipFlop_0.3-input-nand_0.B 0.851043
R33299 D_FlipFlop_0.D.n19 D_FlipFlop_3.Inverter_0.Vin 0.851043
R33300 D_FlipFlop_0.D.n25 D_FlipFlop_3.3-input-nand_0.B 0.851043
R33301 D_FlipFlop_0.D.n33 D_FlipFlop_2.Inverter_0.Vin 0.851043
R33302 D_FlipFlop_0.D.n39 D_FlipFlop_2.3-input-nand_0.B 0.851043
R33303 D_FlipFlop_0.D.n47 D_FlipFlop_1.Inverter_0.Vin 0.851043
R33304 D_FlipFlop_0.D.n53 D_FlipFlop_1.3-input-nand_0.B 0.851043
R33305 D_FlipFlop_0.D.n61 D_FlipFlop_4.Inverter_0.Vin 0.851043
R33306 D_FlipFlop_0.D.n67 D_FlipFlop_4.3-input-nand_0.B 0.851043
R33307 D_FlipFlop_0.D.n88 D_FlipFlop_6.Inverter_0.Vin 0.851043
R33308 D_FlipFlop_0.D.n94 D_FlipFlop_6.3-input-nand_0.B 0.851043
R33309 D_FlipFlop_0.D.n75 D_FlipFlop_7.Inverter_0.Vin 0.851043
R33310 D_FlipFlop_0.D.n81 D_FlipFlop_7.3-input-nand_0.B 0.851043
R33311 D_FlipFlop_0.D.n106 D_FlipFlop_0.D.n105 0.55213
R33312 D_FlipFlop_0.D.n112 D_FlipFlop_0.D.n111 0.55213
R33313 D_FlipFlop_0.D.n9 D_FlipFlop_0.D.n8 0.55213
R33314 D_FlipFlop_0.D.n15 D_FlipFlop_0.D.n14 0.55213
R33315 D_FlipFlop_0.D.n22 D_FlipFlop_0.D.n21 0.55213
R33316 D_FlipFlop_0.D.n28 D_FlipFlop_0.D.n27 0.55213
R33317 D_FlipFlop_0.D.n36 D_FlipFlop_0.D.n35 0.55213
R33318 D_FlipFlop_0.D.n42 D_FlipFlop_0.D.n41 0.55213
R33319 D_FlipFlop_0.D.n50 D_FlipFlop_0.D.n49 0.55213
R33320 D_FlipFlop_0.D.n56 D_FlipFlop_0.D.n55 0.55213
R33321 D_FlipFlop_0.D.n64 D_FlipFlop_0.D.n63 0.55213
R33322 D_FlipFlop_0.D.n70 D_FlipFlop_0.D.n69 0.55213
R33323 D_FlipFlop_0.D.n91 D_FlipFlop_0.D.n90 0.55213
R33324 D_FlipFlop_0.D.n97 D_FlipFlop_0.D.n96 0.55213
R33325 D_FlipFlop_0.D.n78 D_FlipFlop_0.D.n77 0.55213
R33326 D_FlipFlop_0.D.n84 D_FlipFlop_0.D.n83 0.55213
R33327 D_FlipFlop_0.D.n73 D_FlipFlop_0.D.n59 0.515159
R33328 D_FlipFlop_0.D.n106 D_FlipFlop_5.Inverter_0.Vin 0.486828
R33329 D_FlipFlop_0.D.n112 D_FlipFlop_5.3-input-nand_0.B 0.486828
R33330 D_FlipFlop_0.D.n9 D_FlipFlop_0.Inverter_0.Vin 0.486828
R33331 D_FlipFlop_0.D.n15 D_FlipFlop_0.3-input-nand_0.B 0.486828
R33332 D_FlipFlop_0.D.n22 D_FlipFlop_3.Inverter_0.Vin 0.486828
R33333 D_FlipFlop_0.D.n28 D_FlipFlop_3.3-input-nand_0.B 0.486828
R33334 D_FlipFlop_0.D.n36 D_FlipFlop_2.Inverter_0.Vin 0.486828
R33335 D_FlipFlop_0.D.n42 D_FlipFlop_2.3-input-nand_0.B 0.486828
R33336 D_FlipFlop_0.D.n50 D_FlipFlop_1.Inverter_0.Vin 0.486828
R33337 D_FlipFlop_0.D.n56 D_FlipFlop_1.3-input-nand_0.B 0.486828
R33338 D_FlipFlop_0.D.n64 D_FlipFlop_4.Inverter_0.Vin 0.486828
R33339 D_FlipFlop_0.D.n70 D_FlipFlop_4.3-input-nand_0.B 0.486828
R33340 D_FlipFlop_0.D.n91 D_FlipFlop_6.Inverter_0.Vin 0.486828
R33341 D_FlipFlop_0.D.n97 D_FlipFlop_6.3-input-nand_0.B 0.486828
R33342 D_FlipFlop_0.D.n78 D_FlipFlop_7.Inverter_0.Vin 0.486828
R33343 D_FlipFlop_0.D.n84 D_FlipFlop_7.3-input-nand_0.B 0.486828
R33344 D_FlipFlop_0.D.n103 D_FlipFlop_0.D.n102 0.470609
R33345 D_FlipFlop_0.D.n109 D_FlipFlop_0.D.n108 0.470609
R33346 D_FlipFlop_0.D.n6 D_FlipFlop_0.D.n5 0.470609
R33347 D_FlipFlop_0.D.n12 D_FlipFlop_0.D.n11 0.470609
R33348 D_FlipFlop_0.D.n19 D_FlipFlop_0.D.n18 0.470609
R33349 D_FlipFlop_0.D.n25 D_FlipFlop_0.D.n24 0.470609
R33350 D_FlipFlop_0.D.n33 D_FlipFlop_0.D.n32 0.470609
R33351 D_FlipFlop_0.D.n39 D_FlipFlop_0.D.n38 0.470609
R33352 D_FlipFlop_0.D.n47 D_FlipFlop_0.D.n46 0.470609
R33353 D_FlipFlop_0.D.n53 D_FlipFlop_0.D.n52 0.470609
R33354 D_FlipFlop_0.D.n61 D_FlipFlop_0.D.n60 0.470609
R33355 D_FlipFlop_0.D.n67 D_FlipFlop_0.D.n66 0.470609
R33356 D_FlipFlop_0.D.n88 D_FlipFlop_0.D.n87 0.470609
R33357 D_FlipFlop_0.D.n94 D_FlipFlop_0.D.n93 0.470609
R33358 D_FlipFlop_0.D.n75 D_FlipFlop_0.D.n74 0.470609
R33359 D_FlipFlop_0.D.n81 D_FlipFlop_0.D.n80 0.470609
R33360 D_FlipFlop_0.D.n115 D_FlipFlop_0.D.n101 0.3805
R33361 D_FlipFlop_0.D.n4 D_FlipFlop_0.D.n3 0.3805
R33362 D_FlipFlop_0.D.n45 D_FlipFlop_0.D.n31 0.323487
R33363 D_FlipFlop_0.D.n59 D_FlipFlop_0.D.n45 0.323487
R33364 D_FlipFlop_0.D.n101 D_FlipFlop_0.D.n73 0.323487
R33365 D_FlipFlop_0.D.n101 D_FlipFlop_0.D.n100 0.323487
R33366 D_FlipFlop_0.D.n116 D_FlipFlop_0.D.n4 0.280803
R33367 D_FlipFlop_0.D.n102 D_FlipFlop_5.Inverter_0.Vin 0.217464
R33368 D_FlipFlop_0.D.n108 D_FlipFlop_5.3-input-nand_0.B 0.217464
R33369 D_FlipFlop_0.D.n5 D_FlipFlop_0.Inverter_0.Vin 0.217464
R33370 D_FlipFlop_0.D.n11 D_FlipFlop_0.3-input-nand_0.B 0.217464
R33371 D_FlipFlop_0.D.n18 D_FlipFlop_3.Inverter_0.Vin 0.217464
R33372 D_FlipFlop_0.D.n24 D_FlipFlop_3.3-input-nand_0.B 0.217464
R33373 D_FlipFlop_0.D.n32 D_FlipFlop_2.Inverter_0.Vin 0.217464
R33374 D_FlipFlop_0.D.n38 D_FlipFlop_2.3-input-nand_0.B 0.217464
R33375 D_FlipFlop_0.D.n46 D_FlipFlop_1.Inverter_0.Vin 0.217464
R33376 D_FlipFlop_0.D.n52 D_FlipFlop_1.3-input-nand_0.B 0.217464
R33377 D_FlipFlop_0.D.n60 D_FlipFlop_4.Inverter_0.Vin 0.217464
R33378 D_FlipFlop_0.D.n66 D_FlipFlop_4.3-input-nand_0.B 0.217464
R33379 D_FlipFlop_0.D.n87 D_FlipFlop_6.Inverter_0.Vin 0.217464
R33380 D_FlipFlop_0.D.n93 D_FlipFlop_6.3-input-nand_0.B 0.217464
R33381 D_FlipFlop_0.D.n74 D_FlipFlop_7.Inverter_0.Vin 0.217464
R33382 D_FlipFlop_0.D.n80 D_FlipFlop_7.3-input-nand_0.B 0.217464
R33383 D_FlipFlop_0.D.n105 D_FlipFlop_5.Inverter_0.Vin 0.1255
R33384 D_FlipFlop_0.D.n111 D_FlipFlop_5.3-input-nand_0.B 0.1255
R33385 D_FlipFlop_0.D.n8 D_FlipFlop_0.Inverter_0.Vin 0.1255
R33386 D_FlipFlop_0.D.n14 D_FlipFlop_0.3-input-nand_0.B 0.1255
R33387 D_FlipFlop_0.D.n21 D_FlipFlop_3.Inverter_0.Vin 0.1255
R33388 D_FlipFlop_0.D.n27 D_FlipFlop_3.3-input-nand_0.B 0.1255
R33389 D_FlipFlop_0.D.n35 D_FlipFlop_2.Inverter_0.Vin 0.1255
R33390 D_FlipFlop_0.D.n41 D_FlipFlop_2.3-input-nand_0.B 0.1255
R33391 D_FlipFlop_0.D.n49 D_FlipFlop_1.Inverter_0.Vin 0.1255
R33392 D_FlipFlop_0.D.n55 D_FlipFlop_1.3-input-nand_0.B 0.1255
R33393 D_FlipFlop_0.D.n63 D_FlipFlop_4.Inverter_0.Vin 0.1255
R33394 D_FlipFlop_0.D.n69 D_FlipFlop_4.3-input-nand_0.B 0.1255
R33395 D_FlipFlop_0.D.n90 D_FlipFlop_6.Inverter_0.Vin 0.1255
R33396 D_FlipFlop_0.D.n96 D_FlipFlop_6.3-input-nand_0.B 0.1255
R33397 D_FlipFlop_0.D.n77 D_FlipFlop_7.Inverter_0.Vin 0.1255
R33398 D_FlipFlop_0.D.n83 D_FlipFlop_7.3-input-nand_0.B 0.1255
R33399 D_FlipFlop_0.D.n117 D_FlipFlop_0.D.n116 0.105716
R33400 D_FlipFlop_0.D.n3 D_FlipFlop_0.D.t0 0.0856875
R33401 D_FlipFlop_0.D.n107 D_FlipFlop_0.D.n103 0.063
R33402 D_FlipFlop_0.D.n107 D_FlipFlop_0.D.n106 0.063
R33403 D_FlipFlop_0.D.n113 D_FlipFlop_0.D.n109 0.063
R33404 D_FlipFlop_0.D.n113 D_FlipFlop_0.D.n112 0.063
R33405 D_FlipFlop_0.D.n10 D_FlipFlop_0.D.n6 0.063
R33406 D_FlipFlop_0.D.n10 D_FlipFlop_0.D.n9 0.063
R33407 D_FlipFlop_0.D.n16 D_FlipFlop_0.D.n12 0.063
R33408 D_FlipFlop_0.D.n16 D_FlipFlop_0.D.n15 0.063
R33409 D_FlipFlop_0.D.n23 D_FlipFlop_0.D.n19 0.063
R33410 D_FlipFlop_0.D.n23 D_FlipFlop_0.D.n22 0.063
R33411 D_FlipFlop_0.D.n29 D_FlipFlop_0.D.n25 0.063
R33412 D_FlipFlop_0.D.n29 D_FlipFlop_0.D.n28 0.063
R33413 D_FlipFlop_0.D.n37 D_FlipFlop_0.D.n33 0.063
R33414 D_FlipFlop_0.D.n37 D_FlipFlop_0.D.n36 0.063
R33415 D_FlipFlop_0.D.n43 D_FlipFlop_0.D.n39 0.063
R33416 D_FlipFlop_0.D.n43 D_FlipFlop_0.D.n42 0.063
R33417 D_FlipFlop_0.D.n51 D_FlipFlop_0.D.n47 0.063
R33418 D_FlipFlop_0.D.n51 D_FlipFlop_0.D.n50 0.063
R33419 D_FlipFlop_0.D.n57 D_FlipFlop_0.D.n53 0.063
R33420 D_FlipFlop_0.D.n57 D_FlipFlop_0.D.n56 0.063
R33421 D_FlipFlop_0.D.n65 D_FlipFlop_0.D.n61 0.063
R33422 D_FlipFlop_0.D.n65 D_FlipFlop_0.D.n64 0.063
R33423 D_FlipFlop_0.D.n71 D_FlipFlop_0.D.n67 0.063
R33424 D_FlipFlop_0.D.n71 D_FlipFlop_0.D.n70 0.063
R33425 D_FlipFlop_0.D.n92 D_FlipFlop_0.D.n88 0.063
R33426 D_FlipFlop_0.D.n92 D_FlipFlop_0.D.n91 0.063
R33427 D_FlipFlop_0.D.n98 D_FlipFlop_0.D.n94 0.063
R33428 D_FlipFlop_0.D.n98 D_FlipFlop_0.D.n97 0.063
R33429 D_FlipFlop_0.D.n79 D_FlipFlop_0.D.n75 0.063
R33430 D_FlipFlop_0.D.n79 D_FlipFlop_0.D.n78 0.063
R33431 D_FlipFlop_0.D.n85 D_FlipFlop_0.D.n81 0.063
R33432 D_FlipFlop_0.D.n85 D_FlipFlop_0.D.n84 0.063
R33433 Comparator_0.Vout D_FlipFlop_0.D.n117 0.0620344
R33434 D_FlipFlop_0.D.n117 D_FlipFlop_0.D.n0 0.0413995
R33435 D_FlipFlop_0.D.n105 D_FlipFlop_0.D.n104 0.0216397
R33436 D_FlipFlop_0.D.n104 D_FlipFlop_5.Inverter_0.Vin 0.0216397
R33437 D_FlipFlop_0.D.n111 D_FlipFlop_0.D.n110 0.0216397
R33438 D_FlipFlop_0.D.n110 D_FlipFlop_5.3-input-nand_0.B 0.0216397
R33439 D_FlipFlop_0.D.n8 D_FlipFlop_0.D.n7 0.0216397
R33440 D_FlipFlop_0.D.n7 D_FlipFlop_0.Inverter_0.Vin 0.0216397
R33441 D_FlipFlop_0.D.n14 D_FlipFlop_0.D.n13 0.0216397
R33442 D_FlipFlop_0.D.n13 D_FlipFlop_0.3-input-nand_0.B 0.0216397
R33443 D_FlipFlop_0.D.n21 D_FlipFlop_0.D.n20 0.0216397
R33444 D_FlipFlop_0.D.n20 D_FlipFlop_3.Inverter_0.Vin 0.0216397
R33445 D_FlipFlop_0.D.n27 D_FlipFlop_0.D.n26 0.0216397
R33446 D_FlipFlop_0.D.n26 D_FlipFlop_3.3-input-nand_0.B 0.0216397
R33447 D_FlipFlop_0.D.n35 D_FlipFlop_0.D.n34 0.0216397
R33448 D_FlipFlop_0.D.n34 D_FlipFlop_2.Inverter_0.Vin 0.0216397
R33449 D_FlipFlop_0.D.n41 D_FlipFlop_0.D.n40 0.0216397
R33450 D_FlipFlop_0.D.n40 D_FlipFlop_2.3-input-nand_0.B 0.0216397
R33451 D_FlipFlop_0.D.n49 D_FlipFlop_0.D.n48 0.0216397
R33452 D_FlipFlop_0.D.n48 D_FlipFlop_1.Inverter_0.Vin 0.0216397
R33453 D_FlipFlop_0.D.n55 D_FlipFlop_0.D.n54 0.0216397
R33454 D_FlipFlop_0.D.n54 D_FlipFlop_1.3-input-nand_0.B 0.0216397
R33455 D_FlipFlop_0.D.n63 D_FlipFlop_0.D.n62 0.0216397
R33456 D_FlipFlop_0.D.n62 D_FlipFlop_4.Inverter_0.Vin 0.0216397
R33457 D_FlipFlop_0.D.n69 D_FlipFlop_0.D.n68 0.0216397
R33458 D_FlipFlop_0.D.n68 D_FlipFlop_4.3-input-nand_0.B 0.0216397
R33459 D_FlipFlop_0.D.n90 D_FlipFlop_0.D.n89 0.0216397
R33460 D_FlipFlop_0.D.n89 D_FlipFlop_6.Inverter_0.Vin 0.0216397
R33461 D_FlipFlop_0.D.n96 D_FlipFlop_0.D.n95 0.0216397
R33462 D_FlipFlop_0.D.n95 D_FlipFlop_6.3-input-nand_0.B 0.0216397
R33463 D_FlipFlop_0.D.n77 D_FlipFlop_0.D.n76 0.0216397
R33464 D_FlipFlop_0.D.n76 D_FlipFlop_7.Inverter_0.Vin 0.0216397
R33465 D_FlipFlop_0.D.n83 D_FlipFlop_0.D.n82 0.0216397
R33466 D_FlipFlop_0.D.n82 D_FlipFlop_7.3-input-nand_0.B 0.0216397
R33467 D_FlipFlop_0.D.n0 Comparator_0.Vout 0.0131087
R33468 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 169.46
R33469 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 168.089
R33470 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 167.809
R33471 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 150.273
R33472 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 73.6406
R33473 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 60.3809
R33474 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 12.0358
R33475 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 11.4489
R33476 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 1.08746
R33477 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.851043
R33478 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.848156
R33479 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 0.788543
R33480 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 0.682565
R33481 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.65675
R33482 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 0.55213
R33483 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.486828
R33484 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 0.470609
R33485 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 0.262643
R33486 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.217464
R33487 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.1255
R33488 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.1255
R33489 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 0.063
R33490 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 0.063
R33491 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 0.063
R33492 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 0.063
R33493 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 0.063
R33494 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 0.0216397
R33495 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.0216397
R33496 Nand_Gate_0.A.n55 Nand_Gate_0.A.t0 169.46
R33497 Nand_Gate_0.A.n55 Nand_Gate_0.A.t1 167.809
R33498 Nand_Gate_0.A.n57 Nand_Gate_0.A.t3 167.809
R33499 Nand_Gate_0.A Nand_Gate_0.A.t13 158.585
R33500 Nand_Gate_0.A Nand_Gate_0.A.t16 158.581
R33501 Nand_Gate_0.A.n42 Nand_Gate_0.A.t11 150.293
R33502 Nand_Gate_0.A.t16 Nand_Gate_0.A.n38 150.293
R33503 Nand_Gate_0.A.t13 Nand_Gate_0.A.n2 150.293
R33504 Nand_Gate_0.A.n29 Nand_Gate_0.A.t10 150.273
R33505 Nand_Gate_0.A.n23 Nand_Gate_0.A.t17 150.273
R33506 Nand_Gate_0.A.n14 Nand_Gate_0.A.t12 150.273
R33507 Nand_Gate_0.A.n8 Nand_Gate_0.A.t8 150.273
R33508 Nand_Gate_0.A.n27 Nand_Gate_0.A.t6 73.6406
R33509 Nand_Gate_0.A.n21 Nand_Gate_0.A.t15 73.6406
R33510 Nand_Gate_0.A.n12 Nand_Gate_0.A.t7 73.6406
R33511 Nand_Gate_0.A.n6 Nand_Gate_0.A.t14 73.6406
R33512 Nand_Gate_0.A.n44 Nand_Gate_0.A.t4 73.6304
R33513 Nand_Gate_0.A.n36 Nand_Gate_0.A.t5 73.6304
R33514 Nand_Gate_0.A.n0 Nand_Gate_0.A.t9 73.6304
R33515 Nand_Gate_0.A.n48 Nand_Gate_0.A.n41 65.2862
R33516 Nand_Gate_0.A.n4 Nand_Gate_0.A.t2 60.3809
R33517 Nand_Gate_0.A.n33 Nand_Gate_0.A.n26 15.5222
R33518 Nand_Gate_0.A.n56 Nand_Gate_0.A.n55 11.4489
R33519 Nand_Gate_0.A.n48 Nand_Gate_0.A.n47 9.57083
R33520 Nand_Gate_0.A.n34 Nand_Gate_0.A.n33 8.26552
R33521 Nand_Gate_0.A.n58 Nand_Gate_0.A.n57 8.21389
R33522 Nand_Gate_0.A.n18 Nand_Gate_0.A.n11 8.1418
R33523 Nand_Gate_0.A.n49 Nand_Gate_0.A.n48 6.58222
R33524 Nand_Gate_0.A.n20 Nand_Gate_0.A.n19 6.47604
R33525 Nand_Gate_0.A.n19 Nand_Gate_0.A 5.35402
R33526 Nand_Gate_0.A.n52 Nand_Gate_0.A 4.55128
R33527 Nand_Gate_0.A.n33 Nand_Gate_0.A.n32 4.5005
R33528 Nand_Gate_0.A.n18 Nand_Gate_0.A.n17 4.5005
R33529 Nand_Gate_0.A.n38 Nand_Gate_0.A.n37 1.19615
R33530 Nand_Gate_0.A.n2 Nand_Gate_0.A.n1 1.19615
R33531 Nand_Gate_0.A.n5 Nand_Gate_0.A 1.08746
R33532 Nand_Gate_0.A.n20 Nand_Gate_0.A 0.973326
R33533 Nand_Gate_0.A.n13 Nand_Gate_0.A 0.851043
R33534 Nand_Gate_0.A.n7 Nand_Gate_0.A 0.851043
R33535 Nand_Gate_0.A.n4 Nand_Gate_0.A 0.848156
R33536 Nand_Gate_0.A.n28 Nand_Gate_0.A.n27 0.796696
R33537 Nand_Gate_0.A.n22 Nand_Gate_0.A.n21 0.796696
R33538 Nand_Gate_0.A.n54 Nand_Gate_0.A.n53 0.788543
R33539 Nand_Gate_0.A.n43 Nand_Gate_0.A 0.769522
R33540 Nand_Gate_0.A.n51 Nand_Gate_0.A.n50 0.755935
R33541 Nand_Gate_0.A.n34 Nand_Gate_0.A 0.716182
R33542 Nand_Gate_0.A.n5 Nand_Gate_0.A.n4 0.682565
R33543 Nand_Gate_0.A.n53 Nand_Gate_0.A 0.65675
R33544 Nand_Gate_0.A.n35 Nand_Gate_0.A.n34 0.556667
R33545 Nand_Gate_0.A.n43 Nand_Gate_0.A.n42 0.55213
R33546 Nand_Gate_0.A.n16 Nand_Gate_0.A.n15 0.55213
R33547 Nand_Gate_0.A.n10 Nand_Gate_0.A.n9 0.55213
R33548 Nand_Gate_0.A.n28 Nand_Gate_0.A 0.524957
R33549 Nand_Gate_0.A.n22 Nand_Gate_0.A 0.524957
R33550 Nand_Gate_0.A.n16 Nand_Gate_0.A 0.486828
R33551 Nand_Gate_0.A.n10 Nand_Gate_0.A 0.486828
R33552 Nand_Gate_0.A.n50 Nand_Gate_0.A 0.48023
R33553 Nand_Gate_0.A.n46 Nand_Gate_0.A.n45 0.470609
R33554 Nand_Gate_0.A.n13 Nand_Gate_0.A.n12 0.470609
R33555 Nand_Gate_0.A.n7 Nand_Gate_0.A.n6 0.470609
R33556 Nand_Gate_0.A.n42 Nand_Gate_0.A 0.447191
R33557 Nand_Gate_0.A.n38 Nand_Gate_0.A 0.447191
R33558 Nand_Gate_0.A.n2 Nand_Gate_0.A 0.447191
R33559 Nand_Gate_0.A.n46 Nand_Gate_0.A 0.428234
R33560 Nand_Gate_0.A.n58 Nand_Gate_0.A.n3 0.425067
R33561 Nand_Gate_0.A Nand_Gate_0.A.n58 0.39003
R33562 Nand_Gate_0.A.n57 Nand_Gate_0.A.n56 0.280391
R33563 Nand_Gate_0.A.n31 Nand_Gate_0.A 0.252453
R33564 Nand_Gate_0.A.n25 Nand_Gate_0.A 0.252453
R33565 Nand_Gate_0.A.n35 Nand_Gate_0.A 0.231583
R33566 Nand_Gate_0.A.n31 Nand_Gate_0.A.n30 0.226043
R33567 Nand_Gate_0.A.n25 Nand_Gate_0.A.n24 0.226043
R33568 Nand_Gate_0.A.n27 Nand_Gate_0.A 0.217464
R33569 Nand_Gate_0.A.n21 Nand_Gate_0.A 0.217464
R33570 Nand_Gate_0.A.n12 Nand_Gate_0.A 0.217464
R33571 Nand_Gate_0.A.n6 Nand_Gate_0.A 0.217464
R33572 Nand_Gate_0.A.n56 Nand_Gate_0.A 0.200143
R33573 Nand_Gate_0.A.n40 Nand_Gate_0.A.n39 0.168133
R33574 Nand_Gate_0.A.n40 Nand_Gate_0.A 0.135934
R33575 Nand_Gate_0.A.n45 Nand_Gate_0.A 0.1255
R33576 Nand_Gate_0.A.n30 Nand_Gate_0.A 0.1255
R33577 Nand_Gate_0.A.n24 Nand_Gate_0.A 0.1255
R33578 Nand_Gate_0.A.n37 Nand_Gate_0.A 0.1255
R33579 Nand_Gate_0.A.n15 Nand_Gate_0.A 0.1255
R33580 Nand_Gate_0.A.n9 Nand_Gate_0.A 0.1255
R33581 Nand_Gate_0.A.n54 Nand_Gate_0.A 0.1255
R33582 Nand_Gate_0.A.n1 Nand_Gate_0.A 0.1255
R33583 Nand_Gate_0.A.n47 Nand_Gate_0.A.n43 0.063
R33584 Nand_Gate_0.A.n47 Nand_Gate_0.A.n46 0.063
R33585 Nand_Gate_0.A.n32 Nand_Gate_0.A.n28 0.063
R33586 Nand_Gate_0.A.n32 Nand_Gate_0.A.n31 0.063
R33587 Nand_Gate_0.A.n26 Nand_Gate_0.A.n22 0.063
R33588 Nand_Gate_0.A.n26 Nand_Gate_0.A.n25 0.063
R33589 Nand_Gate_0.A.n17 Nand_Gate_0.A.n13 0.063
R33590 Nand_Gate_0.A.n17 Nand_Gate_0.A.n16 0.063
R33591 Nand_Gate_0.A.n11 Nand_Gate_0.A.n7 0.063
R33592 Nand_Gate_0.A.n11 Nand_Gate_0.A.n10 0.063
R33593 Nand_Gate_0.A.n19 Nand_Gate_0.A.n18 0.063
R33594 Nand_Gate_0.A.n49 Nand_Gate_0.A.n20 0.063
R33595 Nand_Gate_0.A.n50 Nand_Gate_0.A.n49 0.063
R33596 Nand_Gate_0.A.n52 Nand_Gate_0.A.n5 0.063
R33597 Nand_Gate_0.A.n53 Nand_Gate_0.A.n52 0.063
R33598 Nand_Gate_0.A Nand_Gate_0.A.n54 0.063
R33599 Nand_Gate_0.A.n41 Nand_Gate_0.A.n35 0.024
R33600 Nand_Gate_0.A.n41 Nand_Gate_0.A.n40 0.024
R33601 Nand_Gate_0.A.n30 Nand_Gate_0.A.n29 0.0216397
R33602 Nand_Gate_0.A.n29 Nand_Gate_0.A 0.0216397
R33603 Nand_Gate_0.A.n24 Nand_Gate_0.A.n23 0.0216397
R33604 Nand_Gate_0.A.n23 Nand_Gate_0.A 0.0216397
R33605 Nand_Gate_0.A.n15 Nand_Gate_0.A.n14 0.0216397
R33606 Nand_Gate_0.A.n14 Nand_Gate_0.A 0.0216397
R33607 Nand_Gate_0.A.n9 Nand_Gate_0.A.n8 0.0216397
R33608 Nand_Gate_0.A.n8 Nand_Gate_0.A 0.0216397
R33609 Nand_Gate_0.A.n51 Nand_Gate_0.A 0.0168043
R33610 Nand_Gate_0.A Nand_Gate_0.A.n51 0.0122188
R33611 Nand_Gate_0.A.n45 Nand_Gate_0.A.n44 0.0107679
R33612 Nand_Gate_0.A.n44 Nand_Gate_0.A 0.0107679
R33613 Nand_Gate_0.A.n37 Nand_Gate_0.A.n36 0.0107679
R33614 Nand_Gate_0.A.n36 Nand_Gate_0.A 0.0107679
R33615 Nand_Gate_0.A.n1 Nand_Gate_0.A.n0 0.0107679
R33616 Nand_Gate_0.A.n0 Nand_Gate_0.A 0.0107679
R33617 Nand_Gate_0.A.n39 Nand_Gate_0.A 0.00441667
R33618 Nand_Gate_0.A.n3 Nand_Gate_0.A 0.00441667
R33619 Nand_Gate_0.A.n39 Nand_Gate_0.A 0.00406061
R33620 Nand_Gate_0.A.n3 Nand_Gate_0.A 0.00406061
R33621 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 316.762
R33622 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 168.108
R33623 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 150.293
R33624 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 150.273
R33625 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 73.6406
R33626 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 73.6304
R33627 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 60.3943
R33628 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 12.0358
R33629 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 1.19615
R33630 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.981478
R33631 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 0.788543
R33632 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.769522
R33633 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 0.682565
R33634 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.580578
R33635 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 0.55213
R33636 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 0.484875
R33637 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 0.470609
R33638 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.447191
R33639 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.428234
R33640 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.217464
R33641 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R33642 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R33643 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.1255
R33644 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 0.063
R33645 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 0.063
R33646 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.063
R33647 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 0.063
R33648 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 0.063
R33649 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 0.0216397
R33650 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.0216397
R33651 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 0.0107679
R33652 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.0107679
R33653 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 179.256
R33654 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 168.089
R33655 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 150.293
R33656 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 73.6304
R33657 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 60.3943
R33658 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 12.0358
R33659 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.981478
R33660 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 0.788543
R33661 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.769522
R33662 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.720633
R33663 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 0.682565
R33664 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.580578
R33665 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 0.55213
R33666 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 0.470609
R33667 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.447191
R33668 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.428234
R33669 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1255
R33670 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1255
R33671 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 0.063
R33672 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 0.063
R33673 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 0.063
R33674 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 0.063
R33675 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 0.063
R33676 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 0.0435206
R33677 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 0.0107679
R33678 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.0107679
R33679 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 169.46
R33680 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 168.089
R33681 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 167.809
R33682 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 150.293
R33683 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 73.6304
R33684 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 60.3943
R33685 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 12.0358
R33686 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 11.4489
R33687 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.981478
R33688 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 0.788543
R33689 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.769522
R33690 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 0.720633
R33691 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 0.682565
R33692 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.580578
R33693 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 0.55213
R33694 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 0.470609
R33695 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.447191
R33696 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.428234
R33697 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.1255
R33698 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.1255
R33699 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 0.063
R33700 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 0.063
R33701 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.063
R33702 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 0.063
R33703 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 0.063
R33704 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 0.0435206
R33705 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 0.0107679
R33706 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.0107679
R33707 Nand_Gate_2.A.n55 Nand_Gate_2.A.t0 169.46
R33708 Nand_Gate_2.A.n55 Nand_Gate_2.A.t3 167.809
R33709 Nand_Gate_2.A.n57 Nand_Gate_2.A.t1 167.809
R33710 Nand_Gate_2.A Nand_Gate_2.A.t11 158.585
R33711 Nand_Gate_2.A Nand_Gate_2.A.t7 158.581
R33712 Nand_Gate_2.A.n42 Nand_Gate_2.A.t14 150.293
R33713 Nand_Gate_2.A.t7 Nand_Gate_2.A.n38 150.293
R33714 Nand_Gate_2.A.t11 Nand_Gate_2.A.n2 150.293
R33715 Nand_Gate_2.A.n29 Nand_Gate_2.A.t5 150.273
R33716 Nand_Gate_2.A.n23 Nand_Gate_2.A.t9 150.273
R33717 Nand_Gate_2.A.n14 Nand_Gate_2.A.t15 150.273
R33718 Nand_Gate_2.A.n8 Nand_Gate_2.A.t17 150.273
R33719 Nand_Gate_2.A.n27 Nand_Gate_2.A.t10 73.6406
R33720 Nand_Gate_2.A.n21 Nand_Gate_2.A.t6 73.6406
R33721 Nand_Gate_2.A.n12 Nand_Gate_2.A.t4 73.6406
R33722 Nand_Gate_2.A.n6 Nand_Gate_2.A.t16 73.6406
R33723 Nand_Gate_2.A.n44 Nand_Gate_2.A.t12 73.6304
R33724 Nand_Gate_2.A.n36 Nand_Gate_2.A.t13 73.6304
R33725 Nand_Gate_2.A.n0 Nand_Gate_2.A.t8 73.6304
R33726 Nand_Gate_2.A.n4 Nand_Gate_2.A.t2 60.3809
R33727 Nand_Gate_2.A.n48 Nand_Gate_2.A.n41 45.1913
R33728 Nand_Gate_2.A.n33 Nand_Gate_2.A.n26 15.5222
R33729 Nand_Gate_2.A.n56 Nand_Gate_2.A.n55 11.4489
R33730 Nand_Gate_2.A.n48 Nand_Gate_2.A.n47 9.57083
R33731 Nand_Gate_2.A.n34 Nand_Gate_2.A.n33 8.26552
R33732 Nand_Gate_2.A.n58 Nand_Gate_2.A.n57 8.21389
R33733 Nand_Gate_2.A.n18 Nand_Gate_2.A.n11 8.1418
R33734 Nand_Gate_2.A.n49 Nand_Gate_2.A.n48 6.58222
R33735 Nand_Gate_2.A.n20 Nand_Gate_2.A.n19 6.47604
R33736 Nand_Gate_2.A.n19 Nand_Gate_2.A 5.35402
R33737 Nand_Gate_2.A.n52 Nand_Gate_2.A 4.55128
R33738 Nand_Gate_2.A.n33 Nand_Gate_2.A.n32 4.5005
R33739 Nand_Gate_2.A.n18 Nand_Gate_2.A.n17 4.5005
R33740 Nand_Gate_2.A.n38 Nand_Gate_2.A.n37 1.19615
R33741 Nand_Gate_2.A.n2 Nand_Gate_2.A.n1 1.19615
R33742 Nand_Gate_2.A.n5 Nand_Gate_2.A 1.08746
R33743 Nand_Gate_2.A.n20 Nand_Gate_2.A 0.973326
R33744 Nand_Gate_2.A.n13 Nand_Gate_2.A 0.851043
R33745 Nand_Gate_2.A.n7 Nand_Gate_2.A 0.851043
R33746 Nand_Gate_2.A.n4 Nand_Gate_2.A 0.848156
R33747 Nand_Gate_2.A.n28 Nand_Gate_2.A.n27 0.796696
R33748 Nand_Gate_2.A.n22 Nand_Gate_2.A.n21 0.796696
R33749 Nand_Gate_2.A.n54 Nand_Gate_2.A.n53 0.788543
R33750 Nand_Gate_2.A.n43 Nand_Gate_2.A 0.769522
R33751 Nand_Gate_2.A.n51 Nand_Gate_2.A.n50 0.755935
R33752 Nand_Gate_2.A.n34 Nand_Gate_2.A 0.716182
R33753 Nand_Gate_2.A.n5 Nand_Gate_2.A.n4 0.682565
R33754 Nand_Gate_2.A.n53 Nand_Gate_2.A 0.65675
R33755 Nand_Gate_2.A.n43 Nand_Gate_2.A.n42 0.55213
R33756 Nand_Gate_2.A.n16 Nand_Gate_2.A.n15 0.55213
R33757 Nand_Gate_2.A.n10 Nand_Gate_2.A.n9 0.55213
R33758 Nand_Gate_2.A.n35 Nand_Gate_2.A.n34 0.549617
R33759 Nand_Gate_2.A.n28 Nand_Gate_2.A 0.524957
R33760 Nand_Gate_2.A.n22 Nand_Gate_2.A 0.524957
R33761 Nand_Gate_2.A.n16 Nand_Gate_2.A 0.486828
R33762 Nand_Gate_2.A.n10 Nand_Gate_2.A 0.486828
R33763 Nand_Gate_2.A.n50 Nand_Gate_2.A 0.48023
R33764 Nand_Gate_2.A.n46 Nand_Gate_2.A.n45 0.470609
R33765 Nand_Gate_2.A.n13 Nand_Gate_2.A.n12 0.470609
R33766 Nand_Gate_2.A.n7 Nand_Gate_2.A.n6 0.470609
R33767 Nand_Gate_2.A.n42 Nand_Gate_2.A 0.447191
R33768 Nand_Gate_2.A.n38 Nand_Gate_2.A 0.447191
R33769 Nand_Gate_2.A.n2 Nand_Gate_2.A 0.447191
R33770 Nand_Gate_2.A.n46 Nand_Gate_2.A 0.428234
R33771 Nand_Gate_2.A.n58 Nand_Gate_2.A.n3 0.425067
R33772 Nand_Gate_2.A Nand_Gate_2.A.n58 0.39003
R33773 Nand_Gate_2.A.n57 Nand_Gate_2.A.n56 0.280391
R33774 Nand_Gate_2.A.n31 Nand_Gate_2.A 0.252453
R33775 Nand_Gate_2.A.n25 Nand_Gate_2.A 0.252453
R33776 Nand_Gate_2.A.n35 Nand_Gate_2.A 0.238633
R33777 Nand_Gate_2.A.n31 Nand_Gate_2.A.n30 0.226043
R33778 Nand_Gate_2.A.n25 Nand_Gate_2.A.n24 0.226043
R33779 Nand_Gate_2.A.n27 Nand_Gate_2.A 0.217464
R33780 Nand_Gate_2.A.n21 Nand_Gate_2.A 0.217464
R33781 Nand_Gate_2.A.n12 Nand_Gate_2.A 0.217464
R33782 Nand_Gate_2.A.n6 Nand_Gate_2.A 0.217464
R33783 Nand_Gate_2.A.n56 Nand_Gate_2.A 0.200143
R33784 Nand_Gate_2.A.n40 Nand_Gate_2.A.n39 0.175183
R33785 Nand_Gate_2.A.n40 Nand_Gate_2.A 0.1415
R33786 Nand_Gate_2.A.n45 Nand_Gate_2.A 0.1255
R33787 Nand_Gate_2.A.n30 Nand_Gate_2.A 0.1255
R33788 Nand_Gate_2.A.n24 Nand_Gate_2.A 0.1255
R33789 Nand_Gate_2.A.n37 Nand_Gate_2.A 0.1255
R33790 Nand_Gate_2.A.n15 Nand_Gate_2.A 0.1255
R33791 Nand_Gate_2.A.n9 Nand_Gate_2.A 0.1255
R33792 Nand_Gate_2.A.n54 Nand_Gate_2.A 0.1255
R33793 Nand_Gate_2.A.n1 Nand_Gate_2.A 0.1255
R33794 Nand_Gate_2.A.n47 Nand_Gate_2.A.n43 0.063
R33795 Nand_Gate_2.A.n47 Nand_Gate_2.A.n46 0.063
R33796 Nand_Gate_2.A.n32 Nand_Gate_2.A.n28 0.063
R33797 Nand_Gate_2.A.n32 Nand_Gate_2.A.n31 0.063
R33798 Nand_Gate_2.A.n26 Nand_Gate_2.A.n22 0.063
R33799 Nand_Gate_2.A.n26 Nand_Gate_2.A.n25 0.063
R33800 Nand_Gate_2.A.n17 Nand_Gate_2.A.n13 0.063
R33801 Nand_Gate_2.A.n17 Nand_Gate_2.A.n16 0.063
R33802 Nand_Gate_2.A.n11 Nand_Gate_2.A.n7 0.063
R33803 Nand_Gate_2.A.n11 Nand_Gate_2.A.n10 0.063
R33804 Nand_Gate_2.A.n19 Nand_Gate_2.A.n18 0.063
R33805 Nand_Gate_2.A.n49 Nand_Gate_2.A.n20 0.063
R33806 Nand_Gate_2.A.n50 Nand_Gate_2.A.n49 0.063
R33807 Nand_Gate_2.A.n52 Nand_Gate_2.A.n5 0.063
R33808 Nand_Gate_2.A.n53 Nand_Gate_2.A.n52 0.063
R33809 Nand_Gate_2.A Nand_Gate_2.A.n54 0.063
R33810 Nand_Gate_2.A.n41 Nand_Gate_2.A.n35 0.024
R33811 Nand_Gate_2.A.n41 Nand_Gate_2.A.n40 0.024
R33812 Nand_Gate_2.A.n30 Nand_Gate_2.A.n29 0.0216397
R33813 Nand_Gate_2.A.n29 Nand_Gate_2.A 0.0216397
R33814 Nand_Gate_2.A.n24 Nand_Gate_2.A.n23 0.0216397
R33815 Nand_Gate_2.A.n23 Nand_Gate_2.A 0.0216397
R33816 Nand_Gate_2.A.n15 Nand_Gate_2.A.n14 0.0216397
R33817 Nand_Gate_2.A.n14 Nand_Gate_2.A 0.0216397
R33818 Nand_Gate_2.A.n9 Nand_Gate_2.A.n8 0.0216397
R33819 Nand_Gate_2.A.n8 Nand_Gate_2.A 0.0216397
R33820 Nand_Gate_2.A.n51 Nand_Gate_2.A 0.0168043
R33821 Nand_Gate_2.A Nand_Gate_2.A.n51 0.0122188
R33822 Nand_Gate_2.A.n45 Nand_Gate_2.A.n44 0.0107679
R33823 Nand_Gate_2.A.n44 Nand_Gate_2.A 0.0107679
R33824 Nand_Gate_2.A.n37 Nand_Gate_2.A.n36 0.0107679
R33825 Nand_Gate_2.A.n36 Nand_Gate_2.A 0.0107679
R33826 Nand_Gate_2.A.n1 Nand_Gate_2.A.n0 0.0107679
R33827 Nand_Gate_2.A.n0 Nand_Gate_2.A 0.0107679
R33828 Nand_Gate_2.A.n39 Nand_Gate_2.A 0.00441667
R33829 Nand_Gate_2.A.n3 Nand_Gate_2.A 0.00441667
R33830 Nand_Gate_2.A.n39 Nand_Gate_2.A 0.00406061
R33831 Nand_Gate_2.A.n3 Nand_Gate_2.A 0.00406061
R33832 And_Gate_1.Vout.n13 And_Gate_1.Vout.t0 168.32
R33833 And_Gate_1.Vout.n4 And_Gate_1.Vout.t3 158.207
R33834 D_FlipFlop_7.CLK And_Gate_1.Vout.t5 158.202
R33835 And_Gate_1.Vout.n6 And_Gate_1.Vout.t4 150.293
R33836 And_Gate_1.Vout.t5 And_Gate_1.Vout.n9 150.293
R33837 And_Gate_1.Vout.t3 And_Gate_1.Vout.n3 150.273
R33838 And_Gate_1.Vout.n13 And_Gate_1.Vout.n12 81.2012
R33839 And_Gate_1.Vout.n1 And_Gate_1.Vout.t6 73.6406
R33840 And_Gate_1.Vout.n8 And_Gate_1.Vout.t2 73.6304
R33841 And_Gate_1.Vout.n7 And_Gate_1.Vout.t7 73.6304
R33842 And_Gate_1.Inverter_0.Vout And_Gate_1.Vout.t1 60.3943
R33843 And_Gate_1.Vout.n8 And_Gate_1.Vout.n7 16.332
R33844 And_Gate_1.Vout.n14 And_Gate_1.Vout.n0 1.62007
R33845 And_Gate_1.Inverter_0.Vout And_Gate_1.Vout.n14 1.25441
R33846 And_Gate_1.Vout.n2 And_Gate_1.Vout.n1 1.19615
R33847 And_Gate_1.Vout.n7 And_Gate_1.Vout.n6 1.1717
R33848 And_Gate_1.Vout.n9 And_Gate_1.Vout.n8 1.1717
R33849 And_Gate_1.Vout.n9 D_FlipFlop_7.3-input-nand_1.C 0.447191
R33850 And_Gate_1.Vout.n6 D_FlipFlop_7.Inverter_1.Vin 0.436162
R33851 And_Gate_1.Vout.n4 D_FlipFlop_7.CLK 0.321667
R33852 And_Gate_1.Vout.n5 D_FlipFlop_7.CLK 0.250383
R33853 And_Gate_1.Vout.n1 D_FlipFlop_7.3-input-nand_0.C 0.217464
R33854 And_Gate_1.Vout.n11 And_Gate_1.Vout.n10 0.186933
R33855 And_Gate_1.Vout.n11 D_FlipFlop_7.CLK 0.150776
R33856 And_Gate_1.Vout.n8 D_FlipFlop_7.3-input-nand_1.C 0.149957
R33857 And_Gate_1.Vout.n2 D_FlipFlop_7.3-input-nand_0.C 0.1255
R33858 And_Gate_1.Vout.n0 And_Gate_1.Inverter_0.Vout 0.1255
R33859 And_Gate_1.Vout.n7 D_FlipFlop_7.Inverter_1.Vin 0.117348
R33860 And_Gate_1.Vout.n5 And_Gate_1.Vout.n4 0.1039
R33861 And_Gate_1.Vout.n0 And_Gate_1.Inverter_0.Vout 0.063
R33862 And_Gate_1.Vout.n14 And_Gate_1.Vout.n13 0.063
R33863 And_Gate_1.Vout.n7 D_FlipFlop_7.Inverter_1.Vin 0.0454219
R33864 And_Gate_1.Vout.n8 D_FlipFlop_7.3-input-nand_1.C 0.0454219
R33865 And_Gate_1.Vout.n12 And_Gate_1.Vout.n5 0.024
R33866 And_Gate_1.Vout.n12 And_Gate_1.Vout.n11 0.024
R33867 And_Gate_1.Vout.n3 And_Gate_1.Vout.n2 0.0216397
R33868 And_Gate_1.Vout.n3 D_FlipFlop_7.3-input-nand_0.C 0.0216397
R33869 And_Gate_1.Vout.n10 D_FlipFlop_7.CLK 0.00441667
R33870 And_Gate_1.Vout.n10 D_FlipFlop_7.CLK 0.00406061
R33871 Nand_Gate_2.B.n31 Nand_Gate_2.B.t0 169.46
R33872 Nand_Gate_2.B.n31 Nand_Gate_2.B.t1 167.809
R33873 Nand_Gate_2.B.n33 Nand_Gate_2.B.t3 167.809
R33874 Nand_Gate_2.B Nand_Gate_2.B.t5 158.585
R33875 Nand_Gate_2.B.t5 Nand_Gate_2.B.n2 150.293
R33876 Nand_Gate_2.B.n24 Nand_Gate_2.B.t11 150.273
R33877 Nand_Gate_2.B.n14 Nand_Gate_2.B.t8 150.273
R33878 Nand_Gate_2.B.n8 Nand_Gate_2.B.t4 150.273
R33879 Nand_Gate_2.B.n12 Nand_Gate_2.B.t6 73.6406
R33880 Nand_Gate_2.B.n6 Nand_Gate_2.B.t7 73.6406
R33881 Nand_Gate_2.B.n21 Nand_Gate_2.B.t9 73.6304
R33882 Nand_Gate_2.B.n0 Nand_Gate_2.B.t10 73.6304
R33883 Nand_Gate_2.B.n4 Nand_Gate_2.B.t2 60.3809
R33884 Nand_Gate_2.B.n25 Nand_Gate_2.B.n24 40.8363
R33885 Nand_Gate_2.B.n32 Nand_Gate_2.B.n31 11.4489
R33886 Nand_Gate_2.B.n34 Nand_Gate_2.B.n33 8.21389
R33887 Nand_Gate_2.B.n18 Nand_Gate_2.B.n11 8.1418
R33888 Nand_Gate_2.B.n20 Nand_Gate_2.B.n19 6.47604
R33889 Nand_Gate_2.B.n19 Nand_Gate_2.B 5.35402
R33890 Nand_Gate_2.B.n28 Nand_Gate_2.B 4.55128
R33891 Nand_Gate_2.B.n18 Nand_Gate_2.B.n17 4.5005
R33892 Nand_Gate_2.B.n2 Nand_Gate_2.B.n1 1.19615
R33893 Nand_Gate_2.B.n23 Nand_Gate_2.B.n22 1.1717
R33894 Nand_Gate_2.B.n5 Nand_Gate_2.B 1.08746
R33895 Nand_Gate_2.B.n20 Nand_Gate_2.B 0.973326
R33896 Nand_Gate_2.B.n23 Nand_Gate_2.B 0.932141
R33897 Nand_Gate_2.B.n13 Nand_Gate_2.B 0.851043
R33898 Nand_Gate_2.B.n7 Nand_Gate_2.B 0.851043
R33899 Nand_Gate_2.B.n4 Nand_Gate_2.B 0.848156
R33900 Nand_Gate_2.B.n30 Nand_Gate_2.B.n29 0.788543
R33901 Nand_Gate_2.B.n27 Nand_Gate_2.B.n26 0.755935
R33902 Nand_Gate_2.B.n5 Nand_Gate_2.B.n4 0.682565
R33903 Nand_Gate_2.B.n29 Nand_Gate_2.B 0.65675
R33904 Nand_Gate_2.B.n16 Nand_Gate_2.B.n15 0.55213
R33905 Nand_Gate_2.B.n10 Nand_Gate_2.B.n9 0.55213
R33906 Nand_Gate_2.B.n16 Nand_Gate_2.B 0.486828
R33907 Nand_Gate_2.B.n10 Nand_Gate_2.B 0.486828
R33908 Nand_Gate_2.B.n26 Nand_Gate_2.B 0.48023
R33909 Nand_Gate_2.B.n13 Nand_Gate_2.B.n12 0.470609
R33910 Nand_Gate_2.B.n7 Nand_Gate_2.B.n6 0.470609
R33911 Nand_Gate_2.B.n2 Nand_Gate_2.B 0.447191
R33912 Nand_Gate_2.B.n34 Nand_Gate_2.B.n3 0.425067
R33913 Nand_Gate_2.B Nand_Gate_2.B.n34 0.39003
R33914 Nand_Gate_2.B.n33 Nand_Gate_2.B.n32 0.280391
R33915 Nand_Gate_2.B.n12 Nand_Gate_2.B 0.217464
R33916 Nand_Gate_2.B.n6 Nand_Gate_2.B 0.217464
R33917 Nand_Gate_2.B.n32 Nand_Gate_2.B 0.200143
R33918 Nand_Gate_2.B.n22 Nand_Gate_2.B 0.1255
R33919 Nand_Gate_2.B.n15 Nand_Gate_2.B 0.1255
R33920 Nand_Gate_2.B.n9 Nand_Gate_2.B 0.1255
R33921 Nand_Gate_2.B.n30 Nand_Gate_2.B 0.1255
R33922 Nand_Gate_2.B.n1 Nand_Gate_2.B 0.1255
R33923 Nand_Gate_2.B.n24 Nand_Gate_2.B.n23 0.063
R33924 Nand_Gate_2.B.n17 Nand_Gate_2.B.n13 0.063
R33925 Nand_Gate_2.B.n17 Nand_Gate_2.B.n16 0.063
R33926 Nand_Gate_2.B.n11 Nand_Gate_2.B.n7 0.063
R33927 Nand_Gate_2.B.n11 Nand_Gate_2.B.n10 0.063
R33928 Nand_Gate_2.B.n19 Nand_Gate_2.B.n18 0.063
R33929 Nand_Gate_2.B.n25 Nand_Gate_2.B.n20 0.063
R33930 Nand_Gate_2.B.n26 Nand_Gate_2.B.n25 0.063
R33931 Nand_Gate_2.B.n28 Nand_Gate_2.B.n5 0.063
R33932 Nand_Gate_2.B.n29 Nand_Gate_2.B.n28 0.063
R33933 Nand_Gate_2.B Nand_Gate_2.B.n30 0.063
R33934 Nand_Gate_2.B.n15 Nand_Gate_2.B.n14 0.0216397
R33935 Nand_Gate_2.B.n14 Nand_Gate_2.B 0.0216397
R33936 Nand_Gate_2.B.n9 Nand_Gate_2.B.n8 0.0216397
R33937 Nand_Gate_2.B.n8 Nand_Gate_2.B 0.0216397
R33938 Nand_Gate_2.B.n27 Nand_Gate_2.B 0.0168043
R33939 Nand_Gate_2.B Nand_Gate_2.B.n27 0.0122188
R33940 Nand_Gate_2.B.n22 Nand_Gate_2.B.n21 0.0107679
R33941 Nand_Gate_2.B.n21 Nand_Gate_2.B 0.0107679
R33942 Nand_Gate_2.B.n1 Nand_Gate_2.B.n0 0.0107679
R33943 Nand_Gate_2.B.n0 Nand_Gate_2.B 0.0107679
R33944 Nand_Gate_2.B.n3 Nand_Gate_2.B 0.00441667
R33945 Nand_Gate_2.B.n3 Nand_Gate_2.B 0.00406061
R33946 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 316.762
R33947 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 168.108
R33948 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 150.293
R33949 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 150.273
R33950 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 73.6406
R33951 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 73.6304
R33952 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 60.4568
R33953 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 12.0358
R33954 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 1.19615
R33955 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.981478
R33956 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 0.788543
R33957 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.769522
R33958 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 0.682565
R33959 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.580578
R33960 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 0.55213
R33961 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 0.484875
R33962 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 0.470609
R33963 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.447191
R33964 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.428234
R33965 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.217464
R33966 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R33967 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R33968 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.1255
R33969 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 0.063
R33970 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 0.063
R33971 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.063
R33972 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 0.063
R33973 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 0.063
R33974 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 0.0216397
R33975 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.0216397
R33976 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 0.0107679
R33977 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.0107679
R33978 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 179.256
R33979 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 168.089
R33980 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 150.293
R33981 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 73.6304
R33982 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 60.4568
R33983 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 12.0358
R33984 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.981478
R33985 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 0.788543
R33986 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.769522
R33987 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 0.720633
R33988 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 0.682565
R33989 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.580578
R33990 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 0.55213
R33991 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 0.470609
R33992 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.447191
R33993 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.428234
R33994 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1255
R33995 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1255
R33996 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 0.063
R33997 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 0.063
R33998 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.063
R33999 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 0.063
R34000 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 0.063
R34001 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 0.0435206
R34002 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 0.0107679
R34003 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.0107679
R34004 And_Gate_4.Vout.n14 And_Gate_4.Vout.t0 168.108
R34005 And_Gate_4.Vout.n5 And_Gate_4.Vout.t6 158.207
R34006 D_FlipFlop_2.CLK And_Gate_4.Vout.t2 158.202
R34007 And_Gate_4.Vout.n7 And_Gate_4.Vout.t7 150.293
R34008 And_Gate_4.Vout.t2 And_Gate_4.Vout.n10 150.293
R34009 And_Gate_4.Vout.t6 And_Gate_4.Vout.n4 150.273
R34010 And_Gate_4.Vout.n2 And_Gate_4.Vout.t5 73.6406
R34011 And_Gate_4.Vout.n9 And_Gate_4.Vout.t4 73.6304
R34012 And_Gate_4.Vout.n8 And_Gate_4.Vout.t3 73.6304
R34013 And_Gate_4.Vout.n12 And_Gate_4.Vout.n11 62.4488
R34014 And_Gate_4.Inverter_0.Vout And_Gate_4.Vout.t1 60.3943
R34015 And_Gate_4.Vout.n9 And_Gate_4.Vout.n8 16.332
R34016 And_Gate_4.Vout.n3 And_Gate_4.Vout.n2 1.19615
R34017 And_Gate_4.Vout.n8 And_Gate_4.Vout.n7 1.1717
R34018 And_Gate_4.Vout.n10 And_Gate_4.Vout.n9 1.1717
R34019 And_Gate_4.Vout.n13 And_Gate_4.Inverter_0.Vout 0.981478
R34020 And_Gate_4.Vout.n14 And_Gate_4.Vout.n13 0.788543
R34021 And_Gate_4.Vout.n1 And_Gate_4.Vout.n0 0.682565
R34022 And_Gate_4.Vout.n1 And_Gate_4.Inverter_0.Vout 0.580578
R34023 And_Gate_4.Inverter_0.Vout And_Gate_4.Vout.n14 0.484875
R34024 And_Gate_4.Vout.n10 D_FlipFlop_2.3-input-nand_1.C 0.447191
R34025 And_Gate_4.Vout.n7 D_FlipFlop_2.Inverter_1.Vin 0.436162
R34026 And_Gate_4.Vout.n5 D_FlipFlop_2.CLK 0.321667
R34027 And_Gate_4.Vout.n6 And_Gate_4.Vout.n5 0.295033
R34028 And_Gate_4.Vout.n2 D_FlipFlop_2.3-input-nand_0.C 0.217464
R34029 And_Gate_4.Vout.n9 D_FlipFlop_2.3-input-nand_1.C 0.149957
R34030 And_Gate_4.Vout.n3 D_FlipFlop_2.3-input-nand_0.C 0.1255
R34031 And_Gate_4.Vout.n0 And_Gate_4.Inverter_0.Vout 0.1255
R34032 And_Gate_4.Vout.n8 D_FlipFlop_2.Inverter_1.Vin 0.117348
R34033 And_Gate_4.Vout.n0 And_Gate_4.Inverter_0.Vout 0.063
R34034 And_Gate_4.Vout.n13 And_Gate_4.Vout.n12 0.063
R34035 And_Gate_4.Vout.n12 And_Gate_4.Vout.n1 0.063
R34036 And_Gate_4.Vout.n6 D_FlipFlop_2.CLK 0.05925
R34037 And_Gate_4.Vout.n8 D_FlipFlop_2.Inverter_1.Vin 0.0454219
R34038 And_Gate_4.Vout.n9 D_FlipFlop_2.3-input-nand_1.C 0.0454219
R34039 And_Gate_4.Vout.n11 And_Gate_4.Vout.n6 0.024
R34040 And_Gate_4.Vout.n11 D_FlipFlop_2.CLK 0.0233816
R34041 And_Gate_4.Vout.n4 And_Gate_4.Vout.n3 0.0216397
R34042 And_Gate_4.Vout.n4 D_FlipFlop_2.3-input-nand_0.C 0.0216397
R34043 And_Gate_7.Vout.n15 And_Gate_7.Vout.t0 168.108
R34044 And_Gate_7.Vout.n3 And_Gate_7.Vout.t6 158.207
R34045 D_FlipFlop_0.CLK And_Gate_7.Vout.t2 158.202
R34046 And_Gate_7.Vout.n5 And_Gate_7.Vout.t7 150.293
R34047 And_Gate_7.Vout.t2 And_Gate_7.Vout.n8 150.293
R34048 And_Gate_7.Vout.t6 And_Gate_7.Vout.n2 150.273
R34049 And_Gate_7.Vout.n0 And_Gate_7.Vout.t3 73.6406
R34050 And_Gate_7.Vout.n7 And_Gate_7.Vout.t5 73.6304
R34051 And_Gate_7.Vout.n6 And_Gate_7.Vout.t4 73.6304
R34052 And_Gate_7.Inverter_0.Vout And_Gate_7.Vout.t1 60.3072
R34053 And_Gate_7.Vout.n12 And_Gate_7.Vout.n11 21.9583
R34054 And_Gate_7.Vout.n7 And_Gate_7.Vout.n6 16.332
R34055 And_Gate_7.Vout.n15 And_Gate_7.Vout.n14 1.62007
R34056 And_Gate_7.Vout.n1 And_Gate_7.Vout.n0 1.19615
R34057 And_Gate_7.Vout.n6 And_Gate_7.Vout.n5 1.1717
R34058 And_Gate_7.Vout.n8 And_Gate_7.Vout.n7 1.1717
R34059 And_Gate_7.Inverter_0.Vout And_Gate_7.Vout.n15 0.484875
R34060 And_Gate_7.Vout.n8 D_FlipFlop_0.3-input-nand_1.C 0.447191
R34061 And_Gate_7.Vout.n5 D_FlipFlop_0.Inverter_1.Vin 0.436162
R34062 And_Gate_7.Vout.n3 D_FlipFlop_0.CLK 0.321667
R34063 And_Gate_7.Vout.n4 And_Gate_7.Vout.n3 0.219833
R34064 And_Gate_7.Vout.n0 D_FlipFlop_0.3-input-nand_0.C 0.217464
R34065 And_Gate_7.Vout.n7 D_FlipFlop_0.3-input-nand_1.C 0.149957
R34066 And_Gate_7.Vout.n14 And_Gate_7.Inverter_0.Vout 0.149957
R34067 And_Gate_7.Vout.n4 D_FlipFlop_0.CLK 0.13445
R34068 And_Gate_7.Vout.n1 D_FlipFlop_0.3-input-nand_0.C 0.1255
R34069 And_Gate_7.Vout.n6 D_FlipFlop_0.Inverter_1.Vin 0.117348
R34070 And_Gate_7.Vout.n13 And_Gate_7.Inverter_0.Vout 0.0903438
R34071 And_Gate_7.Vout.n10 And_Gate_7.Vout.n9 0.071
R34072 And_Gate_7.Vout.n10 D_FlipFlop_0.CLK 0.05925
R34073 And_Gate_7.Vout.n6 D_FlipFlop_0.Inverter_1.Vin 0.0454219
R34074 And_Gate_7.Vout.n7 D_FlipFlop_0.3-input-nand_1.C 0.0454219
R34075 And_Gate_7.Vout.n13 And_Gate_7.Vout.n12 0.027881
R34076 And_Gate_7.Vout.n12 And_Gate_7.Inverter_0.Vout 0.027881
R34077 And_Gate_7.Vout.n11 And_Gate_7.Vout.n4 0.024
R34078 And_Gate_7.Vout.n11 And_Gate_7.Vout.n10 0.024
R34079 And_Gate_7.Vout.n2 And_Gate_7.Vout.n1 0.0216397
R34080 And_Gate_7.Vout.n2 D_FlipFlop_0.3-input-nand_0.C 0.0216397
R34081 And_Gate_7.Vout.n14 And_Gate_7.Vout.n13 0.0180781
R34082 And_Gate_7.Vout.n9 D_FlipFlop_0.CLK 0.00441667
R34083 And_Gate_7.Vout.n9 D_FlipFlop_0.CLK 0.00406061
R34084 And_Gate_3.Vout.n12 And_Gate_3.Vout.t0 168.32
R34085 And_Gate_3.Vout.n4 And_Gate_3.Vout.t3 158.226
R34086 D_FlipFlop_4.CLK And_Gate_3.Vout.t6 158.202
R34087 And_Gate_3.Vout.n5 And_Gate_3.Vout.t4 150.293
R34088 And_Gate_3.Vout.t6 And_Gate_3.Vout.n8 150.293
R34089 And_Gate_3.Vout.t3 And_Gate_3.Vout.n3 150.273
R34090 And_Gate_3.Vout.n1 And_Gate_3.Vout.t5 73.6406
R34091 And_Gate_3.Vout.n7 And_Gate_3.Vout.t2 73.6304
R34092 And_Gate_3.Vout.n6 And_Gate_3.Vout.t7 73.6304
R34093 And_Gate_3.Inverter_0.Vout And_Gate_3.Vout.t1 60.3943
R34094 And_Gate_3.Vout.n12 And_Gate_3.Vout.n11 37.7699
R34095 And_Gate_3.Vout.n7 And_Gate_3.Vout.n6 16.332
R34096 And_Gate_3.Vout.n13 And_Gate_3.Vout.n0 1.62007
R34097 And_Gate_3.Inverter_0.Vout And_Gate_3.Vout.n13 1.25441
R34098 And_Gate_3.Vout.n2 And_Gate_3.Vout.n1 1.19615
R34099 And_Gate_3.Vout.n6 And_Gate_3.Vout.n5 1.1717
R34100 And_Gate_3.Vout.n8 And_Gate_3.Vout.n7 1.1717
R34101 And_Gate_3.Vout.n8 D_FlipFlop_4.3-input-nand_1.C 0.447191
R34102 And_Gate_3.Vout.n5 D_FlipFlop_4.Inverter_1.Vin 0.436162
R34103 And_Gate_3.Vout.n4 D_FlipFlop_4.CLK 0.302439
R34104 And_Gate_3.Vout.n10 And_Gate_3.Vout.n9 0.269183
R34105 And_Gate_3.Vout.n1 D_FlipFlop_4.3-input-nand_0.C 0.217464
R34106 And_Gate_3.Vout.n10 D_FlipFlop_4.CLK 0.215711
R34107 And_Gate_3.Vout.n7 D_FlipFlop_4.3-input-nand_1.C 0.149957
R34108 And_Gate_3.Vout.n2 D_FlipFlop_4.3-input-nand_0.C 0.1255
R34109 And_Gate_3.Vout.n0 And_Gate_3.Inverter_0.Vout 0.1255
R34110 And_Gate_3.Vout.n6 D_FlipFlop_4.Inverter_1.Vin 0.117348
R34111 And_Gate_3.Vout.n0 And_Gate_3.Inverter_0.Vout 0.063
R34112 And_Gate_3.Vout.n13 And_Gate_3.Vout.n12 0.063
R34113 And_Gate_3.Vout.n6 D_FlipFlop_4.Inverter_1.Vin 0.0454219
R34114 And_Gate_3.Vout.n7 D_FlipFlop_4.3-input-nand_1.C 0.0454219
R34115 And_Gate_3.Vout.n11 And_Gate_3.Vout.n4 0.024
R34116 And_Gate_3.Vout.n11 And_Gate_3.Vout.n10 0.024
R34117 And_Gate_3.Vout.n3 And_Gate_3.Vout.n2 0.0216397
R34118 And_Gate_3.Vout.n3 D_FlipFlop_4.3-input-nand_0.C 0.0216397
R34119 And_Gate_3.Vout.n9 D_FlipFlop_4.CLK 0.00441667
R34120 And_Gate_3.Vout.n9 D_FlipFlop_4.CLK 0.00406061
R34121 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 316.762
R34122 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 168.108
R34123 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 150.293
R34124 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 150.273
R34125 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 73.6406
R34126 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 73.6304
R34127 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 60.4568
R34128 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 12.0358
R34129 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 1.19615
R34130 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.981478
R34131 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 0.788543
R34132 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.769522
R34133 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 0.682565
R34134 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.580578
R34135 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 0.55213
R34136 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 0.484875
R34137 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 0.470609
R34138 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.447191
R34139 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.428234
R34140 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.217464
R34141 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R34142 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R34143 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.1255
R34144 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 0.063
R34145 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 0.063
R34146 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.063
R34147 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 0.063
R34148 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 0.063
R34149 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 0.0216397
R34150 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.0216397
R34151 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 0.0107679
R34152 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.0107679
R34153 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t0 169.46
R34154 D_FlipFlop_2.3-input-nand_2.C.n11 D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R34155 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.t3 167.809
R34156 D_FlipFlop_2.3-input-nand_2.C.t6 D_FlipFlop_2.3-input-nand_2.C.n13 167.226
R34157 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C.t4 150.273
R34158 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.t6 150.273
R34159 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C.t7 73.6406
R34160 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C.t5 73.6304
R34161 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C.t1 60.4568
R34162 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C.n7 12.3891
R34163 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.n11 11.4489
R34164 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C 1.68257
R34165 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C.n2 1.38365
R34166 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C.n0 1.19615
R34167 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C.n5 1.1717
R34168 D_FlipFlop_2.3-input-nand_2.C.n3 D_FlipFlop_2.3-input-nand_2.C 1.08448
R34169 D_FlipFlop_2.3-input-nand_2.C.n6 D_FlipFlop_2.3-input-nand_2.C 0.932141
R34170 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C 0.720633
R34171 D_FlipFlop_2.3-input-nand_2.C.n13 D_FlipFlop_2.3-input-nand_2.C.n12 0.280391
R34172 D_FlipFlop_2.3-input-nand_2.C.n0 D_FlipFlop_2.3-input-nand_2.C 0.217464
R34173 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C 0.1255
R34174 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C 0.1255
R34175 D_FlipFlop_2.3-input-nand_2.C.n1 D_FlipFlop_2.3-input-nand_2.C 0.1255
R34176 D_FlipFlop_2.3-input-nand_2.C.n10 D_FlipFlop_2.3-input-nand_2.C.n9 0.0874565
R34177 D_FlipFlop_2.3-input-nand_2.C.n7 D_FlipFlop_2.3-input-nand_2.C.n6 0.063
R34178 D_FlipFlop_2.3-input-nand_2.C.n2 D_FlipFlop_2.3-input-nand_2.C 0.063
R34179 D_FlipFlop_2.3-input-nand_2.C.n9 D_FlipFlop_2.3-input-nand_2.C.n8 0.063
R34180 D_FlipFlop_2.3-input-nand_2.C.n8 D_FlipFlop_2.3-input-nand_2.C.n3 0.063
R34181 D_FlipFlop_2.3-input-nand_2.C.n12 D_FlipFlop_2.3-input-nand_2.C.n10 0.0435206
R34182 D_FlipFlop_2.3-input-nand_2.C.n14 D_FlipFlop_2.3-input-nand_2.C.n1 0.0216397
R34183 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.C.n14 0.0216397
R34184 D_FlipFlop_2.3-input-nand_2.C.n5 D_FlipFlop_2.3-input-nand_2.C.n4 0.0107679
R34185 D_FlipFlop_2.3-input-nand_2.C.n4 D_FlipFlop_2.3-input-nand_2.C 0.0107679
R34186 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.t2 168.553
R34187 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.t0 168.542
R34188 CDAC8_0.switch_9.Z.n0 CDAC8_0.switch_9.Z.t1 60.321
R34189 CDAC8_0.switch_9.Z.n0 CDAC8_0.switch_9.Z.t3 60.321
R34190 CDAC8_0.switch_9.Z.n23 CDAC8_0.switch_9.Z.n22 14.237
R34191 CDAC8_0.switch_9.Z.n36 CDAC8_0.switch_9.Z.n35 11.3711
R34192 CDAC8_0.switch_9.Z.n35 CDAC8_0.switch_9.Z.n5 7.35843
R34193 CDAC8_0.switch_9.Z.n35 CDAC8_0.switch_9.Z.n34 6.87433
R34194 CDAC8_0.switch_9.Z.n2 CDAC8_0.switch_9.Z.n1 1.58202
R34195 CDAC8_0.switch_9.Z.n3 CDAC8_0.switch_9.Z.t25 0.77316
R34196 CDAC8_0.switch_9.Z.n6 CDAC8_0.switch_9.Z.t28 0.77316
R34197 CDAC8_0.switch_9.Z.n8 CDAC8_0.switch_9.Z.t31 0.77316
R34198 CDAC8_0.switch_9.Z.n20 CDAC8_0.switch_9.Z.t29 0.77316
R34199 CDAC8_0.switch_9.Z.n3 CDAC8_0.switch_9.Z.t23 0.611304
R34200 CDAC8_0.switch_9.Z.n4 CDAC8_0.switch_9.Z.t32 0.611304
R34201 CDAC8_0.switch_9.Z.n10 CDAC8_0.switch_9.Z.t30 0.611304
R34202 CDAC8_0.switch_9.Z.n11 CDAC8_0.switch_9.Z.t10 0.611304
R34203 CDAC8_0.switch_9.Z.n12 CDAC8_0.switch_9.Z.t14 0.611304
R34204 CDAC8_0.switch_9.Z.n13 CDAC8_0.switch_9.Z.t13 0.611304
R34205 CDAC8_0.switch_9.Z.n14 CDAC8_0.switch_9.Z.t18 0.611304
R34206 CDAC8_0.switch_9.Z.n15 CDAC8_0.switch_9.Z.t17 0.611304
R34207 CDAC8_0.switch_9.Z.n16 CDAC8_0.switch_9.Z.t34 0.611304
R34208 CDAC8_0.switch_9.Z.n17 CDAC8_0.switch_9.Z.t6 0.611304
R34209 CDAC8_0.switch_9.Z.n18 CDAC8_0.switch_9.Z.t5 0.611304
R34210 CDAC8_0.switch_9.Z.n19 CDAC8_0.switch_9.Z.t9 0.611304
R34211 CDAC8_0.switch_9.Z.n6 CDAC8_0.switch_9.Z.t27 0.611304
R34212 CDAC8_0.switch_9.Z.n7 CDAC8_0.switch_9.Z.t35 0.611304
R34213 CDAC8_0.switch_9.Z.n33 CDAC8_0.switch_9.Z.t33 0.611304
R34214 CDAC8_0.switch_9.Z.n32 CDAC8_0.switch_9.Z.t12 0.611304
R34215 CDAC8_0.switch_9.Z.n31 CDAC8_0.switch_9.Z.t16 0.611304
R34216 CDAC8_0.switch_9.Z.n30 CDAC8_0.switch_9.Z.t15 0.611304
R34217 CDAC8_0.switch_9.Z.n29 CDAC8_0.switch_9.Z.t21 0.611304
R34218 CDAC8_0.switch_9.Z.n28 CDAC8_0.switch_9.Z.t19 0.611304
R34219 CDAC8_0.switch_9.Z.n27 CDAC8_0.switch_9.Z.t4 0.611304
R34220 CDAC8_0.switch_9.Z.n26 CDAC8_0.switch_9.Z.t8 0.611304
R34221 CDAC8_0.switch_9.Z.n25 CDAC8_0.switch_9.Z.t7 0.611304
R34222 CDAC8_0.switch_9.Z.n24 CDAC8_0.switch_9.Z.t11 0.611304
R34223 CDAC8_0.switch_9.Z.n9 CDAC8_0.switch_9.Z.t26 0.611304
R34224 CDAC8_0.switch_9.Z.n8 CDAC8_0.switch_9.Z.t24 0.611304
R34225 CDAC8_0.switch_9.Z.n21 CDAC8_0.switch_9.Z.t22 0.611304
R34226 CDAC8_0.switch_9.Z.n20 CDAC8_0.switch_9.Z.t20 0.611304
R34227 CDAC8_0.switch_9.Z.n1 CDAC8_0.switch_9.Z 0.259656
R34228 CDAC8_0.switch_9.Z.n2 CDAC8_0.switch_9.Z 0.188
R34229 CDAC8_0.switch_9.Z.n7 CDAC8_0.switch_9.Z.n6 0.162356
R34230 CDAC8_0.switch_9.Z.n33 CDAC8_0.switch_9.Z.n32 0.162356
R34231 CDAC8_0.switch_9.Z.n32 CDAC8_0.switch_9.Z.n31 0.162356
R34232 CDAC8_0.switch_9.Z.n31 CDAC8_0.switch_9.Z.n30 0.162356
R34233 CDAC8_0.switch_9.Z.n30 CDAC8_0.switch_9.Z.n29 0.162356
R34234 CDAC8_0.switch_9.Z.n29 CDAC8_0.switch_9.Z.n28 0.162356
R34235 CDAC8_0.switch_9.Z.n28 CDAC8_0.switch_9.Z.n27 0.162356
R34236 CDAC8_0.switch_9.Z.n27 CDAC8_0.switch_9.Z.n26 0.162356
R34237 CDAC8_0.switch_9.Z.n26 CDAC8_0.switch_9.Z.n25 0.162356
R34238 CDAC8_0.switch_9.Z.n25 CDAC8_0.switch_9.Z.n24 0.162356
R34239 CDAC8_0.switch_9.Z.n9 CDAC8_0.switch_9.Z.n8 0.162356
R34240 CDAC8_0.switch_9.Z.n4 CDAC8_0.switch_9.Z.n3 0.162356
R34241 CDAC8_0.switch_9.Z.n11 CDAC8_0.switch_9.Z.n10 0.162356
R34242 CDAC8_0.switch_9.Z.n12 CDAC8_0.switch_9.Z.n11 0.162356
R34243 CDAC8_0.switch_9.Z.n13 CDAC8_0.switch_9.Z.n12 0.162356
R34244 CDAC8_0.switch_9.Z.n14 CDAC8_0.switch_9.Z.n13 0.162356
R34245 CDAC8_0.switch_9.Z.n15 CDAC8_0.switch_9.Z.n14 0.162356
R34246 CDAC8_0.switch_9.Z.n16 CDAC8_0.switch_9.Z.n15 0.162356
R34247 CDAC8_0.switch_9.Z.n17 CDAC8_0.switch_9.Z.n16 0.162356
R34248 CDAC8_0.switch_9.Z.n18 CDAC8_0.switch_9.Z.n17 0.162356
R34249 CDAC8_0.switch_9.Z.n19 CDAC8_0.switch_9.Z.n18 0.162356
R34250 CDAC8_0.switch_9.Z.n21 CDAC8_0.switch_9.Z.n20 0.162356
R34251 CDAC8_0.switch_9.Z.n34 CDAC8_0.switch_9.Z.n33 0.115412
R34252 CDAC8_0.switch_9.Z.n10 CDAC8_0.switch_9.Z.n5 0.115412
R34253 CDAC8_0.switch_9.Z.n23 CDAC8_0.switch_9.Z.n9 0.0845094
R34254 CDAC8_0.switch_9.Z.n22 CDAC8_0.switch_9.Z.n21 0.0845094
R34255 CDAC8_0.switch_9.Z.n24 CDAC8_0.switch_9.Z.n23 0.0783469
R34256 CDAC8_0.switch_9.Z.n22 CDAC8_0.switch_9.Z.n19 0.0783469
R34257 CDAC8_0.switch_9.Z.n36 CDAC8_0.switch_9.Z.n2 0.063
R34258 CDAC8_0.switch_9.Z.n34 CDAC8_0.switch_9.Z.n7 0.0474438
R34259 CDAC8_0.switch_9.Z.n5 CDAC8_0.switch_9.Z.n4 0.0474438
R34260 CDAC8_0.switch_9.Z CDAC8_0.switch_9.Z.n37 0.0454219
R34261 CDAC8_0.switch_9.Z.n37 CDAC8_0.switch_9.Z.n36 0.0278438
R34262 CDAC8_0.switch_9.Z.n1 CDAC8_0.switch_9.Z.n0 0.0188121
R34263 Nand_Gate_5.B.n24 Nand_Gate_5.B.t0 169.46
R34264 Nand_Gate_5.B.n24 Nand_Gate_5.B.t1 167.809
R34265 Nand_Gate_5.B.n26 Nand_Gate_5.B.t2 167.809
R34266 Nand_Gate_5.B Nand_Gate_5.B.t7 158.585
R34267 Nand_Gate_5.B.t7 Nand_Gate_5.B.n20 150.293
R34268 Nand_Gate_5.B.n16 Nand_Gate_5.B.t6 150.273
R34269 Nand_Gate_5.B.n5 Nand_Gate_5.B.t11 150.273
R34270 Nand_Gate_5.B.n0 Nand_Gate_5.B.t9 150.273
R34271 Nand_Gate_5.B.t5 Nand_Gate_5.B.n17 82.5626
R34272 Nand_Gate_5.B Nand_Gate_5.B.t10 81.5603
R34273 Nand_Gate_5.B.n3 Nand_Gate_5.B.t8 73.6406
R34274 Nand_Gate_5.B.t10 Nand_Gate_5.B.n11 73.6406
R34275 Nand_Gate_5.B.n13 Nand_Gate_5.B.t4 73.6304
R34276 Nand_Gate_5.B.n18 Nand_Gate_5.B.t5 73.6304
R34277 Nand_Gate_5.B.n22 Nand_Gate_5.B.t3 60.3809
R34278 Nand_Gate_5.B.n17 Nand_Gate_5.B.n16 32.9078
R34279 Nand_Gate_5.B.n17 Nand_Gate_5.B.n12 25.3147
R34280 Nand_Gate_5.B.n9 Nand_Gate_5.B.n8 12.6418
R34281 Nand_Gate_5.B.n25 Nand_Gate_5.B.n24 11.4489
R34282 Nand_Gate_5.B.n27 Nand_Gate_5.B.n26 8.21389
R34283 Nand_Gate_5.B.n23 Nand_Gate_5.B.n22 1.64452
R34284 Nand_Gate_5.B.n20 Nand_Gate_5.B.n19 1.19615
R34285 Nand_Gate_5.B.n15 Nand_Gate_5.B.n14 1.1717
R34286 Nand_Gate_5.B.n15 Nand_Gate_5.B 0.932141
R34287 Nand_Gate_5.B.n4 Nand_Gate_5.B 0.851043
R34288 Nand_Gate_5.B.n10 Nand_Gate_5.B 0.851043
R34289 Nand_Gate_5.B.n22 Nand_Gate_5.B 0.848156
R34290 Nand_Gate_5.B.n7 Nand_Gate_5.B.n6 0.55213
R34291 Nand_Gate_5.B.n2 Nand_Gate_5.B.n1 0.55213
R34292 Nand_Gate_5.B.n7 Nand_Gate_5.B 0.486828
R34293 Nand_Gate_5.B.n2 Nand_Gate_5.B 0.486828
R34294 Nand_Gate_5.B.n4 Nand_Gate_5.B.n3 0.470609
R34295 Nand_Gate_5.B.n11 Nand_Gate_5.B.n10 0.470609
R34296 Nand_Gate_5.B.n20 Nand_Gate_5.B 0.447191
R34297 Nand_Gate_5.B.n27 Nand_Gate_5.B.n21 0.425067
R34298 Nand_Gate_5.B Nand_Gate_5.B.n27 0.39003
R34299 Nand_Gate_5.B.n26 Nand_Gate_5.B.n25 0.280391
R34300 Nand_Gate_5.B.n3 Nand_Gate_5.B 0.217464
R34301 Nand_Gate_5.B.n11 Nand_Gate_5.B 0.217464
R34302 Nand_Gate_5.B.n25 Nand_Gate_5.B 0.200143
R34303 Nand_Gate_5.B.n23 Nand_Gate_5.B 0.1255
R34304 Nand_Gate_5.B.n14 Nand_Gate_5.B 0.1255
R34305 Nand_Gate_5.B.n6 Nand_Gate_5.B 0.1255
R34306 Nand_Gate_5.B.n1 Nand_Gate_5.B 0.1255
R34307 Nand_Gate_5.B.n19 Nand_Gate_5.B 0.1255
R34308 Nand_Gate_5.B Nand_Gate_5.B.n23 0.063
R34309 Nand_Gate_5.B.n16 Nand_Gate_5.B.n15 0.063
R34310 Nand_Gate_5.B.n8 Nand_Gate_5.B.n4 0.063
R34311 Nand_Gate_5.B.n8 Nand_Gate_5.B.n7 0.063
R34312 Nand_Gate_5.B.n10 Nand_Gate_5.B.n9 0.063
R34313 Nand_Gate_5.B.n9 Nand_Gate_5.B.n2 0.063
R34314 Nand_Gate_5.B.n6 Nand_Gate_5.B.n5 0.0216397
R34315 Nand_Gate_5.B.n5 Nand_Gate_5.B 0.0216397
R34316 Nand_Gate_5.B.n1 Nand_Gate_5.B.n0 0.0216397
R34317 Nand_Gate_5.B.n0 Nand_Gate_5.B 0.0216397
R34318 Nand_Gate_5.B.n14 Nand_Gate_5.B.n13 0.0107679
R34319 Nand_Gate_5.B.n13 Nand_Gate_5.B 0.0107679
R34320 Nand_Gate_5.B.n19 Nand_Gate_5.B.n18 0.0107679
R34321 Nand_Gate_5.B.n18 Nand_Gate_5.B 0.0107679
R34322 Nand_Gate_5.B.n12 Nand_Gate_5.B 0.00441667
R34323 Nand_Gate_5.B.n21 Nand_Gate_5.B 0.00441667
R34324 Nand_Gate_5.B.n12 Nand_Gate_5.B 0.00406061
R34325 Nand_Gate_5.B.n21 Nand_Gate_5.B 0.00406061
R34326 Nand_Gate_6.A.n33 Nand_Gate_6.A.t0 169.46
R34327 Nand_Gate_6.A.n33 Nand_Gate_6.A.t3 167.809
R34328 Nand_Gate_6.A.n35 Nand_Gate_6.A.t2 167.809
R34329 Nand_Gate_6.A Nand_Gate_6.A.t11 158.585
R34330 Nand_Gate_6.A.n21 Nand_Gate_6.A.t9 150.293
R34331 Nand_Gate_6.A.t11 Nand_Gate_6.A.n2 150.293
R34332 Nand_Gate_6.A.n14 Nand_Gate_6.A.t8 150.273
R34333 Nand_Gate_6.A.n8 Nand_Gate_6.A.t10 150.273
R34334 Nand_Gate_6.A.n12 Nand_Gate_6.A.t6 73.6406
R34335 Nand_Gate_6.A.n6 Nand_Gate_6.A.t4 73.6406
R34336 Nand_Gate_6.A.n23 Nand_Gate_6.A.t5 73.6304
R34337 Nand_Gate_6.A.n0 Nand_Gate_6.A.t7 73.6304
R34338 Nand_Gate_6.A.n4 Nand_Gate_6.A.t1 60.3809
R34339 Nand_Gate_6.A.n27 Nand_Gate_6.A.n26 14.3097
R34340 Nand_Gate_6.A.n34 Nand_Gate_6.A.n33 11.4489
R34341 Nand_Gate_6.A.n36 Nand_Gate_6.A.n35 8.21389
R34342 Nand_Gate_6.A.n18 Nand_Gate_6.A.n11 8.1418
R34343 Nand_Gate_6.A.n29 Nand_Gate_6.A.n28 5.61191
R34344 Nand_Gate_6.A.n29 Nand_Gate_6.A 5.35402
R34345 Nand_Gate_6.A.n30 Nand_Gate_6.A.n29 4.563
R34346 Nand_Gate_6.A.n18 Nand_Gate_6.A.n17 4.5005
R34347 Nand_Gate_6.A.n28 Nand_Gate_6.A 1.83746
R34348 Nand_Gate_6.A.n20 Nand_Gate_6.A.n19 1.62007
R34349 Nand_Gate_6.A.n2 Nand_Gate_6.A.n1 1.19615
R34350 Nand_Gate_6.A.n5 Nand_Gate_6.A 1.08746
R34351 Nand_Gate_6.A.n20 Nand_Gate_6.A 1.01739
R34352 Nand_Gate_6.A.n13 Nand_Gate_6.A 0.851043
R34353 Nand_Gate_6.A.n7 Nand_Gate_6.A 0.851043
R34354 Nand_Gate_6.A.n4 Nand_Gate_6.A 0.848156
R34355 Nand_Gate_6.A.n32 Nand_Gate_6.A.n31 0.788543
R34356 Nand_Gate_6.A.n22 Nand_Gate_6.A 0.769522
R34357 Nand_Gate_6.A.n5 Nand_Gate_6.A.n4 0.682565
R34358 Nand_Gate_6.A.n31 Nand_Gate_6.A 0.65675
R34359 Nand_Gate_6.A.n22 Nand_Gate_6.A.n21 0.55213
R34360 Nand_Gate_6.A.n16 Nand_Gate_6.A.n15 0.55213
R34361 Nand_Gate_6.A.n10 Nand_Gate_6.A.n9 0.55213
R34362 Nand_Gate_6.A.n16 Nand_Gate_6.A 0.486828
R34363 Nand_Gate_6.A.n10 Nand_Gate_6.A 0.486828
R34364 Nand_Gate_6.A.n25 Nand_Gate_6.A.n24 0.470609
R34365 Nand_Gate_6.A.n13 Nand_Gate_6.A.n12 0.470609
R34366 Nand_Gate_6.A.n7 Nand_Gate_6.A.n6 0.470609
R34367 Nand_Gate_6.A.n21 Nand_Gate_6.A 0.447191
R34368 Nand_Gate_6.A.n2 Nand_Gate_6.A 0.447191
R34369 Nand_Gate_6.A.n25 Nand_Gate_6.A 0.428234
R34370 Nand_Gate_6.A.n36 Nand_Gate_6.A.n3 0.425067
R34371 Nand_Gate_6.A Nand_Gate_6.A.n36 0.39003
R34372 Nand_Gate_6.A.n35 Nand_Gate_6.A.n34 0.280391
R34373 Nand_Gate_6.A.n34 Nand_Gate_6.A.n32 0.262643
R34374 Nand_Gate_6.A.n12 Nand_Gate_6.A 0.217464
R34375 Nand_Gate_6.A.n6 Nand_Gate_6.A 0.217464
R34376 Nand_Gate_6.A.n24 Nand_Gate_6.A 0.1255
R34377 Nand_Gate_6.A.n15 Nand_Gate_6.A 0.1255
R34378 Nand_Gate_6.A.n9 Nand_Gate_6.A 0.1255
R34379 Nand_Gate_6.A.n32 Nand_Gate_6.A 0.1255
R34380 Nand_Gate_6.A.n1 Nand_Gate_6.A 0.1255
R34381 Nand_Gate_6.A.n26 Nand_Gate_6.A.n22 0.063
R34382 Nand_Gate_6.A.n26 Nand_Gate_6.A.n25 0.063
R34383 Nand_Gate_6.A.n17 Nand_Gate_6.A.n13 0.063
R34384 Nand_Gate_6.A.n17 Nand_Gate_6.A.n16 0.063
R34385 Nand_Gate_6.A.n11 Nand_Gate_6.A.n7 0.063
R34386 Nand_Gate_6.A.n11 Nand_Gate_6.A.n10 0.063
R34387 Nand_Gate_6.A.n28 Nand_Gate_6.A.n27 0.063
R34388 Nand_Gate_6.A.n27 Nand_Gate_6.A.n20 0.063
R34389 Nand_Gate_6.A.n30 Nand_Gate_6.A.n5 0.063
R34390 Nand_Gate_6.A.n31 Nand_Gate_6.A.n30 0.063
R34391 Nand_Gate_6.A.n32 Nand_Gate_6.A 0.063
R34392 Nand_Gate_6.A Nand_Gate_6.A.n18 0.0512812
R34393 Nand_Gate_6.A.n15 Nand_Gate_6.A.n14 0.0216397
R34394 Nand_Gate_6.A.n14 Nand_Gate_6.A 0.0216397
R34395 Nand_Gate_6.A.n9 Nand_Gate_6.A.n8 0.0216397
R34396 Nand_Gate_6.A.n8 Nand_Gate_6.A 0.0216397
R34397 Nand_Gate_6.A.n19 Nand_Gate_6.A 0.0168043
R34398 Nand_Gate_6.A.n19 Nand_Gate_6.A 0.0122188
R34399 Nand_Gate_6.A.n24 Nand_Gate_6.A.n23 0.0107679
R34400 Nand_Gate_6.A.n23 Nand_Gate_6.A 0.0107679
R34401 Nand_Gate_6.A.n1 Nand_Gate_6.A.n0 0.0107679
R34402 Nand_Gate_6.A.n0 Nand_Gate_6.A 0.0107679
R34403 Nand_Gate_6.A.n3 Nand_Gate_6.A 0.00441667
R34404 Nand_Gate_6.A.n3 Nand_Gate_6.A 0.00406061
R34405 FFCLR.n205 FFCLR.t1 169.46
R34406 FFCLR.n207 FFCLR.t3 167.809
R34407 FFCLR.n205 FFCLR.t0 167.809
R34408 FFCLR.n45 FFCLR.t27 158.988
R34409 FFCLR.n84 FFCLR.t7 158.965
R34410 FFCLR.n64 FFCLR.t45 158.965
R34411 FFCLR.n187 FFCLR.t55 158.965
R34412 FFCLR.n165 FFCLR.t5 158.965
R34413 FFCLR.n143 FFCLR.t9 158.965
R34414 FFCLR.n121 FFCLR.t49 158.965
R34415 FFCLR FFCLR.t6 158.585
R34416 FFCLR FFCLR.t44 158.581
R34417 FFCLR.n192 FFCLR.t16 150.293
R34418 FFCLR.n93 FFCLR.t56 150.293
R34419 FFCLR.n87 FFCLR.t24 150.293
R34420 FFCLR.n73 FFCLR.t22 150.293
R34421 FFCLR.n67 FFCLR.t50 150.293
R34422 FFCLR.n53 FFCLR.t8 150.293
R34423 FFCLR.n47 FFCLR.t33 150.293
R34424 FFCLR.n174 FFCLR.t30 150.293
R34425 FFCLR.n168 FFCLR.t58 150.293
R34426 FFCLR.n152 FFCLR.t51 150.293
R34427 FFCLR.n146 FFCLR.t21 150.293
R34428 FFCLR.n130 FFCLR.t36 150.293
R34429 FFCLR.n124 FFCLR.t10 150.293
R34430 FFCLR.n108 FFCLR.t28 150.293
R34431 FFCLR.n102 FFCLR.t54 150.293
R34432 FFCLR.t44 FFCLR.n38 150.293
R34433 FFCLR.t6 FFCLR.n2 150.293
R34434 FFCLR.t7 FFCLR.n83 150.273
R34435 FFCLR.t45 FFCLR.n63 150.273
R34436 FFCLR.t27 FFCLR.n44 150.273
R34437 FFCLR.t55 FFCLR.n186 150.273
R34438 FFCLR.t5 FFCLR.n164 150.273
R34439 FFCLR.t9 FFCLR.n142 150.273
R34440 FFCLR.t49 FFCLR.n120 150.273
R34441 FFCLR.n29 FFCLR.t38 150.273
R34442 FFCLR.n23 FFCLR.t11 150.273
R34443 FFCLR.n14 FFCLR.t40 150.273
R34444 FFCLR.n8 FFCLR.t34 150.273
R34445 FFCLR.n198 FFCLR.n191 88.4503
R34446 FFCLR.n81 FFCLR.t14 73.6406
R34447 FFCLR.n61 FFCLR.t37 73.6406
R34448 FFCLR.n42 FFCLR.t19 73.6406
R34449 FFCLR.n184 FFCLR.t20 73.6406
R34450 FFCLR.n162 FFCLR.t52 73.6406
R34451 FFCLR.n140 FFCLR.t15 73.6406
R34452 FFCLR.n118 FFCLR.t43 73.6406
R34453 FFCLR.n27 FFCLR.t13 73.6406
R34454 FFCLR.n21 FFCLR.t39 73.6406
R34455 FFCLR.n12 FFCLR.t32 73.6406
R34456 FFCLR.n6 FFCLR.t41 73.6406
R34457 FFCLR.n194 FFCLR.t48 73.6304
R34458 FFCLR.n95 FFCLR.t4 73.6304
R34459 FFCLR.n89 FFCLR.t31 73.6304
R34460 FFCLR.n75 FFCLR.t42 73.6304
R34461 FFCLR.n69 FFCLR.t12 73.6304
R34462 FFCLR.n55 FFCLR.t23 73.6304
R34463 FFCLR.n49 FFCLR.t53 73.6304
R34464 FFCLR.n176 FFCLR.t47 73.6304
R34465 FFCLR.n170 FFCLR.t18 73.6304
R34466 FFCLR.n154 FFCLR.t57 73.6304
R34467 FFCLR.n148 FFCLR.t25 73.6304
R34468 FFCLR.n132 FFCLR.t59 73.6304
R34469 FFCLR.n126 FFCLR.t29 73.6304
R34470 FFCLR.n110 FFCLR.t46 73.6304
R34471 FFCLR.n104 FFCLR.t17 73.6304
R34472 FFCLR.n36 FFCLR.t26 73.6304
R34473 FFCLR.n0 FFCLR.t35 73.6304
R34474 FFCLR.n4 FFCLR.t2 60.3809
R34475 FFCLR.n99 FFCLR.n92 15.5222
R34476 FFCLR.n79 FFCLR.n72 15.5222
R34477 FFCLR.n59 FFCLR.n52 15.5222
R34478 FFCLR.n180 FFCLR.n173 15.5222
R34479 FFCLR.n158 FFCLR.n151 15.5222
R34480 FFCLR.n136 FFCLR.n129 15.5222
R34481 FFCLR.n114 FFCLR.n107 15.5222
R34482 FFCLR.n33 FFCLR.n26 15.5222
R34483 FFCLR.n206 FFCLR.n205 11.4489
R34484 FFCLR.n189 FFCLR 10.7094
R34485 FFCLR.n190 FFCLR.n100 9.59712
R34486 FFCLR.n198 FFCLR.n197 9.57083
R34487 FFCLR.n188 FFCLR 9.51957
R34488 FFCLR.n190 FFCLR.n189 9.43184
R34489 FFCLR.n34 FFCLR.n33 8.26552
R34490 FFCLR.n208 FFCLR.n207 8.21389
R34491 FFCLR.n18 FFCLR.n11 8.1418
R34492 FFCLR.n167 FFCLR 7.84808
R34493 FFCLR.n100 FFCLR.n99 7.83713
R34494 FFCLR.n80 FFCLR.n79 7.83713
R34495 FFCLR.n60 FFCLR.n59 7.83713
R34496 FFCLR.n181 FFCLR.n180 7.83713
R34497 FFCLR.n159 FFCLR.n158 7.83713
R34498 FFCLR.n137 FFCLR.n136 7.83713
R34499 FFCLR.n115 FFCLR.n114 7.83713
R34500 FFCLR.n166 FFCLR 6.72777
R34501 FFCLR.n199 FFCLR.n198 6.58222
R34502 FFCLR.n20 FFCLR.n19 6.47604
R34503 FFCLR.n19 FFCLR 5.35402
R34504 FFCLR.n145 FFCLR 5.31008
R34505 FFCLR.n202 FFCLR 4.55128
R34506 FFCLR.n99 FFCLR.n98 4.5005
R34507 FFCLR.n79 FFCLR.n78 4.5005
R34508 FFCLR.n59 FFCLR.n58 4.5005
R34509 FFCLR.n180 FFCLR.n179 4.5005
R34510 FFCLR.n158 FFCLR.n157 4.5005
R34511 FFCLR.n136 FFCLR.n135 4.5005
R34512 FFCLR.n114 FFCLR.n113 4.5005
R34513 FFCLR.n33 FFCLR.n32 4.5005
R34514 FFCLR.n18 FFCLR.n17 4.5005
R34515 FFCLR.n144 FFCLR 3.93597
R34516 FFCLR.n191 FFCLR.n41 3.73088
R34517 FFCLR.n191 FFCLR.n190 3.4105
R34518 FFCLR.n123 FFCLR 2.77208
R34519 FFCLR.n189 FFCLR.n188 2.2612
R34520 FFCLR.n64 FFCLR.n60 1.95257
R34521 FFCLR.n84 FFCLR.n80 1.95257
R34522 FFCLR.n123 FFCLR.n122 1.90557
R34523 FFCLR.n145 FFCLR.n144 1.90557
R34524 FFCLR.n167 FFCLR.n166 1.90557
R34525 FFCLR.n82 FFCLR.n81 1.19615
R34526 FFCLR.n62 FFCLR.n61 1.19615
R34527 FFCLR.n43 FFCLR.n42 1.19615
R34528 FFCLR.n185 FFCLR.n184 1.19615
R34529 FFCLR.n163 FFCLR.n162 1.19615
R34530 FFCLR.n141 FFCLR.n140 1.19615
R34531 FFCLR.n119 FFCLR.n118 1.19615
R34532 FFCLR.n38 FFCLR.n37 1.19615
R34533 FFCLR.n2 FFCLR.n1 1.19615
R34534 FFCLR.n122 FFCLR 1.14417
R34535 FFCLR.n94 FFCLR 1.09561
R34536 FFCLR.n88 FFCLR 1.09561
R34537 FFCLR.n74 FFCLR 1.09561
R34538 FFCLR.n68 FFCLR 1.09561
R34539 FFCLR.n54 FFCLR 1.09561
R34540 FFCLR.n48 FFCLR 1.09561
R34541 FFCLR.n175 FFCLR 1.09561
R34542 FFCLR.n169 FFCLR 1.09561
R34543 FFCLR.n153 FFCLR 1.09561
R34544 FFCLR.n147 FFCLR 1.09561
R34545 FFCLR.n131 FFCLR 1.09561
R34546 FFCLR.n125 FFCLR 1.09561
R34547 FFCLR.n109 FFCLR 1.09561
R34548 FFCLR.n103 FFCLR 1.09561
R34549 FFCLR.n5 FFCLR 1.08746
R34550 FFCLR.n20 FFCLR 0.973326
R34551 FFCLR.n13 FFCLR 0.851043
R34552 FFCLR.n7 FFCLR 0.851043
R34553 FFCLR.n4 FFCLR 0.848156
R34554 FFCLR.n97 FFCLR.n96 0.796696
R34555 FFCLR.n91 FFCLR.n90 0.796696
R34556 FFCLR.n77 FFCLR.n76 0.796696
R34557 FFCLR.n71 FFCLR.n70 0.796696
R34558 FFCLR.n57 FFCLR.n56 0.796696
R34559 FFCLR.n51 FFCLR.n50 0.796696
R34560 FFCLR.n178 FFCLR.n177 0.796696
R34561 FFCLR.n172 FFCLR.n171 0.796696
R34562 FFCLR.n156 FFCLR.n155 0.796696
R34563 FFCLR.n150 FFCLR.n149 0.796696
R34564 FFCLR.n134 FFCLR.n133 0.796696
R34565 FFCLR.n128 FFCLR.n127 0.796696
R34566 FFCLR.n112 FFCLR.n111 0.796696
R34567 FFCLR.n106 FFCLR.n105 0.796696
R34568 FFCLR.n28 FFCLR.n27 0.796696
R34569 FFCLR.n22 FFCLR.n21 0.796696
R34570 FFCLR.n204 FFCLR.n203 0.788543
R34571 FFCLR.n46 FFCLR.n45 0.783833
R34572 FFCLR.n66 FFCLR.n65 0.783833
R34573 FFCLR.n86 FFCLR.n85 0.783833
R34574 FFCLR.n117 FFCLR.n116 0.783833
R34575 FFCLR.n139 FFCLR.n138 0.783833
R34576 FFCLR.n161 FFCLR.n160 0.783833
R34577 FFCLR.n183 FFCLR.n182 0.783833
R34578 FFCLR.n193 FFCLR 0.769522
R34579 FFCLR.n201 FFCLR.n200 0.755935
R34580 FFCLR.n45 FFCLR 0.716182
R34581 FFCLR.n65 FFCLR 0.716182
R34582 FFCLR.n85 FFCLR 0.716182
R34583 FFCLR.n117 FFCLR 0.716182
R34584 FFCLR.n139 FFCLR 0.716182
R34585 FFCLR.n161 FFCLR 0.716182
R34586 FFCLR.n183 FFCLR 0.716182
R34587 FFCLR.n34 FFCLR 0.716182
R34588 FFCLR.n5 FFCLR.n4 0.682565
R34589 FFCLR.n97 FFCLR 0.662609
R34590 FFCLR.n91 FFCLR 0.662609
R34591 FFCLR.n77 FFCLR 0.662609
R34592 FFCLR.n71 FFCLR 0.662609
R34593 FFCLR.n57 FFCLR 0.662609
R34594 FFCLR.n51 FFCLR 0.662609
R34595 FFCLR.n178 FFCLR 0.662609
R34596 FFCLR.n172 FFCLR 0.662609
R34597 FFCLR.n156 FFCLR 0.662609
R34598 FFCLR.n150 FFCLR 0.662609
R34599 FFCLR.n134 FFCLR 0.662609
R34600 FFCLR.n128 FFCLR 0.662609
R34601 FFCLR.n112 FFCLR 0.662609
R34602 FFCLR.n106 FFCLR 0.662609
R34603 FFCLR.n203 FFCLR 0.65675
R34604 FFCLR.n35 FFCLR.n34 0.565283
R34605 FFCLR.n193 FFCLR.n192 0.55213
R34606 FFCLR.n16 FFCLR.n15 0.55213
R34607 FFCLR.n10 FFCLR.n9 0.55213
R34608 FFCLR.n28 FFCLR 0.524957
R34609 FFCLR.n22 FFCLR 0.524957
R34610 FFCLR.n16 FFCLR 0.486828
R34611 FFCLR.n10 FFCLR 0.486828
R34612 FFCLR.n200 FFCLR 0.48023
R34613 FFCLR.n196 FFCLR.n195 0.470609
R34614 FFCLR.n13 FFCLR.n12 0.470609
R34615 FFCLR.n7 FFCLR.n6 0.470609
R34616 FFCLR.n192 FFCLR 0.447191
R34617 FFCLR.n93 FFCLR 0.447191
R34618 FFCLR.n87 FFCLR 0.447191
R34619 FFCLR.n73 FFCLR 0.447191
R34620 FFCLR.n67 FFCLR 0.447191
R34621 FFCLR.n53 FFCLR 0.447191
R34622 FFCLR.n47 FFCLR 0.447191
R34623 FFCLR.n174 FFCLR 0.447191
R34624 FFCLR.n168 FFCLR 0.447191
R34625 FFCLR.n152 FFCLR 0.447191
R34626 FFCLR.n146 FFCLR 0.447191
R34627 FFCLR.n130 FFCLR 0.447191
R34628 FFCLR.n124 FFCLR 0.447191
R34629 FFCLR.n108 FFCLR 0.447191
R34630 FFCLR.n102 FFCLR 0.447191
R34631 FFCLR.n38 FFCLR 0.447191
R34632 FFCLR.n2 FFCLR 0.447191
R34633 FFCLR.n196 FFCLR 0.428234
R34634 FFCLR.n208 FFCLR.n3 0.425067
R34635 FFCLR FFCLR.n208 0.39003
R34636 FFCLR.n207 FFCLR.n206 0.280391
R34637 FFCLR.n101 FFCLR 0.257433
R34638 FFCLR.n31 FFCLR 0.252453
R34639 FFCLR.n25 FFCLR 0.252453
R34640 FFCLR.n101 FFCLR 0.234076
R34641 FFCLR.n94 FFCLR.n93 0.226043
R34642 FFCLR.n88 FFCLR.n87 0.226043
R34643 FFCLR.n74 FFCLR.n73 0.226043
R34644 FFCLR.n68 FFCLR.n67 0.226043
R34645 FFCLR.n54 FFCLR.n53 0.226043
R34646 FFCLR.n48 FFCLR.n47 0.226043
R34647 FFCLR.n175 FFCLR.n174 0.226043
R34648 FFCLR.n169 FFCLR.n168 0.226043
R34649 FFCLR.n153 FFCLR.n152 0.226043
R34650 FFCLR.n147 FFCLR.n146 0.226043
R34651 FFCLR.n131 FFCLR.n130 0.226043
R34652 FFCLR.n125 FFCLR.n124 0.226043
R34653 FFCLR.n109 FFCLR.n108 0.226043
R34654 FFCLR.n103 FFCLR.n102 0.226043
R34655 FFCLR.n31 FFCLR.n30 0.226043
R34656 FFCLR.n25 FFCLR.n24 0.226043
R34657 FFCLR.n35 FFCLR 0.222967
R34658 FFCLR.n81 FFCLR 0.217464
R34659 FFCLR.n61 FFCLR 0.217464
R34660 FFCLR.n42 FFCLR 0.217464
R34661 FFCLR.n184 FFCLR 0.217464
R34662 FFCLR.n162 FFCLR 0.217464
R34663 FFCLR.n140 FFCLR 0.217464
R34664 FFCLR.n118 FFCLR 0.217464
R34665 FFCLR.n27 FFCLR 0.217464
R34666 FFCLR.n21 FFCLR 0.217464
R34667 FFCLR.n12 FFCLR 0.217464
R34668 FFCLR.n6 FFCLR 0.217464
R34669 FFCLR.n206 FFCLR 0.200143
R34670 FFCLR.n40 FFCLR.n39 0.159517
R34671 FFCLR.n40 FFCLR 0.129132
R34672 FFCLR.n195 FFCLR 0.1255
R34673 FFCLR.n96 FFCLR 0.1255
R34674 FFCLR.n90 FFCLR 0.1255
R34675 FFCLR.n82 FFCLR 0.1255
R34676 FFCLR.n76 FFCLR 0.1255
R34677 FFCLR.n70 FFCLR 0.1255
R34678 FFCLR.n62 FFCLR 0.1255
R34679 FFCLR.n56 FFCLR 0.1255
R34680 FFCLR.n50 FFCLR 0.1255
R34681 FFCLR.n43 FFCLR 0.1255
R34682 FFCLR.n185 FFCLR 0.1255
R34683 FFCLR.n177 FFCLR 0.1255
R34684 FFCLR.n171 FFCLR 0.1255
R34685 FFCLR.n163 FFCLR 0.1255
R34686 FFCLR.n155 FFCLR 0.1255
R34687 FFCLR.n149 FFCLR 0.1255
R34688 FFCLR.n141 FFCLR 0.1255
R34689 FFCLR.n133 FFCLR 0.1255
R34690 FFCLR.n127 FFCLR 0.1255
R34691 FFCLR.n119 FFCLR 0.1255
R34692 FFCLR.n111 FFCLR 0.1255
R34693 FFCLR.n105 FFCLR 0.1255
R34694 FFCLR.n30 FFCLR 0.1255
R34695 FFCLR.n24 FFCLR 0.1255
R34696 FFCLR.n37 FFCLR 0.1255
R34697 FFCLR.n15 FFCLR 0.1255
R34698 FFCLR.n9 FFCLR 0.1255
R34699 FFCLR.n204 FFCLR 0.1255
R34700 FFCLR.n1 FFCLR 0.1255
R34701 FFCLR.n197 FFCLR.n193 0.063
R34702 FFCLR.n197 FFCLR.n196 0.063
R34703 FFCLR.n98 FFCLR.n94 0.063
R34704 FFCLR.n98 FFCLR.n97 0.063
R34705 FFCLR.n92 FFCLR.n88 0.063
R34706 FFCLR.n92 FFCLR.n91 0.063
R34707 FFCLR.n78 FFCLR.n74 0.063
R34708 FFCLR.n78 FFCLR.n77 0.063
R34709 FFCLR.n72 FFCLR.n68 0.063
R34710 FFCLR.n72 FFCLR.n71 0.063
R34711 FFCLR.n58 FFCLR.n54 0.063
R34712 FFCLR.n58 FFCLR.n57 0.063
R34713 FFCLR.n52 FFCLR.n48 0.063
R34714 FFCLR.n52 FFCLR.n51 0.063
R34715 FFCLR.n179 FFCLR.n175 0.063
R34716 FFCLR.n179 FFCLR.n178 0.063
R34717 FFCLR.n173 FFCLR.n169 0.063
R34718 FFCLR.n173 FFCLR.n172 0.063
R34719 FFCLR.n157 FFCLR.n153 0.063
R34720 FFCLR.n157 FFCLR.n156 0.063
R34721 FFCLR.n151 FFCLR.n147 0.063
R34722 FFCLR.n151 FFCLR.n150 0.063
R34723 FFCLR.n135 FFCLR.n131 0.063
R34724 FFCLR.n135 FFCLR.n134 0.063
R34725 FFCLR.n129 FFCLR.n125 0.063
R34726 FFCLR.n129 FFCLR.n128 0.063
R34727 FFCLR.n113 FFCLR.n109 0.063
R34728 FFCLR.n113 FFCLR.n112 0.063
R34729 FFCLR.n107 FFCLR.n103 0.063
R34730 FFCLR.n107 FFCLR.n106 0.063
R34731 FFCLR.n32 FFCLR.n28 0.063
R34732 FFCLR.n32 FFCLR.n31 0.063
R34733 FFCLR.n26 FFCLR.n22 0.063
R34734 FFCLR.n26 FFCLR.n25 0.063
R34735 FFCLR.n17 FFCLR.n13 0.063
R34736 FFCLR.n17 FFCLR.n16 0.063
R34737 FFCLR.n11 FFCLR.n7 0.063
R34738 FFCLR.n11 FFCLR.n10 0.063
R34739 FFCLR.n19 FFCLR.n18 0.063
R34740 FFCLR.n199 FFCLR.n20 0.063
R34741 FFCLR.n200 FFCLR.n199 0.063
R34742 FFCLR.n202 FFCLR.n5 0.063
R34743 FFCLR.n203 FFCLR.n202 0.063
R34744 FFCLR FFCLR.n204 0.063
R34745 FFCLR.n65 FFCLR.n64 0.024
R34746 FFCLR.n85 FFCLR.n84 0.024
R34747 FFCLR.n115 FFCLR.n101 0.024
R34748 FFCLR.n122 FFCLR.n121 0.024
R34749 FFCLR.n121 FFCLR.n117 0.024
R34750 FFCLR.n137 FFCLR.n123 0.024
R34751 FFCLR.n144 FFCLR.n143 0.024
R34752 FFCLR.n143 FFCLR.n139 0.024
R34753 FFCLR.n159 FFCLR.n145 0.024
R34754 FFCLR.n166 FFCLR.n165 0.024
R34755 FFCLR.n165 FFCLR.n161 0.024
R34756 FFCLR.n181 FFCLR.n167 0.024
R34757 FFCLR.n188 FFCLR.n187 0.024
R34758 FFCLR.n187 FFCLR.n183 0.024
R34759 FFCLR.n41 FFCLR.n35 0.024
R34760 FFCLR.n41 FFCLR.n40 0.024
R34761 FFCLR.n83 FFCLR.n82 0.0216397
R34762 FFCLR.n83 FFCLR 0.0216397
R34763 FFCLR.n63 FFCLR.n62 0.0216397
R34764 FFCLR.n63 FFCLR 0.0216397
R34765 FFCLR.n44 FFCLR.n43 0.0216397
R34766 FFCLR.n44 FFCLR 0.0216397
R34767 FFCLR.n186 FFCLR.n185 0.0216397
R34768 FFCLR.n186 FFCLR 0.0216397
R34769 FFCLR.n164 FFCLR.n163 0.0216397
R34770 FFCLR.n164 FFCLR 0.0216397
R34771 FFCLR.n142 FFCLR.n141 0.0216397
R34772 FFCLR.n142 FFCLR 0.0216397
R34773 FFCLR.n120 FFCLR.n119 0.0216397
R34774 FFCLR.n120 FFCLR 0.0216397
R34775 FFCLR.n30 FFCLR.n29 0.0216397
R34776 FFCLR.n29 FFCLR 0.0216397
R34777 FFCLR.n24 FFCLR.n23 0.0216397
R34778 FFCLR.n23 FFCLR 0.0216397
R34779 FFCLR.n15 FFCLR.n14 0.0216397
R34780 FFCLR.n14 FFCLR 0.0216397
R34781 FFCLR.n9 FFCLR.n8 0.0216397
R34782 FFCLR.n8 FFCLR 0.0216397
R34783 FFCLR.n60 FFCLR 0.0204394
R34784 FFCLR.n80 FFCLR 0.0204394
R34785 FFCLR.n100 FFCLR 0.0204394
R34786 FFCLR FFCLR.n115 0.0204394
R34787 FFCLR FFCLR.n137 0.0204394
R34788 FFCLR FFCLR.n159 0.0204394
R34789 FFCLR FFCLR.n181 0.0204394
R34790 FFCLR.n201 FFCLR 0.0168043
R34791 FFCLR FFCLR.n201 0.0122188
R34792 FFCLR.n195 FFCLR.n194 0.0107679
R34793 FFCLR.n194 FFCLR 0.0107679
R34794 FFCLR.n96 FFCLR.n95 0.0107679
R34795 FFCLR.n95 FFCLR 0.0107679
R34796 FFCLR.n90 FFCLR.n89 0.0107679
R34797 FFCLR.n89 FFCLR 0.0107679
R34798 FFCLR.n76 FFCLR.n75 0.0107679
R34799 FFCLR.n75 FFCLR 0.0107679
R34800 FFCLR.n70 FFCLR.n69 0.0107679
R34801 FFCLR.n69 FFCLR 0.0107679
R34802 FFCLR.n56 FFCLR.n55 0.0107679
R34803 FFCLR.n55 FFCLR 0.0107679
R34804 FFCLR.n50 FFCLR.n49 0.0107679
R34805 FFCLR.n49 FFCLR 0.0107679
R34806 FFCLR.n177 FFCLR.n176 0.0107679
R34807 FFCLR.n176 FFCLR 0.0107679
R34808 FFCLR.n171 FFCLR.n170 0.0107679
R34809 FFCLR.n170 FFCLR 0.0107679
R34810 FFCLR.n155 FFCLR.n154 0.0107679
R34811 FFCLR.n154 FFCLR 0.0107679
R34812 FFCLR.n149 FFCLR.n148 0.0107679
R34813 FFCLR.n148 FFCLR 0.0107679
R34814 FFCLR.n133 FFCLR.n132 0.0107679
R34815 FFCLR.n132 FFCLR 0.0107679
R34816 FFCLR.n127 FFCLR.n126 0.0107679
R34817 FFCLR.n126 FFCLR 0.0107679
R34818 FFCLR.n111 FFCLR.n110 0.0107679
R34819 FFCLR.n110 FFCLR 0.0107679
R34820 FFCLR.n105 FFCLR.n104 0.0107679
R34821 FFCLR.n104 FFCLR 0.0107679
R34822 FFCLR.n37 FFCLR.n36 0.0107679
R34823 FFCLR.n36 FFCLR 0.0107679
R34824 FFCLR.n1 FFCLR.n0 0.0107679
R34825 FFCLR.n0 FFCLR 0.0107679
R34826 FFCLR.n46 FFCLR 0.00441667
R34827 FFCLR.n66 FFCLR 0.00441667
R34828 FFCLR.n86 FFCLR 0.00441667
R34829 FFCLR.n116 FFCLR 0.00441667
R34830 FFCLR.n138 FFCLR 0.00441667
R34831 FFCLR.n160 FFCLR 0.00441667
R34832 FFCLR.n182 FFCLR 0.00441667
R34833 FFCLR.n39 FFCLR 0.00441667
R34834 FFCLR.n3 FFCLR 0.00441667
R34835 FFCLR FFCLR.n46 0.00406061
R34836 FFCLR FFCLR.n66 0.00406061
R34837 FFCLR FFCLR.n86 0.00406061
R34838 FFCLR.n116 FFCLR 0.00406061
R34839 FFCLR.n138 FFCLR 0.00406061
R34840 FFCLR.n160 FFCLR 0.00406061
R34841 FFCLR.n182 FFCLR 0.00406061
R34842 FFCLR.n39 FFCLR 0.00406061
R34843 FFCLR.n3 FFCLR 0.00406061
R34844 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 316.762
R34845 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 168.108
R34846 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 150.293
R34847 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 150.273
R34848 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 73.6406
R34849 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 73.6304
R34850 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 60.3943
R34851 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 12.0358
R34852 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 1.19615
R34853 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.981478
R34854 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 0.788543
R34855 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.769522
R34856 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 0.682565
R34857 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.580578
R34858 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 0.55213
R34859 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 0.484875
R34860 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 0.470609
R34861 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.447191
R34862 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.428234
R34863 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.217464
R34864 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R34865 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R34866 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.1255
R34867 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 0.063
R34868 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 0.063
R34869 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.063
R34870 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 0.063
R34871 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 0.063
R34872 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 0.0216397
R34873 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.0216397
R34874 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 0.0107679
R34875 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.0107679
R34876 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 179.256
R34877 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 168.089
R34878 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 150.293
R34879 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 73.6304
R34880 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 60.3943
R34881 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 12.0358
R34882 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.981478
R34883 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 0.788543
R34884 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.769522
R34885 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 0.720633
R34886 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 0.682565
R34887 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.580578
R34888 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 0.55213
R34889 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 0.470609
R34890 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.447191
R34891 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.428234
R34892 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1255
R34893 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1255
R34894 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 0.063
R34895 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 0.063
R34896 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.063
R34897 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 0.063
R34898 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 0.063
R34899 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 0.0435206
R34900 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 0.0107679
R34901 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.0107679
R34902 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 316.762
R34903 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 168.108
R34904 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 150.293
R34905 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 150.273
R34906 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 73.6406
R34907 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 73.6304
R34908 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 60.4568
R34909 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 12.0358
R34910 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 1.19615
R34911 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.981478
R34912 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 0.788543
R34913 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.769522
R34914 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 0.682565
R34915 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.580578
R34916 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 0.55213
R34917 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 0.484875
R34918 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 0.470609
R34919 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.447191
R34920 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.428234
R34921 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.217464
R34922 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R34923 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R34924 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.1255
R34925 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 0.063
R34926 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 0.063
R34927 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.063
R34928 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 0.063
R34929 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 0.063
R34930 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 0.0216397
R34931 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.0216397
R34932 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 0.0107679
R34933 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.0107679
R34934 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 179.256
R34935 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 168.089
R34936 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 150.293
R34937 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 73.6304
R34938 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 60.4568
R34939 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 12.0358
R34940 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.981478
R34941 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 0.788543
R34942 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.769522
R34943 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 0.720633
R34944 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 0.682565
R34945 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.580578
R34946 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 0.55213
R34947 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 0.470609
R34948 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.447191
R34949 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.428234
R34950 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1255
R34951 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1255
R34952 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 0.063
R34953 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 0.063
R34954 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.063
R34955 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 0.063
R34956 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 0.063
R34957 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 0.0435206
R34958 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 0.0107679
R34959 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.0107679
R34960 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 169.46
R34961 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 167.809
R34962 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 167.809
R34963 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 167.226
R34964 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 150.273
R34965 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 150.273
R34966 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 73.6406
R34967 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 73.6304
R34968 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 60.3943
R34969 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 12.3891
R34970 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 11.4489
R34971 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 1.68257
R34972 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 1.38365
R34973 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 1.19615
R34974 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 1.1717
R34975 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 1.08448
R34976 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.932141
R34977 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.720633
R34978 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 0.280391
R34979 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.217464
R34980 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R34981 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R34982 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.1255
R34983 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 0.0874565
R34984 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 0.063
R34985 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.063
R34986 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 0.063
R34987 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 0.063
R34988 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 0.0435206
R34989 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 0.0216397
R34990 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 0.0216397
R34991 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 0.0107679
R34992 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.0107679
R34993 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 316.762
R34994 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 168.108
R34995 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 150.293
R34996 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 150.273
R34997 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 73.6406
R34998 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 73.6304
R34999 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 60.4568
R35000 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 12.0358
R35001 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 1.19615
R35002 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.981478
R35003 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 0.788543
R35004 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.769522
R35005 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 0.682565
R35006 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.580578
R35007 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 0.55213
R35008 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 0.484875
R35009 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 0.470609
R35010 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.447191
R35011 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.428234
R35012 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.217464
R35013 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R35014 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R35015 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.1255
R35016 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 0.063
R35017 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 0.063
R35018 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.063
R35019 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 0.063
R35020 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 0.063
R35021 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 0.0216397
R35022 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.0216397
R35023 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 0.0107679
R35024 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.0107679
R35025 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 169.46
R35026 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 168.089
R35027 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 167.809
R35028 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 150.293
R35029 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 73.6304
R35030 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 60.4568
R35031 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 12.0358
R35032 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 11.4489
R35033 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.981478
R35034 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 0.788543
R35035 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.769522
R35036 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 0.720633
R35037 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 0.682565
R35038 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.580578
R35039 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 0.55213
R35040 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 0.470609
R35041 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.447191
R35042 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.428234
R35043 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.1255
R35044 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.1255
R35045 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 0.063
R35046 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 0.063
R35047 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.063
R35048 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 0.063
R35049 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 0.063
R35050 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 0.0435206
R35051 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 0.0107679
R35052 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.0107679
R35053 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 169.46
R35054 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 167.809
R35055 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 167.809
R35056 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 167.226
R35057 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 150.273
R35058 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 150.273
R35059 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 73.6406
R35060 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 73.6304
R35061 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 60.3943
R35062 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 12.3891
R35063 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 11.4489
R35064 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 1.68257
R35065 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 1.38365
R35066 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 1.19615
R35067 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 1.1717
R35068 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 1.08448
R35069 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.932141
R35070 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.720633
R35071 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 0.280391
R35072 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.217464
R35073 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R35074 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R35075 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.1255
R35076 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 0.0874565
R35077 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 0.063
R35078 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 0.063
R35079 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 0.063
R35080 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 0.063
R35081 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 0.0435206
R35082 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 0.0216397
R35083 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.0216397
R35084 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 0.0107679
R35085 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.0107679
R35086 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 169.46
R35087 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 167.809
R35088 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 167.809
R35089 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 167.227
R35090 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 150.293
R35091 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 150.273
R35092 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 73.6406
R35093 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 73.6304
R35094 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 60.3809
R35095 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 12.3891
R35096 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 11.4489
R35097 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 1.38365
R35098 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 1.19615
R35099 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 1.1717
R35100 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.848156
R35101 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 0.447191
R35102 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R35103 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 0.280391
R35104 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.217464
R35105 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.200143
R35106 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R35107 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R35108 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R35109 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R35110 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 0.0874565
R35111 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 0.063
R35112 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 0.063
R35113 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 0.063
R35114 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R35115 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 0.0107679
R35116 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0107679
R35117 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 169.46
R35118 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 167.809
R35119 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 167.809
R35120 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 167.226
R35121 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 150.273
R35122 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 150.273
R35123 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 73.6406
R35124 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 73.6304
R35125 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 60.3943
R35126 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 12.3891
R35127 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 11.4489
R35128 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 1.68257
R35129 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 1.38365
R35130 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 1.19615
R35131 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 1.1717
R35132 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 1.08448
R35133 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.932141
R35134 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.720633
R35135 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 0.280391
R35136 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.217464
R35137 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R35138 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R35139 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.1255
R35140 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 0.0874565
R35141 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 0.063
R35142 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 0.063
R35143 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 0.063
R35144 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 0.063
R35145 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 0.0435206
R35146 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 0.0216397
R35147 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.0216397
R35148 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 0.0107679
R35149 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.0107679
R35150 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 169.46
R35151 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 167.809
R35152 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 167.809
R35153 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 167.226
R35154 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 150.273
R35155 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 150.273
R35156 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 73.6406
R35157 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 73.6304
R35158 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 60.3943
R35159 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 12.3891
R35160 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 11.4489
R35161 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 1.68257
R35162 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 1.38365
R35163 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 1.19615
R35164 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 1.1717
R35165 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 1.08448
R35166 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.932141
R35167 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.720633
R35168 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 0.280391
R35169 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.217464
R35170 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R35171 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R35172 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.1255
R35173 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 0.0874565
R35174 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 0.063
R35175 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.063
R35176 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 0.063
R35177 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 0.063
R35178 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 0.0435206
R35179 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 0.0216397
R35180 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 0.0216397
R35181 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 0.0107679
R35182 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.0107679
R35183 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 169.46
R35184 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 167.809
R35185 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 167.809
R35186 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 167.227
R35187 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 150.293
R35188 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 150.273
R35189 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 73.6406
R35190 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 73.6304
R35191 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 60.3809
R35192 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 12.3891
R35193 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 11.4489
R35194 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 1.38365
R35195 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 1.19615
R35196 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 1.1717
R35197 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.848156
R35198 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 0.447191
R35199 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R35200 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 0.280391
R35201 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.217464
R35202 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.200143
R35203 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R35204 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R35205 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R35206 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R35207 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 0.0874565
R35208 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 0.063
R35209 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 0.063
R35210 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 0.063
R35211 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R35212 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 0.0107679
R35213 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0107679
R35214 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 169.46
R35215 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 167.809
R35216 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 167.809
R35217 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 167.226
R35218 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 150.273
R35219 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 150.273
R35220 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 73.6406
R35221 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 73.6304
R35222 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 60.4568
R35223 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 12.3891
R35224 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 11.4489
R35225 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.68257
R35226 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 1.38365
R35227 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 1.19615
R35228 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 1.1717
R35229 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.08448
R35230 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.932141
R35231 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.720633
R35232 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 0.280391
R35233 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.217464
R35234 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R35235 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R35236 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.1255
R35237 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 0.0874565
R35238 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 0.063
R35239 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 0.063
R35240 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 0.063
R35241 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 0.063
R35242 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 0.0435206
R35243 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 0.0216397
R35244 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.0216397
R35245 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 0.0107679
R35246 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.0107679
R35247 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 169.46
R35248 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 167.809
R35249 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 167.809
R35250 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 167.227
R35251 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 150.293
R35252 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 150.273
R35253 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 73.6406
R35254 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 73.6304
R35255 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 60.3809
R35256 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 12.3891
R35257 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 11.4489
R35258 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 1.38365
R35259 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 1.19615
R35260 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 1.1717
R35261 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.848156
R35262 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 0.447191
R35263 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.38637
R35264 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 0.280391
R35265 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 0.262643
R35266 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.217464
R35267 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.152844
R35268 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.149957
R35269 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.1255
R35270 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.1255
R35271 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 0.0874565
R35272 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 0.063
R35273 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 0.063
R35274 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.063
R35275 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.0454219
R35276 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 0.0107679
R35277 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.0107679
R35278 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t3 169.46
R35279 D_FlipFlop_0.3-input-nand_2.Vout.n9 D_FlipFlop_0.3-input-nand_2.Vout.t2 167.809
R35280 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.t0 167.809
R35281 D_FlipFlop_0.3-input-nand_2.Vout.t4 D_FlipFlop_0.3-input-nand_2.Vout.n11 167.227
R35282 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.t4 150.293
R35283 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.t7 150.273
R35284 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout.t5 73.6406
R35285 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout.t6 73.6304
R35286 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout.t1 60.3809
R35287 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n5 12.3891
R35288 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout.n9 11.4489
R35289 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout.n2 1.38365
R35290 D_FlipFlop_0.3-input-nand_2.Vout.n12 D_FlipFlop_0.3-input-nand_2.Vout.n1 1.19615
R35291 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout.n4 1.1717
R35292 D_FlipFlop_0.3-input-nand_2.Vout.n2 D_FlipFlop_0.3-input-nand_2.Vout 0.848156
R35293 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.Vout.n12 0.447191
R35294 D_FlipFlop_0.3-input-nand_2.Vout.n3 D_FlipFlop_0.3-input-nand_2.Vout 0.38637
R35295 D_FlipFlop_0.3-input-nand_2.Vout.n11 D_FlipFlop_0.3-input-nand_2.Vout.n10 0.280391
R35296 D_FlipFlop_0.3-input-nand_2.Vout.n10 D_FlipFlop_0.3-input-nand_2.Vout.n8 0.262643
R35297 D_FlipFlop_0.3-input-nand_2.Vout.n4 D_FlipFlop_0.3-input-nand_2.Vout 0.217464
R35298 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout 0.152844
R35299 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.149957
R35300 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R35301 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout 0.1255
R35302 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout.n7 0.0874565
R35303 D_FlipFlop_0.3-input-nand_2.Vout.n6 D_FlipFlop_0.3-input-nand_2.Vout.n3 0.063
R35304 D_FlipFlop_0.3-input-nand_2.Vout.n7 D_FlipFlop_0.3-input-nand_2.Vout.n6 0.063
R35305 D_FlipFlop_0.3-input-nand_2.Vout.n8 D_FlipFlop_0.3-input-nand_2.Vout 0.063
R35306 D_FlipFlop_0.3-input-nand_2.Vout.n5 D_FlipFlop_0.3-input-nand_2.Vout 0.0454219
R35307 D_FlipFlop_0.3-input-nand_2.Vout.n1 D_FlipFlop_0.3-input-nand_2.Vout.n0 0.0107679
R35308 D_FlipFlop_0.3-input-nand_2.Vout.n0 D_FlipFlop_0.3-input-nand_2.Vout 0.0107679
R35309 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 169.46
R35310 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 167.809
R35311 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 167.809
R35312 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 167.227
R35313 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 150.293
R35314 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 150.273
R35315 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 73.6406
R35316 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 73.6304
R35317 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 60.3809
R35318 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 12.3891
R35319 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 11.4489
R35320 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 1.38365
R35321 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 1.19615
R35322 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 1.1717
R35323 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.848156
R35324 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 0.447191
R35325 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.38637
R35326 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 0.280391
R35327 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 0.262643
R35328 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.217464
R35329 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.152844
R35330 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.149957
R35331 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.1255
R35332 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.1255
R35333 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 0.0874565
R35334 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 0.063
R35335 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 0.063
R35336 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.063
R35337 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.0454219
R35338 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 0.0107679
R35339 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.0107679
R35340 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 169.46
R35341 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 167.809
R35342 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 167.809
R35343 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 167.226
R35344 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 150.273
R35345 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 150.273
R35346 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 73.6406
R35347 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 73.6304
R35348 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 60.4568
R35349 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 12.3891
R35350 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 11.4489
R35351 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.68257
R35352 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 1.38365
R35353 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 1.19615
R35354 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 1.1717
R35355 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.08448
R35356 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.932141
R35357 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.720633
R35358 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 0.280391
R35359 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.217464
R35360 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R35361 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R35362 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.1255
R35363 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 0.0874565
R35364 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 0.063
R35365 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 0.063
R35366 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 0.063
R35367 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 0.063
R35368 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 0.0435206
R35369 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 0.0216397
R35370 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.0216397
R35371 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 0.0107679
R35372 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.0107679
R35373 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 169.46
R35374 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 167.809
R35375 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 167.809
R35376 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 167.227
R35377 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 150.293
R35378 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 150.273
R35379 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 73.6406
R35380 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 73.6304
R35381 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 60.3809
R35382 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 12.3891
R35383 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 11.4489
R35384 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 1.38365
R35385 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 1.19615
R35386 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 1.1717
R35387 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.848156
R35388 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 0.447191
R35389 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.38637
R35390 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 0.280391
R35391 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 0.262643
R35392 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.217464
R35393 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.152844
R35394 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.149957
R35395 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.1255
R35396 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.1255
R35397 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 0.0874565
R35398 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 0.063
R35399 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 0.063
R35400 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.063
R35401 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.0454219
R35402 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 0.0107679
R35403 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.0107679
R35404 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 169.46
R35405 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 167.809
R35406 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 167.809
R35407 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 167.226
R35408 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 150.273
R35409 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 150.273
R35410 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 73.6406
R35411 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 73.6304
R35412 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 60.4568
R35413 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 12.3891
R35414 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 11.4489
R35415 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.68257
R35416 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 1.38365
R35417 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 1.19615
R35418 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 1.1717
R35419 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.08448
R35420 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.932141
R35421 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.720633
R35422 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 0.280391
R35423 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.217464
R35424 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R35425 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R35426 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.1255
R35427 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 0.0874565
R35428 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 0.063
R35429 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 0.063
R35430 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 0.063
R35431 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 0.063
R35432 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 0.0435206
R35433 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 0.0216397
R35434 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.0216397
R35435 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 0.0107679
R35436 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.0107679
R35437 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 316.762
R35438 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 168.108
R35439 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 150.293
R35440 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 150.273
R35441 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 73.6406
R35442 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 73.6304
R35443 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 60.3943
R35444 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 12.0358
R35445 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 1.19615
R35446 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.981478
R35447 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 0.788543
R35448 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.769522
R35449 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 0.682565
R35450 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.580578
R35451 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 0.55213
R35452 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 0.484875
R35453 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 0.470609
R35454 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.447191
R35455 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.428234
R35456 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.217464
R35457 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R35458 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R35459 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.1255
R35460 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 0.063
R35461 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 0.063
R35462 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.063
R35463 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 0.063
R35464 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 0.063
R35465 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 0.0216397
R35466 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.0216397
R35467 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 0.0107679
R35468 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.0107679
R35469 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 169.46
R35470 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 167.809
R35471 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 167.809
R35472 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 167.227
R35473 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 150.293
R35474 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 150.273
R35475 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 73.6406
R35476 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 73.6304
R35477 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 60.3809
R35478 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 12.3891
R35479 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 11.4489
R35480 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 1.38365
R35481 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 1.19615
R35482 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 1.1717
R35483 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.848156
R35484 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 0.447191
R35485 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R35486 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 0.280391
R35487 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.217464
R35488 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.200143
R35489 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R35490 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R35491 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R35492 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R35493 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 0.0874565
R35494 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 0.063
R35495 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 0.063
R35496 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 0.063
R35497 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R35498 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 0.0107679
R35499 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0107679
R35500 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C.t3 169.46
R35501 D_FlipFlop_5.3-input-nand_2.C.n4 D_FlipFlop_5.3-input-nand_2.C.t2 167.809
R35502 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C.t1 167.809
R35503 D_FlipFlop_5.3-input-nand_2.C.n3 D_FlipFlop_5.3-input-nand_2.C.t6 167.226
R35504 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.t7 150.273
R35505 D_FlipFlop_5.3-input-nand_2.C.t6 D_FlipFlop_5.3-input-nand_2.C.n2 150.273
R35506 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C.t5 73.6406
R35507 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C.t4 73.6304
R35508 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.t0 60.4568
R35509 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n11 12.3891
R35510 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C.n4 11.4489
R35511 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C 1.68257
R35512 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C.n13 1.38365
R35513 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C.n0 1.19615
R35514 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C.n9 1.1717
R35515 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C 1.08448
R35516 D_FlipFlop_5.3-input-nand_2.C.n10 D_FlipFlop_5.3-input-nand_2.C 0.932141
R35517 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C 0.720633
R35518 D_FlipFlop_5.3-input-nand_2.C.n5 D_FlipFlop_5.3-input-nand_2.C.n3 0.280391
R35519 D_FlipFlop_5.3-input-nand_2.C.n0 D_FlipFlop_5.3-input-nand_2.C 0.217464
R35520 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C 0.1255
R35521 D_FlipFlop_5.3-input-nand_2.C.n1 D_FlipFlop_5.3-input-nand_2.C 0.1255
R35522 D_FlipFlop_5.3-input-nand_2.C.n14 D_FlipFlop_5.3-input-nand_2.C 0.1255
R35523 D_FlipFlop_5.3-input-nand_2.C.n7 D_FlipFlop_5.3-input-nand_2.C.n6 0.0874565
R35524 D_FlipFlop_5.3-input-nand_2.C.n11 D_FlipFlop_5.3-input-nand_2.C.n10 0.063
R35525 D_FlipFlop_5.3-input-nand_2.C.n12 D_FlipFlop_5.3-input-nand_2.C.n7 0.063
R35526 D_FlipFlop_5.3-input-nand_2.C.n13 D_FlipFlop_5.3-input-nand_2.C.n12 0.063
R35527 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.C.n14 0.063
R35528 D_FlipFlop_5.3-input-nand_2.C.n6 D_FlipFlop_5.3-input-nand_2.C.n5 0.0435206
R35529 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C.n1 0.0216397
R35530 D_FlipFlop_5.3-input-nand_2.C.n2 D_FlipFlop_5.3-input-nand_2.C 0.0216397
R35531 D_FlipFlop_5.3-input-nand_2.C.n9 D_FlipFlop_5.3-input-nand_2.C.n8 0.0107679
R35532 D_FlipFlop_5.3-input-nand_2.C.n8 D_FlipFlop_5.3-input-nand_2.C 0.0107679
R35533 Q6.n2 Q6.t1 169.46
R35534 Q6.n4 Q6.t2 167.809
R35535 Q6.n2 Q6.t0 167.809
R35536 Q6 Q6.t6 158.585
R35537 Q6 Q6.t7 154.823
R35538 Q6.n14 Q6.t9 150.869
R35539 Q6.t7 Q6.n15 150.869
R35540 Q6.t6 Q6.n9 150.293
R35541 Q6.n16 Q6.n13 137.644
R35542 Q6.n13 Q6 85.5731
R35543 Q6.n15 Q6.t4 74.1352
R35544 Q6.n14 Q6.t5 74.1352
R35545 Q6.n7 Q6.t8 73.6304
R35546 Q6.n0 Q6.t3 60.3809
R35547 Q6.n3 Q6.n2 11.4489
R35548 Q6.n5 Q6.n4 8.21389
R35549 Q6.n13 Q6.n12 3.473
R35550 Q6.n15 Q6.n14 1.66898
R35551 Q6.n1 Q6.n0 1.64452
R35552 Q6.n9 Q6.n8 1.19615
R35553 Q6.n0 Q6 0.848156
R35554 Q6.n9 Q6 0.447191
R35555 Q6.n5 Q6 0.39003
R35556 Q6.n4 Q6.n3 0.280391
R35557 Q6.n3 Q6.n1 0.262643
R35558 Q6.n6 Q6 0.2167
R35559 Q6.n6 Q6.n5 0.212783
R35560 Q6.n11 Q6.n10 0.161083
R35561 Q6.n11 Q6 0.150045
R35562 Q6.n1 Q6 0.1255
R35563 Q6.n8 Q6 0.1255
R35564 Q6.n14 Q6 0.063
R35565 Q6.n1 Q6 0.063
R35566 Q6.n12 Q6.n6 0.024
R35567 Q6.n12 Q6.n11 0.024
R35568 Q6 Q6.n16 0.0168043
R35569 Q6.n16 Q6 0.0122188
R35570 Q6.n8 Q6.n7 0.0107679
R35571 Q6.n7 Q6 0.0107679
R35572 Q6.n10 Q6 0.00441667
R35573 Q6.n10 Q6 0.00406061
R35574 CDAC8_0.switch_2.Z.n0 CDAC8_0.switch_2.Z.t1 168.548
R35575 CDAC8_0.switch_2.Z.n0 CDAC8_0.switch_2.Z.t2 168.548
R35576 CDAC8_0.switch_2.Z.n4 CDAC8_0.switch_2.Z.t3 60.321
R35577 CDAC8_0.switch_2.Z.n4 CDAC8_0.switch_2.Z.t0 60.321
R35578 CDAC8_0.switch_2.Z.n2 CDAC8_0.switch_2.Z.n1 11.3205
R35579 CDAC8_0.switch_2.Z.n1 CDAC8_0.switch_2.Z.t5 3.64361
R35580 CDAC8_0.switch_2.Z.n1 CDAC8_0.switch_2.Z.t4 3.16265
R35581 CDAC8_0.switch_2.Z.n5 CDAC8_0.switch_2.Z.n3 1.59289
R35582 CDAC8_0.switch_2.Z CDAC8_0.switch_2.Z.n5 0.259656
R35583 CDAC8_0.switch_2.Z.n3 CDAC8_0.switch_2.Z 0.17713
R35584 CDAC8_0.switch_2.Z.n3 CDAC8_0.switch_2.Z.n2 0.063
R35585 CDAC8_0.switch_2.Z.n0 CDAC8_0.switch_2.Z 0.0454219
R35586 CDAC8_0.switch_2.Z.n2 CDAC8_0.switch_2.Z.n0 0.0200312
R35587 CDAC8_0.switch_2.Z.n5 CDAC8_0.switch_2.Z.n4 0.0188121
R35588 Q3.n5 Q3.t0 169.46
R35589 Q3.n7 Q3.t2 167.809
R35590 Q3.n5 Q3.t3 167.809
R35591 Q3.n11 Q3.t5 155.12
R35592 Q3.n14 Q3.t6 150.869
R35593 Q3.n13 Q3.t7 150.869
R35594 Q3.t5 Q3.n2 150.293
R35595 Q3.n15 Q3.n12 137.644
R35596 Q3 Q3.t9 78.1811
R35597 Q3.n13 Q3.t4 74.1352
R35598 Q3.t9 Q3.n14 74.1352
R35599 Q3.n0 Q3.t8 73.6304
R35600 Q3.n3 Q3.t1 60.3809
R35601 Q3.n12 Q3 36.8166
R35602 Q3.n6 Q3.n5 11.4489
R35603 Q3.n8 Q3.n7 8.21389
R35604 Q3.n11 Q3.n10 1.6986
R35605 Q3.n14 Q3.n13 1.66898
R35606 Q3.n4 Q3.n3 1.64452
R35607 Q3.n2 Q3.n1 1.19615
R35608 Q3.n3 Q3 0.848156
R35609 Q3.n2 Q3 0.447191
R35610 Q3.n8 Q3 0.39003
R35611 Q3.n9 Q3.n8 0.3483
R35612 Q3.n7 Q3.n6 0.280391
R35613 Q3.n6 Q3.n4 0.262643
R35614 Q3.n4 Q3 0.1255
R35615 Q3.n1 Q3 0.1255
R35616 Q3.n9 Q3 0.0811833
R35617 Q3.n13 Q3 0.063
R35618 Q3.n4 Q3 0.063
R35619 Q3.n10 Q3.n9 0.0491718
R35620 Q3.n12 Q3.n11 0.0273895
R35621 Q3.n10 Q3 0.025816
R35622 Q3 Q3.n15 0.0168043
R35623 Q3.n15 Q3 0.0122188
R35624 Q3.n1 Q3.n0 0.0107679
R35625 Q3.n0 Q3 0.0107679
R35626 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.t3 168.609
R35627 CDAC8_0.switch_5.Z CDAC8_0.switch_5.Z.t0 168.565
R35628 CDAC8_0.switch_5.Z.n0 CDAC8_0.switch_5.Z.t1 60.321
R35629 CDAC8_0.switch_5.Z.n0 CDAC8_0.switch_5.Z.t2 60.321
R35630 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.n10 11.3205
R35631 CDAC8_0.switch_5.Z.n6 CDAC8_0.switch_5.Z.n5 5.49497
R35632 CDAC8_0.switch_5.Z.n10 CDAC8_0.switch_5.Z.n2 2.98587
R35633 CDAC8_0.switch_5.Z.n10 CDAC8_0.switch_5.Z.n9 2.5049
R35634 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z.n1 1.60376
R35635 CDAC8_0.switch_5.Z.n9 CDAC8_0.switch_5.Z.t10 0.726216
R35636 CDAC8_0.switch_5.Z.n2 CDAC8_0.switch_5.Z.t6 0.726216
R35637 CDAC8_0.switch_5.Z.n5 CDAC8_0.switch_5.Z.t9 0.658247
R35638 CDAC8_0.switch_5.Z.n6 CDAC8_0.switch_5.Z.t5 0.658247
R35639 CDAC8_0.switch_5.Z.n7 CDAC8_0.switch_5.Z.t8 0.611304
R35640 CDAC8_0.switch_5.Z.n8 CDAC8_0.switch_5.Z.t11 0.611304
R35641 CDAC8_0.switch_5.Z.n4 CDAC8_0.switch_5.Z.t4 0.611304
R35642 CDAC8_0.switch_5.Z.n3 CDAC8_0.switch_5.Z.t7 0.611304
R35643 CDAC8_0.switch_5.Z.n1 CDAC8_0.switch_5.Z 0.259656
R35644 CDAC8_0.switch_5.Z.n11 CDAC8_0.switch_5.Z 0.166261
R35645 CDAC8_0.switch_5.Z.n8 CDAC8_0.switch_5.Z.n7 0.162356
R35646 CDAC8_0.switch_5.Z.n4 CDAC8_0.switch_5.Z.n3 0.162356
R35647 CDAC8_0.switch_5.Z.n7 CDAC8_0.switch_5.Z.n6 0.115412
R35648 CDAC8_0.switch_5.Z.n5 CDAC8_0.switch_5.Z.n4 0.115412
R35649 CDAC8_0.switch_5.Z.n9 CDAC8_0.switch_5.Z.n8 0.0474438
R35650 CDAC8_0.switch_5.Z.n3 CDAC8_0.switch_5.Z.n2 0.0474438
R35651 CDAC8_0.switch_5.Z CDAC8_0.switch_5.Z.n11 0.0454219
R35652 CDAC8_0.switch_5.Z.n1 CDAC8_0.switch_5.Z.n0 0.0188121
R35653 Nand_Gate_5.Vout.n10 Nand_Gate_5.Vout.t0 179.256
R35654 Nand_Gate_5.Vout.n10 Nand_Gate_5.Vout.t1 168.089
R35655 Nand_Gate_5.Vout.n2 Nand_Gate_5.Vout.t3 150.293
R35656 Nand_Gate_5.Vout.n4 Nand_Gate_5.Vout.t4 73.6304
R35657 Nand_Gate_5.Vout Nand_Gate_5.Vout.t2 60.3943
R35658 Nand_Gate_5.Vout.n8 Nand_Gate_5.Vout.n7 35.6663
R35659 Nand_Gate_5.Vout.n9 Nand_Gate_5.Vout 0.981478
R35660 Nand_Gate_5.Vout.n11 Nand_Gate_5.Vout.n9 0.788543
R35661 Nand_Gate_5.Vout.n3 Nand_Gate_5.Vout 0.769522
R35662 Nand_Gate_5.Vout Nand_Gate_5.Vout.n11 0.720633
R35663 Nand_Gate_5.Vout.n1 Nand_Gate_5.Vout.n0 0.682565
R35664 Nand_Gate_5.Vout.n1 Nand_Gate_5.Vout 0.580578
R35665 Nand_Gate_5.Vout.n3 Nand_Gate_5.Vout.n2 0.55213
R35666 Nand_Gate_5.Vout.n6 Nand_Gate_5.Vout.n5 0.470609
R35667 Nand_Gate_5.Vout.n2 Nand_Gate_5.Vout 0.447191
R35668 Nand_Gate_5.Vout.n6 Nand_Gate_5.Vout 0.428234
R35669 Nand_Gate_5.Vout.n5 Nand_Gate_5.Vout 0.1255
R35670 Nand_Gate_5.Vout.n0 Nand_Gate_5.Vout 0.1255
R35671 Nand_Gate_5.Vout.n7 Nand_Gate_5.Vout.n3 0.063
R35672 Nand_Gate_5.Vout.n7 Nand_Gate_5.Vout.n6 0.063
R35673 Nand_Gate_5.Vout.n0 Nand_Gate_5.Vout 0.063
R35674 Nand_Gate_5.Vout.n9 Nand_Gate_5.Vout.n8 0.063
R35675 Nand_Gate_5.Vout.n8 Nand_Gate_5.Vout.n1 0.063
R35676 Nand_Gate_5.Vout.n11 Nand_Gate_5.Vout.n10 0.0435206
R35677 Nand_Gate_5.Vout.n5 Nand_Gate_5.Vout.n4 0.0107679
R35678 Nand_Gate_5.Vout.n4 Nand_Gate_5.Vout 0.0107679
R35679 Nand_Gate_6.B.n51 Nand_Gate_6.B.t0 169.46
R35680 Nand_Gate_6.B.n51 Nand_Gate_6.B.t1 167.809
R35681 Nand_Gate_6.B.n53 Nand_Gate_6.B.t3 167.809
R35682 Nand_Gate_6.B Nand_Gate_6.B.t5 158.585
R35683 Nand_Gate_6.B Nand_Gate_6.B.t9 158.581
R35684 Nand_Gate_6.B.n42 Nand_Gate_6.B.t8 150.293
R35685 Nand_Gate_6.B.t9 Nand_Gate_6.B.n38 150.293
R35686 Nand_Gate_6.B.t5 Nand_Gate_6.B.n2 150.293
R35687 Nand_Gate_6.B.n29 Nand_Gate_6.B.t7 150.273
R35688 Nand_Gate_6.B.n23 Nand_Gate_6.B.t12 150.273
R35689 Nand_Gate_6.B.n14 Nand_Gate_6.B.t11 150.273
R35690 Nand_Gate_6.B.n8 Nand_Gate_6.B.t17 150.273
R35691 Nand_Gate_6.B.n27 Nand_Gate_6.B.t13 73.6406
R35692 Nand_Gate_6.B.n21 Nand_Gate_6.B.t6 73.6406
R35693 Nand_Gate_6.B.n12 Nand_Gate_6.B.t15 73.6406
R35694 Nand_Gate_6.B.n6 Nand_Gate_6.B.t10 73.6406
R35695 Nand_Gate_6.B.n43 Nand_Gate_6.B.t14 73.6304
R35696 Nand_Gate_6.B.n36 Nand_Gate_6.B.t4 73.6304
R35697 Nand_Gate_6.B.n0 Nand_Gate_6.B.t16 73.6304
R35698 Nand_Gate_6.B.n4 Nand_Gate_6.B.t2 60.3809
R35699 Nand_Gate_6.B.n44 Nand_Gate_6.B.n41 47.1622
R35700 Nand_Gate_6.B.n44 Nand_Gate_6.B.n43 34.7148
R35701 Nand_Gate_6.B.n33 Nand_Gate_6.B.n26 15.5222
R35702 Nand_Gate_6.B.n52 Nand_Gate_6.B.n51 11.4489
R35703 Nand_Gate_6.B.n34 Nand_Gate_6.B.n33 8.26552
R35704 Nand_Gate_6.B.n54 Nand_Gate_6.B.n53 8.21389
R35705 Nand_Gate_6.B.n18 Nand_Gate_6.B.n11 8.1418
R35706 Nand_Gate_6.B.n47 Nand_Gate_6.B.n46 5.61191
R35707 Nand_Gate_6.B.n47 Nand_Gate_6.B 5.35402
R35708 Nand_Gate_6.B.n45 Nand_Gate_6.B.n44 4.81893
R35709 Nand_Gate_6.B.n48 Nand_Gate_6.B.n47 4.563
R35710 Nand_Gate_6.B.n33 Nand_Gate_6.B.n32 4.5005
R35711 Nand_Gate_6.B.n18 Nand_Gate_6.B.n17 4.5005
R35712 Nand_Gate_6.B.n46 Nand_Gate_6.B 1.83746
R35713 Nand_Gate_6.B.n20 Nand_Gate_6.B.n19 1.62007
R35714 Nand_Gate_6.B.n38 Nand_Gate_6.B.n37 1.19615
R35715 Nand_Gate_6.B.n2 Nand_Gate_6.B.n1 1.19615
R35716 Nand_Gate_6.B.n43 Nand_Gate_6.B.n42 1.1717
R35717 Nand_Gate_6.B.n5 Nand_Gate_6.B 1.08746
R35718 Nand_Gate_6.B.n20 Nand_Gate_6.B 1.01739
R35719 Nand_Gate_6.B.n13 Nand_Gate_6.B 0.851043
R35720 Nand_Gate_6.B.n7 Nand_Gate_6.B 0.851043
R35721 Nand_Gate_6.B.n4 Nand_Gate_6.B 0.848156
R35722 Nand_Gate_6.B.n28 Nand_Gate_6.B.n27 0.796696
R35723 Nand_Gate_6.B.n22 Nand_Gate_6.B.n21 0.796696
R35724 Nand_Gate_6.B.n50 Nand_Gate_6.B.n49 0.788543
R35725 Nand_Gate_6.B.n34 Nand_Gate_6.B 0.716182
R35726 Nand_Gate_6.B.n5 Nand_Gate_6.B.n4 0.682565
R35727 Nand_Gate_6.B.n49 Nand_Gate_6.B 0.65675
R35728 Nand_Gate_6.B.n16 Nand_Gate_6.B.n15 0.55213
R35729 Nand_Gate_6.B.n10 Nand_Gate_6.B.n9 0.55213
R35730 Nand_Gate_6.B.n28 Nand_Gate_6.B 0.524957
R35731 Nand_Gate_6.B.n22 Nand_Gate_6.B 0.524957
R35732 Nand_Gate_6.B.n16 Nand_Gate_6.B 0.486828
R35733 Nand_Gate_6.B.n10 Nand_Gate_6.B 0.486828
R35734 Nand_Gate_6.B.n35 Nand_Gate_6.B 0.4846
R35735 Nand_Gate_6.B.n13 Nand_Gate_6.B.n12 0.470609
R35736 Nand_Gate_6.B.n7 Nand_Gate_6.B.n6 0.470609
R35737 Nand_Gate_6.B.n42 Nand_Gate_6.B 0.447191
R35738 Nand_Gate_6.B.n38 Nand_Gate_6.B 0.447191
R35739 Nand_Gate_6.B.n2 Nand_Gate_6.B 0.447191
R35740 Nand_Gate_6.B.n54 Nand_Gate_6.B.n3 0.425067
R35741 Nand_Gate_6.B.n40 Nand_Gate_6.B.n39 0.42115
R35742 Nand_Gate_6.B Nand_Gate_6.B.n54 0.39003
R35743 Nand_Gate_6.B.n40 Nand_Gate_6.B 0.335684
R35744 Nand_Gate_6.B.n35 Nand_Gate_6.B.n34 0.30365
R35745 Nand_Gate_6.B.n53 Nand_Gate_6.B.n52 0.280391
R35746 Nand_Gate_6.B.n52 Nand_Gate_6.B.n50 0.262643
R35747 Nand_Gate_6.B.n31 Nand_Gate_6.B 0.252453
R35748 Nand_Gate_6.B.n25 Nand_Gate_6.B 0.252453
R35749 Nand_Gate_6.B.n31 Nand_Gate_6.B.n30 0.226043
R35750 Nand_Gate_6.B.n25 Nand_Gate_6.B.n24 0.226043
R35751 Nand_Gate_6.B.n27 Nand_Gate_6.B 0.217464
R35752 Nand_Gate_6.B.n21 Nand_Gate_6.B 0.217464
R35753 Nand_Gate_6.B.n12 Nand_Gate_6.B 0.217464
R35754 Nand_Gate_6.B.n6 Nand_Gate_6.B 0.217464
R35755 Nand_Gate_6.B.n43 Nand_Gate_6.B 0.149957
R35756 Nand_Gate_6.B.n30 Nand_Gate_6.B 0.1255
R35757 Nand_Gate_6.B.n24 Nand_Gate_6.B 0.1255
R35758 Nand_Gate_6.B.n37 Nand_Gate_6.B 0.1255
R35759 Nand_Gate_6.B.n15 Nand_Gate_6.B 0.1255
R35760 Nand_Gate_6.B.n9 Nand_Gate_6.B 0.1255
R35761 Nand_Gate_6.B.n50 Nand_Gate_6.B 0.1255
R35762 Nand_Gate_6.B.n1 Nand_Gate_6.B 0.1255
R35763 Nand_Gate_6.B.n32 Nand_Gate_6.B.n28 0.063
R35764 Nand_Gate_6.B.n32 Nand_Gate_6.B.n31 0.063
R35765 Nand_Gate_6.B.n26 Nand_Gate_6.B.n22 0.063
R35766 Nand_Gate_6.B.n26 Nand_Gate_6.B.n25 0.063
R35767 Nand_Gate_6.B.n17 Nand_Gate_6.B.n13 0.063
R35768 Nand_Gate_6.B.n17 Nand_Gate_6.B.n16 0.063
R35769 Nand_Gate_6.B.n11 Nand_Gate_6.B.n7 0.063
R35770 Nand_Gate_6.B.n11 Nand_Gate_6.B.n10 0.063
R35771 Nand_Gate_6.B.n46 Nand_Gate_6.B.n45 0.063
R35772 Nand_Gate_6.B.n45 Nand_Gate_6.B.n20 0.063
R35773 Nand_Gate_6.B.n48 Nand_Gate_6.B.n5 0.063
R35774 Nand_Gate_6.B.n49 Nand_Gate_6.B.n48 0.063
R35775 Nand_Gate_6.B.n50 Nand_Gate_6.B 0.063
R35776 Nand_Gate_6.B Nand_Gate_6.B.n18 0.0512812
R35777 Nand_Gate_6.B.n43 Nand_Gate_6.B 0.0454219
R35778 Nand_Gate_6.B.n41 Nand_Gate_6.B.n35 0.024
R35779 Nand_Gate_6.B.n41 Nand_Gate_6.B.n40 0.024
R35780 Nand_Gate_6.B.n30 Nand_Gate_6.B.n29 0.0216397
R35781 Nand_Gate_6.B.n29 Nand_Gate_6.B 0.0216397
R35782 Nand_Gate_6.B.n24 Nand_Gate_6.B.n23 0.0216397
R35783 Nand_Gate_6.B.n23 Nand_Gate_6.B 0.0216397
R35784 Nand_Gate_6.B.n15 Nand_Gate_6.B.n14 0.0216397
R35785 Nand_Gate_6.B.n14 Nand_Gate_6.B 0.0216397
R35786 Nand_Gate_6.B.n9 Nand_Gate_6.B.n8 0.0216397
R35787 Nand_Gate_6.B.n8 Nand_Gate_6.B 0.0216397
R35788 Nand_Gate_6.B.n19 Nand_Gate_6.B 0.0168043
R35789 Nand_Gate_6.B.n19 Nand_Gate_6.B 0.0122188
R35790 Nand_Gate_6.B.n37 Nand_Gate_6.B.n36 0.0107679
R35791 Nand_Gate_6.B.n36 Nand_Gate_6.B 0.0107679
R35792 Nand_Gate_6.B.n1 Nand_Gate_6.B.n0 0.0107679
R35793 Nand_Gate_6.B.n0 Nand_Gate_6.B 0.0107679
R35794 Nand_Gate_6.B.n39 Nand_Gate_6.B 0.00441667
R35795 Nand_Gate_6.B.n3 Nand_Gate_6.B 0.00441667
R35796 Nand_Gate_6.B.n39 Nand_Gate_6.B 0.00406061
R35797 Nand_Gate_6.B.n3 Nand_Gate_6.B 0.00406061
R35798 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 169.46
R35799 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 168.089
R35800 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 167.809
R35801 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 150.273
R35802 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 73.6406
R35803 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 60.3809
R35804 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 12.0358
R35805 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 11.4489
R35806 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 1.08746
R35807 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.851043
R35808 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.848156
R35809 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 0.788543
R35810 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 0.682565
R35811 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.65675
R35812 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 0.55213
R35813 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.486828
R35814 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 0.470609
R35815 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 0.262643
R35816 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.217464
R35817 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.1255
R35818 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.1255
R35819 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 0.063
R35820 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 0.063
R35821 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 0.063
R35822 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 0.063
R35823 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 0.063
R35824 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 0.0216397
R35825 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0216397
R35826 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 179.256
R35827 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 168.089
R35828 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 150.293
R35829 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 73.6304
R35830 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 60.3943
R35831 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 12.0358
R35832 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.981478
R35833 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 0.788543
R35834 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.769522
R35835 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.720633
R35836 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 0.682565
R35837 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.580578
R35838 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 0.55213
R35839 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 0.470609
R35840 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.447191
R35841 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.428234
R35842 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1255
R35843 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1255
R35844 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 0.063
R35845 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 0.063
R35846 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 0.063
R35847 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 0.063
R35848 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 0.063
R35849 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 0.0435206
R35850 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 0.0107679
R35851 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.0107679
R35852 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 316.762
R35853 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 168.108
R35854 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 150.293
R35855 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 150.273
R35856 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 73.6406
R35857 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 73.6304
R35858 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 60.3943
R35859 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 12.0358
R35860 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 1.19615
R35861 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.981478
R35862 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 0.788543
R35863 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.769522
R35864 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 0.682565
R35865 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.580578
R35866 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 0.55213
R35867 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 0.484875
R35868 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 0.470609
R35869 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.447191
R35870 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.428234
R35871 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.217464
R35872 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R35873 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R35874 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.1255
R35875 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 0.063
R35876 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 0.063
R35877 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.063
R35878 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 0.063
R35879 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 0.063
R35880 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 0.0216397
R35881 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.0216397
R35882 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 0.0107679
R35883 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.0107679
R35884 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 316.762
R35885 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 168.108
R35886 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 150.293
R35887 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 150.273
R35888 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 73.6406
R35889 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 73.6304
R35890 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 60.4568
R35891 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 12.0358
R35892 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 1.19615
R35893 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.981478
R35894 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 0.788543
R35895 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.769522
R35896 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 0.682565
R35897 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.580578
R35898 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 0.55213
R35899 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 0.484875
R35900 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 0.470609
R35901 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.447191
R35902 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.428234
R35903 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.217464
R35904 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R35905 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R35906 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.1255
R35907 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 0.063
R35908 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 0.063
R35909 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.063
R35910 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 0.063
R35911 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 0.063
R35912 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 0.0216397
R35913 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.0216397
R35914 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 0.0107679
R35915 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.0107679
R35916 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 179.256
R35917 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 168.089
R35918 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 150.293
R35919 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 73.6304
R35920 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 60.4568
R35921 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 12.0358
R35922 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.981478
R35923 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 0.788543
R35924 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.769522
R35925 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 0.720633
R35926 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 0.682565
R35927 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.580578
R35928 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 0.55213
R35929 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 0.470609
R35930 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.447191
R35931 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.428234
R35932 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1255
R35933 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1255
R35934 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 0.063
R35935 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 0.063
R35936 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.063
R35937 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 0.063
R35938 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 0.063
R35939 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 0.0435206
R35940 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 0.0107679
R35941 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.0107679
R35942 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 169.46
R35943 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 168.089
R35944 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 167.809
R35945 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 150.273
R35946 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 73.6406
R35947 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 60.3809
R35948 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 12.0358
R35949 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 11.4489
R35950 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 1.08746
R35951 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.851043
R35952 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.848156
R35953 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 0.788543
R35954 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 0.682565
R35955 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.65675
R35956 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 0.55213
R35957 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.486828
R35958 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 0.470609
R35959 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 0.262643
R35960 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.217464
R35961 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.1255
R35962 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.1255
R35963 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 0.063
R35964 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 0.063
R35965 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 0.063
R35966 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 0.063
R35967 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 0.063
R35968 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 0.0216397
R35969 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.0216397
R35970 Nand_Gate_5.A.n55 Nand_Gate_5.A.t0 169.46
R35971 Nand_Gate_5.A.n55 Nand_Gate_5.A.t1 167.809
R35972 Nand_Gate_5.A.n57 Nand_Gate_5.A.t2 167.809
R35973 Nand_Gate_5.A Nand_Gate_5.A.t7 158.585
R35974 Nand_Gate_5.A Nand_Gate_5.A.t17 158.581
R35975 Nand_Gate_5.A.n42 Nand_Gate_5.A.t9 150.293
R35976 Nand_Gate_5.A.t17 Nand_Gate_5.A.n38 150.293
R35977 Nand_Gate_5.A.t7 Nand_Gate_5.A.n2 150.293
R35978 Nand_Gate_5.A.n29 Nand_Gate_5.A.t14 150.273
R35979 Nand_Gate_5.A.n23 Nand_Gate_5.A.t5 150.273
R35980 Nand_Gate_5.A.n14 Nand_Gate_5.A.t11 150.273
R35981 Nand_Gate_5.A.n8 Nand_Gate_5.A.t12 150.273
R35982 Nand_Gate_5.A.n27 Nand_Gate_5.A.t6 73.6406
R35983 Nand_Gate_5.A.n21 Nand_Gate_5.A.t15 73.6406
R35984 Nand_Gate_5.A.n12 Nand_Gate_5.A.t13 73.6406
R35985 Nand_Gate_5.A.n6 Nand_Gate_5.A.t8 73.6406
R35986 Nand_Gate_5.A.n44 Nand_Gate_5.A.t4 73.6304
R35987 Nand_Gate_5.A.n36 Nand_Gate_5.A.t10 73.6304
R35988 Nand_Gate_5.A.n0 Nand_Gate_5.A.t16 73.6304
R35989 Nand_Gate_5.A.n4 Nand_Gate_5.A.t3 60.3809
R35990 Nand_Gate_5.A.n48 Nand_Gate_5.A.n41 25.1004
R35991 Nand_Gate_5.A.n33 Nand_Gate_5.A.n26 15.5222
R35992 Nand_Gate_5.A.n56 Nand_Gate_5.A.n55 11.4489
R35993 Nand_Gate_5.A.n48 Nand_Gate_5.A.n47 9.57083
R35994 Nand_Gate_5.A.n34 Nand_Gate_5.A.n33 8.26552
R35995 Nand_Gate_5.A.n58 Nand_Gate_5.A.n57 8.21389
R35996 Nand_Gate_5.A.n18 Nand_Gate_5.A.n11 8.1418
R35997 Nand_Gate_5.A.n49 Nand_Gate_5.A.n48 6.58222
R35998 Nand_Gate_5.A.n20 Nand_Gate_5.A.n19 6.47604
R35999 Nand_Gate_5.A.n19 Nand_Gate_5.A 5.35402
R36000 Nand_Gate_5.A.n52 Nand_Gate_5.A 4.55128
R36001 Nand_Gate_5.A.n33 Nand_Gate_5.A.n32 4.5005
R36002 Nand_Gate_5.A.n18 Nand_Gate_5.A.n17 4.5005
R36003 Nand_Gate_5.A.n38 Nand_Gate_5.A.n37 1.19615
R36004 Nand_Gate_5.A.n2 Nand_Gate_5.A.n1 1.19615
R36005 Nand_Gate_5.A.n5 Nand_Gate_5.A 1.08746
R36006 Nand_Gate_5.A.n20 Nand_Gate_5.A 0.973326
R36007 Nand_Gate_5.A.n13 Nand_Gate_5.A 0.851043
R36008 Nand_Gate_5.A.n7 Nand_Gate_5.A 0.851043
R36009 Nand_Gate_5.A.n4 Nand_Gate_5.A 0.848156
R36010 Nand_Gate_5.A.n28 Nand_Gate_5.A.n27 0.796696
R36011 Nand_Gate_5.A.n22 Nand_Gate_5.A.n21 0.796696
R36012 Nand_Gate_5.A.n54 Nand_Gate_5.A.n53 0.788543
R36013 Nand_Gate_5.A.n43 Nand_Gate_5.A 0.769522
R36014 Nand_Gate_5.A.n51 Nand_Gate_5.A.n50 0.755935
R36015 Nand_Gate_5.A.n34 Nand_Gate_5.A 0.716182
R36016 Nand_Gate_5.A.n5 Nand_Gate_5.A.n4 0.682565
R36017 Nand_Gate_5.A.n53 Nand_Gate_5.A 0.65675
R36018 Nand_Gate_5.A.n43 Nand_Gate_5.A.n42 0.55213
R36019 Nand_Gate_5.A.n16 Nand_Gate_5.A.n15 0.55213
R36020 Nand_Gate_5.A.n10 Nand_Gate_5.A.n9 0.55213
R36021 Nand_Gate_5.A.n35 Nand_Gate_5.A.n34 0.546483
R36022 Nand_Gate_5.A.n28 Nand_Gate_5.A 0.524957
R36023 Nand_Gate_5.A.n22 Nand_Gate_5.A 0.524957
R36024 Nand_Gate_5.A.n16 Nand_Gate_5.A 0.486828
R36025 Nand_Gate_5.A.n10 Nand_Gate_5.A 0.486828
R36026 Nand_Gate_5.A.n50 Nand_Gate_5.A 0.48023
R36027 Nand_Gate_5.A.n46 Nand_Gate_5.A.n45 0.470609
R36028 Nand_Gate_5.A.n13 Nand_Gate_5.A.n12 0.470609
R36029 Nand_Gate_5.A.n7 Nand_Gate_5.A.n6 0.470609
R36030 Nand_Gate_5.A.n42 Nand_Gate_5.A 0.447191
R36031 Nand_Gate_5.A.n38 Nand_Gate_5.A 0.447191
R36032 Nand_Gate_5.A.n2 Nand_Gate_5.A 0.447191
R36033 Nand_Gate_5.A.n46 Nand_Gate_5.A 0.428234
R36034 Nand_Gate_5.A.n58 Nand_Gate_5.A.n3 0.425067
R36035 Nand_Gate_5.A Nand_Gate_5.A.n58 0.39003
R36036 Nand_Gate_5.A.n57 Nand_Gate_5.A.n56 0.280391
R36037 Nand_Gate_5.A.n31 Nand_Gate_5.A 0.252453
R36038 Nand_Gate_5.A.n25 Nand_Gate_5.A 0.252453
R36039 Nand_Gate_5.A.n35 Nand_Gate_5.A 0.241767
R36040 Nand_Gate_5.A.n31 Nand_Gate_5.A.n30 0.226043
R36041 Nand_Gate_5.A.n25 Nand_Gate_5.A.n24 0.226043
R36042 Nand_Gate_5.A.n27 Nand_Gate_5.A 0.217464
R36043 Nand_Gate_5.A.n21 Nand_Gate_5.A 0.217464
R36044 Nand_Gate_5.A.n12 Nand_Gate_5.A 0.217464
R36045 Nand_Gate_5.A.n6 Nand_Gate_5.A 0.217464
R36046 Nand_Gate_5.A.n56 Nand_Gate_5.A 0.200143
R36047 Nand_Gate_5.A.n40 Nand_Gate_5.A.n39 0.178317
R36048 Nand_Gate_5.A.n40 Nand_Gate_5.A 0.143974
R36049 Nand_Gate_5.A.n45 Nand_Gate_5.A 0.1255
R36050 Nand_Gate_5.A.n30 Nand_Gate_5.A 0.1255
R36051 Nand_Gate_5.A.n24 Nand_Gate_5.A 0.1255
R36052 Nand_Gate_5.A.n37 Nand_Gate_5.A 0.1255
R36053 Nand_Gate_5.A.n15 Nand_Gate_5.A 0.1255
R36054 Nand_Gate_5.A.n9 Nand_Gate_5.A 0.1255
R36055 Nand_Gate_5.A.n54 Nand_Gate_5.A 0.1255
R36056 Nand_Gate_5.A.n1 Nand_Gate_5.A 0.1255
R36057 Nand_Gate_5.A.n47 Nand_Gate_5.A.n43 0.063
R36058 Nand_Gate_5.A.n47 Nand_Gate_5.A.n46 0.063
R36059 Nand_Gate_5.A.n32 Nand_Gate_5.A.n28 0.063
R36060 Nand_Gate_5.A.n32 Nand_Gate_5.A.n31 0.063
R36061 Nand_Gate_5.A.n26 Nand_Gate_5.A.n22 0.063
R36062 Nand_Gate_5.A.n26 Nand_Gate_5.A.n25 0.063
R36063 Nand_Gate_5.A.n17 Nand_Gate_5.A.n13 0.063
R36064 Nand_Gate_5.A.n17 Nand_Gate_5.A.n16 0.063
R36065 Nand_Gate_5.A.n11 Nand_Gate_5.A.n7 0.063
R36066 Nand_Gate_5.A.n11 Nand_Gate_5.A.n10 0.063
R36067 Nand_Gate_5.A.n19 Nand_Gate_5.A.n18 0.063
R36068 Nand_Gate_5.A.n49 Nand_Gate_5.A.n20 0.063
R36069 Nand_Gate_5.A.n50 Nand_Gate_5.A.n49 0.063
R36070 Nand_Gate_5.A.n52 Nand_Gate_5.A.n5 0.063
R36071 Nand_Gate_5.A.n53 Nand_Gate_5.A.n52 0.063
R36072 Nand_Gate_5.A Nand_Gate_5.A.n54 0.063
R36073 Nand_Gate_5.A.n41 Nand_Gate_5.A.n35 0.024
R36074 Nand_Gate_5.A.n41 Nand_Gate_5.A.n40 0.024
R36075 Nand_Gate_5.A.n30 Nand_Gate_5.A.n29 0.0216397
R36076 Nand_Gate_5.A.n29 Nand_Gate_5.A 0.0216397
R36077 Nand_Gate_5.A.n24 Nand_Gate_5.A.n23 0.0216397
R36078 Nand_Gate_5.A.n23 Nand_Gate_5.A 0.0216397
R36079 Nand_Gate_5.A.n15 Nand_Gate_5.A.n14 0.0216397
R36080 Nand_Gate_5.A.n14 Nand_Gate_5.A 0.0216397
R36081 Nand_Gate_5.A.n9 Nand_Gate_5.A.n8 0.0216397
R36082 Nand_Gate_5.A.n8 Nand_Gate_5.A 0.0216397
R36083 Nand_Gate_5.A.n51 Nand_Gate_5.A 0.0168043
R36084 Nand_Gate_5.A Nand_Gate_5.A.n51 0.0122188
R36085 Nand_Gate_5.A.n45 Nand_Gate_5.A.n44 0.0107679
R36086 Nand_Gate_5.A.n44 Nand_Gate_5.A 0.0107679
R36087 Nand_Gate_5.A.n37 Nand_Gate_5.A.n36 0.0107679
R36088 Nand_Gate_5.A.n36 Nand_Gate_5.A 0.0107679
R36089 Nand_Gate_5.A.n1 Nand_Gate_5.A.n0 0.0107679
R36090 Nand_Gate_5.A.n0 Nand_Gate_5.A 0.0107679
R36091 Nand_Gate_5.A.n39 Nand_Gate_5.A 0.00441667
R36092 Nand_Gate_5.A.n3 Nand_Gate_5.A 0.00441667
R36093 Nand_Gate_5.A.n39 Nand_Gate_5.A 0.00406061
R36094 Nand_Gate_5.A.n3 Nand_Gate_5.A 0.00406061
R36095 Nand_Gate_4.B.n51 Nand_Gate_4.B.t1 169.46
R36096 Nand_Gate_4.B.n53 Nand_Gate_4.B.t3 167.809
R36097 Nand_Gate_4.B.n51 Nand_Gate_4.B.t0 167.809
R36098 Nand_Gate_4.B Nand_Gate_4.B.t17 158.585
R36099 Nand_Gate_4.B Nand_Gate_4.B.t7 158.581
R36100 Nand_Gate_4.B.n42 Nand_Gate_4.B.t10 150.293
R36101 Nand_Gate_4.B.t7 Nand_Gate_4.B.n38 150.293
R36102 Nand_Gate_4.B.t17 Nand_Gate_4.B.n2 150.293
R36103 Nand_Gate_4.B.n29 Nand_Gate_4.B.t4 150.273
R36104 Nand_Gate_4.B.n23 Nand_Gate_4.B.t11 150.273
R36105 Nand_Gate_4.B.n14 Nand_Gate_4.B.t6 150.273
R36106 Nand_Gate_4.B.n8 Nand_Gate_4.B.t16 150.273
R36107 Nand_Gate_4.B.n44 Nand_Gate_4.B.n41 76.0985
R36108 Nand_Gate_4.B.n27 Nand_Gate_4.B.t12 73.6406
R36109 Nand_Gate_4.B.n21 Nand_Gate_4.B.t5 73.6406
R36110 Nand_Gate_4.B.n12 Nand_Gate_4.B.t14 73.6406
R36111 Nand_Gate_4.B.n6 Nand_Gate_4.B.t13 73.6406
R36112 Nand_Gate_4.B.n43 Nand_Gate_4.B.t8 73.6304
R36113 Nand_Gate_4.B.n36 Nand_Gate_4.B.t15 73.6304
R36114 Nand_Gate_4.B.n0 Nand_Gate_4.B.t9 73.6304
R36115 Nand_Gate_4.B.n4 Nand_Gate_4.B.t2 60.3809
R36116 Nand_Gate_4.B.n44 Nand_Gate_4.B.n43 34.7148
R36117 Nand_Gate_4.B.n33 Nand_Gate_4.B.n26 15.5222
R36118 Nand_Gate_4.B.n52 Nand_Gate_4.B.n51 11.4489
R36119 Nand_Gate_4.B.n34 Nand_Gate_4.B.n33 8.26552
R36120 Nand_Gate_4.B.n54 Nand_Gate_4.B.n53 8.21389
R36121 Nand_Gate_4.B.n18 Nand_Gate_4.B.n11 8.1418
R36122 Nand_Gate_4.B.n47 Nand_Gate_4.B.n46 5.61191
R36123 Nand_Gate_4.B.n47 Nand_Gate_4.B 5.35402
R36124 Nand_Gate_4.B.n45 Nand_Gate_4.B.n44 4.81893
R36125 Nand_Gate_4.B.n48 Nand_Gate_4.B.n47 4.563
R36126 Nand_Gate_4.B.n33 Nand_Gate_4.B.n32 4.5005
R36127 Nand_Gate_4.B.n18 Nand_Gate_4.B.n17 4.5005
R36128 Nand_Gate_4.B.n46 Nand_Gate_4.B 1.83746
R36129 Nand_Gate_4.B.n20 Nand_Gate_4.B.n19 1.62007
R36130 Nand_Gate_4.B.n38 Nand_Gate_4.B.n37 1.19615
R36131 Nand_Gate_4.B.n2 Nand_Gate_4.B.n1 1.19615
R36132 Nand_Gate_4.B.n43 Nand_Gate_4.B.n42 1.1717
R36133 Nand_Gate_4.B.n5 Nand_Gate_4.B 1.08746
R36134 Nand_Gate_4.B.n20 Nand_Gate_4.B 1.01739
R36135 Nand_Gate_4.B.n13 Nand_Gate_4.B 0.851043
R36136 Nand_Gate_4.B.n7 Nand_Gate_4.B 0.851043
R36137 Nand_Gate_4.B.n4 Nand_Gate_4.B 0.848156
R36138 Nand_Gate_4.B.n28 Nand_Gate_4.B.n27 0.796696
R36139 Nand_Gate_4.B.n22 Nand_Gate_4.B.n21 0.796696
R36140 Nand_Gate_4.B.n50 Nand_Gate_4.B.n49 0.788543
R36141 Nand_Gate_4.B.n34 Nand_Gate_4.B 0.716182
R36142 Nand_Gate_4.B.n5 Nand_Gate_4.B.n4 0.682565
R36143 Nand_Gate_4.B.n49 Nand_Gate_4.B 0.65675
R36144 Nand_Gate_4.B.n16 Nand_Gate_4.B.n15 0.55213
R36145 Nand_Gate_4.B.n10 Nand_Gate_4.B.n9 0.55213
R36146 Nand_Gate_4.B.n28 Nand_Gate_4.B 0.524957
R36147 Nand_Gate_4.B.n22 Nand_Gate_4.B 0.524957
R36148 Nand_Gate_4.B.n16 Nand_Gate_4.B 0.486828
R36149 Nand_Gate_4.B.n10 Nand_Gate_4.B 0.486828
R36150 Nand_Gate_4.B.n13 Nand_Gate_4.B.n12 0.470609
R36151 Nand_Gate_4.B.n7 Nand_Gate_4.B.n6 0.470609
R36152 Nand_Gate_4.B.n42 Nand_Gate_4.B 0.447191
R36153 Nand_Gate_4.B.n38 Nand_Gate_4.B 0.447191
R36154 Nand_Gate_4.B.n2 Nand_Gate_4.B 0.447191
R36155 Nand_Gate_4.B.n54 Nand_Gate_4.B.n3 0.425067
R36156 Nand_Gate_4.B.n35 Nand_Gate_4.B 0.412533
R36157 Nand_Gate_4.B Nand_Gate_4.B.n54 0.39003
R36158 Nand_Gate_4.B.n35 Nand_Gate_4.B.n34 0.375717
R36159 Nand_Gate_4.B.n40 Nand_Gate_4.B.n39 0.349083
R36160 Nand_Gate_4.B.n53 Nand_Gate_4.B.n52 0.280391
R36161 Nand_Gate_4.B.n40 Nand_Gate_4.B 0.278789
R36162 Nand_Gate_4.B.n52 Nand_Gate_4.B.n50 0.262643
R36163 Nand_Gate_4.B.n31 Nand_Gate_4.B 0.252453
R36164 Nand_Gate_4.B.n25 Nand_Gate_4.B 0.252453
R36165 Nand_Gate_4.B.n31 Nand_Gate_4.B.n30 0.226043
R36166 Nand_Gate_4.B.n25 Nand_Gate_4.B.n24 0.226043
R36167 Nand_Gate_4.B.n27 Nand_Gate_4.B 0.217464
R36168 Nand_Gate_4.B.n21 Nand_Gate_4.B 0.217464
R36169 Nand_Gate_4.B.n12 Nand_Gate_4.B 0.217464
R36170 Nand_Gate_4.B.n6 Nand_Gate_4.B 0.217464
R36171 Nand_Gate_4.B.n43 Nand_Gate_4.B 0.149957
R36172 Nand_Gate_4.B.n30 Nand_Gate_4.B 0.1255
R36173 Nand_Gate_4.B.n24 Nand_Gate_4.B 0.1255
R36174 Nand_Gate_4.B.n37 Nand_Gate_4.B 0.1255
R36175 Nand_Gate_4.B.n15 Nand_Gate_4.B 0.1255
R36176 Nand_Gate_4.B.n9 Nand_Gate_4.B 0.1255
R36177 Nand_Gate_4.B.n50 Nand_Gate_4.B 0.1255
R36178 Nand_Gate_4.B.n1 Nand_Gate_4.B 0.1255
R36179 Nand_Gate_4.B.n32 Nand_Gate_4.B.n28 0.063
R36180 Nand_Gate_4.B.n32 Nand_Gate_4.B.n31 0.063
R36181 Nand_Gate_4.B.n26 Nand_Gate_4.B.n22 0.063
R36182 Nand_Gate_4.B.n26 Nand_Gate_4.B.n25 0.063
R36183 Nand_Gate_4.B.n17 Nand_Gate_4.B.n13 0.063
R36184 Nand_Gate_4.B.n17 Nand_Gate_4.B.n16 0.063
R36185 Nand_Gate_4.B.n11 Nand_Gate_4.B.n7 0.063
R36186 Nand_Gate_4.B.n11 Nand_Gate_4.B.n10 0.063
R36187 Nand_Gate_4.B.n46 Nand_Gate_4.B.n45 0.063
R36188 Nand_Gate_4.B.n45 Nand_Gate_4.B.n20 0.063
R36189 Nand_Gate_4.B.n48 Nand_Gate_4.B.n5 0.063
R36190 Nand_Gate_4.B.n49 Nand_Gate_4.B.n48 0.063
R36191 Nand_Gate_4.B.n50 Nand_Gate_4.B 0.063
R36192 Nand_Gate_4.B Nand_Gate_4.B.n18 0.0512812
R36193 Nand_Gate_4.B.n43 Nand_Gate_4.B 0.0454219
R36194 Nand_Gate_4.B.n41 Nand_Gate_4.B.n35 0.024
R36195 Nand_Gate_4.B.n41 Nand_Gate_4.B.n40 0.024
R36196 Nand_Gate_4.B.n30 Nand_Gate_4.B.n29 0.0216397
R36197 Nand_Gate_4.B.n29 Nand_Gate_4.B 0.0216397
R36198 Nand_Gate_4.B.n24 Nand_Gate_4.B.n23 0.0216397
R36199 Nand_Gate_4.B.n23 Nand_Gate_4.B 0.0216397
R36200 Nand_Gate_4.B.n15 Nand_Gate_4.B.n14 0.0216397
R36201 Nand_Gate_4.B.n14 Nand_Gate_4.B 0.0216397
R36202 Nand_Gate_4.B.n9 Nand_Gate_4.B.n8 0.0216397
R36203 Nand_Gate_4.B.n8 Nand_Gate_4.B 0.0216397
R36204 Nand_Gate_4.B.n19 Nand_Gate_4.B 0.0168043
R36205 Nand_Gate_4.B.n19 Nand_Gate_4.B 0.0122188
R36206 Nand_Gate_4.B.n37 Nand_Gate_4.B.n36 0.0107679
R36207 Nand_Gate_4.B.n36 Nand_Gate_4.B 0.0107679
R36208 Nand_Gate_4.B.n1 Nand_Gate_4.B.n0 0.0107679
R36209 Nand_Gate_4.B.n0 Nand_Gate_4.B 0.0107679
R36210 Nand_Gate_4.B.n39 Nand_Gate_4.B 0.00441667
R36211 Nand_Gate_4.B.n3 Nand_Gate_4.B 0.00441667
R36212 Nand_Gate_4.B.n39 Nand_Gate_4.B 0.00406061
R36213 Nand_Gate_4.B.n3 Nand_Gate_4.B 0.00406061
R36214 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t2 169.46
R36215 D_FlipFlop_3.3-input-nand_2.Vout.n9 D_FlipFlop_3.3-input-nand_2.Vout.t3 167.809
R36216 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.t0 167.809
R36217 D_FlipFlop_3.3-input-nand_2.Vout.t6 D_FlipFlop_3.3-input-nand_2.Vout.n11 167.227
R36218 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.t6 150.293
R36219 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.t5 150.273
R36220 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout.t7 73.6406
R36221 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout.t4 73.6304
R36222 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout.t1 60.3809
R36223 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n5 12.3891
R36224 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout.n9 11.4489
R36225 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout.n2 1.38365
R36226 D_FlipFlop_3.3-input-nand_2.Vout.n12 D_FlipFlop_3.3-input-nand_2.Vout.n1 1.19615
R36227 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout.n4 1.1717
R36228 D_FlipFlop_3.3-input-nand_2.Vout.n2 D_FlipFlop_3.3-input-nand_2.Vout 0.848156
R36229 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.Vout.n12 0.447191
R36230 D_FlipFlop_3.3-input-nand_2.Vout.n3 D_FlipFlop_3.3-input-nand_2.Vout 0.38637
R36231 D_FlipFlop_3.3-input-nand_2.Vout.n11 D_FlipFlop_3.3-input-nand_2.Vout.n10 0.280391
R36232 D_FlipFlop_3.3-input-nand_2.Vout.n10 D_FlipFlop_3.3-input-nand_2.Vout.n8 0.262643
R36233 D_FlipFlop_3.3-input-nand_2.Vout.n4 D_FlipFlop_3.3-input-nand_2.Vout 0.217464
R36234 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout 0.152844
R36235 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.149957
R36236 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R36237 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout 0.1255
R36238 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout.n7 0.0874565
R36239 D_FlipFlop_3.3-input-nand_2.Vout.n6 D_FlipFlop_3.3-input-nand_2.Vout.n3 0.063
R36240 D_FlipFlop_3.3-input-nand_2.Vout.n7 D_FlipFlop_3.3-input-nand_2.Vout.n6 0.063
R36241 D_FlipFlop_3.3-input-nand_2.Vout.n8 D_FlipFlop_3.3-input-nand_2.Vout 0.063
R36242 D_FlipFlop_3.3-input-nand_2.Vout.n5 D_FlipFlop_3.3-input-nand_2.Vout 0.0454219
R36243 D_FlipFlop_3.3-input-nand_2.Vout.n1 D_FlipFlop_3.3-input-nand_2.Vout.n0 0.0107679
R36244 D_FlipFlop_3.3-input-nand_2.Vout.n0 D_FlipFlop_3.3-input-nand_2.Vout 0.0107679
R36245 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t3 169.46
R36246 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.t1 167.809
R36247 D_FlipFlop_3.3-input-nand_2.C.n11 D_FlipFlop_3.3-input-nand_2.C.t0 167.809
R36248 D_FlipFlop_3.3-input-nand_2.C.t4 D_FlipFlop_3.3-input-nand_2.C.n13 167.226
R36249 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.t5 150.273
R36250 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.t4 150.273
R36251 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C.t7 73.6406
R36252 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C.t6 73.6304
R36253 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C.t2 60.4568
R36254 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n7 12.3891
R36255 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n11 11.4489
R36256 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C 1.68257
R36257 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C.n2 1.38365
R36258 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C.n0 1.19615
R36259 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C.n5 1.1717
R36260 D_FlipFlop_3.3-input-nand_2.C.n3 D_FlipFlop_3.3-input-nand_2.C 1.08448
R36261 D_FlipFlop_3.3-input-nand_2.C.n6 D_FlipFlop_3.3-input-nand_2.C 0.932141
R36262 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C 0.720633
R36263 D_FlipFlop_3.3-input-nand_2.C.n13 D_FlipFlop_3.3-input-nand_2.C.n12 0.280391
R36264 D_FlipFlop_3.3-input-nand_2.C.n0 D_FlipFlop_3.3-input-nand_2.C 0.217464
R36265 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C 0.1255
R36266 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.1255
R36267 D_FlipFlop_3.3-input-nand_2.C.n1 D_FlipFlop_3.3-input-nand_2.C 0.1255
R36268 D_FlipFlop_3.3-input-nand_2.C.n10 D_FlipFlop_3.3-input-nand_2.C.n9 0.0874565
R36269 D_FlipFlop_3.3-input-nand_2.C.n7 D_FlipFlop_3.3-input-nand_2.C.n6 0.063
R36270 D_FlipFlop_3.3-input-nand_2.C.n2 D_FlipFlop_3.3-input-nand_2.C 0.063
R36271 D_FlipFlop_3.3-input-nand_2.C.n9 D_FlipFlop_3.3-input-nand_2.C.n8 0.063
R36272 D_FlipFlop_3.3-input-nand_2.C.n8 D_FlipFlop_3.3-input-nand_2.C.n3 0.063
R36273 D_FlipFlop_3.3-input-nand_2.C.n12 D_FlipFlop_3.3-input-nand_2.C.n10 0.0435206
R36274 D_FlipFlop_3.3-input-nand_2.C.n14 D_FlipFlop_3.3-input-nand_2.C.n1 0.0216397
R36275 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.C.n14 0.0216397
R36276 D_FlipFlop_3.3-input-nand_2.C.n5 D_FlipFlop_3.3-input-nand_2.C.n4 0.0107679
R36277 D_FlipFlop_3.3-input-nand_2.C.n4 D_FlipFlop_3.3-input-nand_2.C 0.0107679
R36278 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C.t3 169.46
R36279 D_FlipFlop_0.3-input-nand_2.C.n4 D_FlipFlop_0.3-input-nand_2.C.t2 167.809
R36280 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C.t1 167.809
R36281 D_FlipFlop_0.3-input-nand_2.C.n3 D_FlipFlop_0.3-input-nand_2.C.t7 167.226
R36282 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.t4 150.273
R36283 D_FlipFlop_0.3-input-nand_2.C.t7 D_FlipFlop_0.3-input-nand_2.C.n2 150.273
R36284 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C.t6 73.6406
R36285 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C.t5 73.6304
R36286 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.t0 60.4568
R36287 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n11 12.3891
R36288 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C.n4 11.4489
R36289 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C 1.68257
R36290 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C.n13 1.38365
R36291 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C.n0 1.19615
R36292 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C.n9 1.1717
R36293 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C 1.08448
R36294 D_FlipFlop_0.3-input-nand_2.C.n10 D_FlipFlop_0.3-input-nand_2.C 0.932141
R36295 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C 0.720633
R36296 D_FlipFlop_0.3-input-nand_2.C.n5 D_FlipFlop_0.3-input-nand_2.C.n3 0.280391
R36297 D_FlipFlop_0.3-input-nand_2.C.n0 D_FlipFlop_0.3-input-nand_2.C 0.217464
R36298 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C 0.1255
R36299 D_FlipFlop_0.3-input-nand_2.C.n1 D_FlipFlop_0.3-input-nand_2.C 0.1255
R36300 D_FlipFlop_0.3-input-nand_2.C.n14 D_FlipFlop_0.3-input-nand_2.C 0.1255
R36301 D_FlipFlop_0.3-input-nand_2.C.n7 D_FlipFlop_0.3-input-nand_2.C.n6 0.0874565
R36302 D_FlipFlop_0.3-input-nand_2.C.n11 D_FlipFlop_0.3-input-nand_2.C.n10 0.063
R36303 D_FlipFlop_0.3-input-nand_2.C.n12 D_FlipFlop_0.3-input-nand_2.C.n7 0.063
R36304 D_FlipFlop_0.3-input-nand_2.C.n13 D_FlipFlop_0.3-input-nand_2.C.n12 0.063
R36305 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_2.C.n14 0.063
R36306 D_FlipFlop_0.3-input-nand_2.C.n6 D_FlipFlop_0.3-input-nand_2.C.n5 0.0435206
R36307 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C.n1 0.0216397
R36308 D_FlipFlop_0.3-input-nand_2.C.n2 D_FlipFlop_0.3-input-nand_2.C 0.0216397
R36309 D_FlipFlop_0.3-input-nand_2.C.n9 D_FlipFlop_0.3-input-nand_2.C.n8 0.0107679
R36310 D_FlipFlop_0.3-input-nand_2.C.n8 D_FlipFlop_0.3-input-nand_2.C 0.0107679
R36311 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 169.46
R36312 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 168.089
R36313 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 167.809
R36314 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 150.293
R36315 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 73.6304
R36316 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 60.3943
R36317 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 12.0358
R36318 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 11.4489
R36319 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.981478
R36320 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 0.788543
R36321 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.769522
R36322 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 0.720633
R36323 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 0.682565
R36324 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.580578
R36325 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 0.55213
R36326 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 0.470609
R36327 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.447191
R36328 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.428234
R36329 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.1255
R36330 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.1255
R36331 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 0.063
R36332 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 0.063
R36333 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.063
R36334 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 0.063
R36335 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 0.063
R36336 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 0.0435206
R36337 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 0.0107679
R36338 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.0107679
R36339 a_139496_37417.n0 a_139496_37417.t3 1306.95
R36340 a_139496_37417.n0 a_139496_37417.t0 1305.57
R36341 a_139496_37417.n1 a_139496_37417.t2 24.4157
R36342 a_139496_37417.t1 a_139496_37417.n1 22.6645
R36343 a_139496_37417.n1 a_139496_37417.n0 0.301808
R36344 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 169.46
R36345 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 168.089
R36346 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 167.809
R36347 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 150.293
R36348 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 73.6304
R36349 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 60.4568
R36350 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 12.0358
R36351 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 11.4489
R36352 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.981478
R36353 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 0.788543
R36354 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.769522
R36355 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 0.720633
R36356 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 0.682565
R36357 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.580578
R36358 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 0.55213
R36359 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 0.470609
R36360 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.447191
R36361 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.428234
R36362 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.1255
R36363 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.1255
R36364 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 0.063
R36365 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 0.063
R36366 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.063
R36367 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 0.063
R36368 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 0.063
R36369 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 0.0435206
R36370 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 0.0107679
R36371 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.0107679
R36372 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 169.46
R36373 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 168.089
R36374 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 167.809
R36375 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 150.273
R36376 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 73.6406
R36377 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 60.3809
R36378 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 12.0358
R36379 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 11.4489
R36380 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 1.08746
R36381 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.851043
R36382 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.848156
R36383 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 0.788543
R36384 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 0.682565
R36385 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.65675
R36386 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 0.55213
R36387 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.486828
R36388 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 0.470609
R36389 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.217464
R36390 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 0.200143
R36391 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.1255
R36392 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.1255
R36393 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 0.063
R36394 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 0.063
R36395 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 0.063
R36396 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 0.063
R36397 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 0.063
R36398 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 0.0216397
R36399 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.0216397
R36400 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 169.46
R36401 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 167.809
R36402 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 167.809
R36403 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 167.226
R36404 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 150.273
R36405 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 150.273
R36406 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 73.6406
R36407 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 73.6304
R36408 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 60.4568
R36409 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 12.3891
R36410 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 11.4489
R36411 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.68257
R36412 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 1.38365
R36413 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 1.19615
R36414 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 1.1717
R36415 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.08448
R36416 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.932141
R36417 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.720633
R36418 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 0.280391
R36419 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.217464
R36420 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R36421 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R36422 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.1255
R36423 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 0.0874565
R36424 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 0.063
R36425 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 0.063
R36426 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 0.063
R36427 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 0.063
R36428 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 0.0435206
R36429 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 0.0216397
R36430 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.0216397
R36431 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 0.0107679
R36432 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.0107679
R36433 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 169.46
R36434 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 167.809
R36435 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 167.809
R36436 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 167.227
R36437 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 150.293
R36438 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 150.273
R36439 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 73.6406
R36440 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 73.6304
R36441 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 60.3809
R36442 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 12.3891
R36443 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 11.4489
R36444 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 1.38365
R36445 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 1.19615
R36446 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 1.1717
R36447 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.848156
R36448 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 0.447191
R36449 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.38637
R36450 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 0.280391
R36451 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 0.262643
R36452 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.217464
R36453 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.152844
R36454 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.149957
R36455 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.1255
R36456 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.1255
R36457 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 0.0874565
R36458 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 0.063
R36459 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 0.063
R36460 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.063
R36461 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.0454219
R36462 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 0.0107679
R36463 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.0107679
R36464 Nand_Gate_7.B.n51 Nand_Gate_7.B.t0 169.46
R36465 Nand_Gate_7.B.n51 Nand_Gate_7.B.t1 167.809
R36466 Nand_Gate_7.B.n53 Nand_Gate_7.B.t3 167.809
R36467 Nand_Gate_7.B Nand_Gate_7.B.t15 158.585
R36468 Nand_Gate_7.B Nand_Gate_7.B.t8 158.581
R36469 Nand_Gate_7.B.n42 Nand_Gate_7.B.t16 150.293
R36470 Nand_Gate_7.B.t8 Nand_Gate_7.B.n38 150.293
R36471 Nand_Gate_7.B.t15 Nand_Gate_7.B.n2 150.293
R36472 Nand_Gate_7.B.n29 Nand_Gate_7.B.t7 150.273
R36473 Nand_Gate_7.B.n23 Nand_Gate_7.B.t17 150.273
R36474 Nand_Gate_7.B.n14 Nand_Gate_7.B.t11 150.273
R36475 Nand_Gate_7.B.n8 Nand_Gate_7.B.t14 150.273
R36476 Nand_Gate_7.B.n27 Nand_Gate_7.B.t6 73.6406
R36477 Nand_Gate_7.B.n21 Nand_Gate_7.B.t12 73.6406
R36478 Nand_Gate_7.B.n12 Nand_Gate_7.B.t13 73.6406
R36479 Nand_Gate_7.B.n6 Nand_Gate_7.B.t10 73.6406
R36480 Nand_Gate_7.B.n43 Nand_Gate_7.B.t9 73.6304
R36481 Nand_Gate_7.B.n36 Nand_Gate_7.B.t4 73.6304
R36482 Nand_Gate_7.B.n0 Nand_Gate_7.B.t5 73.6304
R36483 Nand_Gate_7.B.n44 Nand_Gate_7.B.n41 61.6632
R36484 Nand_Gate_7.B.n4 Nand_Gate_7.B.t2 60.3809
R36485 Nand_Gate_7.B.n44 Nand_Gate_7.B.n43 34.7148
R36486 Nand_Gate_7.B.n33 Nand_Gate_7.B.n26 15.5222
R36487 Nand_Gate_7.B.n52 Nand_Gate_7.B.n51 11.4489
R36488 Nand_Gate_7.B.n34 Nand_Gate_7.B.n33 8.26552
R36489 Nand_Gate_7.B.n54 Nand_Gate_7.B.n53 8.21389
R36490 Nand_Gate_7.B.n18 Nand_Gate_7.B.n11 8.1418
R36491 Nand_Gate_7.B.n47 Nand_Gate_7.B.n46 5.61191
R36492 Nand_Gate_7.B.n47 Nand_Gate_7.B 5.35402
R36493 Nand_Gate_7.B.n45 Nand_Gate_7.B.n44 4.81893
R36494 Nand_Gate_7.B.n48 Nand_Gate_7.B.n47 4.563
R36495 Nand_Gate_7.B.n33 Nand_Gate_7.B.n32 4.5005
R36496 Nand_Gate_7.B.n18 Nand_Gate_7.B.n17 4.5005
R36497 Nand_Gate_7.B.n46 Nand_Gate_7.B 1.83746
R36498 Nand_Gate_7.B.n20 Nand_Gate_7.B.n19 1.62007
R36499 Nand_Gate_7.B.n38 Nand_Gate_7.B.n37 1.19615
R36500 Nand_Gate_7.B.n2 Nand_Gate_7.B.n1 1.19615
R36501 Nand_Gate_7.B.n43 Nand_Gate_7.B.n42 1.1717
R36502 Nand_Gate_7.B.n5 Nand_Gate_7.B 1.08746
R36503 Nand_Gate_7.B.n20 Nand_Gate_7.B 1.01739
R36504 Nand_Gate_7.B.n13 Nand_Gate_7.B 0.851043
R36505 Nand_Gate_7.B.n7 Nand_Gate_7.B 0.851043
R36506 Nand_Gate_7.B.n4 Nand_Gate_7.B 0.848156
R36507 Nand_Gate_7.B.n28 Nand_Gate_7.B.n27 0.796696
R36508 Nand_Gate_7.B.n22 Nand_Gate_7.B.n21 0.796696
R36509 Nand_Gate_7.B.n50 Nand_Gate_7.B.n49 0.788543
R36510 Nand_Gate_7.B.n34 Nand_Gate_7.B 0.716182
R36511 Nand_Gate_7.B.n5 Nand_Gate_7.B.n4 0.682565
R36512 Nand_Gate_7.B.n49 Nand_Gate_7.B 0.65675
R36513 Nand_Gate_7.B.n16 Nand_Gate_7.B.n15 0.55213
R36514 Nand_Gate_7.B.n10 Nand_Gate_7.B.n9 0.55213
R36515 Nand_Gate_7.B.n28 Nand_Gate_7.B 0.524957
R36516 Nand_Gate_7.B.n22 Nand_Gate_7.B 0.524957
R36517 Nand_Gate_7.B.n16 Nand_Gate_7.B 0.486828
R36518 Nand_Gate_7.B.n10 Nand_Gate_7.B 0.486828
R36519 Nand_Gate_7.B.n35 Nand_Gate_7.B 0.481467
R36520 Nand_Gate_7.B.n13 Nand_Gate_7.B.n12 0.470609
R36521 Nand_Gate_7.B.n7 Nand_Gate_7.B.n6 0.470609
R36522 Nand_Gate_7.B.n42 Nand_Gate_7.B 0.447191
R36523 Nand_Gate_7.B.n38 Nand_Gate_7.B 0.447191
R36524 Nand_Gate_7.B.n2 Nand_Gate_7.B 0.447191
R36525 Nand_Gate_7.B.n54 Nand_Gate_7.B.n3 0.425067
R36526 Nand_Gate_7.B.n40 Nand_Gate_7.B.n39 0.418017
R36527 Nand_Gate_7.B Nand_Gate_7.B.n54 0.39003
R36528 Nand_Gate_7.B.n40 Nand_Gate_7.B 0.333211
R36529 Nand_Gate_7.B.n35 Nand_Gate_7.B.n34 0.306783
R36530 Nand_Gate_7.B.n53 Nand_Gate_7.B.n52 0.280391
R36531 Nand_Gate_7.B.n52 Nand_Gate_7.B.n50 0.262643
R36532 Nand_Gate_7.B.n31 Nand_Gate_7.B 0.252453
R36533 Nand_Gate_7.B.n25 Nand_Gate_7.B 0.252453
R36534 Nand_Gate_7.B.n31 Nand_Gate_7.B.n30 0.226043
R36535 Nand_Gate_7.B.n25 Nand_Gate_7.B.n24 0.226043
R36536 Nand_Gate_7.B.n27 Nand_Gate_7.B 0.217464
R36537 Nand_Gate_7.B.n21 Nand_Gate_7.B 0.217464
R36538 Nand_Gate_7.B.n12 Nand_Gate_7.B 0.217464
R36539 Nand_Gate_7.B.n6 Nand_Gate_7.B 0.217464
R36540 Nand_Gate_7.B.n43 Nand_Gate_7.B 0.149957
R36541 Nand_Gate_7.B.n30 Nand_Gate_7.B 0.1255
R36542 Nand_Gate_7.B.n24 Nand_Gate_7.B 0.1255
R36543 Nand_Gate_7.B.n37 Nand_Gate_7.B 0.1255
R36544 Nand_Gate_7.B.n15 Nand_Gate_7.B 0.1255
R36545 Nand_Gate_7.B.n9 Nand_Gate_7.B 0.1255
R36546 Nand_Gate_7.B.n50 Nand_Gate_7.B 0.1255
R36547 Nand_Gate_7.B.n1 Nand_Gate_7.B 0.1255
R36548 Nand_Gate_7.B.n32 Nand_Gate_7.B.n28 0.063
R36549 Nand_Gate_7.B.n32 Nand_Gate_7.B.n31 0.063
R36550 Nand_Gate_7.B.n26 Nand_Gate_7.B.n22 0.063
R36551 Nand_Gate_7.B.n26 Nand_Gate_7.B.n25 0.063
R36552 Nand_Gate_7.B.n17 Nand_Gate_7.B.n13 0.063
R36553 Nand_Gate_7.B.n17 Nand_Gate_7.B.n16 0.063
R36554 Nand_Gate_7.B.n11 Nand_Gate_7.B.n7 0.063
R36555 Nand_Gate_7.B.n11 Nand_Gate_7.B.n10 0.063
R36556 Nand_Gate_7.B.n46 Nand_Gate_7.B.n45 0.063
R36557 Nand_Gate_7.B.n45 Nand_Gate_7.B.n20 0.063
R36558 Nand_Gate_7.B.n48 Nand_Gate_7.B.n5 0.063
R36559 Nand_Gate_7.B.n49 Nand_Gate_7.B.n48 0.063
R36560 Nand_Gate_7.B.n50 Nand_Gate_7.B 0.063
R36561 Nand_Gate_7.B Nand_Gate_7.B.n18 0.0512812
R36562 Nand_Gate_7.B.n43 Nand_Gate_7.B 0.0454219
R36563 Nand_Gate_7.B.n41 Nand_Gate_7.B.n35 0.024
R36564 Nand_Gate_7.B.n41 Nand_Gate_7.B.n40 0.024
R36565 Nand_Gate_7.B.n30 Nand_Gate_7.B.n29 0.0216397
R36566 Nand_Gate_7.B.n29 Nand_Gate_7.B 0.0216397
R36567 Nand_Gate_7.B.n24 Nand_Gate_7.B.n23 0.0216397
R36568 Nand_Gate_7.B.n23 Nand_Gate_7.B 0.0216397
R36569 Nand_Gate_7.B.n15 Nand_Gate_7.B.n14 0.0216397
R36570 Nand_Gate_7.B.n14 Nand_Gate_7.B 0.0216397
R36571 Nand_Gate_7.B.n9 Nand_Gate_7.B.n8 0.0216397
R36572 Nand_Gate_7.B.n8 Nand_Gate_7.B 0.0216397
R36573 Nand_Gate_7.B.n19 Nand_Gate_7.B 0.0168043
R36574 Nand_Gate_7.B.n19 Nand_Gate_7.B 0.0122188
R36575 Nand_Gate_7.B.n37 Nand_Gate_7.B.n36 0.0107679
R36576 Nand_Gate_7.B.n36 Nand_Gate_7.B 0.0107679
R36577 Nand_Gate_7.B.n1 Nand_Gate_7.B.n0 0.0107679
R36578 Nand_Gate_7.B.n0 Nand_Gate_7.B 0.0107679
R36579 Nand_Gate_7.B.n39 Nand_Gate_7.B 0.00441667
R36580 Nand_Gate_7.B.n3 Nand_Gate_7.B 0.00441667
R36581 Nand_Gate_7.B.n39 Nand_Gate_7.B 0.00406061
R36582 Nand_Gate_7.B.n3 Nand_Gate_7.B 0.00406061
R36583 Q1.n5 Q1.t1 169.46
R36584 Q1.n7 Q1.t2 167.809
R36585 Q1.n5 Q1.t0 167.809
R36586 Q1.n11 Q1.t4 155.124
R36587 Q1.n14 Q1.t7 150.869
R36588 Q1.n13 Q1.t9 150.869
R36589 Q1.t4 Q1.n2 150.293
R36590 Q1.n15 Q1.n12 137.644
R36591 Q1 Q1.t5 78.1811
R36592 Q1.n13 Q1.t6 74.1352
R36593 Q1.t5 Q1.n14 74.1352
R36594 Q1.n0 Q1.t8 73.6304
R36595 Q1.n3 Q1.t3 60.3809
R36596 Q1.n12 Q1 41.1198
R36597 Q1.n6 Q1.n5 11.4489
R36598 Q1.n8 Q1.n7 8.21389
R36599 Q1.n11 Q1.n10 1.70176
R36600 Q1.n14 Q1.n13 1.66898
R36601 Q1.n4 Q1.n3 1.64452
R36602 Q1.n2 Q1.n1 1.19615
R36603 Q1.n3 Q1 0.848156
R36604 Q1.n2 Q1 0.447191
R36605 Q1.n8 Q1 0.39003
R36606 Q1.n9 Q1.n8 0.3624
R36607 Q1.n7 Q1.n6 0.280391
R36608 Q1.n6 Q1.n4 0.262643
R36609 Q1.n4 Q1 0.1255
R36610 Q1.n1 Q1 0.1255
R36611 Q1.n9 Q1 0.0670833
R36612 Q1.n13 Q1 0.063
R36613 Q1.n4 Q1 0.063
R36614 Q1.n10 Q1.n9 0.0428618
R36615 Q1.n12 Q1.n11 0.0305325
R36616 Q1.n10 Q1 0.0194691
R36617 Q1 Q1.n15 0.0168043
R36618 Q1.n15 Q1 0.0122188
R36619 Q1.n1 Q1.n0 0.0107679
R36620 Q1.n0 Q1 0.0107679
R36621 Vin Vin.t0 467.378
R36622 a_138366_35417.n0 a_138366_35417.t3 1546.57
R36623 a_138366_35417.t0 a_138366_35417.n1 27.6313
R36624 a_138366_35417.n1 a_138366_35417.t1 21.1653
R36625 a_138366_35417.n0 a_138366_35417.t2 11.1233
R36626 a_138366_35417.n1 a_138366_35417.n0 6.05452
R36627 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 169.46
R36628 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 167.809
R36629 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 167.809
R36630 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 167.227
R36631 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 150.293
R36632 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 150.273
R36633 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 73.6406
R36634 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 73.6304
R36635 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 60.3809
R36636 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 12.3891
R36637 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 11.4489
R36638 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 1.38365
R36639 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 1.19615
R36640 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 1.1717
R36641 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.848156
R36642 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 0.447191
R36643 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.38637
R36644 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 0.280391
R36645 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 0.262643
R36646 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.217464
R36647 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.152844
R36648 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.149957
R36649 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.1255
R36650 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.1255
R36651 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 0.0874565
R36652 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 0.063
R36653 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 0.063
R36654 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.063
R36655 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.0454219
R36656 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 0.0107679
R36657 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.0107679
R36658 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 169.46
R36659 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 167.809
R36660 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 167.809
R36661 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 167.226
R36662 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 150.273
R36663 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 150.273
R36664 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 73.6406
R36665 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 73.6304
R36666 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 60.4568
R36667 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 12.3891
R36668 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 11.4489
R36669 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.68257
R36670 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 1.38365
R36671 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 1.19615
R36672 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 1.1717
R36673 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.08448
R36674 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.932141
R36675 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 0.720633
R36676 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 0.280391
R36677 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.217464
R36678 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R36679 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R36680 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.1255
R36681 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 0.0874565
R36682 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 0.063
R36683 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.063
R36684 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 0.063
R36685 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 0.063
R36686 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 0.0435206
R36687 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 0.0216397
R36688 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.0216397
R36689 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 0.0107679
R36690 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.0107679
R36691 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 169.46
R36692 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 167.809
R36693 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 167.809
R36694 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 167.227
R36695 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 150.293
R36696 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 150.273
R36697 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 73.6406
R36698 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 73.6304
R36699 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 60.3809
R36700 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 12.3891
R36701 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 11.4489
R36702 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 1.38365
R36703 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 1.19615
R36704 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 1.1717
R36705 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.848156
R36706 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 0.447191
R36707 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.38637
R36708 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 0.280391
R36709 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.217464
R36710 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.200143
R36711 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.152844
R36712 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.149957
R36713 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.1255
R36714 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.1255
R36715 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 0.0874565
R36716 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 0.063
R36717 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 0.063
R36718 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 0.063
R36719 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0454219
R36720 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 0.0107679
R36721 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0107679
R36722 CDAC8_0.switch_1.Z.n4 CDAC8_0.switch_1.Z.t3 168.075
R36723 CDAC8_0.switch_1.Z.n4 CDAC8_0.switch_1.Z.t0 168.075
R36724 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z.t2 60.6851
R36725 CDAC8_0.switch_1.Z CDAC8_0.switch_1.Z.t1 60.6226
R36726 CDAC8_0.switch_1.Z.n2 CDAC8_0.switch_1.Z.t4 14.5332
R36727 CDAC8_0.switch_1.Z.n5 CDAC8_0.switch_1.Z.n3 1.29126
R36728 CDAC8_0.switch_1.Z.n3 CDAC8_0.switch_1.Z 0.478761
R36729 CDAC8_0.switch_1.Z.n1 CDAC8_0.switch_1.Z 0.21925
R36730 CDAC8_0.switch_1.Z.n1 CDAC8_0.switch_1.Z.n0 0.179848
R36731 CDAC8_0.switch_1.Z CDAC8_0.switch_1.Z.n5 0.178175
R36732 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z 0.1255
R36733 CDAC8_0.switch_1.Z.n0 CDAC8_0.switch_1.Z 0.063
R36734 CDAC8_0.switch_1.Z.n3 CDAC8_0.switch_1.Z.n2 0.063
R36735 CDAC8_0.switch_1.Z.n2 CDAC8_0.switch_1.Z.n1 0.063
R36736 CDAC8_0.switch_1.Z.n5 CDAC8_0.switch_1.Z.n4 0.0130546
R36737 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 169.46
R36738 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 167.809
R36739 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 167.809
R36740 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 167.227
R36741 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 150.293
R36742 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 150.273
R36743 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 73.6406
R36744 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 73.6304
R36745 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 60.3809
R36746 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 12.3891
R36747 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 11.4489
R36748 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 1.38365
R36749 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 1.19615
R36750 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 1.1717
R36751 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.848156
R36752 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 0.447191
R36753 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R36754 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 0.280391
R36755 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.217464
R36756 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.200143
R36757 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R36758 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R36759 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R36760 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R36761 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 0.0874565
R36762 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 0.063
R36763 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 0.063
R36764 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 0.063
R36765 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R36766 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 0.0107679
R36767 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0107679
R36768 Nand_Gate_2.Vout.n10 Nand_Gate_2.Vout.t0 179.256
R36769 Nand_Gate_2.Vout.n10 Nand_Gate_2.Vout.t1 168.089
R36770 Nand_Gate_2.Vout.n2 Nand_Gate_2.Vout.t4 150.293
R36771 Nand_Gate_2.Vout.n4 Nand_Gate_2.Vout.t3 73.6304
R36772 Nand_Gate_2.Vout Nand_Gate_2.Vout.t2 60.3943
R36773 Nand_Gate_2.Vout.n8 Nand_Gate_2.Vout.n7 35.6663
R36774 Nand_Gate_2.Vout.n9 Nand_Gate_2.Vout 0.981478
R36775 Nand_Gate_2.Vout.n11 Nand_Gate_2.Vout.n9 0.788543
R36776 Nand_Gate_2.Vout.n3 Nand_Gate_2.Vout 0.769522
R36777 Nand_Gate_2.Vout Nand_Gate_2.Vout.n11 0.720633
R36778 Nand_Gate_2.Vout.n1 Nand_Gate_2.Vout.n0 0.682565
R36779 Nand_Gate_2.Vout.n1 Nand_Gate_2.Vout 0.580578
R36780 Nand_Gate_2.Vout.n3 Nand_Gate_2.Vout.n2 0.55213
R36781 Nand_Gate_2.Vout.n6 Nand_Gate_2.Vout.n5 0.470609
R36782 Nand_Gate_2.Vout.n2 Nand_Gate_2.Vout 0.447191
R36783 Nand_Gate_2.Vout.n6 Nand_Gate_2.Vout 0.428234
R36784 Nand_Gate_2.Vout.n5 Nand_Gate_2.Vout 0.1255
R36785 Nand_Gate_2.Vout.n0 Nand_Gate_2.Vout 0.1255
R36786 Nand_Gate_2.Vout.n7 Nand_Gate_2.Vout.n3 0.063
R36787 Nand_Gate_2.Vout.n7 Nand_Gate_2.Vout.n6 0.063
R36788 Nand_Gate_2.Vout.n0 Nand_Gate_2.Vout 0.063
R36789 Nand_Gate_2.Vout.n9 Nand_Gate_2.Vout.n8 0.063
R36790 Nand_Gate_2.Vout.n8 Nand_Gate_2.Vout.n1 0.063
R36791 Nand_Gate_2.Vout.n11 Nand_Gate_2.Vout.n10 0.0435206
R36792 Nand_Gate_2.Vout.n5 Nand_Gate_2.Vout.n4 0.0107679
R36793 Nand_Gate_2.Vout.n4 Nand_Gate_2.Vout 0.0107679
R36794 Nand_Gate_3.B.n31 Nand_Gate_3.B.t0 169.46
R36795 Nand_Gate_3.B.n31 Nand_Gate_3.B.t1 167.809
R36796 Nand_Gate_3.B.n33 Nand_Gate_3.B.t3 167.809
R36797 Nand_Gate_3.B Nand_Gate_3.B.t7 158.585
R36798 Nand_Gate_3.B.t7 Nand_Gate_3.B.n2 150.293
R36799 Nand_Gate_3.B.n24 Nand_Gate_3.B.t6 150.273
R36800 Nand_Gate_3.B.n14 Nand_Gate_3.B.t10 150.273
R36801 Nand_Gate_3.B.n8 Nand_Gate_3.B.t5 150.273
R36802 Nand_Gate_3.B.n12 Nand_Gate_3.B.t4 73.6406
R36803 Nand_Gate_3.B.n6 Nand_Gate_3.B.t11 73.6406
R36804 Nand_Gate_3.B.n21 Nand_Gate_3.B.t8 73.6304
R36805 Nand_Gate_3.B.n0 Nand_Gate_3.B.t9 73.6304
R36806 Nand_Gate_3.B.n4 Nand_Gate_3.B.t2 60.3809
R36807 Nand_Gate_3.B.n25 Nand_Gate_3.B.n24 40.8363
R36808 Nand_Gate_3.B.n32 Nand_Gate_3.B.n31 11.4489
R36809 Nand_Gate_3.B.n34 Nand_Gate_3.B.n33 8.21389
R36810 Nand_Gate_3.B.n18 Nand_Gate_3.B.n11 8.1418
R36811 Nand_Gate_3.B.n20 Nand_Gate_3.B.n19 6.47604
R36812 Nand_Gate_3.B.n19 Nand_Gate_3.B 5.35402
R36813 Nand_Gate_3.B.n28 Nand_Gate_3.B 4.55128
R36814 Nand_Gate_3.B.n18 Nand_Gate_3.B.n17 4.5005
R36815 Nand_Gate_3.B.n2 Nand_Gate_3.B.n1 1.19615
R36816 Nand_Gate_3.B.n23 Nand_Gate_3.B.n22 1.1717
R36817 Nand_Gate_3.B.n5 Nand_Gate_3.B 1.08746
R36818 Nand_Gate_3.B.n20 Nand_Gate_3.B 0.973326
R36819 Nand_Gate_3.B.n23 Nand_Gate_3.B 0.932141
R36820 Nand_Gate_3.B.n13 Nand_Gate_3.B 0.851043
R36821 Nand_Gate_3.B.n7 Nand_Gate_3.B 0.851043
R36822 Nand_Gate_3.B.n4 Nand_Gate_3.B 0.848156
R36823 Nand_Gate_3.B.n30 Nand_Gate_3.B.n29 0.788543
R36824 Nand_Gate_3.B.n27 Nand_Gate_3.B.n26 0.755935
R36825 Nand_Gate_3.B.n5 Nand_Gate_3.B.n4 0.682565
R36826 Nand_Gate_3.B.n29 Nand_Gate_3.B 0.65675
R36827 Nand_Gate_3.B.n16 Nand_Gate_3.B.n15 0.55213
R36828 Nand_Gate_3.B.n10 Nand_Gate_3.B.n9 0.55213
R36829 Nand_Gate_3.B.n16 Nand_Gate_3.B 0.486828
R36830 Nand_Gate_3.B.n10 Nand_Gate_3.B 0.486828
R36831 Nand_Gate_3.B.n26 Nand_Gate_3.B 0.48023
R36832 Nand_Gate_3.B.n13 Nand_Gate_3.B.n12 0.470609
R36833 Nand_Gate_3.B.n7 Nand_Gate_3.B.n6 0.470609
R36834 Nand_Gate_3.B.n2 Nand_Gate_3.B 0.447191
R36835 Nand_Gate_3.B.n34 Nand_Gate_3.B.n3 0.425067
R36836 Nand_Gate_3.B Nand_Gate_3.B.n34 0.39003
R36837 Nand_Gate_3.B.n33 Nand_Gate_3.B.n32 0.280391
R36838 Nand_Gate_3.B.n12 Nand_Gate_3.B 0.217464
R36839 Nand_Gate_3.B.n6 Nand_Gate_3.B 0.217464
R36840 Nand_Gate_3.B.n32 Nand_Gate_3.B 0.200143
R36841 Nand_Gate_3.B.n22 Nand_Gate_3.B 0.1255
R36842 Nand_Gate_3.B.n15 Nand_Gate_3.B 0.1255
R36843 Nand_Gate_3.B.n9 Nand_Gate_3.B 0.1255
R36844 Nand_Gate_3.B.n30 Nand_Gate_3.B 0.1255
R36845 Nand_Gate_3.B.n1 Nand_Gate_3.B 0.1255
R36846 Nand_Gate_3.B.n24 Nand_Gate_3.B.n23 0.063
R36847 Nand_Gate_3.B.n17 Nand_Gate_3.B.n13 0.063
R36848 Nand_Gate_3.B.n17 Nand_Gate_3.B.n16 0.063
R36849 Nand_Gate_3.B.n11 Nand_Gate_3.B.n7 0.063
R36850 Nand_Gate_3.B.n11 Nand_Gate_3.B.n10 0.063
R36851 Nand_Gate_3.B.n19 Nand_Gate_3.B.n18 0.063
R36852 Nand_Gate_3.B.n25 Nand_Gate_3.B.n20 0.063
R36853 Nand_Gate_3.B.n26 Nand_Gate_3.B.n25 0.063
R36854 Nand_Gate_3.B.n28 Nand_Gate_3.B.n5 0.063
R36855 Nand_Gate_3.B.n29 Nand_Gate_3.B.n28 0.063
R36856 Nand_Gate_3.B Nand_Gate_3.B.n30 0.063
R36857 Nand_Gate_3.B.n15 Nand_Gate_3.B.n14 0.0216397
R36858 Nand_Gate_3.B.n14 Nand_Gate_3.B 0.0216397
R36859 Nand_Gate_3.B.n9 Nand_Gate_3.B.n8 0.0216397
R36860 Nand_Gate_3.B.n8 Nand_Gate_3.B 0.0216397
R36861 Nand_Gate_3.B.n27 Nand_Gate_3.B 0.0168043
R36862 Nand_Gate_3.B Nand_Gate_3.B.n27 0.0122188
R36863 Nand_Gate_3.B.n22 Nand_Gate_3.B.n21 0.0107679
R36864 Nand_Gate_3.B.n21 Nand_Gate_3.B 0.0107679
R36865 Nand_Gate_3.B.n1 Nand_Gate_3.B.n0 0.0107679
R36866 Nand_Gate_3.B.n0 Nand_Gate_3.B 0.0107679
R36867 Nand_Gate_3.B.n3 Nand_Gate_3.B 0.00441667
R36868 Nand_Gate_3.B.n3 Nand_Gate_3.B 0.00406061
R36869 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 316.762
R36870 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 168.108
R36871 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 150.293
R36872 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 150.273
R36873 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 73.6406
R36874 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 73.6304
R36875 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 60.4568
R36876 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 12.0358
R36877 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 1.19615
R36878 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.981478
R36879 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 0.788543
R36880 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.769522
R36881 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 0.682565
R36882 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.580578
R36883 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 0.55213
R36884 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 0.484875
R36885 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 0.470609
R36886 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.447191
R36887 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.428234
R36888 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.217464
R36889 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R36890 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R36891 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.1255
R36892 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 0.063
R36893 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 0.063
R36894 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.063
R36895 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 0.063
R36896 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 0.063
R36897 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 0.0216397
R36898 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.0216397
R36899 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 0.0107679
R36900 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.0107679
R36901 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 169.46
R36902 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 167.809
R36903 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 167.809
R36904 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 167.227
R36905 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 150.293
R36906 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 150.273
R36907 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 73.6406
R36908 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 73.6304
R36909 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 60.3809
R36910 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 12.3891
R36911 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 11.4489
R36912 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 1.38365
R36913 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 1.19615
R36914 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 1.1717
R36915 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.848156
R36916 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 0.447191
R36917 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R36918 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 0.280391
R36919 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.217464
R36920 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.200143
R36921 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R36922 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R36923 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R36924 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R36925 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 0.0874565
R36926 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 0.063
R36927 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 0.063
R36928 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 0.063
R36929 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R36930 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 0.0107679
R36931 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0107679
R36932 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 316.762
R36933 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 168.108
R36934 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 150.293
R36935 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 150.273
R36936 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 73.6406
R36937 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 73.6304
R36938 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 60.3943
R36939 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 12.0358
R36940 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 1.19615
R36941 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.981478
R36942 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 0.788543
R36943 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.769522
R36944 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 0.682565
R36945 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.580578
R36946 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 0.55213
R36947 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 0.484875
R36948 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 0.470609
R36949 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.447191
R36950 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.428234
R36951 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.217464
R36952 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R36953 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R36954 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.1255
R36955 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 0.063
R36956 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 0.063
R36957 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.063
R36958 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 0.063
R36959 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 0.063
R36960 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 0.0216397
R36961 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.0216397
R36962 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 0.0107679
R36963 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.0107679
R36964 Nand_Gate_1.B.n51 Nand_Gate_1.B.t0 169.46
R36965 Nand_Gate_1.B.n51 Nand_Gate_1.B.t3 167.809
R36966 Nand_Gate_1.B.n53 Nand_Gate_1.B.t2 167.809
R36967 Nand_Gate_1.B Nand_Gate_1.B.t16 158.585
R36968 Nand_Gate_1.B Nand_Gate_1.B.t9 158.581
R36969 Nand_Gate_1.B.n42 Nand_Gate_1.B.t4 150.293
R36970 Nand_Gate_1.B.t9 Nand_Gate_1.B.n38 150.293
R36971 Nand_Gate_1.B.t16 Nand_Gate_1.B.n2 150.293
R36972 Nand_Gate_1.B.n29 Nand_Gate_1.B.t7 150.273
R36973 Nand_Gate_1.B.n23 Nand_Gate_1.B.t14 150.273
R36974 Nand_Gate_1.B.n14 Nand_Gate_1.B.t11 150.273
R36975 Nand_Gate_1.B.n8 Nand_Gate_1.B.t6 150.273
R36976 Nand_Gate_1.B.n27 Nand_Gate_1.B.t8 73.6406
R36977 Nand_Gate_1.B.n21 Nand_Gate_1.B.t15 73.6406
R36978 Nand_Gate_1.B.n12 Nand_Gate_1.B.t5 73.6406
R36979 Nand_Gate_1.B.n6 Nand_Gate_1.B.t10 73.6406
R36980 Nand_Gate_1.B.n43 Nand_Gate_1.B.t12 73.6304
R36981 Nand_Gate_1.B.n36 Nand_Gate_1.B.t17 73.6304
R36982 Nand_Gate_1.B.n0 Nand_Gate_1.B.t13 73.6304
R36983 Nand_Gate_1.B.n4 Nand_Gate_1.B.t1 60.3809
R36984 Nand_Gate_1.B.n44 Nand_Gate_1.B.n43 34.7148
R36985 Nand_Gate_1.B.n44 Nand_Gate_1.B.n41 32.6611
R36986 Nand_Gate_1.B.n33 Nand_Gate_1.B.n26 15.5222
R36987 Nand_Gate_1.B.n52 Nand_Gate_1.B.n51 11.4489
R36988 Nand_Gate_1.B.n34 Nand_Gate_1.B.n33 8.26552
R36989 Nand_Gate_1.B.n54 Nand_Gate_1.B.n53 8.21389
R36990 Nand_Gate_1.B.n18 Nand_Gate_1.B.n11 8.1418
R36991 Nand_Gate_1.B.n47 Nand_Gate_1.B.n46 5.61191
R36992 Nand_Gate_1.B.n47 Nand_Gate_1.B 5.35402
R36993 Nand_Gate_1.B.n45 Nand_Gate_1.B.n44 4.81893
R36994 Nand_Gate_1.B.n48 Nand_Gate_1.B.n47 4.563
R36995 Nand_Gate_1.B.n33 Nand_Gate_1.B.n32 4.5005
R36996 Nand_Gate_1.B.n18 Nand_Gate_1.B.n17 4.5005
R36997 Nand_Gate_1.B.n46 Nand_Gate_1.B 1.83746
R36998 Nand_Gate_1.B.n20 Nand_Gate_1.B.n19 1.62007
R36999 Nand_Gate_1.B.n38 Nand_Gate_1.B.n37 1.19615
R37000 Nand_Gate_1.B.n2 Nand_Gate_1.B.n1 1.19615
R37001 Nand_Gate_1.B.n43 Nand_Gate_1.B.n42 1.1717
R37002 Nand_Gate_1.B.n5 Nand_Gate_1.B 1.08746
R37003 Nand_Gate_1.B.n20 Nand_Gate_1.B 1.01739
R37004 Nand_Gate_1.B.n13 Nand_Gate_1.B 0.851043
R37005 Nand_Gate_1.B.n7 Nand_Gate_1.B 0.851043
R37006 Nand_Gate_1.B.n4 Nand_Gate_1.B 0.848156
R37007 Nand_Gate_1.B.n28 Nand_Gate_1.B.n27 0.796696
R37008 Nand_Gate_1.B.n22 Nand_Gate_1.B.n21 0.796696
R37009 Nand_Gate_1.B.n50 Nand_Gate_1.B.n49 0.788543
R37010 Nand_Gate_1.B.n34 Nand_Gate_1.B 0.716182
R37011 Nand_Gate_1.B.n5 Nand_Gate_1.B.n4 0.682565
R37012 Nand_Gate_1.B.n49 Nand_Gate_1.B 0.65675
R37013 Nand_Gate_1.B.n16 Nand_Gate_1.B.n15 0.55213
R37014 Nand_Gate_1.B.n10 Nand_Gate_1.B.n9 0.55213
R37015 Nand_Gate_1.B.n28 Nand_Gate_1.B 0.524957
R37016 Nand_Gate_1.B.n22 Nand_Gate_1.B 0.524957
R37017 Nand_Gate_1.B.n35 Nand_Gate_1.B 0.487733
R37018 Nand_Gate_1.B.n16 Nand_Gate_1.B 0.486828
R37019 Nand_Gate_1.B.n10 Nand_Gate_1.B 0.486828
R37020 Nand_Gate_1.B.n13 Nand_Gate_1.B.n12 0.470609
R37021 Nand_Gate_1.B.n7 Nand_Gate_1.B.n6 0.470609
R37022 Nand_Gate_1.B.n42 Nand_Gate_1.B 0.447191
R37023 Nand_Gate_1.B.n38 Nand_Gate_1.B 0.447191
R37024 Nand_Gate_1.B.n2 Nand_Gate_1.B 0.447191
R37025 Nand_Gate_1.B.n54 Nand_Gate_1.B.n3 0.425067
R37026 Nand_Gate_1.B.n40 Nand_Gate_1.B.n39 0.424283
R37027 Nand_Gate_1.B Nand_Gate_1.B.n54 0.39003
R37028 Nand_Gate_1.B.n40 Nand_Gate_1.B 0.338158
R37029 Nand_Gate_1.B.n35 Nand_Gate_1.B.n34 0.300517
R37030 Nand_Gate_1.B.n53 Nand_Gate_1.B.n52 0.280391
R37031 Nand_Gate_1.B.n52 Nand_Gate_1.B.n50 0.262643
R37032 Nand_Gate_1.B.n31 Nand_Gate_1.B 0.252453
R37033 Nand_Gate_1.B.n25 Nand_Gate_1.B 0.252453
R37034 Nand_Gate_1.B.n31 Nand_Gate_1.B.n30 0.226043
R37035 Nand_Gate_1.B.n25 Nand_Gate_1.B.n24 0.226043
R37036 Nand_Gate_1.B.n27 Nand_Gate_1.B 0.217464
R37037 Nand_Gate_1.B.n21 Nand_Gate_1.B 0.217464
R37038 Nand_Gate_1.B.n12 Nand_Gate_1.B 0.217464
R37039 Nand_Gate_1.B.n6 Nand_Gate_1.B 0.217464
R37040 Nand_Gate_1.B.n43 Nand_Gate_1.B 0.149957
R37041 Nand_Gate_1.B.n30 Nand_Gate_1.B 0.1255
R37042 Nand_Gate_1.B.n24 Nand_Gate_1.B 0.1255
R37043 Nand_Gate_1.B.n37 Nand_Gate_1.B 0.1255
R37044 Nand_Gate_1.B.n15 Nand_Gate_1.B 0.1255
R37045 Nand_Gate_1.B.n9 Nand_Gate_1.B 0.1255
R37046 Nand_Gate_1.B.n50 Nand_Gate_1.B 0.1255
R37047 Nand_Gate_1.B.n1 Nand_Gate_1.B 0.1255
R37048 Nand_Gate_1.B.n32 Nand_Gate_1.B.n28 0.063
R37049 Nand_Gate_1.B.n32 Nand_Gate_1.B.n31 0.063
R37050 Nand_Gate_1.B.n26 Nand_Gate_1.B.n22 0.063
R37051 Nand_Gate_1.B.n26 Nand_Gate_1.B.n25 0.063
R37052 Nand_Gate_1.B.n17 Nand_Gate_1.B.n13 0.063
R37053 Nand_Gate_1.B.n17 Nand_Gate_1.B.n16 0.063
R37054 Nand_Gate_1.B.n11 Nand_Gate_1.B.n7 0.063
R37055 Nand_Gate_1.B.n11 Nand_Gate_1.B.n10 0.063
R37056 Nand_Gate_1.B.n46 Nand_Gate_1.B.n45 0.063
R37057 Nand_Gate_1.B.n45 Nand_Gate_1.B.n20 0.063
R37058 Nand_Gate_1.B.n48 Nand_Gate_1.B.n5 0.063
R37059 Nand_Gate_1.B.n49 Nand_Gate_1.B.n48 0.063
R37060 Nand_Gate_1.B.n50 Nand_Gate_1.B 0.063
R37061 Nand_Gate_1.B Nand_Gate_1.B.n18 0.0512812
R37062 Nand_Gate_1.B.n43 Nand_Gate_1.B 0.0454219
R37063 Nand_Gate_1.B.n41 Nand_Gate_1.B.n35 0.024
R37064 Nand_Gate_1.B.n41 Nand_Gate_1.B.n40 0.024
R37065 Nand_Gate_1.B.n30 Nand_Gate_1.B.n29 0.0216397
R37066 Nand_Gate_1.B.n29 Nand_Gate_1.B 0.0216397
R37067 Nand_Gate_1.B.n24 Nand_Gate_1.B.n23 0.0216397
R37068 Nand_Gate_1.B.n23 Nand_Gate_1.B 0.0216397
R37069 Nand_Gate_1.B.n15 Nand_Gate_1.B.n14 0.0216397
R37070 Nand_Gate_1.B.n14 Nand_Gate_1.B 0.0216397
R37071 Nand_Gate_1.B.n9 Nand_Gate_1.B.n8 0.0216397
R37072 Nand_Gate_1.B.n8 Nand_Gate_1.B 0.0216397
R37073 Nand_Gate_1.B.n19 Nand_Gate_1.B 0.0168043
R37074 Nand_Gate_1.B.n19 Nand_Gate_1.B 0.0122188
R37075 Nand_Gate_1.B.n37 Nand_Gate_1.B.n36 0.0107679
R37076 Nand_Gate_1.B.n36 Nand_Gate_1.B 0.0107679
R37077 Nand_Gate_1.B.n1 Nand_Gate_1.B.n0 0.0107679
R37078 Nand_Gate_1.B.n0 Nand_Gate_1.B 0.0107679
R37079 Nand_Gate_1.B.n39 Nand_Gate_1.B 0.00441667
R37080 Nand_Gate_1.B.n3 Nand_Gate_1.B 0.00441667
R37081 Nand_Gate_1.B.n39 Nand_Gate_1.B 0.00406061
R37082 Nand_Gate_1.B.n3 Nand_Gate_1.B 0.00406061
R37083 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 169.46
R37084 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 168.089
R37085 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 167.809
R37086 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 150.293
R37087 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 73.6304
R37088 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 60.3943
R37089 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 12.0358
R37090 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 11.4489
R37091 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.981478
R37092 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 0.788543
R37093 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.769522
R37094 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 0.720633
R37095 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 0.682565
R37096 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.580578
R37097 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 0.55213
R37098 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 0.470609
R37099 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.447191
R37100 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.428234
R37101 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.1255
R37102 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.1255
R37103 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 0.063
R37104 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 0.063
R37105 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.063
R37106 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 0.063
R37107 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 0.063
R37108 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 0.0435206
R37109 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 0.0107679
R37110 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.0107679
R37111 Q7.n2 Q7.t3 169.46
R37112 Q7.n4 Q7.t1 167.809
R37113 Q7.n2 Q7.t2 167.809
R37114 Q7 Q7.t6 158.585
R37115 Q7 Q7.t9 154.823
R37116 Q7.n14 Q7.t4 150.869
R37117 Q7.t9 Q7.n15 150.869
R37118 Q7.t6 Q7.n9 150.293
R37119 Q7.n16 Q7.n13 137.644
R37120 Q7.n13 Q7 85.5731
R37121 Q7.n15 Q7.t7 74.1352
R37122 Q7.n14 Q7.t8 74.1352
R37123 Q7.n7 Q7.t5 73.6304
R37124 Q7.n0 Q7.t0 60.3809
R37125 Q7.n3 Q7.n2 11.4489
R37126 Q7.n5 Q7.n4 8.21389
R37127 Q7.n13 Q7.n12 3.473
R37128 Q7.n15 Q7.n14 1.66898
R37129 Q7.n1 Q7.n0 1.64452
R37130 Q7.n9 Q7.n8 1.19615
R37131 Q7.n0 Q7 0.848156
R37132 Q7.n9 Q7 0.447191
R37133 Q7.n5 Q7 0.39003
R37134 Q7.n4 Q7.n3 0.280391
R37135 Q7.n3 Q7.n1 0.262643
R37136 Q7.n6 Q7.n5 0.224533
R37137 Q7.n6 Q7 0.20495
R37138 Q7.n11 Q7.n10 0.149333
R37139 Q7.n11 Q7 0.139364
R37140 Q7.n1 Q7 0.1255
R37141 Q7.n8 Q7 0.1255
R37142 Q7.n14 Q7 0.063
R37143 Q7.n1 Q7 0.063
R37144 Q7.n12 Q7.n6 0.024
R37145 Q7.n12 Q7.n11 0.024
R37146 Q7 Q7.n16 0.0168043
R37147 Q7.n16 Q7 0.0122188
R37148 Q7.n8 Q7.n7 0.0107679
R37149 Q7.n7 Q7 0.0107679
R37150 Q7.n10 Q7 0.00441667
R37151 Q7.n10 Q7 0.00406061
R37152 And_Gate_5.Vout.n15 And_Gate_5.Vout.t0 168.108
R37153 And_Gate_5.Vout.n5 And_Gate_5.Vout.t6 158.207
R37154 D_FlipFlop_1.CLK And_Gate_5.Vout.t2 158.202
R37155 And_Gate_5.Vout.n7 And_Gate_5.Vout.t7 150.293
R37156 And_Gate_5.Vout.t2 And_Gate_5.Vout.n10 150.293
R37157 And_Gate_5.Vout.t6 And_Gate_5.Vout.n4 150.273
R37158 And_Gate_5.Vout.n13 And_Gate_5.Vout.n12 89.3276
R37159 And_Gate_5.Vout.n2 And_Gate_5.Vout.t3 73.6406
R37160 And_Gate_5.Vout.n9 And_Gate_5.Vout.t5 73.6304
R37161 And_Gate_5.Vout.n8 And_Gate_5.Vout.t4 73.6304
R37162 And_Gate_5.Inverter_0.Vout And_Gate_5.Vout.t1 60.3943
R37163 And_Gate_5.Vout.n9 And_Gate_5.Vout.n8 16.332
R37164 And_Gate_5.Vout.n3 And_Gate_5.Vout.n2 1.19615
R37165 And_Gate_5.Vout.n8 And_Gate_5.Vout.n7 1.1717
R37166 And_Gate_5.Vout.n10 And_Gate_5.Vout.n9 1.1717
R37167 And_Gate_5.Vout.n14 And_Gate_5.Inverter_0.Vout 0.981478
R37168 And_Gate_5.Vout.n15 And_Gate_5.Vout.n14 0.788543
R37169 And_Gate_5.Vout.n1 And_Gate_5.Vout.n0 0.682565
R37170 And_Gate_5.Vout.n1 And_Gate_5.Inverter_0.Vout 0.580578
R37171 And_Gate_5.Inverter_0.Vout And_Gate_5.Vout.n15 0.484875
R37172 And_Gate_5.Vout.n10 D_FlipFlop_1.3-input-nand_1.C 0.447191
R37173 And_Gate_5.Vout.n7 D_FlipFlop_1.Inverter_1.Vin 0.436162
R37174 And_Gate_5.Vout.n5 D_FlipFlop_1.CLK 0.321667
R37175 And_Gate_5.Vout.n6 And_Gate_5.Vout.n5 0.283283
R37176 And_Gate_5.Vout.n2 D_FlipFlop_1.3-input-nand_0.C 0.217464
R37177 And_Gate_5.Vout.n9 D_FlipFlop_1.3-input-nand_1.C 0.149957
R37178 And_Gate_5.Vout.n3 D_FlipFlop_1.3-input-nand_0.C 0.1255
R37179 And_Gate_5.Vout.n0 And_Gate_5.Inverter_0.Vout 0.1255
R37180 And_Gate_5.Vout.n8 D_FlipFlop_1.Inverter_1.Vin 0.117348
R37181 And_Gate_5.Vout.n6 D_FlipFlop_1.CLK 0.071
R37182 And_Gate_5.Vout.n0 And_Gate_5.Inverter_0.Vout 0.063
R37183 And_Gate_5.Vout.n14 And_Gate_5.Vout.n13 0.063
R37184 And_Gate_5.Vout.n13 And_Gate_5.Vout.n1 0.063
R37185 And_Gate_5.Vout.n8 D_FlipFlop_1.Inverter_1.Vin 0.0454219
R37186 And_Gate_5.Vout.n9 D_FlipFlop_1.3-input-nand_1.C 0.0454219
R37187 And_Gate_5.Vout.n12 And_Gate_5.Vout.n6 0.024
R37188 And_Gate_5.Vout.n12 And_Gate_5.Vout.n11 0.024
R37189 And_Gate_5.Vout.n4 And_Gate_5.Vout.n3 0.0216397
R37190 And_Gate_5.Vout.n4 D_FlipFlop_1.3-input-nand_0.C 0.0216397
R37191 And_Gate_5.Vout.n11 D_FlipFlop_1.CLK 0.0104697
R37192 And_Gate_5.Vout.n11 D_FlipFlop_1.CLK 0.0091579
R37193 Q5.n2 Q5.t3 169.46
R37194 Q5.n4 Q5.t1 167.809
R37195 Q5.n2 Q5.t2 167.809
R37196 Q5 Q5.t9 158.585
R37197 Q5 Q5.t4 154.823
R37198 Q5.n14 Q5.t5 150.869
R37199 Q5.t4 Q5.n15 150.869
R37200 Q5.t9 Q5.n9 150.293
R37201 Q5.n16 Q5.n13 137.644
R37202 Q5.n13 Q5 85.5731
R37203 Q5.n15 Q5.t6 74.1352
R37204 Q5.n14 Q5.t7 74.1352
R37205 Q5.n7 Q5.t8 73.6304
R37206 Q5.n0 Q5.t0 60.3809
R37207 Q5.n3 Q5.n2 11.4489
R37208 Q5.n5 Q5.n4 8.21389
R37209 Q5.n13 Q5.n12 3.473
R37210 Q5.n15 Q5.n14 1.66898
R37211 Q5.n1 Q5.n0 1.64452
R37212 Q5.n9 Q5.n8 1.19615
R37213 Q5.n0 Q5 0.848156
R37214 Q5.n9 Q5 0.447191
R37215 Q5.n5 Q5 0.39003
R37216 Q5.n4 Q5.n3 0.280391
R37217 Q5.n3 Q5.n1 0.262643
R37218 Q5.n6 Q5 0.222967
R37219 Q5.n6 Q5.n5 0.206517
R37220 Q5.n11 Q5.n10 0.16735
R37221 Q5.n11 Q5 0.155742
R37222 Q5.n1 Q5 0.1255
R37223 Q5.n8 Q5 0.1255
R37224 Q5.n14 Q5 0.063
R37225 Q5.n1 Q5 0.063
R37226 Q5.n12 Q5.n6 0.024
R37227 Q5.n12 Q5.n11 0.024
R37228 Q5 Q5.n16 0.0168043
R37229 Q5.n16 Q5 0.0122188
R37230 Q5.n8 Q5.n7 0.0107679
R37231 Q5.n7 Q5 0.0107679
R37232 Q5.n10 Q5 0.00441667
R37233 Q5.n10 Q5 0.00406061
R37234 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t3 169.46
R37235 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.t2 167.809
R37236 D_FlipFlop_7.3-input-nand_2.C.n11 D_FlipFlop_7.3-input-nand_2.C.t0 167.809
R37237 D_FlipFlop_7.3-input-nand_2.C.t4 D_FlipFlop_7.3-input-nand_2.C.n13 167.226
R37238 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C.t5 150.273
R37239 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.t4 150.273
R37240 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C.t7 73.6406
R37241 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C.t6 73.6304
R37242 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C.t1 60.4568
R37243 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C.n7 12.3891
R37244 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.n11 11.4489
R37245 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C 1.68257
R37246 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C.n2 1.38365
R37247 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C.n0 1.19615
R37248 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C.n5 1.1717
R37249 D_FlipFlop_7.3-input-nand_2.C.n3 D_FlipFlop_7.3-input-nand_2.C 1.08448
R37250 D_FlipFlop_7.3-input-nand_2.C.n6 D_FlipFlop_7.3-input-nand_2.C 0.932141
R37251 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C 0.720633
R37252 D_FlipFlop_7.3-input-nand_2.C.n13 D_FlipFlop_7.3-input-nand_2.C.n12 0.280391
R37253 D_FlipFlop_7.3-input-nand_2.C.n0 D_FlipFlop_7.3-input-nand_2.C 0.217464
R37254 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C 0.1255
R37255 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C 0.1255
R37256 D_FlipFlop_7.3-input-nand_2.C.n1 D_FlipFlop_7.3-input-nand_2.C 0.1255
R37257 D_FlipFlop_7.3-input-nand_2.C.n10 D_FlipFlop_7.3-input-nand_2.C.n9 0.0874565
R37258 D_FlipFlop_7.3-input-nand_2.C.n7 D_FlipFlop_7.3-input-nand_2.C.n6 0.063
R37259 D_FlipFlop_7.3-input-nand_2.C.n2 D_FlipFlop_7.3-input-nand_2.C 0.063
R37260 D_FlipFlop_7.3-input-nand_2.C.n9 D_FlipFlop_7.3-input-nand_2.C.n8 0.063
R37261 D_FlipFlop_7.3-input-nand_2.C.n8 D_FlipFlop_7.3-input-nand_2.C.n3 0.063
R37262 D_FlipFlop_7.3-input-nand_2.C.n12 D_FlipFlop_7.3-input-nand_2.C.n10 0.0435206
R37263 D_FlipFlop_7.3-input-nand_2.C.n14 D_FlipFlop_7.3-input-nand_2.C.n1 0.0216397
R37264 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.C.n14 0.0216397
R37265 D_FlipFlop_7.3-input-nand_2.C.n5 D_FlipFlop_7.3-input-nand_2.C.n4 0.0107679
R37266 D_FlipFlop_7.3-input-nand_2.C.n4 D_FlipFlop_7.3-input-nand_2.C 0.0107679
R37267 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t1 169.46
R37268 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.t3 167.809
R37269 D_FlipFlop_7.3-input-nand_2.Vout.n9 D_FlipFlop_7.3-input-nand_2.Vout.t0 167.809
R37270 D_FlipFlop_7.3-input-nand_2.Vout.t6 D_FlipFlop_7.3-input-nand_2.Vout.n11 167.227
R37271 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.t6 150.293
R37272 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.t5 150.273
R37273 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout.t7 73.6406
R37274 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout.t4 73.6304
R37275 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout.t2 60.3809
R37276 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n5 12.3891
R37277 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout.n9 11.4489
R37278 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout.n2 1.38365
R37279 D_FlipFlop_7.3-input-nand_2.Vout.n12 D_FlipFlop_7.3-input-nand_2.Vout.n1 1.19615
R37280 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout.n4 1.1717
R37281 D_FlipFlop_7.3-input-nand_2.Vout.n2 D_FlipFlop_7.3-input-nand_2.Vout 0.848156
R37282 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.Vout.n12 0.447191
R37283 D_FlipFlop_7.3-input-nand_2.Vout.n3 D_FlipFlop_7.3-input-nand_2.Vout 0.38637
R37284 D_FlipFlop_7.3-input-nand_2.Vout.n11 D_FlipFlop_7.3-input-nand_2.Vout.n10 0.280391
R37285 D_FlipFlop_7.3-input-nand_2.Vout.n10 D_FlipFlop_7.3-input-nand_2.Vout.n8 0.262643
R37286 D_FlipFlop_7.3-input-nand_2.Vout.n4 D_FlipFlop_7.3-input-nand_2.Vout 0.217464
R37287 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout 0.152844
R37288 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.149957
R37289 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R37290 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout 0.1255
R37291 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout.n7 0.0874565
R37292 D_FlipFlop_7.3-input-nand_2.Vout.n6 D_FlipFlop_7.3-input-nand_2.Vout.n3 0.063
R37293 D_FlipFlop_7.3-input-nand_2.Vout.n7 D_FlipFlop_7.3-input-nand_2.Vout.n6 0.063
R37294 D_FlipFlop_7.3-input-nand_2.Vout.n8 D_FlipFlop_7.3-input-nand_2.Vout 0.063
R37295 D_FlipFlop_7.3-input-nand_2.Vout.n5 D_FlipFlop_7.3-input-nand_2.Vout 0.0454219
R37296 D_FlipFlop_7.3-input-nand_2.Vout.n1 D_FlipFlop_7.3-input-nand_2.Vout.n0 0.0107679
R37297 D_FlipFlop_7.3-input-nand_2.Vout.n0 D_FlipFlop_7.3-input-nand_2.Vout 0.0107679
R37298 Nand_Gate_1.Vout.n0 Nand_Gate_1.Vout.t2 179.256
R37299 Nand_Gate_1.Vout.n0 Nand_Gate_1.Vout.t1 168.089
R37300 Nand_Gate_1.Vout.n3 Nand_Gate_1.Vout.t4 150.293
R37301 Nand_Gate_1.Vout.n5 Nand_Gate_1.Vout.t3 73.6304
R37302 Nand_Gate_1.Vout Nand_Gate_1.Vout.t0 60.3943
R37303 Nand_Gate_1.Vout.n9 Nand_Gate_1.Vout.n8 37.3347
R37304 Nand_Gate_1.Vout.n2 Nand_Gate_1.Vout 0.981478
R37305 Nand_Gate_1.Vout.n2 Nand_Gate_1.Vout.n1 0.788543
R37306 Nand_Gate_1.Vout.n4 Nand_Gate_1.Vout 0.769522
R37307 Nand_Gate_1.Vout.n1 Nand_Gate_1.Vout 0.720633
R37308 Nand_Gate_1.Vout.n11 Nand_Gate_1.Vout.n10 0.682565
R37309 Nand_Gate_1.Vout.n10 Nand_Gate_1.Vout 0.580578
R37310 Nand_Gate_1.Vout.n4 Nand_Gate_1.Vout.n3 0.55213
R37311 Nand_Gate_1.Vout.n7 Nand_Gate_1.Vout.n6 0.470609
R37312 Nand_Gate_1.Vout.n3 Nand_Gate_1.Vout 0.447191
R37313 Nand_Gate_1.Vout.n7 Nand_Gate_1.Vout 0.428234
R37314 Nand_Gate_1.Vout.n6 Nand_Gate_1.Vout 0.1255
R37315 Nand_Gate_1.Vout.n11 Nand_Gate_1.Vout 0.1255
R37316 Nand_Gate_1.Vout.n8 Nand_Gate_1.Vout.n4 0.063
R37317 Nand_Gate_1.Vout.n8 Nand_Gate_1.Vout.n7 0.063
R37318 Nand_Gate_1.Vout.n9 Nand_Gate_1.Vout.n2 0.063
R37319 Nand_Gate_1.Vout.n10 Nand_Gate_1.Vout.n9 0.063
R37320 Nand_Gate_1.Vout Nand_Gate_1.Vout.n11 0.063
R37321 Nand_Gate_1.Vout.n1 Nand_Gate_1.Vout.n0 0.0435206
R37322 Nand_Gate_1.Vout.n6 Nand_Gate_1.Vout.n5 0.0107679
R37323 Nand_Gate_1.Vout.n5 Nand_Gate_1.Vout 0.0107679
R37324 Nand_Gate_7.A.n32 Nand_Gate_7.A.t0 169.46
R37325 Nand_Gate_7.A.n32 Nand_Gate_7.A.t3 167.809
R37326 Nand_Gate_7.A.n34 Nand_Gate_7.A.t1 167.809
R37327 Nand_Gate_7.A Nand_Gate_7.A.t6 158.585
R37328 Nand_Gate_7.A.n20 Nand_Gate_7.A.t9 150.293
R37329 Nand_Gate_7.A.t6 Nand_Gate_7.A.n2 150.293
R37330 Nand_Gate_7.A.n14 Nand_Gate_7.A.t8 150.273
R37331 Nand_Gate_7.A.n8 Nand_Gate_7.A.t5 150.273
R37332 Nand_Gate_7.A.n12 Nand_Gate_7.A.t4 73.6406
R37333 Nand_Gate_7.A.n6 Nand_Gate_7.A.t7 73.6406
R37334 Nand_Gate_7.A.n22 Nand_Gate_7.A.t11 73.6304
R37335 Nand_Gate_7.A.n0 Nand_Gate_7.A.t10 73.6304
R37336 Nand_Gate_7.A.n4 Nand_Gate_7.A.t2 60.3809
R37337 Nand_Gate_7.A.n26 Nand_Gate_7.A.n25 14.3097
R37338 Nand_Gate_7.A.n33 Nand_Gate_7.A.n32 11.4489
R37339 Nand_Gate_7.A.n35 Nand_Gate_7.A.n34 8.21389
R37340 Nand_Gate_7.A.n18 Nand_Gate_7.A.n11 8.1418
R37341 Nand_Gate_7.A.n28 Nand_Gate_7.A.n27 5.61191
R37342 Nand_Gate_7.A.n28 Nand_Gate_7.A 5.3423
R37343 Nand_Gate_7.A.n29 Nand_Gate_7.A.n28 4.563
R37344 Nand_Gate_7.A.n18 Nand_Gate_7.A.n17 4.5005
R37345 Nand_Gate_7.A.n27 Nand_Gate_7.A 1.82115
R37346 Nand_Gate_7.A.n19 Nand_Gate_7.A 1.62007
R37347 Nand_Gate_7.A.n2 Nand_Gate_7.A.n1 1.19615
R37348 Nand_Gate_7.A.n5 Nand_Gate_7.A 1.08746
R37349 Nand_Gate_7.A.n19 Nand_Gate_7.A 1.00726
R37350 Nand_Gate_7.A.n13 Nand_Gate_7.A 0.851043
R37351 Nand_Gate_7.A.n7 Nand_Gate_7.A 0.851043
R37352 Nand_Gate_7.A.n4 Nand_Gate_7.A 0.848156
R37353 Nand_Gate_7.A.n31 Nand_Gate_7.A.n30 0.788543
R37354 Nand_Gate_7.A.n21 Nand_Gate_7.A 0.769522
R37355 Nand_Gate_7.A.n5 Nand_Gate_7.A.n4 0.682565
R37356 Nand_Gate_7.A.n30 Nand_Gate_7.A 0.65675
R37357 Nand_Gate_7.A.n21 Nand_Gate_7.A.n20 0.55213
R37358 Nand_Gate_7.A.n16 Nand_Gate_7.A.n15 0.55213
R37359 Nand_Gate_7.A.n10 Nand_Gate_7.A.n9 0.55213
R37360 Nand_Gate_7.A.n16 Nand_Gate_7.A 0.486828
R37361 Nand_Gate_7.A.n10 Nand_Gate_7.A 0.486828
R37362 Nand_Gate_7.A.n24 Nand_Gate_7.A.n23 0.470609
R37363 Nand_Gate_7.A.n13 Nand_Gate_7.A.n12 0.470609
R37364 Nand_Gate_7.A.n7 Nand_Gate_7.A.n6 0.470609
R37365 Nand_Gate_7.A.n20 Nand_Gate_7.A 0.447191
R37366 Nand_Gate_7.A.n2 Nand_Gate_7.A 0.447191
R37367 Nand_Gate_7.A.n24 Nand_Gate_7.A 0.428234
R37368 Nand_Gate_7.A.n35 Nand_Gate_7.A.n3 0.425067
R37369 Nand_Gate_7.A Nand_Gate_7.A.n35 0.39003
R37370 Nand_Gate_7.A.n34 Nand_Gate_7.A.n33 0.280391
R37371 Nand_Gate_7.A.n33 Nand_Gate_7.A.n31 0.262643
R37372 Nand_Gate_7.A.n12 Nand_Gate_7.A 0.217464
R37373 Nand_Gate_7.A.n6 Nand_Gate_7.A 0.217464
R37374 Nand_Gate_7.A.n23 Nand_Gate_7.A 0.1255
R37375 Nand_Gate_7.A.n15 Nand_Gate_7.A 0.1255
R37376 Nand_Gate_7.A.n9 Nand_Gate_7.A 0.1255
R37377 Nand_Gate_7.A.n31 Nand_Gate_7.A 0.1255
R37378 Nand_Gate_7.A.n1 Nand_Gate_7.A 0.1255
R37379 Nand_Gate_7.A.n25 Nand_Gate_7.A.n21 0.063
R37380 Nand_Gate_7.A.n25 Nand_Gate_7.A.n24 0.063
R37381 Nand_Gate_7.A.n17 Nand_Gate_7.A.n13 0.063
R37382 Nand_Gate_7.A.n17 Nand_Gate_7.A.n16 0.063
R37383 Nand_Gate_7.A.n11 Nand_Gate_7.A.n7 0.063
R37384 Nand_Gate_7.A.n11 Nand_Gate_7.A.n10 0.063
R37385 Nand_Gate_7.A Nand_Gate_7.A.n18 0.063
R37386 Nand_Gate_7.A.n27 Nand_Gate_7.A.n26 0.063
R37387 Nand_Gate_7.A.n26 Nand_Gate_7.A.n19 0.063
R37388 Nand_Gate_7.A.n29 Nand_Gate_7.A.n5 0.063
R37389 Nand_Gate_7.A.n30 Nand_Gate_7.A.n29 0.063
R37390 Nand_Gate_7.A.n31 Nand_Gate_7.A 0.063
R37391 Nand_Gate_7.A.n15 Nand_Gate_7.A.n14 0.0216397
R37392 Nand_Gate_7.A.n14 Nand_Gate_7.A 0.0216397
R37393 Nand_Gate_7.A.n9 Nand_Gate_7.A.n8 0.0216397
R37394 Nand_Gate_7.A.n8 Nand_Gate_7.A 0.0216397
R37395 Nand_Gate_7.A.n23 Nand_Gate_7.A.n22 0.0107679
R37396 Nand_Gate_7.A.n22 Nand_Gate_7.A 0.0107679
R37397 Nand_Gate_7.A.n1 Nand_Gate_7.A.n0 0.0107679
R37398 Nand_Gate_7.A.n0 Nand_Gate_7.A 0.0107679
R37399 Nand_Gate_7.A.n3 Nand_Gate_7.A 0.00441667
R37400 Nand_Gate_7.A.n3 Nand_Gate_7.A 0.00406061
R37401 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.t0 169.46
R37402 D_FlipFlop_5.3-input-nand_2.Vout.n9 D_FlipFlop_5.3-input-nand_2.Vout.t3 167.809
R37403 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout.t2 167.809
R37404 D_FlipFlop_5.3-input-nand_2.Vout.t6 D_FlipFlop_5.3-input-nand_2.Vout.n11 167.227
R37405 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.t6 150.293
R37406 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.t5 150.273
R37407 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout.t7 73.6406
R37408 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout.t4 73.6304
R37409 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout.t1 60.3809
R37410 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout.n5 12.3891
R37411 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n9 11.4489
R37412 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout.n2 1.38365
R37413 D_FlipFlop_5.3-input-nand_2.Vout.n12 D_FlipFlop_5.3-input-nand_2.Vout.n1 1.19615
R37414 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout.n4 1.1717
R37415 D_FlipFlop_5.3-input-nand_2.Vout.n2 D_FlipFlop_5.3-input-nand_2.Vout 0.848156
R37416 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.Vout.n12 0.447191
R37417 D_FlipFlop_5.3-input-nand_2.Vout.n3 D_FlipFlop_5.3-input-nand_2.Vout 0.38637
R37418 D_FlipFlop_5.3-input-nand_2.Vout.n11 D_FlipFlop_5.3-input-nand_2.Vout.n10 0.280391
R37419 D_FlipFlop_5.3-input-nand_2.Vout.n10 D_FlipFlop_5.3-input-nand_2.Vout.n8 0.262643
R37420 D_FlipFlop_5.3-input-nand_2.Vout.n4 D_FlipFlop_5.3-input-nand_2.Vout 0.217464
R37421 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout 0.152844
R37422 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout 0.149957
R37423 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R37424 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout 0.1255
R37425 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout.n7 0.0874565
R37426 D_FlipFlop_5.3-input-nand_2.Vout.n6 D_FlipFlop_5.3-input-nand_2.Vout.n3 0.063
R37427 D_FlipFlop_5.3-input-nand_2.Vout.n7 D_FlipFlop_5.3-input-nand_2.Vout.n6 0.063
R37428 D_FlipFlop_5.3-input-nand_2.Vout.n8 D_FlipFlop_5.3-input-nand_2.Vout 0.063
R37429 D_FlipFlop_5.3-input-nand_2.Vout.n5 D_FlipFlop_5.3-input-nand_2.Vout 0.0454219
R37430 D_FlipFlop_5.3-input-nand_2.Vout.n1 D_FlipFlop_5.3-input-nand_2.Vout.n0 0.0107679
R37431 D_FlipFlop_5.3-input-nand_2.Vout.n0 D_FlipFlop_5.3-input-nand_2.Vout 0.0107679
R37432 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 169.46
R37433 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 168.089
R37434 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 167.809
R37435 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 150.293
R37436 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 73.6304
R37437 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 60.4568
R37438 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 12.0358
R37439 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 11.4489
R37440 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.981478
R37441 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 0.788543
R37442 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.769522
R37443 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 0.720633
R37444 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 0.682565
R37445 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.580578
R37446 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 0.55213
R37447 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 0.470609
R37448 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.447191
R37449 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.428234
R37450 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.1255
R37451 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.1255
R37452 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 0.063
R37453 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 0.063
R37454 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.063
R37455 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 0.063
R37456 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 0.063
R37457 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 0.0435206
R37458 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 0.0107679
R37459 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.0107679
R37460 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 169.46
R37461 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 167.809
R37462 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 167.809
R37463 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 167.227
R37464 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 150.293
R37465 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 150.273
R37466 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 73.6406
R37467 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 73.6304
R37468 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 60.3809
R37469 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 12.3891
R37470 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 11.4489
R37471 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 1.38365
R37472 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 1.19615
R37473 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 1.1717
R37474 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.848156
R37475 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 0.447191
R37476 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.38637
R37477 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 0.280391
R37478 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 0.262643
R37479 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.217464
R37480 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.152844
R37481 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.149957
R37482 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.1255
R37483 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.1255
R37484 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 0.0874565
R37485 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 0.063
R37486 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 0.063
R37487 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.063
R37488 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.0454219
R37489 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 0.0107679
R37490 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.0107679
R37491 And_Gate_2.Vout.n12 And_Gate_2.Vout.t0 168.32
R37492 And_Gate_2.Vout.n4 And_Gate_2.Vout.t4 158.23
R37493 D_FlipFlop_5.CLK And_Gate_2.Vout.t6 158.202
R37494 And_Gate_2.Vout.n5 And_Gate_2.Vout.t5 150.293
R37495 And_Gate_2.Vout.t6 And_Gate_2.Vout.n8 150.293
R37496 And_Gate_2.Vout.t4 And_Gate_2.Vout.n3 150.273
R37497 And_Gate_2.Vout.n1 And_Gate_2.Vout.t7 73.6406
R37498 And_Gate_2.Vout.n7 And_Gate_2.Vout.t3 73.6304
R37499 And_Gate_2.Vout.n6 And_Gate_2.Vout.t2 73.6304
R37500 And_Gate_2.Inverter_0.Vout And_Gate_2.Vout.t1 60.3943
R37501 And_Gate_2.Vout.n12 And_Gate_2.Vout.n11 52.2702
R37502 And_Gate_2.Vout.n7 And_Gate_2.Vout.n6 16.332
R37503 And_Gate_2.Vout.n13 And_Gate_2.Vout.n0 1.62007
R37504 And_Gate_2.Inverter_0.Vout And_Gate_2.Vout.n13 1.25441
R37505 And_Gate_2.Vout.n2 And_Gate_2.Vout.n1 1.19615
R37506 And_Gate_2.Vout.n6 And_Gate_2.Vout.n5 1.1717
R37507 And_Gate_2.Vout.n8 And_Gate_2.Vout.n7 1.1717
R37508 And_Gate_2.Vout.n8 D_FlipFlop_5.3-input-nand_1.C 0.447191
R37509 And_Gate_2.Vout.n5 D_FlipFlop_5.Inverter_1.Vin 0.436162
R37510 And_Gate_2.Vout.n4 D_FlipFlop_5.CLK 0.298879
R37511 And_Gate_2.Vout.n10 And_Gate_2.Vout.n9 0.265267
R37512 And_Gate_2.Vout.n1 D_FlipFlop_5.3-input-nand_0.C 0.217464
R37513 And_Gate_2.Vout.n10 D_FlipFlop_5.CLK 0.212618
R37514 And_Gate_2.Vout.n7 D_FlipFlop_5.3-input-nand_1.C 0.149957
R37515 And_Gate_2.Vout.n2 D_FlipFlop_5.3-input-nand_0.C 0.1255
R37516 And_Gate_2.Vout.n0 And_Gate_2.Inverter_0.Vout 0.1255
R37517 And_Gate_2.Vout.n6 D_FlipFlop_5.Inverter_1.Vin 0.117348
R37518 And_Gate_2.Vout.n0 And_Gate_2.Inverter_0.Vout 0.063
R37519 And_Gate_2.Vout.n13 And_Gate_2.Vout.n12 0.063
R37520 And_Gate_2.Vout.n6 D_FlipFlop_5.Inverter_1.Vin 0.0454219
R37521 And_Gate_2.Vout.n7 D_FlipFlop_5.3-input-nand_1.C 0.0454219
R37522 And_Gate_2.Vout.n11 And_Gate_2.Vout.n4 0.024
R37523 And_Gate_2.Vout.n11 And_Gate_2.Vout.n10 0.024
R37524 And_Gate_2.Vout.n3 And_Gate_2.Vout.n2 0.0216397
R37525 And_Gate_2.Vout.n3 D_FlipFlop_5.3-input-nand_0.C 0.0216397
R37526 And_Gate_2.Vout.n9 D_FlipFlop_5.CLK 0.00441667
R37527 And_Gate_2.Vout.n9 D_FlipFlop_5.CLK 0.00406061
R37528 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 169.46
R37529 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 168.089
R37530 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 167.809
R37531 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 150.293
R37532 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 73.6304
R37533 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 60.3943
R37534 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 12.0358
R37535 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 11.4489
R37536 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.981478
R37537 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 0.788543
R37538 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.769522
R37539 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 0.720633
R37540 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 0.682565
R37541 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.580578
R37542 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 0.55213
R37543 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 0.470609
R37544 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.447191
R37545 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.428234
R37546 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.1255
R37547 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.1255
R37548 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 0.063
R37549 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 0.063
R37550 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.063
R37551 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 0.063
R37552 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 0.063
R37553 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 0.0435206
R37554 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 0.0107679
R37555 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.0107679
R37556 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 169.46
R37557 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 168.089
R37558 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 167.809
R37559 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 150.293
R37560 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 73.6304
R37561 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 60.4568
R37562 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 12.0358
R37563 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 11.4489
R37564 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.981478
R37565 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 0.788543
R37566 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.769522
R37567 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 0.720633
R37568 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 0.682565
R37569 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.580578
R37570 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 0.55213
R37571 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 0.470609
R37572 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.447191
R37573 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.428234
R37574 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.1255
R37575 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.1255
R37576 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 0.063
R37577 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 0.063
R37578 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.063
R37579 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 0.063
R37580 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 0.063
R37581 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 0.0435206
R37582 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 0.0107679
R37583 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.0107679
R37584 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 169.46
R37585 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 167.809
R37586 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 167.809
R37587 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 167.226
R37588 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 150.273
R37589 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 150.273
R37590 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 73.6406
R37591 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 73.6304
R37592 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 60.3943
R37593 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 12.3891
R37594 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 11.4489
R37595 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 1.68257
R37596 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 1.38365
R37597 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 1.19615
R37598 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 1.1717
R37599 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 1.08448
R37600 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.932141
R37601 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.720633
R37602 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 0.280391
R37603 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.217464
R37604 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R37605 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R37606 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.1255
R37607 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 0.0874565
R37608 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 0.063
R37609 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 0.063
R37610 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 0.063
R37611 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 0.063
R37612 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 0.0435206
R37613 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 0.0216397
R37614 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.0216397
R37615 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 0.0107679
R37616 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.0107679
R37617 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 179.256
R37618 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 168.089
R37619 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 150.293
R37620 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 73.6304
R37621 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 60.3943
R37622 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 12.0358
R37623 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.981478
R37624 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 0.788543
R37625 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.769522
R37626 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 0.720633
R37627 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 0.682565
R37628 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.580578
R37629 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 0.55213
R37630 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 0.470609
R37631 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.447191
R37632 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.428234
R37633 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1255
R37634 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1255
R37635 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 0.063
R37636 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 0.063
R37637 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.063
R37638 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 0.063
R37639 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 0.063
R37640 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 0.0435206
R37641 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 0.0107679
R37642 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.0107679
R37643 And_Gate_4.A.n0 And_Gate_4.A.t1 179.256
R37644 And_Gate_4.A.n0 And_Gate_4.A.t2 168.089
R37645 And_Gate_4.A.n3 And_Gate_4.A.t3 150.293
R37646 And_Gate_4.A.n5 And_Gate_4.A.t4 73.6304
R37647 Nand_Gate_0.Vout And_Gate_4.A.t0 60.3943
R37648 And_Gate_4.A.n9 And_Gate_4.A.n8 35.6663
R37649 And_Gate_4.A.n2 Nand_Gate_0.Vout 0.981478
R37650 And_Gate_4.A.n2 And_Gate_4.A.n1 0.788543
R37651 And_Gate_4.A.n4 And_Gate_4.Nand_Gate_0.A 0.769522
R37652 And_Gate_4.A.n1 Nand_Gate_0.Vout 0.720633
R37653 And_Gate_4.A.n11 And_Gate_4.A.n10 0.682565
R37654 And_Gate_4.A.n10 Nand_Gate_0.Vout 0.580578
R37655 And_Gate_4.A.n4 And_Gate_4.A.n3 0.55213
R37656 And_Gate_4.A.n7 And_Gate_4.A.n6 0.470609
R37657 And_Gate_4.A.n3 And_Gate_4.Nand_Gate_0.A 0.447191
R37658 And_Gate_4.A.n7 And_Gate_4.Nand_Gate_0.A 0.428234
R37659 And_Gate_4.A.n6 And_Gate_4.Nand_Gate_0.A 0.1255
R37660 And_Gate_4.A.n11 Nand_Gate_0.Vout 0.1255
R37661 And_Gate_4.A.n8 And_Gate_4.A.n4 0.063
R37662 And_Gate_4.A.n8 And_Gate_4.A.n7 0.063
R37663 And_Gate_4.A.n9 And_Gate_4.A.n2 0.063
R37664 And_Gate_4.A.n10 And_Gate_4.A.n9 0.063
R37665 Nand_Gate_0.Vout And_Gate_4.A.n11 0.063
R37666 And_Gate_4.A.n1 And_Gate_4.A.n0 0.0435206
R37667 And_Gate_4.A.n6 And_Gate_4.A.n5 0.0107679
R37668 And_Gate_4.A.n5 And_Gate_4.Nand_Gate_0.A 0.0107679
R37669 Q2.n5 Q2.t0 169.46
R37670 Q2.n7 Q2.t2 167.809
R37671 Q2.n5 Q2.t3 167.809
R37672 Q2.n11 Q2.t8 155.121
R37673 Q2.n14 Q2.t4 150.869
R37674 Q2.n13 Q2.t5 150.869
R37675 Q2.t8 Q2.n2 150.293
R37676 Q2.n15 Q2.n12 137.644
R37677 Q2 Q2.t6 78.1811
R37678 Q2.n13 Q2.t7 74.1352
R37679 Q2.t6 Q2.n14 74.1352
R37680 Q2.n0 Q2.t9 73.6304
R37681 Q2.n3 Q2.t1 60.3809
R37682 Q2.n12 Q2 38.8494
R37683 Q2.n6 Q2.n5 11.4489
R37684 Q2.n8 Q2.n7 8.21389
R37685 Q2.n11 Q2.n10 1.70018
R37686 Q2.n14 Q2.n13 1.66898
R37687 Q2.n4 Q2.n3 1.64452
R37688 Q2.n2 Q2.n1 1.19615
R37689 Q2.n3 Q2 0.848156
R37690 Q2.n2 Q2 0.447191
R37691 Q2.n8 Q2 0.39003
R37692 Q2.n9 Q2.n8 0.35535
R37693 Q2.n7 Q2.n6 0.280391
R37694 Q2.n6 Q2.n4 0.262643
R37695 Q2.n4 Q2 0.1255
R37696 Q2.n1 Q2 0.1255
R37697 Q2.n9 Q2 0.0741333
R37698 Q2.n13 Q2 0.063
R37699 Q2.n4 Q2 0.063
R37700 Q2.n10 Q2.n9 0.0460197
R37701 Q2.n12 Q2.n11 0.0288742
R37702 Q2.n10 Q2 0.0226455
R37703 Q2 Q2.n15 0.0168043
R37704 Q2.n15 Q2 0.0122188
R37705 Q2.n1 Q2.n0 0.0107679
R37706 Q2.n0 Q2 0.0107679
R37707 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 179.256
R37708 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 168.089
R37709 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 150.293
R37710 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 73.6304
R37711 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 60.4568
R37712 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 12.0358
R37713 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.981478
R37714 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 0.788543
R37715 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.769522
R37716 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 0.720633
R37717 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 0.682565
R37718 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.580578
R37719 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 0.55213
R37720 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 0.470609
R37721 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.447191
R37722 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.428234
R37723 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1255
R37724 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1255
R37725 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 0.063
R37726 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 0.063
R37727 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.063
R37728 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 0.063
R37729 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 0.063
R37730 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 0.0435206
R37731 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 0.0107679
R37732 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.0107679
R37733 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 179.256
R37734 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 168.089
R37735 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 150.293
R37736 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 73.6304
R37737 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 60.4568
R37738 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 12.0358
R37739 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.981478
R37740 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 0.788543
R37741 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.769522
R37742 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 0.720633
R37743 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 0.682565
R37744 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.580578
R37745 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 0.55213
R37746 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 0.470609
R37747 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.447191
R37748 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.428234
R37749 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1255
R37750 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1255
R37751 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 0.063
R37752 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 0.063
R37753 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.063
R37754 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 0.063
R37755 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 0.063
R37756 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 0.0435206
R37757 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 0.0107679
R37758 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.0107679
R37759 Nand_Gate_1.A.n33 Nand_Gate_1.A.t0 169.46
R37760 Nand_Gate_1.A.n33 Nand_Gate_1.A.t1 167.809
R37761 Nand_Gate_1.A.n35 Nand_Gate_1.A.t3 167.809
R37762 Nand_Gate_1.A Nand_Gate_1.A.t6 158.585
R37763 Nand_Gate_1.A.n21 Nand_Gate_1.A.t5 150.293
R37764 Nand_Gate_1.A.t6 Nand_Gate_1.A.n2 150.293
R37765 Nand_Gate_1.A.n14 Nand_Gate_1.A.t4 150.273
R37766 Nand_Gate_1.A.n8 Nand_Gate_1.A.t11 150.273
R37767 Nand_Gate_1.A.n12 Nand_Gate_1.A.t9 73.6406
R37768 Nand_Gate_1.A.n6 Nand_Gate_1.A.t7 73.6406
R37769 Nand_Gate_1.A.n23 Nand_Gate_1.A.t8 73.6304
R37770 Nand_Gate_1.A.n0 Nand_Gate_1.A.t10 73.6304
R37771 Nand_Gate_1.A.n4 Nand_Gate_1.A.t2 60.3809
R37772 Nand_Gate_1.A.n27 Nand_Gate_1.A.n26 14.3097
R37773 Nand_Gate_1.A.n34 Nand_Gate_1.A.n33 11.4489
R37774 Nand_Gate_1.A.n36 Nand_Gate_1.A.n35 8.21389
R37775 Nand_Gate_1.A.n18 Nand_Gate_1.A.n11 8.1418
R37776 Nand_Gate_1.A.n29 Nand_Gate_1.A.n28 5.61191
R37777 Nand_Gate_1.A.n29 Nand_Gate_1.A 5.35402
R37778 Nand_Gate_1.A.n30 Nand_Gate_1.A.n29 4.563
R37779 Nand_Gate_1.A.n18 Nand_Gate_1.A.n17 4.5005
R37780 Nand_Gate_1.A.n28 Nand_Gate_1.A 1.83746
R37781 Nand_Gate_1.A.n20 Nand_Gate_1.A.n19 1.62007
R37782 Nand_Gate_1.A.n2 Nand_Gate_1.A.n1 1.19615
R37783 Nand_Gate_1.A.n5 Nand_Gate_1.A 1.08746
R37784 Nand_Gate_1.A.n20 Nand_Gate_1.A 1.01739
R37785 Nand_Gate_1.A.n13 Nand_Gate_1.A 0.851043
R37786 Nand_Gate_1.A.n7 Nand_Gate_1.A 0.851043
R37787 Nand_Gate_1.A.n4 Nand_Gate_1.A 0.848156
R37788 Nand_Gate_1.A.n32 Nand_Gate_1.A.n31 0.788543
R37789 Nand_Gate_1.A.n22 Nand_Gate_1.A 0.769522
R37790 Nand_Gate_1.A.n5 Nand_Gate_1.A.n4 0.682565
R37791 Nand_Gate_1.A.n31 Nand_Gate_1.A 0.65675
R37792 Nand_Gate_1.A.n22 Nand_Gate_1.A.n21 0.55213
R37793 Nand_Gate_1.A.n16 Nand_Gate_1.A.n15 0.55213
R37794 Nand_Gate_1.A.n10 Nand_Gate_1.A.n9 0.55213
R37795 Nand_Gate_1.A.n16 Nand_Gate_1.A 0.486828
R37796 Nand_Gate_1.A.n10 Nand_Gate_1.A 0.486828
R37797 Nand_Gate_1.A.n25 Nand_Gate_1.A.n24 0.470609
R37798 Nand_Gate_1.A.n13 Nand_Gate_1.A.n12 0.470609
R37799 Nand_Gate_1.A.n7 Nand_Gate_1.A.n6 0.470609
R37800 Nand_Gate_1.A.n21 Nand_Gate_1.A 0.447191
R37801 Nand_Gate_1.A.n2 Nand_Gate_1.A 0.447191
R37802 Nand_Gate_1.A.n25 Nand_Gate_1.A 0.428234
R37803 Nand_Gate_1.A.n36 Nand_Gate_1.A.n3 0.425067
R37804 Nand_Gate_1.A Nand_Gate_1.A.n36 0.39003
R37805 Nand_Gate_1.A.n35 Nand_Gate_1.A.n34 0.280391
R37806 Nand_Gate_1.A.n34 Nand_Gate_1.A.n32 0.262643
R37807 Nand_Gate_1.A.n12 Nand_Gate_1.A 0.217464
R37808 Nand_Gate_1.A.n6 Nand_Gate_1.A 0.217464
R37809 Nand_Gate_1.A.n24 Nand_Gate_1.A 0.1255
R37810 Nand_Gate_1.A.n15 Nand_Gate_1.A 0.1255
R37811 Nand_Gate_1.A.n9 Nand_Gate_1.A 0.1255
R37812 Nand_Gate_1.A.n32 Nand_Gate_1.A 0.1255
R37813 Nand_Gate_1.A.n1 Nand_Gate_1.A 0.1255
R37814 Nand_Gate_1.A.n26 Nand_Gate_1.A.n22 0.063
R37815 Nand_Gate_1.A.n26 Nand_Gate_1.A.n25 0.063
R37816 Nand_Gate_1.A.n17 Nand_Gate_1.A.n13 0.063
R37817 Nand_Gate_1.A.n17 Nand_Gate_1.A.n16 0.063
R37818 Nand_Gate_1.A.n11 Nand_Gate_1.A.n7 0.063
R37819 Nand_Gate_1.A.n11 Nand_Gate_1.A.n10 0.063
R37820 Nand_Gate_1.A.n28 Nand_Gate_1.A.n27 0.063
R37821 Nand_Gate_1.A.n27 Nand_Gate_1.A.n20 0.063
R37822 Nand_Gate_1.A.n30 Nand_Gate_1.A.n5 0.063
R37823 Nand_Gate_1.A.n31 Nand_Gate_1.A.n30 0.063
R37824 Nand_Gate_1.A.n32 Nand_Gate_1.A 0.063
R37825 Nand_Gate_1.A Nand_Gate_1.A.n18 0.0512812
R37826 Nand_Gate_1.A.n15 Nand_Gate_1.A.n14 0.0216397
R37827 Nand_Gate_1.A.n14 Nand_Gate_1.A 0.0216397
R37828 Nand_Gate_1.A.n9 Nand_Gate_1.A.n8 0.0216397
R37829 Nand_Gate_1.A.n8 Nand_Gate_1.A 0.0216397
R37830 Nand_Gate_1.A.n19 Nand_Gate_1.A 0.0168043
R37831 Nand_Gate_1.A.n19 Nand_Gate_1.A 0.0122188
R37832 Nand_Gate_1.A.n24 Nand_Gate_1.A.n23 0.0107679
R37833 Nand_Gate_1.A.n23 Nand_Gate_1.A 0.0107679
R37834 Nand_Gate_1.A.n1 Nand_Gate_1.A.n0 0.0107679
R37835 Nand_Gate_1.A.n0 Nand_Gate_1.A 0.0107679
R37836 Nand_Gate_1.A.n3 Nand_Gate_1.A 0.00441667
R37837 Nand_Gate_1.A.n3 Nand_Gate_1.A 0.00406061
R37838 Q4.n2 Q4.t3 169.46
R37839 Q4.n4 Q4.t2 167.809
R37840 Q4.n2 Q4.t0 167.809
R37841 Q4 Q4.t9 158.585
R37842 Q4.n15 Q4.t8 150.869
R37843 Q4.t9 Q4.n9 150.293
R37844 Q4.n17 Q4.t7 150.273
R37845 Q4.n14 Q4.n13 137.644
R37846 Q4.n13 Q4 85.5731
R37847 Q4.n16 Q4.t4 74.1352
R37848 Q4.n15 Q4.t6 74.1352
R37849 Q4.n7 Q4.t5 73.6304
R37850 Q4.n0 Q4.t1 60.3809
R37851 Q4.n3 Q4.n2 11.4489
R37852 Q4.n5 Q4.n4 8.21389
R37853 Q4 Q4.n17 4.54933
R37854 Q4.n13 Q4.n12 3.473
R37855 Q4.n16 Q4.n15 1.66898
R37856 Q4.n1 Q4.n0 1.64452
R37857 Q4.n9 Q4.n8 1.19615
R37858 Q4.n0 Q4 0.848156
R37859 Q4.n17 Q4.n16 0.55213
R37860 Q4.n9 Q4 0.447191
R37861 Q4.n5 Q4 0.39003
R37862 Q4.n4 Q4.n3 0.280391
R37863 Q4.n3 Q4.n1 0.262643
R37864 Q4.n6 Q4.n5 0.219833
R37865 Q4.n6 Q4 0.20965
R37866 Q4.n11 Q4.n10 0.154033
R37867 Q4.n11 Q4 0.143636
R37868 Q4.n1 Q4 0.1255
R37869 Q4.n8 Q4 0.1255
R37870 Q4.n15 Q4 0.063
R37871 Q4.n1 Q4 0.063
R37872 Q4.n12 Q4.n6 0.024
R37873 Q4.n12 Q4.n11 0.024
R37874 Q4.n14 Q4 0.0168043
R37875 Q4 Q4.n14 0.0122188
R37876 Q4.n8 Q4.n7 0.0107679
R37877 Q4.n7 Q4 0.0107679
R37878 Q4.n10 Q4 0.00441667
R37879 Q4.n10 Q4 0.00406061
R37880 And_Gate_6.Vout.n14 And_Gate_6.Vout.t0 168.108
R37881 And_Gate_6.Vout.n5 And_Gate_6.Vout.t2 158.207
R37882 D_FlipFlop_3.CLK And_Gate_6.Vout.t4 158.202
R37883 And_Gate_6.Vout.n7 And_Gate_6.Vout.t3 150.293
R37884 And_Gate_6.Vout.t4 And_Gate_6.Vout.n10 150.293
R37885 And_Gate_6.Vout.t2 And_Gate_6.Vout.n4 150.273
R37886 And_Gate_6.Vout.n2 And_Gate_6.Vout.t5 73.6406
R37887 And_Gate_6.Vout.n9 And_Gate_6.Vout.t7 73.6304
R37888 And_Gate_6.Vout.n8 And_Gate_6.Vout.t6 73.6304
R37889 And_Gate_6.Inverter_0.Vout And_Gate_6.Vout.t1 60.3943
R37890 And_Gate_6.Vout.n12 And_Gate_6.Vout.n11 42.3602
R37891 And_Gate_6.Vout.n9 And_Gate_6.Vout.n8 16.332
R37892 And_Gate_6.Vout.n3 And_Gate_6.Vout.n2 1.19615
R37893 And_Gate_6.Vout.n8 And_Gate_6.Vout.n7 1.1717
R37894 And_Gate_6.Vout.n10 And_Gate_6.Vout.n9 1.1717
R37895 And_Gate_6.Vout.n13 And_Gate_6.Inverter_0.Vout 0.981478
R37896 And_Gate_6.Vout.n14 And_Gate_6.Vout.n13 0.788543
R37897 And_Gate_6.Vout.n1 And_Gate_6.Vout.n0 0.682565
R37898 And_Gate_6.Vout.n1 And_Gate_6.Inverter_0.Vout 0.580578
R37899 And_Gate_6.Inverter_0.Vout And_Gate_6.Vout.n14 0.484875
R37900 And_Gate_6.Vout.n10 D_FlipFlop_3.3-input-nand_1.C 0.447191
R37901 And_Gate_6.Vout.n7 D_FlipFlop_3.Inverter_1.Vin 0.436162
R37902 And_Gate_6.Vout.n5 D_FlipFlop_3.CLK 0.321667
R37903 And_Gate_6.Vout.n6 And_Gate_6.Vout.n5 0.29425
R37904 And_Gate_6.Vout.n2 D_FlipFlop_3.3-input-nand_0.C 0.217464
R37905 And_Gate_6.Vout.n9 D_FlipFlop_3.3-input-nand_1.C 0.149957
R37906 And_Gate_6.Vout.n3 D_FlipFlop_3.3-input-nand_0.C 0.1255
R37907 And_Gate_6.Vout.n0 And_Gate_6.Inverter_0.Vout 0.1255
R37908 And_Gate_6.Vout.n8 D_FlipFlop_3.Inverter_1.Vin 0.117348
R37909 And_Gate_6.Vout.n0 And_Gate_6.Inverter_0.Vout 0.063
R37910 And_Gate_6.Vout.n13 And_Gate_6.Vout.n12 0.063
R37911 And_Gate_6.Vout.n12 And_Gate_6.Vout.n1 0.063
R37912 And_Gate_6.Vout.n6 D_FlipFlop_3.CLK 0.0600333
R37913 And_Gate_6.Vout.n8 D_FlipFlop_3.Inverter_1.Vin 0.0454219
R37914 And_Gate_6.Vout.n9 D_FlipFlop_3.3-input-nand_1.C 0.0454219
R37915 And_Gate_6.Vout.n11 And_Gate_6.Vout.n6 0.024
R37916 And_Gate_6.Vout.n11 D_FlipFlop_3.CLK 0.024
R37917 And_Gate_6.Vout.n4 And_Gate_6.Vout.n3 0.0216397
R37918 And_Gate_6.Vout.n4 D_FlipFlop_3.3-input-nand_0.C 0.0216397
R37919 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 169.46
R37920 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 168.089
R37921 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 167.809
R37922 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 150.273
R37923 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 73.6406
R37924 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 60.3809
R37925 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 12.0358
R37926 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 11.4489
R37927 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 1.08746
R37928 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.851043
R37929 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.848156
R37930 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 0.788543
R37931 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 0.682565
R37932 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.65675
R37933 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 0.55213
R37934 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.486828
R37935 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 0.470609
R37936 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 0.262643
R37937 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.217464
R37938 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.1255
R37939 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.1255
R37940 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 0.063
R37941 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 0.063
R37942 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 0.063
R37943 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 0.063
R37944 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 0.063
R37945 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 0.0216397
R37946 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0216397
R37947 And_Gate_0.Vout.n12 And_Gate_0.Vout.t0 168.32
R37948 And_Gate_0.Vout.n4 And_Gate_0.Vout.t5 158.246
R37949 D_FlipFlop_6.CLK And_Gate_0.Vout.t7 158.202
R37950 And_Gate_0.Vout.n5 And_Gate_0.Vout.t6 150.293
R37951 And_Gate_0.Vout.t7 And_Gate_0.Vout.n8 150.293
R37952 And_Gate_0.Vout.t5 And_Gate_0.Vout.n3 150.273
R37953 And_Gate_0.Vout.n1 And_Gate_0.Vout.t4 73.6406
R37954 And_Gate_0.Vout.n7 And_Gate_0.Vout.t3 73.6304
R37955 And_Gate_0.Vout.n6 And_Gate_0.Vout.t2 73.6304
R37956 And_Gate_0.Vout.n12 And_Gate_0.Vout.n11 66.7548
R37957 And_Gate_0.Inverter_0.Vout And_Gate_0.Vout.t1 60.3943
R37958 And_Gate_0.Vout.n7 And_Gate_0.Vout.n6 16.332
R37959 And_Gate_0.Vout.n13 And_Gate_0.Vout.n0 1.62007
R37960 And_Gate_0.Inverter_0.Vout And_Gate_0.Vout.n13 1.25441
R37961 And_Gate_0.Vout.n2 And_Gate_0.Vout.n1 1.19615
R37962 And_Gate_0.Vout.n6 And_Gate_0.Vout.n5 1.1717
R37963 And_Gate_0.Vout.n8 And_Gate_0.Vout.n7 1.1717
R37964 And_Gate_0.Vout.n8 D_FlipFlop_6.3-input-nand_1.C 0.447191
R37965 And_Gate_0.Vout.n5 D_FlipFlop_6.Inverter_1.Vin 0.436162
R37966 And_Gate_0.Vout.n4 D_FlipFlop_6.CLK 0.281076
R37967 And_Gate_0.Vout.n10 And_Gate_0.Vout.n9 0.245683
R37968 And_Gate_0.Vout.n1 D_FlipFlop_6.3-input-nand_0.C 0.217464
R37969 And_Gate_0.Vout.n10 D_FlipFlop_6.CLK 0.197158
R37970 And_Gate_0.Vout.n7 D_FlipFlop_6.3-input-nand_1.C 0.149957
R37971 And_Gate_0.Vout.n2 D_FlipFlop_6.3-input-nand_0.C 0.1255
R37972 And_Gate_0.Vout.n0 And_Gate_0.Inverter_0.Vout 0.1255
R37973 And_Gate_0.Vout.n6 D_FlipFlop_6.Inverter_1.Vin 0.117348
R37974 And_Gate_0.Vout.n0 And_Gate_0.Inverter_0.Vout 0.063
R37975 And_Gate_0.Vout.n13 And_Gate_0.Vout.n12 0.063
R37976 And_Gate_0.Vout.n6 D_FlipFlop_6.Inverter_1.Vin 0.0454219
R37977 And_Gate_0.Vout.n7 D_FlipFlop_6.3-input-nand_1.C 0.0454219
R37978 And_Gate_0.Vout.n11 And_Gate_0.Vout.n4 0.024
R37979 And_Gate_0.Vout.n11 And_Gate_0.Vout.n10 0.024
R37980 And_Gate_0.Vout.n3 And_Gate_0.Vout.n2 0.0216397
R37981 And_Gate_0.Vout.n3 D_FlipFlop_6.3-input-nand_0.C 0.0216397
R37982 And_Gate_0.Vout.n9 D_FlipFlop_6.CLK 0.00441667
R37983 And_Gate_0.Vout.n9 D_FlipFlop_6.CLK 0.00406061
R37984 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 169.46
R37985 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 167.809
R37986 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 167.809
R37987 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 167.226
R37988 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 150.273
R37989 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 150.273
R37990 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 73.6406
R37991 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 73.6304
R37992 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 60.4568
R37993 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 12.3891
R37994 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 11.4489
R37995 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.68257
R37996 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 1.38365
R37997 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 1.19615
R37998 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 1.1717
R37999 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.08448
R38000 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.932141
R38001 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.720633
R38002 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 0.280391
R38003 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.217464
R38004 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R38005 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R38006 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.1255
R38007 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 0.0874565
R38008 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 0.063
R38009 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 0.063
R38010 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 0.063
R38011 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 0.063
R38012 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 0.0435206
R38013 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 0.0216397
R38014 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.0216397
R38015 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 0.0107679
R38016 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.0107679
R38017 And_Gate_5.A.n0 And_Gate_5.A.t2 179.256
R38018 And_Gate_5.A.n0 And_Gate_5.A.t1 168.089
R38019 And_Gate_5.A.n3 And_Gate_5.A.t4 150.293
R38020 And_Gate_5.A.n5 And_Gate_5.A.t3 73.6304
R38021 Nand_Gate_3.Vout And_Gate_5.A.t0 60.3943
R38022 And_Gate_5.A.n9 And_Gate_5.A.n8 35.6663
R38023 And_Gate_5.A.n2 Nand_Gate_3.Vout 0.981478
R38024 And_Gate_5.A.n2 And_Gate_5.A.n1 0.788543
R38025 And_Gate_5.A.n4 And_Gate_5.Nand_Gate_0.A 0.769522
R38026 And_Gate_5.A.n1 Nand_Gate_3.Vout 0.720633
R38027 And_Gate_5.A.n11 And_Gate_5.A.n10 0.682565
R38028 And_Gate_5.A.n10 Nand_Gate_3.Vout 0.580578
R38029 And_Gate_5.A.n4 And_Gate_5.A.n3 0.55213
R38030 And_Gate_5.A.n7 And_Gate_5.A.n6 0.470609
R38031 And_Gate_5.A.n3 And_Gate_5.Nand_Gate_0.A 0.447191
R38032 And_Gate_5.A.n7 And_Gate_5.Nand_Gate_0.A 0.428234
R38033 And_Gate_5.A.n6 And_Gate_5.Nand_Gate_0.A 0.1255
R38034 And_Gate_5.A.n11 Nand_Gate_3.Vout 0.1255
R38035 And_Gate_5.A.n8 And_Gate_5.A.n4 0.063
R38036 And_Gate_5.A.n8 And_Gate_5.A.n7 0.063
R38037 And_Gate_5.A.n9 And_Gate_5.A.n2 0.063
R38038 And_Gate_5.A.n10 And_Gate_5.A.n9 0.063
R38039 Nand_Gate_3.Vout And_Gate_5.A.n11 0.063
R38040 And_Gate_5.A.n1 And_Gate_5.A.n0 0.0435206
R38041 And_Gate_5.A.n6 And_Gate_5.A.n5 0.0107679
R38042 And_Gate_5.A.n5 And_Gate_5.Nand_Gate_0.A 0.0107679
R38043 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 169.46
R38044 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 168.089
R38045 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 167.809
R38046 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 150.273
R38047 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 73.6406
R38048 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 60.3809
R38049 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 12.0358
R38050 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 11.4489
R38051 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 1.08746
R38052 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.851043
R38053 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.848156
R38054 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 0.788543
R38055 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 0.682565
R38056 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.65675
R38057 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 0.55213
R38058 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.486828
R38059 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 0.470609
R38060 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 0.262643
R38061 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.217464
R38062 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.1255
R38063 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.1255
R38064 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 0.063
R38065 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 0.063
R38066 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 0.063
R38067 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 0.063
R38068 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 0.063
R38069 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 0.0216397
R38070 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0216397
R38071 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 169.46
R38072 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 168.089
R38073 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 167.809
R38074 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 150.273
R38075 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 73.6406
R38076 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 60.3809
R38077 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 12.0358
R38078 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 11.4489
R38079 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 1.08746
R38080 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.851043
R38081 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.848156
R38082 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 0.788543
R38083 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 0.682565
R38084 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.65675
R38085 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 0.55213
R38086 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.486828
R38087 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 0.470609
R38088 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 0.262643
R38089 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.217464
R38090 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.1255
R38091 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.1255
R38092 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 0.063
R38093 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 0.063
R38094 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 0.063
R38095 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 0.063
R38096 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 0.063
R38097 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 0.0216397
R38098 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.0216397
R38099 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 169.46
R38100 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 168.089
R38101 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 167.809
R38102 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 150.293
R38103 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 73.6304
R38104 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 60.3943
R38105 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 12.0358
R38106 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 11.4489
R38107 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.981478
R38108 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 0.788543
R38109 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.769522
R38110 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 0.720633
R38111 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 0.682565
R38112 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.580578
R38113 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 0.55213
R38114 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 0.470609
R38115 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.447191
R38116 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.428234
R38117 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.1255
R38118 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.1255
R38119 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 0.063
R38120 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 0.063
R38121 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.063
R38122 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 0.063
R38123 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 0.063
R38124 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 0.0435206
R38125 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 0.0107679
R38126 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.0107679
R38127 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t0 169.46
R38128 D_FlipFlop_4.3-input-nand_2.Vout.n9 D_FlipFlop_4.3-input-nand_2.Vout.t1 167.809
R38129 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.t2 167.809
R38130 D_FlipFlop_4.3-input-nand_2.Vout.t7 D_FlipFlop_4.3-input-nand_2.Vout.n11 167.227
R38131 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.t7 150.293
R38132 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.t5 150.273
R38133 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6406
R38134 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout.t4 73.6304
R38135 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout.t3 60.3809
R38136 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n5 12.3891
R38137 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout.n9 11.4489
R38138 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout.n2 1.38365
R38139 D_FlipFlop_4.3-input-nand_2.Vout.n12 D_FlipFlop_4.3-input-nand_2.Vout.n1 1.19615
R38140 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout.n4 1.1717
R38141 D_FlipFlop_4.3-input-nand_2.Vout.n2 D_FlipFlop_4.3-input-nand_2.Vout 0.848156
R38142 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.Vout.n12 0.447191
R38143 D_FlipFlop_4.3-input-nand_2.Vout.n3 D_FlipFlop_4.3-input-nand_2.Vout 0.38637
R38144 D_FlipFlop_4.3-input-nand_2.Vout.n11 D_FlipFlop_4.3-input-nand_2.Vout.n10 0.280391
R38145 D_FlipFlop_4.3-input-nand_2.Vout.n10 D_FlipFlop_4.3-input-nand_2.Vout.n8 0.262643
R38146 D_FlipFlop_4.3-input-nand_2.Vout.n4 D_FlipFlop_4.3-input-nand_2.Vout 0.217464
R38147 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R38148 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R38149 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R38150 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R38151 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout.n7 0.0874565
R38152 D_FlipFlop_4.3-input-nand_2.Vout.n6 D_FlipFlop_4.3-input-nand_2.Vout.n3 0.063
R38153 D_FlipFlop_4.3-input-nand_2.Vout.n7 D_FlipFlop_4.3-input-nand_2.Vout.n6 0.063
R38154 D_FlipFlop_4.3-input-nand_2.Vout.n8 D_FlipFlop_4.3-input-nand_2.Vout 0.063
R38155 D_FlipFlop_4.3-input-nand_2.Vout.n5 D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R38156 D_FlipFlop_4.3-input-nand_2.Vout.n1 D_FlipFlop_4.3-input-nand_2.Vout.n0 0.0107679
R38157 D_FlipFlop_4.3-input-nand_2.Vout.n0 D_FlipFlop_4.3-input-nand_2.Vout 0.0107679
R38158 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C.t3 169.46
R38159 D_FlipFlop_4.3-input-nand_2.C.n4 D_FlipFlop_4.3-input-nand_2.C.t2 167.809
R38160 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C.t1 167.809
R38161 D_FlipFlop_4.3-input-nand_2.C.n3 D_FlipFlop_4.3-input-nand_2.C.t4 167.226
R38162 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.t6 150.273
R38163 D_FlipFlop_4.3-input-nand_2.C.t4 D_FlipFlop_4.3-input-nand_2.C.n2 150.273
R38164 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C.t5 73.6406
R38165 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C.t7 73.6304
R38166 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.t0 60.4568
R38167 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.n11 12.3891
R38168 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C.n4 11.4489
R38169 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C 1.68257
R38170 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C.n13 1.38365
R38171 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C.n0 1.19615
R38172 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C.n9 1.1717
R38173 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C 1.08448
R38174 D_FlipFlop_4.3-input-nand_2.C.n10 D_FlipFlop_4.3-input-nand_2.C 0.932141
R38175 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C 0.720633
R38176 D_FlipFlop_4.3-input-nand_2.C.n5 D_FlipFlop_4.3-input-nand_2.C.n3 0.280391
R38177 D_FlipFlop_4.3-input-nand_2.C.n0 D_FlipFlop_4.3-input-nand_2.C 0.217464
R38178 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C 0.1255
R38179 D_FlipFlop_4.3-input-nand_2.C.n1 D_FlipFlop_4.3-input-nand_2.C 0.1255
R38180 D_FlipFlop_4.3-input-nand_2.C.n14 D_FlipFlop_4.3-input-nand_2.C 0.1255
R38181 D_FlipFlop_4.3-input-nand_2.C.n7 D_FlipFlop_4.3-input-nand_2.C.n6 0.0874565
R38182 D_FlipFlop_4.3-input-nand_2.C.n11 D_FlipFlop_4.3-input-nand_2.C.n10 0.063
R38183 D_FlipFlop_4.3-input-nand_2.C.n12 D_FlipFlop_4.3-input-nand_2.C.n7 0.063
R38184 D_FlipFlop_4.3-input-nand_2.C.n13 D_FlipFlop_4.3-input-nand_2.C.n12 0.063
R38185 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_2.C.n14 0.063
R38186 D_FlipFlop_4.3-input-nand_2.C.n6 D_FlipFlop_4.3-input-nand_2.C.n5 0.0435206
R38187 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C.n1 0.0216397
R38188 D_FlipFlop_4.3-input-nand_2.C.n2 D_FlipFlop_4.3-input-nand_2.C 0.0216397
R38189 D_FlipFlop_4.3-input-nand_2.C.n9 D_FlipFlop_4.3-input-nand_2.C.n8 0.0107679
R38190 D_FlipFlop_4.3-input-nand_2.C.n8 D_FlipFlop_4.3-input-nand_2.C 0.0107679
R38191 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 179.256
R38192 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 168.089
R38193 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 150.293
R38194 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 73.6304
R38195 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 60.4568
R38196 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 12.0358
R38197 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.981478
R38198 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 0.788543
R38199 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.769522
R38200 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.720633
R38201 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 0.682565
R38202 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.580578
R38203 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 0.55213
R38204 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 0.470609
R38205 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.447191
R38206 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.428234
R38207 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1255
R38208 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1255
R38209 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 0.063
R38210 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 0.063
R38211 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 0.063
R38212 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 0.063
R38213 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 0.063
R38214 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 0.0435206
R38215 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 0.0107679
R38216 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.0107679
R38217 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z.t1 168.609
R38218 CDAC8_0.switch_0.Z CDAC8_0.switch_0.Z.t2 168.565
R38219 CDAC8_0.switch_0.Z.n6 CDAC8_0.switch_0.Z.t3 60.321
R38220 CDAC8_0.switch_0.Z.n6 CDAC8_0.switch_0.Z.t0 60.321
R38221 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z.n4 11.3205
R38222 CDAC8_0.switch_0.Z.n2 CDAC8_0.switch_0.Z.n1 5.58885
R38223 CDAC8_0.switch_0.Z.n4 CDAC8_0.switch_0.Z.n0 2.98587
R38224 CDAC8_0.switch_0.Z.n4 CDAC8_0.switch_0.Z.n3 2.5049
R38225 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z.n5 1.60376
R38226 CDAC8_0.switch_0.Z.n0 CDAC8_0.switch_0.Z.t5 0.658247
R38227 CDAC8_0.switch_0.Z.n3 CDAC8_0.switch_0.Z.t7 0.658247
R38228 CDAC8_0.switch_0.Z.n1 CDAC8_0.switch_0.Z.t6 0.611304
R38229 CDAC8_0.switch_0.Z.n2 CDAC8_0.switch_0.Z.t4 0.611304
R38230 CDAC8_0.switch_0.Z CDAC8_0.switch_0.Z.n7 0.259656
R38231 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z 0.166261
R38232 CDAC8_0.switch_0.Z.n3 CDAC8_0.switch_0.Z.n2 0.115412
R38233 CDAC8_0.switch_0.Z.n1 CDAC8_0.switch_0.Z.n0 0.115412
R38234 CDAC8_0.switch_0.Z.n5 CDAC8_0.switch_0.Z 0.0454219
R38235 CDAC8_0.switch_0.Z.n7 CDAC8_0.switch_0.Z.n6 0.0188121
R38236 RingCounter_0.D_FlipFlop_16.Q.n19 RingCounter_0.D_FlipFlop_16.Q.t0 169.46
R38237 RingCounter_0.D_FlipFlop_16.Q.n19 RingCounter_0.D_FlipFlop_16.Q.t3 167.809
R38238 RingCounter_0.D_FlipFlop_16.Q.n21 RingCounter_0.D_FlipFlop_16.Q.t2 167.809
R38239 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Q.t8 158.585
R38240 RingCounter_0.D_FlipFlop_16.Q.t8 RingCounter_0.D_FlipFlop_16.Q.n2 150.293
R38241 RingCounter_0.D_FlipFlop_16.Q.n12 RingCounter_0.D_FlipFlop_16.Q.t7 150.273
R38242 RingCounter_0.D_FlipFlop_16.Q.n6 RingCounter_0.D_FlipFlop_16.Q.t6 150.273
R38243 RingCounter_0.D_FlipFlop_16.Q.n10 RingCounter_0.D_FlipFlop_16.Q.t9 73.6406
R38244 RingCounter_0.D_FlipFlop_16.Q.n4 RingCounter_0.D_FlipFlop_16.Q.t4 73.6406
R38245 RingCounter_0.D_FlipFlop_16.Q.n0 RingCounter_0.D_FlipFlop_16.Q.t5 73.6304
R38246 RingCounter_0.D_FlipFlop_16.Q.n22 RingCounter_0.D_FlipFlop_16.Q.n16 62.8776
R38247 RingCounter_0.D_FlipFlop_16.Q.n17 RingCounter_0.D_FlipFlop_16.Q.t1 60.3809
R38248 RingCounter_0.D_FlipFlop_16.Q.n20 RingCounter_0.D_FlipFlop_16.Q.n19 11.4489
R38249 RingCounter_0.D_FlipFlop_16.Q.n22 RingCounter_0.D_FlipFlop_16.Q.n21 8.19039
R38250 RingCounter_0.D_FlipFlop_16.Q.n16 RingCounter_0.D_FlipFlop_16.Q.n9 8.1418
R38251 RingCounter_0.D_FlipFlop_16.Q.n16 RingCounter_0.D_FlipFlop_16.Q.n15 4.5005
R38252 RingCounter_0.D_FlipFlop_16.Q.n18 RingCounter_0.D_FlipFlop_16.Q.n17 1.64452
R38253 RingCounter_0.D_FlipFlop_16.Q.n2 RingCounter_0.D_FlipFlop_16.Q.n1 1.19615
R38254 RingCounter_0.D_FlipFlop_16.Q.n11 RingCounter_0.D_FlipFlop_16.Q 0.851043
R38255 RingCounter_0.D_FlipFlop_16.Q.n5 RingCounter_0.D_FlipFlop_16.Q 0.851043
R38256 RingCounter_0.D_FlipFlop_16.Q.n17 RingCounter_0.D_FlipFlop_16.Q 0.848156
R38257 RingCounter_0.D_FlipFlop_16.Q.n14 RingCounter_0.D_FlipFlop_16.Q.n13 0.55213
R38258 RingCounter_0.D_FlipFlop_16.Q.n8 RingCounter_0.D_FlipFlop_16.Q.n7 0.55213
R38259 RingCounter_0.D_FlipFlop_16.Q.n14 RingCounter_0.D_FlipFlop_16.Q 0.486828
R38260 RingCounter_0.D_FlipFlop_16.Q.n8 RingCounter_0.D_FlipFlop_16.Q 0.486828
R38261 RingCounter_0.D_FlipFlop_16.Q.n11 RingCounter_0.D_FlipFlop_16.Q.n10 0.470609
R38262 RingCounter_0.D_FlipFlop_16.Q.n5 RingCounter_0.D_FlipFlop_16.Q.n4 0.470609
R38263 RingCounter_0.D_FlipFlop_16.Q.n2 RingCounter_0.D_FlipFlop_16.Q 0.447191
R38264 RingCounter_0.D_FlipFlop_16.Q.n23 RingCounter_0.D_FlipFlop_16.Q.n3 0.425067
R38265 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Q.n23 0.39003
R38266 RingCounter_0.D_FlipFlop_16.Q.n21 RingCounter_0.D_FlipFlop_16.Q.n20 0.280391
R38267 RingCounter_0.D_FlipFlop_16.Q.n20 RingCounter_0.D_FlipFlop_16.Q.n18 0.262643
R38268 RingCounter_0.D_FlipFlop_16.Q.n10 RingCounter_0.D_FlipFlop_16.Q 0.217464
R38269 RingCounter_0.D_FlipFlop_16.Q.n4 RingCounter_0.D_FlipFlop_16.Q 0.217464
R38270 RingCounter_0.D_FlipFlop_16.Q.n18 RingCounter_0.D_FlipFlop_16.Q 0.1255
R38271 RingCounter_0.D_FlipFlop_16.Q.n13 RingCounter_0.D_FlipFlop_16.Q 0.1255
R38272 RingCounter_0.D_FlipFlop_16.Q.n7 RingCounter_0.D_FlipFlop_16.Q 0.1255
R38273 RingCounter_0.D_FlipFlop_16.Q.n1 RingCounter_0.D_FlipFlop_16.Q 0.1255
R38274 RingCounter_0.D_FlipFlop_16.Q.n18 RingCounter_0.D_FlipFlop_16.Q 0.063
R38275 RingCounter_0.D_FlipFlop_16.Q.n15 RingCounter_0.D_FlipFlop_16.Q.n11 0.063
R38276 RingCounter_0.D_FlipFlop_16.Q.n15 RingCounter_0.D_FlipFlop_16.Q.n14 0.063
R38277 RingCounter_0.D_FlipFlop_16.Q.n9 RingCounter_0.D_FlipFlop_16.Q.n5 0.063
R38278 RingCounter_0.D_FlipFlop_16.Q.n9 RingCounter_0.D_FlipFlop_16.Q.n8 0.063
R38279 RingCounter_0.D_FlipFlop_16.Q.n23 RingCounter_0.D_FlipFlop_16.Q.n22 0.024
R38280 RingCounter_0.D_FlipFlop_16.Q.n13 RingCounter_0.D_FlipFlop_16.Q.n12 0.0216397
R38281 RingCounter_0.D_FlipFlop_16.Q.n12 RingCounter_0.D_FlipFlop_16.Q 0.0216397
R38282 RingCounter_0.D_FlipFlop_16.Q.n7 RingCounter_0.D_FlipFlop_16.Q.n6 0.0216397
R38283 RingCounter_0.D_FlipFlop_16.Q.n6 RingCounter_0.D_FlipFlop_16.Q 0.0216397
R38284 RingCounter_0.D_FlipFlop_16.Q.n1 RingCounter_0.D_FlipFlop_16.Q.n0 0.0107679
R38285 RingCounter_0.D_FlipFlop_16.Q.n0 RingCounter_0.D_FlipFlop_16.Q 0.0107679
R38286 RingCounter_0.D_FlipFlop_16.Q.n3 RingCounter_0.D_FlipFlop_16.Q 0.00441667
R38287 RingCounter_0.D_FlipFlop_16.Q.n3 RingCounter_0.D_FlipFlop_16.Q 0.00406061
R38288 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 316.762
R38289 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 168.108
R38290 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 150.293
R38291 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 150.273
R38292 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 73.6406
R38293 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 73.6304
R38294 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 60.3943
R38295 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 12.0358
R38296 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 1.19615
R38297 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.981478
R38298 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 0.788543
R38299 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.769522
R38300 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 0.682565
R38301 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.580578
R38302 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 0.55213
R38303 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 0.484875
R38304 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 0.470609
R38305 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.447191
R38306 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.428234
R38307 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.217464
R38308 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R38309 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R38310 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.1255
R38311 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 0.063
R38312 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 0.063
R38313 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.063
R38314 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 0.063
R38315 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 0.063
R38316 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 0.0216397
R38317 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.0216397
R38318 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 0.0107679
R38319 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.0107679
R38320 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 179.256
R38321 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 168.089
R38322 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 150.273
R38323 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 73.6406
R38324 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 60.3809
R38325 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 12.0358
R38326 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 1.08746
R38327 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.851043
R38328 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.848156
R38329 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 0.788543
R38330 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 0.682565
R38331 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.65675
R38332 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 0.55213
R38333 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.486828
R38334 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 0.470609
R38335 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.217464
R38336 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 0.200143
R38337 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.1255
R38338 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.1255
R38339 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 0.063
R38340 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 0.063
R38341 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 0.063
R38342 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 0.063
R38343 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 0.063
R38344 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 0.0216397
R38345 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.0216397
R38346 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 316.762
R38347 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 168.108
R38348 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 150.293
R38349 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 150.273
R38350 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 73.6406
R38351 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 73.6304
R38352 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 60.3943
R38353 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 12.0358
R38354 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 1.19615
R38355 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.981478
R38356 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 0.788543
R38357 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.769522
R38358 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 0.682565
R38359 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.580578
R38360 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 0.55213
R38361 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 0.484875
R38362 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 0.470609
R38363 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.447191
R38364 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.428234
R38365 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.217464
R38366 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R38367 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R38368 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.1255
R38369 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 0.063
R38370 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 0.063
R38371 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.063
R38372 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 0.063
R38373 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 0.063
R38374 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 0.0216397
R38375 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.0216397
R38376 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 0.0107679
R38377 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.0107679
R38378 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 169.46
R38379 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 167.809
R38380 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 167.809
R38381 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 167.226
R38382 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 150.273
R38383 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 150.273
R38384 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 73.6406
R38385 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 73.6304
R38386 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 60.4568
R38387 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 12.3891
R38388 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 11.4489
R38389 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.68257
R38390 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 1.38365
R38391 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 1.19615
R38392 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 1.1717
R38393 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.08448
R38394 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.932141
R38395 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.720633
R38396 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 0.280391
R38397 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.217464
R38398 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R38399 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R38400 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.1255
R38401 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 0.0874565
R38402 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 0.063
R38403 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.063
R38404 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 0.063
R38405 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 0.063
R38406 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 0.0435206
R38407 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 0.0216397
R38408 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 0.0216397
R38409 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 0.0107679
R38410 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.0107679
R38411 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 169.46
R38412 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 168.089
R38413 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 167.809
R38414 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 150.293
R38415 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 73.6304
R38416 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 60.3943
R38417 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 12.0358
R38418 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 11.4489
R38419 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.981478
R38420 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 0.788543
R38421 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.769522
R38422 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 0.720633
R38423 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 0.682565
R38424 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.580578
R38425 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 0.55213
R38426 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 0.470609
R38427 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.447191
R38428 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.428234
R38429 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.1255
R38430 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.1255
R38431 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 0.063
R38432 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 0.063
R38433 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.063
R38434 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 0.063
R38435 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 0.063
R38436 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 0.0435206
R38437 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 0.0107679
R38438 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.0107679
R38439 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 169.46
R38440 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 168.089
R38441 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 167.809
R38442 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 150.293
R38443 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 73.6304
R38444 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 60.4568
R38445 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 12.0358
R38446 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 11.4489
R38447 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.981478
R38448 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 0.788543
R38449 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.769522
R38450 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 0.720633
R38451 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 0.682565
R38452 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.580578
R38453 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 0.55213
R38454 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 0.470609
R38455 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.447191
R38456 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.428234
R38457 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.1255
R38458 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.1255
R38459 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 0.063
R38460 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 0.063
R38461 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.063
R38462 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 0.063
R38463 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 0.063
R38464 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 0.0435206
R38465 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 0.0107679
R38466 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.0107679
R38467 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 169.46
R38468 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 167.809
R38469 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 167.809
R38470 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 167.226
R38471 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 150.273
R38472 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 150.273
R38473 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 73.6406
R38474 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 73.6304
R38475 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 60.4568
R38476 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 12.3891
R38477 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 11.4489
R38478 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.68257
R38479 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 1.38365
R38480 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 1.19615
R38481 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 1.1717
R38482 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.08448
R38483 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.932141
R38484 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.720633
R38485 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 0.280391
R38486 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.217464
R38487 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R38488 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R38489 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.1255
R38490 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 0.0874565
R38491 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 0.063
R38492 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.063
R38493 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 0.063
R38494 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 0.063
R38495 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 0.0435206
R38496 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 0.0216397
R38497 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 0.0216397
R38498 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 0.0107679
R38499 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.0107679
R38500 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 179.256
R38501 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 168.089
R38502 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 150.293
R38503 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 73.6304
R38504 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 60.4568
R38505 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 12.0358
R38506 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.981478
R38507 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 0.788543
R38508 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.769522
R38509 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 0.720633
R38510 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 0.682565
R38511 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.580578
R38512 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 0.55213
R38513 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 0.470609
R38514 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.447191
R38515 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.428234
R38516 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1255
R38517 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1255
R38518 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 0.063
R38519 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 0.063
R38520 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.063
R38521 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 0.063
R38522 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 0.063
R38523 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 0.0435206
R38524 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 0.0107679
R38525 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.0107679
R38526 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 316.762
R38527 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 168.108
R38528 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 150.293
R38529 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 150.273
R38530 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 73.6406
R38531 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 73.6304
R38532 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 60.4568
R38533 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 12.0358
R38534 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 1.19615
R38535 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.981478
R38536 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 0.788543
R38537 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.769522
R38538 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 0.682565
R38539 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.580578
R38540 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 0.55213
R38541 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 0.484875
R38542 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 0.470609
R38543 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.447191
R38544 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.428234
R38545 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.217464
R38546 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R38547 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R38548 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.1255
R38549 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 0.063
R38550 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 0.063
R38551 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.063
R38552 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 0.063
R38553 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 0.063
R38554 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 0.0216397
R38555 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.0216397
R38556 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 0.0107679
R38557 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.0107679
R38558 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 169.46
R38559 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 167.809
R38560 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 167.809
R38561 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 167.227
R38562 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 150.293
R38563 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 150.273
R38564 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 73.6406
R38565 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 73.6304
R38566 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 60.3809
R38567 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 12.3891
R38568 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 11.4489
R38569 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 1.38365
R38570 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 1.19615
R38571 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 1.1717
R38572 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.848156
R38573 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 0.447191
R38574 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.38637
R38575 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 0.280391
R38576 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.217464
R38577 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.200143
R38578 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.152844
R38579 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.149957
R38580 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R38581 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.1255
R38582 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 0.0874565
R38583 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 0.063
R38584 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 0.063
R38585 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 0.063
R38586 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0454219
R38587 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 0.0107679
R38588 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0107679
R38589 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 169.46
R38590 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 167.809
R38591 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 167.809
R38592 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 167.226
R38593 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 150.273
R38594 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 150.273
R38595 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 73.6406
R38596 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 73.6304
R38597 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 60.4568
R38598 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 12.3891
R38599 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 11.4489
R38600 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.68257
R38601 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 1.38365
R38602 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 1.19615
R38603 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 1.1717
R38604 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.08448
R38605 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.932141
R38606 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 0.720633
R38607 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 0.280391
R38608 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.217464
R38609 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R38610 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R38611 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.1255
R38612 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 0.0874565
R38613 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 0.063
R38614 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.063
R38615 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 0.063
R38616 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 0.063
R38617 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 0.0435206
R38618 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 0.0216397
R38619 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.0216397
R38620 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 0.0107679
R38621 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.0107679
R38622 And_Gate_1.B.n10 And_Gate_1.B.t0 179.256
R38623 And_Gate_1.B.n10 And_Gate_1.B.t2 168.089
R38624 And_Gate_1.B.n2 And_Gate_1.B.t3 150.293
R38625 And_Gate_1.B.n4 And_Gate_1.B.t4 73.6304
R38626 Nand_Gate_4.Vout And_Gate_1.B.t1 60.3943
R38627 And_Gate_1.B.n8 And_Gate_1.B.n7 37.3347
R38628 And_Gate_1.B.n9 Nand_Gate_4.Vout 0.981478
R38629 And_Gate_1.B.n11 And_Gate_1.B.n9 0.788543
R38630 And_Gate_1.B.n3 And_Gate_1.Nand_Gate_0.B 0.769522
R38631 Nand_Gate_4.Vout And_Gate_1.B.n11 0.720633
R38632 And_Gate_1.B.n1 And_Gate_1.B.n0 0.682565
R38633 And_Gate_1.B.n1 Nand_Gate_4.Vout 0.580578
R38634 And_Gate_1.B.n3 And_Gate_1.B.n2 0.55213
R38635 And_Gate_1.B.n6 And_Gate_1.B.n5 0.470609
R38636 And_Gate_1.B.n2 And_Gate_1.Nand_Gate_0.B 0.447191
R38637 And_Gate_1.B.n6 And_Gate_1.Nand_Gate_0.B 0.428234
R38638 And_Gate_1.B.n5 And_Gate_1.Nand_Gate_0.B 0.1255
R38639 And_Gate_1.B.n0 Nand_Gate_4.Vout 0.1255
R38640 And_Gate_1.B.n7 And_Gate_1.B.n3 0.063
R38641 And_Gate_1.B.n7 And_Gate_1.B.n6 0.063
R38642 And_Gate_1.B.n0 Nand_Gate_4.Vout 0.063
R38643 And_Gate_1.B.n9 And_Gate_1.B.n8 0.063
R38644 And_Gate_1.B.n8 And_Gate_1.B.n1 0.063
R38645 And_Gate_1.B.n11 And_Gate_1.B.n10 0.0435206
R38646 And_Gate_1.B.n5 And_Gate_1.B.n4 0.0107679
R38647 And_Gate_1.B.n4 And_Gate_1.Nand_Gate_0.B 0.0107679
R38648 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 179.256
R38649 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 168.089
R38650 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 150.293
R38651 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 73.6304
R38652 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 60.3943
R38653 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 12.0358
R38654 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.981478
R38655 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 0.788543
R38656 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.769522
R38657 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.720633
R38658 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 0.682565
R38659 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.580578
R38660 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 0.55213
R38661 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 0.470609
R38662 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.447191
R38663 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.428234
R38664 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1255
R38665 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1255
R38666 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 0.063
R38667 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 0.063
R38668 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 0.063
R38669 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 0.063
R38670 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 0.063
R38671 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 0.0435206
R38672 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 0.0107679
R38673 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.0107679
R38674 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.t3 169.46
R38675 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout.t1 167.809
R38676 D_FlipFlop_2.3-input-nand_2.Vout.n9 D_FlipFlop_2.3-input-nand_2.Vout.t0 167.809
R38677 D_FlipFlop_2.3-input-nand_2.Vout.t7 D_FlipFlop_2.3-input-nand_2.Vout.n11 167.227
R38678 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.t7 150.293
R38679 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.t6 150.273
R38680 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout.t4 73.6406
R38681 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout.t5 73.6304
R38682 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout.t2 60.3809
R38683 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout.n5 12.3891
R38684 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout.n9 11.4489
R38685 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout.n2 1.38365
R38686 D_FlipFlop_2.3-input-nand_2.Vout.n12 D_FlipFlop_2.3-input-nand_2.Vout.n1 1.19615
R38687 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout.n4 1.1717
R38688 D_FlipFlop_2.3-input-nand_2.Vout.n2 D_FlipFlop_2.3-input-nand_2.Vout 0.848156
R38689 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.Vout.n12 0.447191
R38690 D_FlipFlop_2.3-input-nand_2.Vout.n3 D_FlipFlop_2.3-input-nand_2.Vout 0.38637
R38691 D_FlipFlop_2.3-input-nand_2.Vout.n11 D_FlipFlop_2.3-input-nand_2.Vout.n10 0.280391
R38692 D_FlipFlop_2.3-input-nand_2.Vout.n10 D_FlipFlop_2.3-input-nand_2.Vout.n8 0.262643
R38693 D_FlipFlop_2.3-input-nand_2.Vout.n4 D_FlipFlop_2.3-input-nand_2.Vout 0.217464
R38694 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout 0.152844
R38695 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout 0.149957
R38696 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R38697 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout 0.1255
R38698 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout.n7 0.0874565
R38699 D_FlipFlop_2.3-input-nand_2.Vout.n6 D_FlipFlop_2.3-input-nand_2.Vout.n3 0.063
R38700 D_FlipFlop_2.3-input-nand_2.Vout.n7 D_FlipFlop_2.3-input-nand_2.Vout.n6 0.063
R38701 D_FlipFlop_2.3-input-nand_2.Vout.n8 D_FlipFlop_2.3-input-nand_2.Vout 0.063
R38702 D_FlipFlop_2.3-input-nand_2.Vout.n5 D_FlipFlop_2.3-input-nand_2.Vout 0.0454219
R38703 D_FlipFlop_2.3-input-nand_2.Vout.n1 D_FlipFlop_2.3-input-nand_2.Vout.n0 0.0107679
R38704 D_FlipFlop_2.3-input-nand_2.Vout.n0 D_FlipFlop_2.3-input-nand_2.Vout 0.0107679
R38705 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 179.256
R38706 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 168.089
R38707 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 150.293
R38708 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 73.6304
R38709 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 60.3943
R38710 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 12.0358
R38711 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.981478
R38712 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 0.788543
R38713 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.769522
R38714 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 0.720633
R38715 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 0.682565
R38716 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.580578
R38717 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 0.55213
R38718 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 0.470609
R38719 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.447191
R38720 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.428234
R38721 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1255
R38722 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1255
R38723 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 0.063
R38724 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 0.063
R38725 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.063
R38726 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 0.063
R38727 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 0.063
R38728 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 0.0435206
R38729 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 0.0107679
R38730 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.0107679
R38731 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout.t3 169.46
R38732 D_FlipFlop_6.3-input-nand_2.Vout.n4 D_FlipFlop_6.3-input-nand_2.Vout.t2 167.809
R38733 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout.t1 167.809
R38734 D_FlipFlop_6.3-input-nand_2.Vout.n3 D_FlipFlop_6.3-input-nand_2.Vout.t7 167.227
R38735 D_FlipFlop_6.3-input-nand_2.Vout.t7 D_FlipFlop_6.3-input-nand_2.Vout.n2 150.293
R38736 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.t6 150.273
R38737 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout.t4 73.6406
R38738 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout.t5 73.6304
R38739 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.t0 60.3809
R38740 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout.n9 12.3891
R38741 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.n4 11.4489
R38742 D_FlipFlop_6.3-input-nand_2.Vout.n12 D_FlipFlop_6.3-input-nand_2.Vout.n11 1.38365
R38743 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout.n1 1.19615
R38744 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout.n8 1.1717
R38745 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.Vout.n12 0.848156
R38746 D_FlipFlop_6.3-input-nand_2.Vout.n2 D_FlipFlop_6.3-input-nand_2.Vout 0.447191
R38747 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout 0.38637
R38748 D_FlipFlop_6.3-input-nand_2.Vout.n5 D_FlipFlop_6.3-input-nand_2.Vout.n3 0.280391
R38749 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout.n5 0.262643
R38750 D_FlipFlop_6.3-input-nand_2.Vout.n8 D_FlipFlop_6.3-input-nand_2.Vout 0.217464
R38751 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout 0.152844
R38752 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout 0.149957
R38753 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R38754 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout 0.1255
R38755 D_FlipFlop_6.3-input-nand_2.Vout.n7 D_FlipFlop_6.3-input-nand_2.Vout.n6 0.0874565
R38756 D_FlipFlop_6.3-input-nand_2.Vout.n6 D_FlipFlop_6.3-input-nand_2.Vout 0.063
R38757 D_FlipFlop_6.3-input-nand_2.Vout.n11 D_FlipFlop_6.3-input-nand_2.Vout.n10 0.063
R38758 D_FlipFlop_6.3-input-nand_2.Vout.n10 D_FlipFlop_6.3-input-nand_2.Vout.n7 0.063
R38759 D_FlipFlop_6.3-input-nand_2.Vout.n9 D_FlipFlop_6.3-input-nand_2.Vout 0.0454219
R38760 D_FlipFlop_6.3-input-nand_2.Vout.n1 D_FlipFlop_6.3-input-nand_2.Vout.n0 0.0107679
R38761 D_FlipFlop_6.3-input-nand_2.Vout.n0 D_FlipFlop_6.3-input-nand_2.Vout 0.0107679
R38762 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 316.762
R38763 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 168.108
R38764 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 150.293
R38765 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 150.273
R38766 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 73.6406
R38767 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 73.6304
R38768 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 60.4568
R38769 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 12.0358
R38770 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 1.19615
R38771 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.981478
R38772 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 0.788543
R38773 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.769522
R38774 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 0.682565
R38775 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.580578
R38776 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 0.55213
R38777 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 0.484875
R38778 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 0.470609
R38779 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.447191
R38780 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.428234
R38781 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.217464
R38782 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R38783 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R38784 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.1255
R38785 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 0.063
R38786 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 0.063
R38787 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.063
R38788 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 0.063
R38789 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 0.063
R38790 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 0.0216397
R38791 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.0216397
R38792 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 0.0107679
R38793 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.0107679
R38794 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 169.46
R38795 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 167.809
R38796 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 167.809
R38797 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 167.227
R38798 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 150.293
R38799 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 150.273
R38800 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 73.6406
R38801 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 73.6304
R38802 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 60.3809
R38803 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 12.3891
R38804 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 11.4489
R38805 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 1.38365
R38806 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 1.19615
R38807 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 1.1717
R38808 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.848156
R38809 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 0.447191
R38810 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.38637
R38811 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 0.280391
R38812 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 0.262643
R38813 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.217464
R38814 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.152844
R38815 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.149957
R38816 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.1255
R38817 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.1255
R38818 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 0.0874565
R38819 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 0.063
R38820 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 0.063
R38821 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.063
R38822 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.0454219
R38823 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 0.0107679
R38824 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.0107679
R38825 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 169.46
R38826 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 167.809
R38827 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 167.809
R38828 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 167.227
R38829 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 150.293
R38830 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 150.273
R38831 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 73.6406
R38832 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 73.6304
R38833 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 60.3809
R38834 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 12.3891
R38835 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 11.4489
R38836 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 1.38365
R38837 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 1.19615
R38838 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 1.1717
R38839 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.848156
R38840 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 0.447191
R38841 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.38637
R38842 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 0.280391
R38843 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 0.262643
R38844 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.217464
R38845 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.152844
R38846 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.149957
R38847 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.1255
R38848 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.1255
R38849 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 0.0874565
R38850 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 0.063
R38851 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 0.063
R38852 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.063
R38853 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.0454219
R38854 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 0.0107679
R38855 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.0107679
R38856 Nand_Gate_6.Vout.n0 Nand_Gate_6.Vout.t2 179.256
R38857 Nand_Gate_6.Vout.n0 Nand_Gate_6.Vout.t1 168.089
R38858 Nand_Gate_6.Vout.n3 Nand_Gate_6.Vout.t3 150.293
R38859 Nand_Gate_6.Vout.n5 Nand_Gate_6.Vout.t4 73.6304
R38860 Nand_Gate_6.Vout Nand_Gate_6.Vout.t0 60.3943
R38861 Nand_Gate_6.Vout.n9 Nand_Gate_6.Vout.n8 37.3347
R38862 Nand_Gate_6.Vout.n2 Nand_Gate_6.Vout 0.981478
R38863 Nand_Gate_6.Vout.n2 Nand_Gate_6.Vout.n1 0.788543
R38864 Nand_Gate_6.Vout.n4 Nand_Gate_6.Vout 0.769522
R38865 Nand_Gate_6.Vout.n1 Nand_Gate_6.Vout 0.720633
R38866 Nand_Gate_6.Vout.n11 Nand_Gate_6.Vout.n10 0.682565
R38867 Nand_Gate_6.Vout.n10 Nand_Gate_6.Vout 0.580578
R38868 Nand_Gate_6.Vout.n4 Nand_Gate_6.Vout.n3 0.55213
R38869 Nand_Gate_6.Vout.n7 Nand_Gate_6.Vout.n6 0.470609
R38870 Nand_Gate_6.Vout.n3 Nand_Gate_6.Vout 0.447191
R38871 Nand_Gate_6.Vout.n7 Nand_Gate_6.Vout 0.428234
R38872 Nand_Gate_6.Vout.n6 Nand_Gate_6.Vout 0.1255
R38873 Nand_Gate_6.Vout.n11 Nand_Gate_6.Vout 0.1255
R38874 Nand_Gate_6.Vout.n8 Nand_Gate_6.Vout.n4 0.063
R38875 Nand_Gate_6.Vout.n8 Nand_Gate_6.Vout.n7 0.063
R38876 Nand_Gate_6.Vout.n9 Nand_Gate_6.Vout.n2 0.063
R38877 Nand_Gate_6.Vout.n10 Nand_Gate_6.Vout.n9 0.063
R38878 Nand_Gate_6.Vout Nand_Gate_6.Vout.n11 0.063
R38879 Nand_Gate_6.Vout.n1 Nand_Gate_6.Vout.n0 0.0435206
R38880 Nand_Gate_6.Vout.n6 Nand_Gate_6.Vout.n5 0.0107679
R38881 Nand_Gate_6.Vout.n5 Nand_Gate_6.Vout 0.0107679
R38882 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 169.46
R38883 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 167.809
R38884 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 167.809
R38885 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 167.227
R38886 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 150.293
R38887 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 150.273
R38888 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 73.6406
R38889 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 73.6304
R38890 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 60.3809
R38891 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 12.3891
R38892 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 11.4489
R38893 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 1.38365
R38894 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 1.19615
R38895 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 1.1717
R38896 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.848156
R38897 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 0.447191
R38898 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.38637
R38899 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 0.280391
R38900 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 0.262643
R38901 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.217464
R38902 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.152844
R38903 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.149957
R38904 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.1255
R38905 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.1255
R38906 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 0.0874565
R38907 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 0.063
R38908 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 0.063
R38909 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.063
R38910 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.0454219
R38911 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 0.0107679
R38912 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.0107679
R38913 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 169.46
R38914 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 167.809
R38915 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 167.809
R38916 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 167.227
R38917 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 150.293
R38918 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 150.273
R38919 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 73.6406
R38920 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 73.6304
R38921 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 60.3809
R38922 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 12.3891
R38923 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 11.4489
R38924 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 1.38365
R38925 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 1.19615
R38926 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 1.1717
R38927 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.848156
R38928 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 0.447191
R38929 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.38637
R38930 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 0.280391
R38931 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.217464
R38932 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.200143
R38933 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.152844
R38934 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.149957
R38935 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R38936 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.1255
R38937 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 0.0874565
R38938 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 0.063
R38939 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 0.063
R38940 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 0.063
R38941 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0454219
R38942 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 0.0107679
R38943 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0107679
R38944 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 316.762
R38945 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 168.108
R38946 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 150.293
R38947 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 150.273
R38948 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 73.6406
R38949 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 73.6304
R38950 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 60.3943
R38951 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 12.0358
R38952 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 1.19615
R38953 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.981478
R38954 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 0.788543
R38955 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.769522
R38956 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 0.682565
R38957 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.580578
R38958 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 0.55213
R38959 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 0.484875
R38960 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 0.470609
R38961 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.447191
R38962 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.428234
R38963 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.217464
R38964 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R38965 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R38966 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.1255
R38967 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 0.063
R38968 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 0.063
R38969 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.063
R38970 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 0.063
R38971 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 0.063
R38972 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 0.0216397
R38973 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.0216397
R38974 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 0.0107679
R38975 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.0107679
R38976 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 316.762
R38977 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 168.108
R38978 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 150.293
R38979 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 150.273
R38980 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 73.6406
R38981 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 73.6304
R38982 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 60.4568
R38983 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 12.0358
R38984 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 1.19615
R38985 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.981478
R38986 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 0.788543
R38987 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.769522
R38988 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 0.682565
R38989 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.580578
R38990 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 0.55213
R38991 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 0.484875
R38992 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 0.470609
R38993 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.447191
R38994 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.428234
R38995 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.217464
R38996 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R38997 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R38998 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.1255
R38999 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 0.063
R39000 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 0.063
R39001 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.063
R39002 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 0.063
R39003 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 0.063
R39004 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 0.0216397
R39005 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.0216397
R39006 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 0.0107679
R39007 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.0107679
R39008 Q0.n7 Q0.t1 169.46
R39009 Q0.n9 Q0.t2 167.809
R39010 Q0.n7 Q0.t0 167.809
R39011 Q0 Q0.t9 158.585
R39012 Q0.n13 Q0.t7 150.869
R39013 Q0.n12 Q0.t8 150.869
R39014 Q0.t9 Q0.n2 150.293
R39015 Q0.n14 Q0.n11 137.644
R39016 Q0 Q0.t4 78.1811
R39017 Q0.n12 Q0.t5 74.1352
R39018 Q0.t4 Q0.n13 74.1352
R39019 Q0.n0 Q0.t6 73.6304
R39020 Q0.n5 Q0.t3 60.3809
R39021 Q0.n11 Q0 41.1198
R39022 Q0.n8 Q0.n7 11.4489
R39023 Q0.n10 Q0.n9 4.78039
R39024 Q0.n10 Q0.n4 1.74412
R39025 Q0.n13 Q0.n12 1.66898
R39026 Q0.n6 Q0.n5 1.64452
R39027 Q0.n2 Q0.n1 1.19615
R39028 Q0.n5 Q0 0.848156
R39029 Q0.n2 Q0 0.447191
R39030 Q0.n4 Q0.n3 0.3624
R39031 Q0.n4 Q0 0.333061
R39032 Q0.n9 Q0.n8 0.280391
R39033 Q0.n8 Q0.n6 0.262643
R39034 Q0.n6 Q0 0.1255
R39035 Q0.n1 Q0 0.1255
R39036 Q0.n12 Q0 0.063
R39037 Q0.n6 Q0 0.063
R39038 Q0.n11 Q0.n10 0.0305325
R39039 Q0 Q0.n14 0.0168043
R39040 Q0.n14 Q0 0.0122188
R39041 Q0.n1 Q0.n0 0.0107679
R39042 Q0.n0 Q0 0.0107679
R39043 Q0.n3 Q0 0.00441667
R39044 Q0.n3 Q0 0.00406061
R39045 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 179.256
R39046 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 168.089
R39047 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 150.293
R39048 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 73.6304
R39049 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 60.4568
R39050 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 12.0358
R39051 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.981478
R39052 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 0.788543
R39053 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.769522
R39054 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 0.720633
R39055 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 0.682565
R39056 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.580578
R39057 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 0.55213
R39058 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 0.470609
R39059 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.447191
R39060 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.428234
R39061 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1255
R39062 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1255
R39063 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 0.063
R39064 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 0.063
R39065 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.063
R39066 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 0.063
R39067 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 0.063
R39068 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 0.0435206
R39069 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 0.0107679
R39070 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.0107679
R39071 Nand_Gate_0.B.n31 Nand_Gate_0.B.t0 169.46
R39072 Nand_Gate_0.B.n31 Nand_Gate_0.B.t1 167.809
R39073 Nand_Gate_0.B.n33 Nand_Gate_0.B.t2 167.809
R39074 Nand_Gate_0.B Nand_Gate_0.B.t5 158.585
R39075 Nand_Gate_0.B.t5 Nand_Gate_0.B.n2 150.293
R39076 Nand_Gate_0.B.n24 Nand_Gate_0.B.t4 150.273
R39077 Nand_Gate_0.B.n14 Nand_Gate_0.B.t7 150.273
R39078 Nand_Gate_0.B.n8 Nand_Gate_0.B.t10 150.273
R39079 Nand_Gate_0.B.n12 Nand_Gate_0.B.t6 73.6406
R39080 Nand_Gate_0.B.n6 Nand_Gate_0.B.t9 73.6406
R39081 Nand_Gate_0.B.n21 Nand_Gate_0.B.t8 73.6304
R39082 Nand_Gate_0.B.n0 Nand_Gate_0.B.t11 73.6304
R39083 Nand_Gate_0.B.n4 Nand_Gate_0.B.t3 60.3809
R39084 Nand_Gate_0.B.n25 Nand_Gate_0.B.n24 40.8363
R39085 Nand_Gate_0.B.n32 Nand_Gate_0.B.n31 11.4489
R39086 Nand_Gate_0.B.n34 Nand_Gate_0.B.n33 8.21389
R39087 Nand_Gate_0.B.n18 Nand_Gate_0.B.n11 8.1418
R39088 Nand_Gate_0.B.n20 Nand_Gate_0.B.n19 6.47604
R39089 Nand_Gate_0.B.n19 Nand_Gate_0.B 5.35402
R39090 Nand_Gate_0.B.n28 Nand_Gate_0.B 4.55128
R39091 Nand_Gate_0.B.n18 Nand_Gate_0.B.n17 4.5005
R39092 Nand_Gate_0.B.n2 Nand_Gate_0.B.n1 1.19615
R39093 Nand_Gate_0.B.n23 Nand_Gate_0.B.n22 1.1717
R39094 Nand_Gate_0.B.n5 Nand_Gate_0.B 1.08746
R39095 Nand_Gate_0.B.n20 Nand_Gate_0.B 0.973326
R39096 Nand_Gate_0.B.n23 Nand_Gate_0.B 0.932141
R39097 Nand_Gate_0.B.n13 Nand_Gate_0.B 0.851043
R39098 Nand_Gate_0.B.n7 Nand_Gate_0.B 0.851043
R39099 Nand_Gate_0.B.n4 Nand_Gate_0.B 0.848156
R39100 Nand_Gate_0.B.n30 Nand_Gate_0.B.n29 0.788543
R39101 Nand_Gate_0.B.n27 Nand_Gate_0.B.n26 0.755935
R39102 Nand_Gate_0.B.n5 Nand_Gate_0.B.n4 0.682565
R39103 Nand_Gate_0.B.n29 Nand_Gate_0.B 0.65675
R39104 Nand_Gate_0.B.n16 Nand_Gate_0.B.n15 0.55213
R39105 Nand_Gate_0.B.n10 Nand_Gate_0.B.n9 0.55213
R39106 Nand_Gate_0.B.n16 Nand_Gate_0.B 0.486828
R39107 Nand_Gate_0.B.n10 Nand_Gate_0.B 0.486828
R39108 Nand_Gate_0.B.n26 Nand_Gate_0.B 0.48023
R39109 Nand_Gate_0.B.n13 Nand_Gate_0.B.n12 0.470609
R39110 Nand_Gate_0.B.n7 Nand_Gate_0.B.n6 0.470609
R39111 Nand_Gate_0.B.n2 Nand_Gate_0.B 0.447191
R39112 Nand_Gate_0.B.n34 Nand_Gate_0.B.n3 0.425067
R39113 Nand_Gate_0.B Nand_Gate_0.B.n34 0.39003
R39114 Nand_Gate_0.B.n33 Nand_Gate_0.B.n32 0.280391
R39115 Nand_Gate_0.B.n12 Nand_Gate_0.B 0.217464
R39116 Nand_Gate_0.B.n6 Nand_Gate_0.B 0.217464
R39117 Nand_Gate_0.B.n32 Nand_Gate_0.B 0.200143
R39118 Nand_Gate_0.B.n22 Nand_Gate_0.B 0.1255
R39119 Nand_Gate_0.B.n15 Nand_Gate_0.B 0.1255
R39120 Nand_Gate_0.B.n9 Nand_Gate_0.B 0.1255
R39121 Nand_Gate_0.B.n30 Nand_Gate_0.B 0.1255
R39122 Nand_Gate_0.B.n1 Nand_Gate_0.B 0.1255
R39123 Nand_Gate_0.B.n24 Nand_Gate_0.B.n23 0.063
R39124 Nand_Gate_0.B.n17 Nand_Gate_0.B.n13 0.063
R39125 Nand_Gate_0.B.n17 Nand_Gate_0.B.n16 0.063
R39126 Nand_Gate_0.B.n11 Nand_Gate_0.B.n7 0.063
R39127 Nand_Gate_0.B.n11 Nand_Gate_0.B.n10 0.063
R39128 Nand_Gate_0.B.n19 Nand_Gate_0.B.n18 0.063
R39129 Nand_Gate_0.B.n25 Nand_Gate_0.B.n20 0.063
R39130 Nand_Gate_0.B.n26 Nand_Gate_0.B.n25 0.063
R39131 Nand_Gate_0.B.n28 Nand_Gate_0.B.n5 0.063
R39132 Nand_Gate_0.B.n29 Nand_Gate_0.B.n28 0.063
R39133 Nand_Gate_0.B Nand_Gate_0.B.n30 0.063
R39134 Nand_Gate_0.B.n15 Nand_Gate_0.B.n14 0.0216397
R39135 Nand_Gate_0.B.n14 Nand_Gate_0.B 0.0216397
R39136 Nand_Gate_0.B.n9 Nand_Gate_0.B.n8 0.0216397
R39137 Nand_Gate_0.B.n8 Nand_Gate_0.B 0.0216397
R39138 Nand_Gate_0.B.n27 Nand_Gate_0.B 0.0168043
R39139 Nand_Gate_0.B Nand_Gate_0.B.n27 0.0122188
R39140 Nand_Gate_0.B.n22 Nand_Gate_0.B.n21 0.0107679
R39141 Nand_Gate_0.B.n21 Nand_Gate_0.B 0.0107679
R39142 Nand_Gate_0.B.n1 Nand_Gate_0.B.n0 0.0107679
R39143 Nand_Gate_0.B.n0 Nand_Gate_0.B 0.0107679
R39144 Nand_Gate_0.B.n3 Nand_Gate_0.B 0.00441667
R39145 Nand_Gate_0.B.n3 Nand_Gate_0.B 0.00406061
R39146 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 169.46
R39147 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 168.089
R39148 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 167.809
R39149 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 150.293
R39150 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 73.6304
R39151 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 60.3943
R39152 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 12.0358
R39153 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 11.4489
R39154 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.981478
R39155 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 0.788543
R39156 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.769522
R39157 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 0.720633
R39158 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 0.682565
R39159 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.580578
R39160 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 0.55213
R39161 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 0.470609
R39162 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.447191
R39163 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.428234
R39164 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.1255
R39165 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.1255
R39166 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 0.063
R39167 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 0.063
R39168 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.063
R39169 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 0.063
R39170 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 0.063
R39171 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 0.0435206
R39172 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 0.0107679
R39173 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.0107679
R39174 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 169.46
R39175 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 168.089
R39176 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 167.809
R39177 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 150.293
R39178 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 73.6304
R39179 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 60.4568
R39180 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 12.0358
R39181 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 11.4489
R39182 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.981478
R39183 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 0.788543
R39184 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.769522
R39185 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 0.720633
R39186 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 0.682565
R39187 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.580578
R39188 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 0.55213
R39189 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 0.470609
R39190 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.447191
R39191 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.428234
R39192 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.1255
R39193 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.1255
R39194 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 0.063
R39195 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 0.063
R39196 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.063
R39197 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 0.063
R39198 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 0.063
R39199 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 0.0435206
R39200 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 0.0107679
R39201 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.0107679
R39202 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 169.46
R39203 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 168.089
R39204 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 167.809
R39205 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 150.273
R39206 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 73.6406
R39207 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 60.3809
R39208 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 12.0358
R39209 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 11.4489
R39210 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 1.08746
R39211 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.851043
R39212 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.848156
R39213 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 0.788543
R39214 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 0.682565
R39215 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.65675
R39216 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 0.55213
R39217 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.486828
R39218 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 0.470609
R39219 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 0.262643
R39220 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.217464
R39221 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.1255
R39222 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.1255
R39223 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 0.063
R39224 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 0.063
R39225 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 0.063
R39226 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 0.063
R39227 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 0.063
R39228 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 0.0216397
R39229 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.0216397
R39230 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 169.46
R39231 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 168.089
R39232 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 167.809
R39233 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 150.293
R39234 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 73.6304
R39235 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 60.4568
R39236 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 12.0358
R39237 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 11.4489
R39238 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.981478
R39239 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 0.788543
R39240 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.769522
R39241 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 0.720633
R39242 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 0.682565
R39243 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.580578
R39244 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 0.55213
R39245 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 0.470609
R39246 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.447191
R39247 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.428234
R39248 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.1255
R39249 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.1255
R39250 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 0.063
R39251 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 0.063
R39252 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.063
R39253 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 0.063
R39254 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 0.063
R39255 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 0.0435206
R39256 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 0.0107679
R39257 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.0107679
R39258 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 169.46
R39259 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 168.089
R39260 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 167.809
R39261 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 150.273
R39262 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 73.6406
R39263 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 60.3809
R39264 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 12.0358
R39265 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 11.4489
R39266 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 1.08746
R39267 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.851043
R39268 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.848156
R39269 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 0.788543
R39270 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 0.682565
R39271 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.65675
R39272 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 0.55213
R39273 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.486828
R39274 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 0.470609
R39275 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 0.262643
R39276 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.217464
R39277 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.1255
R39278 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.1255
R39279 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 0.063
R39280 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 0.063
R39281 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 0.063
R39282 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 0.063
R39283 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 0.063
R39284 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 0.0216397
R39285 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0216397
R39286 And_Gate_0.B.n10 And_Gate_0.B.t0 179.256
R39287 And_Gate_0.B.n10 And_Gate_0.B.t2 168.089
R39288 And_Gate_0.B.n2 And_Gate_0.B.t3 150.293
R39289 And_Gate_0.B.n4 And_Gate_0.B.t4 73.6304
R39290 Nand_Gate_7.Vout And_Gate_0.B.t1 60.3943
R39291 And_Gate_0.B.n8 And_Gate_0.B.n7 37.3347
R39292 And_Gate_0.B.n9 Nand_Gate_7.Vout 0.981478
R39293 And_Gate_0.B.n11 And_Gate_0.B.n9 0.788543
R39294 And_Gate_0.B.n3 And_Gate_0.Nand_Gate_0.B 0.769522
R39295 Nand_Gate_7.Vout And_Gate_0.B.n11 0.720633
R39296 And_Gate_0.B.n1 And_Gate_0.B.n0 0.682565
R39297 And_Gate_0.B.n1 Nand_Gate_7.Vout 0.580578
R39298 And_Gate_0.B.n3 And_Gate_0.B.n2 0.55213
R39299 And_Gate_0.B.n6 And_Gate_0.B.n5 0.470609
R39300 And_Gate_0.B.n2 And_Gate_0.Nand_Gate_0.B 0.447191
R39301 And_Gate_0.B.n6 And_Gate_0.Nand_Gate_0.B 0.428234
R39302 And_Gate_0.B.n5 And_Gate_0.Nand_Gate_0.B 0.1255
R39303 And_Gate_0.B.n0 Nand_Gate_7.Vout 0.1255
R39304 And_Gate_0.B.n7 And_Gate_0.B.n3 0.063
R39305 And_Gate_0.B.n7 And_Gate_0.B.n6 0.063
R39306 And_Gate_0.B.n0 Nand_Gate_7.Vout 0.063
R39307 And_Gate_0.B.n9 And_Gate_0.B.n8 0.063
R39308 And_Gate_0.B.n8 And_Gate_0.B.n1 0.063
R39309 And_Gate_0.B.n11 And_Gate_0.B.n10 0.0435206
R39310 And_Gate_0.B.n5 And_Gate_0.B.n4 0.0107679
R39311 And_Gate_0.B.n4 And_Gate_0.Nand_Gate_0.B 0.0107679
R39312 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 169.46
R39313 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 167.809
R39314 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 167.809
R39315 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 167.226
R39316 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 150.273
R39317 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 150.273
R39318 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 73.6406
R39319 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 73.6304
R39320 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 60.3943
R39321 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 12.3891
R39322 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 11.4489
R39323 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 1.68257
R39324 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 1.38365
R39325 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 1.19615
R39326 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 1.1717
R39327 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 1.08448
R39328 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.932141
R39329 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.720633
R39330 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 0.280391
R39331 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.217464
R39332 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R39333 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R39334 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.1255
R39335 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 0.0874565
R39336 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 0.063
R39337 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 0.063
R39338 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 0.063
R39339 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 0.063
R39340 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 0.0435206
R39341 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 0.0216397
R39342 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.0216397
R39343 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 0.0107679
R39344 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.0107679
R39345 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 179.256
R39346 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 168.089
R39347 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 150.293
R39348 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 73.6304
R39349 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 60.3943
R39350 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 12.0358
R39351 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.981478
R39352 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 0.788543
R39353 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.769522
R39354 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 0.720633
R39355 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 0.682565
R39356 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.580578
R39357 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 0.55213
R39358 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 0.470609
R39359 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.447191
R39360 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.428234
R39361 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1255
R39362 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1255
R39363 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 0.063
R39364 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 0.063
R39365 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.063
R39366 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 0.063
R39367 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 0.063
R39368 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 0.0435206
R39369 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 0.0107679
R39370 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.0107679
R39371 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 169.46
R39372 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 167.809
R39373 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 167.809
R39374 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 167.226
R39375 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 150.273
R39376 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 150.273
R39377 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 73.6406
R39378 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 73.6304
R39379 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 60.3943
R39380 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 12.3891
R39381 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 11.4489
R39382 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 1.68257
R39383 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 1.38365
R39384 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 1.19615
R39385 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 1.1717
R39386 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 1.08448
R39387 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.932141
R39388 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 0.720633
R39389 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 0.280391
R39390 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.217464
R39391 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R39392 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R39393 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.1255
R39394 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 0.0874565
R39395 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 0.063
R39396 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.063
R39397 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 0.063
R39398 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 0.063
R39399 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 0.0435206
R39400 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 0.0216397
R39401 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.0216397
R39402 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 0.0107679
R39403 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.0107679
C0 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.16429f
C1 RingCounter_0.D_FlipFlop_15.Q' RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.11654f
C2 CDAC8_0.switch_1.Z EN 0.15062f
C3 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.30154f
C4 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.06445f
C5 FFCLR a_134283_33443# 0.01803f
C6 a_62409_15797# VDD 0.01571f
C7 RingCounter_0.D_FlipFlop_16.Q' a_28675_13083# 0.06113f
C8 a_128237_23350# VDD 0.02521f
C9 a_128237_23350# a_128851_23350# 0.05935f
C10 a_79625_52572# a_80239_52572# 0.05935f
C11 D_FlipFlop_2.Q' a_128237_37007# 0.06113f
C12 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.0846f
C13 a_90535_15797# VDD 0.06072f
C14 D_FlipFlop_5.Inverter_0.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.0857f
C15 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout a_106699_49858# 0.04995f
C16 a_85233_49858# EN 0.01149f
C17 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout CLK 0.27362f
C18 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout VDD 1.56255f
C19 a_87949_13083# CLK 0.03129f
C20 a_62539_49858# a_63153_49858# 0.05935f
C21 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_2.C 0.1486f
C22 a_134283_30478# VDD 0.02521f
C23 a_72835_15797# VDD 0.02906f
C24 Nand_Gate_0.A a_132925_39721# 0.04682f
C25 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.Inverter_1.Vout 0.25963f
C26 D_FlipFlop_2.Inverter_0.Vout a_134283_37007# 0.04443f
C27 a_128237_26914# a_128851_26914# 0.05935f
C28 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 0.25579f
C29 a_123041_13083# a_123655_13083# 0.05935f
C30 a_107313_49858# VDD 0.0325f
C31 a_128237_33443# VDD 0.02521f
C32 D_FlipFlop_6.3-input-nand_1.Vout D_FlipFlop_7.3-input-nand_0.Vout 0.01418f
C33 Nand_Gate_5.Vout a_115177_47663# 0.05964f
C34 FFCLR D_FlipFlop_1.Q' 0.0683f
C35 a_106699_52572# VDD 0.0564f
C36 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout VDD 2.88547f
C37 FFCLR D_FlipFlop_0.Inverter_1.Vout 0.56808f
C38 D_FlipFlop_6.Nand_Gate_1.Vout a_128237_20636# 0.04444f
C39 Nand_Gate_2.A Nand_Gate_2.Vout 0.11161f
C40 a_128851_26914# VDD 0.01186f
C41 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout VDD 2.73332f
C42 a_134283_40571# a_134897_40571# 0.05935f
C43 Nand_Gate_5.A D_FlipFlop_0.Nand_Gate_0.Vout 0.64617f
C44 D_FlipFlop_0.Inverter_1.Vout a_130209_44135# 0.04995f
C45 RingCounter_0.D_FlipFlop_13.Q' a_73449_13083# 0.01335f
C46 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout a_96273_49858# 0.04443f
C47 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_90665_49858# 0.04995f
C48 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.04109f
C49 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.06445f
C50 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.3-input-nand_2.C 0.25579f
C51 Nand_Gate_4.A RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.08377f
C52 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 1.09975f
C53 Nand_Gate_5.Vout EN 0.10962f
C54 RingCounter_0.D_FlipFlop_3.Q' Nand_Gate_0.B 1.10693f
C55 D_FlipFlop_6.Q' Nand_Gate_7.B 0.03706f
C56 a_56801_13083# VDD 0.02865f
C57 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.48392f
C58 CDAC8_0.switch_6.Z Q2 0.74768f
C59 Nand_Gate_7.A a_59977_16975# 0.0476f
C60 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.30154f
C61 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.3-input-nand_2.C 0.25579f
C62 And_Gate_3.Inverter_0.Vin Q0 0.05258f
C63 D_FlipFlop_5.Nand_Gate_1.Vout a_128237_24200# 0.04444f
C64 a_132925_37007# VDD 0.01186f
C65 RingCounter_0.D_FlipFlop_16.Q a_41073_52572# 0.04443f
C66 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout CLK 0.23464f
C67 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout a_98245_49858# 0.04443f
C68 a_108671_52572# a_109285_52572# 0.05935f
C69 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout VDD 2.8604f
C70 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.30154f
C71 a_41073_49858# EN 0.01767f
C72 a_77523_15797# EN 0.045f
C73 a_130209_23350# VDD 0.02521f
C74 a_101575_13083# EN 0.0452f
C75 D_FlipFlop_5.Q' Nand_Gate_6.B 0.03561f
C76 RingCounter_0.D_FlipFlop_8.Q' a_39715_15797# 0.04443f
C77 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_86591_49858# 0.01335f
C78 a_43789_13083# CLK 0.03129f
C79 a_40459_49858# a_41073_49858# 0.05935f
C80 D_FlipFlop_1.Inverter_0.Vout VDD 1.37367f
C81 a_78267_52572# RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.05964f
C82 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout a_111387_49858# 0.04995f
C83 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout EN 0.09127f
C84 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 1.09946f
C85 And_Gate_3.Inverter_0.Vin EN 0.02316f
C86 a_95659_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.01335f
C87 a_63153_49858# VDD 0.0325f
C88 a_100961_13083# a_101575_13083# 0.05935f
C89 D_FlipFlop_3.Nand_Gate_1.Vout Q5 0.06503f
C90 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout VDD 2.07373f
C91 a_123655_13083# VDD 0.01327f
C92 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout VDD 2.08141f
C93 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout EN 0.24889f
C94 a_116995_15797# RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.04444f
C95 a_121683_15797# VDD 0.03339f
C96 RingCounter_0.D_FlipFlop_3.Q' RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.11654f
C97 Nand_Gate_6.B Q0 0.06521f
C98 FFCLR a_134897_23350# 0.08419f
C99 a_134897_40571# VDD 0.01186f
C100 D_FlipFlop_7.Nand_Gate_1.Vout a_130209_17072# 0.05964f
C101 a_63767_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.04443f
C102 CDAC8_0.switch_7.Z Q4 1.28022f
C103 D_FlipFlop_3.3-input-nand_2.Vout a_132311_43285# 0.05964f
C104 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout EN 0.61894f
C105 a_53471_52572# EN 0.045f
C106 a_128851_46849# Q4 0.01335f
C107 a_128237_23350# D_FlipFlop_6.Nand_Gate_0.Vout 0.04444f
C108 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_80239_52572# 0.04444f
C109 D_FlipFlop_1.3-input-nand_2.C a_132925_33443# 0.01335f
C110 a_75898_42964# CDAC8_0.switch_9.Z 0.29215f
C111 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.0857f
C112 a_128851_33443# EN 0.05028f
C113 a_109285_52572# VDD 0.02521f
C114 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_76165_49858# 0.05964f
C115 a_110643_13083# CLK 0.03129f
C116 CDAC8_0.switch_9.Z Q3 0.36261f
C117 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_95529_15797# 0.04995f
C118 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 1.09975f
C119 Nand_Gate_2.A a_132925_43285# 0.04684f
C120 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_46375_13083# 0.01335f
C121 Nand_Gate_6.B EN 1.25083f
C122 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_89921_15797# 0.05964f
C123 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.06445f
C124 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout VDD 1.56255f
C125 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_0.Vout 1.00121f
C126 a_128237_26914# D_FlipFlop_5.Nand_Gate_0.Vout 0.04444f
C127 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout VDD 2.88547f
C128 D_FlipFlop_1.3-input-nand_1.Vout VDD 1.7803f
C129 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout CLK 0.29644f
C130 CDAC8_0.switch_9.Z VDD 12.5515f
C131 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout a_52727_13083# 0.04995f
C132 a_57415_13083# EN 0.0452f
C133 FFCLR a_128851_36157# 0.04623f
C134 Nand_Gate_2.A RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.08377f
C135 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.30154f
C136 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout VDD 1.76876f
C137 a_134283_30478# a_134897_30478# 0.05935f
C138 a_91279_52572# Nand_Gate_2.A 0.06113f
C139 RingCounter_0.D_FlipFlop_5.Q' a_101705_49858# 0.01335f
C140 D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.48313f
C141 a_72835_15797# RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.04444f
C142 a_33363_15797# VDD 0.02954f
C143 CDAC8_0.switch_9.Z CDAC8_0.switch_1.Z 0.14339f
C144 Nand_Gate_2.B EN 0.99738f
C145 a_78881_13083# a_79495_13083# 0.05935f
C146 Nand_Gate_6.B a_90535_15797# 0.04995f
C147 a_79495_13083# VDD 0.01327f
C148 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_99603_13083# 0.01335f
C149 a_128851_23350# Nand_Gate_7.B 0.04723f
C150 Nand_Gate_7.B VDD 8.0573f
C151 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout VDD 2.13993f
C152 a_75898_28676# Q3 0.49857f
C153 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.0857f
C154 a_128237_33443# a_128851_33443# 0.05935f
C155 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_98245_52572# 0.04444f
C156 CLK Q7 0.1175f
C157 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout CLK 0.70923f
C158 Nand_Gate_7.B CDAC8_0.switch_1.Z 0.33175f
C159 D_FlipFlop_7.Q' VDD 1.89473f
C160 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout VDD 2.07373f
C161 D_FlipFlop_7.3-input-nand_0.Vout a_134283_19786# 0.05964f
C162 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout VDD 1.48368f
C163 a_75898_28676# VDD 1.30969f
C164 a_106699_52572# a_107313_52572# 0.05935f
C165 Nand_Gate_6.A RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.08377f
C166 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.30154f
C167 a_128237_19786# Q0 0.06113f
C168 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout CLK 0.20785f
C169 a_128851_26914# Nand_Gate_6.B 0.04727f
C170 a_66483_13083# CLK 0.03129f
C171 D_FlipFlop_6.Nand_Gate_0.Vout a_130209_23350# 0.05964f
C172 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout VDD 2.46653f
C173 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.30154f
C174 a_86591_49858# VDD 0.06071f
C175 Comparator_0.Vinm a_75898_21528# 0.04177f
C176 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.06594f
C177 a_28675_15797# RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.04444f
C178 a_53471_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.01335f
C179 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121069_15797# 0.05964f
C180 RingCounter_0.D_FlipFlop_15.Q' a_50755_15797# 0.04443f
C181 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_90665_52572# 0.04995f
C182 D_FlipFlop_3.Nand_Gate_1.Vout D_FlipFlop_2.Nand_Gate_0.Vout 0.01681f
C183 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C EN 0.07732f
C184 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_57415_13083# 0.01335f
C185 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_52727_13083# 0.05964f
C186 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_95659_49858# 0.01335f
C187 a_51499_52572# VDD 0.0564f
C188 RingCounter_0.D_FlipFlop_7.Q' RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.11654f
C189 a_134897_17072# VDD 0.01186f
C190 Nand_Gate_2.B a_106699_52572# 0.04995f
C191 D_FlipFlop_5.Nand_Gate_0.Vout a_130209_26914# 0.05964f
C192 D_FlipFlop_4.Q' D_FlipFlop_4.Nand_Gate_0.Vout 0.06632f
C193 Comparator_0.Vinm Q7 0.7705f
C194 RingCounter_0.D_FlipFlop_3.Q' VDD 1.96503f
C195 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout a_117739_49858# 0.04995f
C196 a_128237_27764# Q3 0.04443f
C197 D_FlipFlop_0.Nand_Gate_0.Vout Q4 0.11443f
C198 a_56801_13083# a_57415_13083# 0.05935f
C199 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_106569_15797# 0.04995f
C200 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout EN 0.97349f
C201 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout CLK 0.23464f
C202 a_78267_52572# RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.04443f
C203 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_52113_49858# 0.05964f
C204 D_FlipFlop_2.Q' D_FlipFlop_2.Nand_Gate_1.Vout 0.11654f
C205 a_35335_13083# VDD 0.01327f
C206 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_45147_49858# 0.05964f
C207 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_99603_15797# 0.01335f
C208 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_40459_49858# 0.01335f
C209 D_FlipFlop_5.3-input-nand_2.Vout VDD 2.77266f
C210 D_FlipFlop_0.Nand_Gate_1.Vout a_128237_44135# 0.04444f
C211 RingCounter_0.D_FlipFlop_8.Q' VDD 1.95446f
C212 D_FlipFlop_0.Q' VDD 1.89794f
C213 a_128237_27764# VDD 0.02521f
C214 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_0.Vout 1.00205f
C215 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout VDD 2.73618f
C216 a_92725_16975# CLK 0.04479f
C217 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.06503f
C218 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.06445f
C219 FFCLR D_FlipFlop_3.3-input-nand_2.Vout 0.06105f
C220 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout a_107927_15797# 0.04443f
C221 D_FlipFlop_1.Nand_Gate_1.Vout VDD 1.46545f
C222 D_FlipFlop_2.Q' Q6 1.06174f
C223 FFCLR D_FlipFlop_5.Inverter_0.Vout 0.43823f
C224 FFCLR D_FlipFlop_1.Nand_Gate_0.Vout 0.64823f
C225 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_76909_15797# 0.05964f
C226 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.25579f
C227 D_FlipFlop_4.3-input-nand_2.C a_132311_27764# 0.05964f
C228 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_3.3-input-nand_2.Vout 0.01194f
C229 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.C 0.01194f
C230 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_17.Inverter_0.Vout 0.29368f
C231 D_FlipFlop_7.Inverter_1.Vout VDD 1.73058f
C232 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.16429f
C233 a_42431_49858# VDD 0.01186f
C234 a_134283_17072# a_134897_17072# 0.05935f
C235 a_78881_15797# VDD 0.03119f
C236 Nand_Gate_2.A CLK 0.63966f
C237 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_108671_52572# 0.04995f
C238 a_105955_13083# VDD 0.02521f
C239 D_FlipFlop_7.3-input-nand_1.Vout a_132925_17072# 0.04543f
C240 a_130209_23350# D_FlipFlop_6.3-input-nand_2.Vout 0.04443f
C241 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_65869_13083# 0.05964f
C242 CDAC8_0.switch_5.Z EN 1.03162f
C243 a_110643_15797# VDD 0.03339f
C244 FFCLR D_FlipFlop_4.Q' 0.03748f
C245 D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_7.B 0.67495f
C246 a_80239_52572# RingCounter_0.D_FlipFlop_3.Q' 0.04443f
C247 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_54829_13083# 0.04443f
C248 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.04107f
C249 Nand_Gate_5.B Q6 0.06203f
C250 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout VDD 2.04843f
C251 a_34721_13083# a_35335_13083# 0.05935f
C252 a_101705_52572# VDD 0.01186f
C253 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout CLK 0.03574f
C254 a_128851_19786# VDD 0.01186f
C255 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_97631_49858# 0.01335f
C256 a_130209_26914# D_FlipFlop_5.3-input-nand_2.Vout 0.04443f
C257 a_89921_13083# CLK 0.04619f
C258 D_FlipFlop_4.Inverter_0.Vout VDD 1.37371f
C259 a_54085_52572# VDD 0.02521f
C260 CDAC8_0.switch_7.Z Q2 1.5084f
C261 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.1182f
C262 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Inverter_1.Vout 0.25963f
C263 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout a_122427_49858# 0.04995f
C264 D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_6.B 0.67535f
C265 D_FlipFlop_6.3-input-nand_2.C VDD 2.74431f
C266 Nand_Gate_6.A a_82057_16975# 0.0476f
C267 a_109285_49858# VDD 0.0301f
C268 Nand_Gate_6.Vout CLK 2.60401f
C269 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.0857f
C270 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout m3_125329_49141# 0.01611f
C271 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout VDD 2.01342f
C272 a_130209_33443# VDD 0.02521f
C273 a_45147_52572# RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.05964f
C274 a_75898_18814# Nand_Gate_4.B 0.03201f
C275 CDAC8_0.switch_0.Z CLK 0.16657f
C276 FFCLR D_FlipFlop_5.3-input-nand_1.Vout 0.95389f
C277 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_32749_15797# 0.05964f
C278 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_56187_49858# 0.05964f
C279 Nand_Gate_2.A Comparator_0.Vinm 4.04825f
C280 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout VDD 1.86552f
C281 D_FlipFlop_6.Nand_Gate_1.Vout a_130209_20636# 0.05964f
C282 Nand_Gate_6.B Nand_Gate_7.B 0.05683f
C283 Nand_Gate_1.B a_134897_27764# 0.04544f
C284 D_FlipFlop_1.Inverter_1.Vout a_130209_36157# 0.04443f
C285 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout CLK 0.155f
C286 FFCLR a_128851_20636# 0.04443f
C287 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout VDD 1.76876f
C288 Nand_Gate_2.B RingCounter_0.D_FlipFlop_7.Inverter_0.Vout 0.29368f
C289 D_FlipFlop_4.Nand_Gate_0.Vout a_128851_30478# 0.04995f
C290 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.06465f
C291 a_139696_27690# Vin 0.49f
C292 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_0.Vout 0.06594f
C293 CDAC8_0.switch_8.Z Q6 0.24676f
C294 a_96273_49858# CLK 0.04619f
C295 a_61795_13083# VDD 0.02521f
C296 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C VDD 3.56545f
C297 D_FlipFlop_5.Nand_Gate_1.Vout a_130209_24200# 0.05964f
C298 a_134897_37007# VDD 0.01186f
C299 a_51369_15797# EN 0.04443f
C300 a_109285_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.04443f
C301 D_FlipFlop_4.3-input-nand_1.Vout VDD 1.78032f
C302 Comparator_0.Vinm CDAC8_0.switch_0.Z 25.94f
C303 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout VDD 2.16362f
C304 Nand_Gate_4.B Q0 1.41224f
C305 FFCLR D_FlipFlop_4.Inverter_1.Vout 0.56808f
C306 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_2.Vout 0.92942f
C307 a_56801_15797# CLK 0.04619f
C308 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_89307_49858# 0.04443f
C309 a_45761_13083# CLK 0.04619f
C310 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.16429f
C311 a_128237_43285# VDD 0.02521f
C312 CDAC8_0.switch_6.Z Q3 0.78009f
C313 a_128851_39721# Q6 0.01335f
C314 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.0846f
C315 a_65125_49858# VDD 0.0301f
C316 a_43789_15797# a_44403_15797# 0.05935f
C317 FFCLR a_48937_47663# 0.04705f
C318 a_123655_15797# VDD 0.05687f
C319 Nand_Gate_2.Vout CLK 2.32087f
C320 Nand_Gate_4.B EN 1.52428f
C321 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout CLK 0.29759f
C322 CDAC8_0.switch_6.Z VDD 13.0121f
C323 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_2.Vout 0.92857f
C324 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout EN 0.1313f
C325 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C EN 0.07732f
C326 a_61795_15797# a_62409_15797# 0.05935f
C327 a_48565_16975# VDD 0.02521f
C328 RingCounter_0.D_FlipFlop_7.Q' a_113359_49858# 0.06113f
C329 D_FlipFlop_1.Nand_Gate_1.Vout a_128851_33443# 0.04995f
C330 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_55443_15797# 0.04995f
C331 a_52727_15797# VDD 0.02906f
C332 FFCLR D_FlipFlop_0.3-input-nand_1.Vout 0.95389f
C333 D_FlipFlop_7.Nand_Gate_1.Vout Q0 0.06503f
C334 a_132311_26914# VDD 0.02521f
C335 a_52113_49858# CLK 0.04619f
C336 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout VDD 1.48392f
C337 D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.48313f
C338 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_1.Vout 0.08671f
C339 a_87949_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.04444f
C340 a_132925_23350# VDD 0.01186f
C341 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout CLK 0.12047f
C342 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout VDD 2.8604f
C343 D_FlipFlop_7.Q' a_128237_19786# 0.04443f
C344 FFCLR D_FlipFlop_5.Nand_Gate_1.Vout 0.60828f
C345 Nand_Gate_2.Vout Comparator_0.Vinm 0.04618f
C346 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.08671f
C347 a_53471_52572# a_54085_52572# 0.05935f
C348 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_43789_13083# 0.05964f
C349 a_35335_15797# VDD 0.06072f
C350 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.3-input-nand_2.Vout 0.16429f
C351 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C CLK 0.30966f
C352 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout CLK 0.70923f
C353 CDAC8_0.switch_9.Z CDAC8_0.switch_5.Z 1.1471f
C354 Nand_Gate_6.B RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0839f
C355 a_119711_49858# CLK 0.02953f
C356 a_84489_13083# VDD 0.0563f
C357 D_FlipFlop_3.3-input-nand_0.Vout a_132925_43285# 0.04995f
C358 a_108671_49858# a_109285_49858# 0.05935f
C359 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.0857f
C360 a_120325_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.05964f
C361 D_FlipFlop_4.Nand_Gate_1.Vout Q3 0.06503f
C362 a_45147_52572# RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.04443f
C363 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout a_78267_52572# 0.04443f
C364 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Nand_Gate_1.Vout 0.04109f
C365 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.08671f
C366 Nand_Gate_2.A Q4 0.06203f
C367 Nand_Gate_0.A Nand_Gate_0.B 0.07727f
C368 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 0.25579f
C369 a_75551_52572# EN 0.045f
C370 D_FlipFlop_0.Inverter_0.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.0857f
C371 a_75898_46095# VDD 1.30093f
C372 RingCounter_0.D_FlipFlop_14.Q' RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.11654f
C373 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.25963f
C374 a_107313_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.05964f
C375 D_FlipFlop_4.Nand_Gate_1.Vout VDD 1.46545f
C376 D_FlipFlop_4.Inverter_1.Vout a_130209_30478# 0.04443f
C377 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_65869_15797# 0.04443f
C378 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout EN 0.24886f
C379 a_101705_52572# Nand_Gate_2.B 0.01335f
C380 a_110029_15797# VDD 0.03178f
C381 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout CLK 0.03479f
C382 a_89307_49858# VDD 0.04111f
C383 Nand_Gate_5.B Q0 0.06203f
C384 D_FlipFlop_2.Nand_Gate_0.Vout Q6 0.11443f
C385 a_75898_28676# CDAC8_0.switch_5.Z 0.29583f
C386 D_FlipFlop_6.3-input-nand_1.Vout a_132925_20636# 0.04543f
C387 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 1.09975f
C388 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.04109f
C389 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout EN 0.78734f
C390 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.06503f
C391 Nand_Gate_5.B a_115177_47663# 0.04443f
C392 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout CLK 0.29644f
C393 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Q' 0.06632f
C394 FFCLR D_FlipFlop_2.3-input-nand_2.Vout 0.06399f
C395 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_97631_49858# 0.04543f
C396 Nand_Gate_2.B RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.08377f
C397 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.C 1.09975f
C398 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout VDD 1.86552f
C399 D_FlipFlop_1.Q' Q6 0.01194f
C400 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout CLK 0.23464f
C401 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout a_85847_15797# 0.04443f
C402 Nand_Gate_5.B EN 0.57932f
C403 a_75551_49858# CLK 0.03129f
C404 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_54085_49858# 0.04444f
C405 FFCLR D_FlipFlop_0.Nand_Gate_1.Vout 0.60828f
C406 a_40329_13083# VDD 0.0563f
C407 D_FlipFlop_5.3-input-nand_1.Vout a_132925_24200# 0.04543f
C408 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_47119_49858# 0.04444f
C409 a_86591_49858# a_87205_49858# 0.05935f
C410 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout VDD 2.07373f
C411 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_42431_49858# 0.04543f
C412 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout CLK 0.03574f
C413 D_FlipFlop_0.Nand_Gate_1.Vout a_130209_44135# 0.05964f
C414 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_2.Vout 0.88509f
C415 a_130209_27764# VDD 0.02521f
C416 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.C 1.09975f
C417 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.Nand_Gate_1.Vout 0.1541f
C418 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.1541f
C419 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout EN 0.24889f
C420 a_114805_16975# CLK 0.06046f
C421 a_134283_37007# a_134897_37007# 0.05935f
C422 a_66483_15797# VDD 0.03339f
C423 D_FlipFlop_6.3-input-nand_0.Vout VDD 1.77946f
C424 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_63767_15797# 0.05964f
C425 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.30154f
C426 D_FlipFlop_3.Inverter_1.Vout VDD 1.73058f
C427 D_FlipFlop_0.Q' a_128237_46849# 0.04443f
C428 a_128237_19786# a_128851_19786# 0.05935f
C429 CDAC8_0.switch_6.Z Nand_Gate_6.B 4.08114f
C430 a_45761_15797# CLK 0.04619f
C431 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Q' 1.05791f
C432 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout VDD 2.31704f
C433 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_109285_49858# 0.05964f
C434 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout a_78881_13083# 0.04443f
C435 RingCounter_0.D_FlipFlop_17.Q' a_46505_49858# 0.01335f
C436 a_45147_49858# VDD 0.04055f
C437 a_51499_52572# a_52113_52572# 0.05935f
C438 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.3-input-nand_2.C 0.25579f
C439 a_59605_47663# CLK 0.04443f
C440 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout VDD 2.46653f
C441 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout VDD 1.70415f
C442 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.C 0.06594f
C443 CDAC8_0.switch_9.Z Nand_Gate_4.B 1.76363f
C444 a_107927_13083# VDD 0.02578f
C445 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.06465f
C446 a_76909_15797# VDD 0.03178f
C447 D_FlipFlop_7.3-input-nand_1.Vout a_134897_17072# 0.01335f
C448 CDAC8_0.switch_8.Z EN 1.97671f
C449 Nand_Gate_1.B CLK 0.66757f
C450 a_112615_15797# VDD 0.06072f
C451 And_Gate_4.Inverter_0.Vin EN 0.0623f
C452 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout VDD 1.56255f
C453 D_FlipFlop_1.3-input-nand_1.Vout a_132311_33443# 0.04444f
C454 RingCounter_0.D_FlipFlop_9.Q' RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.06632f
C455 D_FlipFlop_7.3-input-nand_2.C a_132311_17072# 0.05964f
C456 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout EN 0.97489f
C457 a_73579_52572# VDD 0.0564f
C458 Nand_Gate_5.A a_117739_52572# 0.04995f
C459 FFCLR D_FlipFlop_0.3-input-nand_2.C 0.76213f
C460 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout a_45761_13083# 0.04443f
C461 a_130209_19786# VDD 0.02521f
C462 RingCounter_0.D_FlipFlop_5.Q' VDD 1.96503f
C463 Nand_Gate_7.B Nand_Gate_4.B 0.0623f
C464 D_FlipFlop_0.3-input-nand_2.C a_130209_44135# 0.04443f
C465 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_100347_49858# 0.04443f
C466 a_64511_49858# a_65125_49858# 0.05935f
C467 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_101705_49858# 0.04995f
C468 RingCounter_0.D_FlipFlop_8.Q' a_39715_13083# 0.06113f
C469 EN Q5 0.2481f
C470 D_FlipFlop_0.3-input-nand_2.Vout a_132311_46849# 0.05964f
C471 a_65125_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.05964f
C472 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout Nand_Gate_2.B 0.12214f
C473 a_112745_49858# VDD 0.06015f
C474 a_132925_33443# VDD 0.01186f
C475 D_FlipFlop_7.Q' Nand_Gate_4.B 0.06645f
C476 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_58159_49858# 0.04444f
C477 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout a_123655_13083# 0.04995f
C478 a_128237_27764# a_128851_27764# 0.05935f
C479 D_FlipFlop_2.3-input-nand_2.Vout a_132311_39721# 0.05964f
C480 RingCounter_0.D_FlipFlop_16.Q VDD 3.43364f
C481 a_123041_15797# a_123655_15797# 0.05935f
C482 FFCLR a_134897_19786# 0.08419f
C483 a_121069_15797# a_121683_15797# 0.05935f
C484 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.04109f
C485 Nand_Gate_1.B Comparator_0.Vinm 1.25742f
C486 a_75898_39392# CDAC8_0.switch_6.Z 0.29045f
C487 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout VDD 2.07373f
C488 D_FlipFlop_6.3-input-nand_2.Vout a_132925_23350# 0.01335f
C489 a_128237_39721# VDD 0.02521f
C490 RingCounter_0.D_FlipFlop_6.Q' a_124399_49858# 0.06113f
C491 CDAC8_0.switch_7.Z Q3 1.50848f
C492 D_FlipFlop_4.Nand_Gate_0.Vout a_130209_30478# 0.05964f
C493 RingCounter_0.D_FlipFlop_13.Q' VDD 1.95446f
C494 RingCounter_0.D_FlipFlop_16.Q a_28675_15797# 0.07417f
C495 a_98245_49858# CLK 0.03129f
C496 a_63767_13083# VDD 0.02578f
C497 Nand_Gate_5.A CLK 0.88296f
C498 D_FlipFlop_3.Q' a_128237_43285# 0.04443f
C499 FFCLR D_FlipFlop_0.Inverter_0.Vout 0.43576f
C500 Nand_Gate_4.B a_134897_17072# 0.04583f
C501 Nand_Gate_0.A VDD 8.23952f
C502 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_118967_13083# 0.04443f
C503 CDAC8_0.switch_7.Z VDD 26.5647f
C504 RingCounter_0.D_FlipFlop_12.Q' a_84489_13083# 0.01335f
C505 Nand_Gate_5.B RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.07174f
C506 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.30154f
C507 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout CLK 0.30735f
C508 a_128851_46849# VDD 0.01186f
C509 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_53471_52572# 0.04995f
C510 D_FlipFlop_7.Q' D_FlipFlop_7.Nand_Gate_1.Vout 0.11654f
C511 D_FlipFlop_5.3-input-nand_2.Vout a_132925_26914# 0.01335f
C512 D_FlipFlop_0.3-input-nand_2.Vout a_132311_44135# 0.04443f
C513 D_FlipFlop_0.3-input-nand_0.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.04107f
C514 And_Gate_7.Inverter_0.Vin VDD 1.43162f
C515 a_46505_49858# EN 0.04443f
C516 FFCLR D_FlipFlop_3.3-input-nand_1.Vout 0.95389f
C517 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout EN 0.97489f
C518 a_123785_52572# VDD 0.01186f
C519 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout CLK 0.15609f
C520 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout EN 0.13192f
C521 a_42431_49858# a_43045_49858# 0.05935f
C522 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.0846f
C523 a_128237_19786# D_FlipFlop_7.Nand_Gate_0.Vout 0.04444f
C524 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout EN 0.24889f
C525 a_76165_52572# VDD 0.02521f
C526 a_78881_15797# a_79495_15797# 0.05935f
C527 Nand_Gate_4.A CLK 0.20423f
C528 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout CLK 0.03479f
C529 a_76909_15797# a_77523_15797# 0.05935f
C530 a_68585_49858# VDD 0.06015f
C531 a_105955_13083# a_106569_13083# 0.05935f
C532 RingCounter_0.D_FlipFlop_1.Q' RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.11654f
C533 Comparator_0.Vinm CLK 2.97464f
C534 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout VDD 2.73332f
C535 a_68585_52572# EN 0.04443f
C536 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_45761_15797# 0.05964f
C537 Nand_Gate_5.A Comparator_0.Vinm 1.94937f
C538 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout VDD 2.01968f
C539 D_FlipFlop_6.3-input-nand_2.C a_132311_23350# 0.04443f
C540 Nand_Gate_1.Vout a_104137_16975# 0.05964f
C541 Nand_Gate_7.B a_59977_16975# 0.04443f
C542 a_70645_16975# VDD 0.02521f
C543 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.Inverter_1.Vout 0.25963f
C544 Nand_Gate_4.B D_FlipFlop_7.Inverter_1.Vout 0.16546f
C545 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout CLK 0.155f
C546 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_57415_15797# 0.01335f
C547 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout VDD 1.76876f
C548 Nand_Gate_5.A RingCounter_0.D_FlipFlop_6.Inverter_0.Vout 0.29368f
C549 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout a_42431_52572# 0.04995f
C550 a_54085_49858# CLK 0.03129f
C551 CDAC8_0.switch_6.Z CDAC8_0.switch_5.Z 3.08882f
C552 D_FlipFlop_0.3-input-nand_1.Vout a_132925_44135# 0.04543f
C553 CDAC8_0.switch_0.Z Q2 0.50649f
C554 D_FlipFlop_5.3-input-nand_2.C a_132311_26914# 0.04443f
C555 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.16429f
C556 Nand_Gate_6.A a_84489_15797# 0.01335f
C557 RingCounter_0.D_FlipFlop_10.Q' RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.06632f
C558 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.3-input-nand_2.C 0.25579f
C559 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C EN 0.07664f
C560 a_134283_23350# VDD 0.02521f
C561 D_FlipFlop_2.Nand_Gate_1.Vout D_FlipFlop_1.Nand_Gate_0.Vout 0.01681f
C562 Nand_Gate_5.B Nand_Gate_7.B 0.06463f
C563 a_101705_52572# a_102319_52572# 0.05935f
C564 RingCounter_0.D_FlipFlop_9.Q' CLK 0.09276f
C565 a_128851_19786# Nand_Gate_4.B 0.04685f
C566 a_34721_15797# a_35335_15797# 0.05935f
C567 a_32749_15797# a_33363_15797# 0.05935f
C568 RingCounter_0.D_FlipFlop_15.Q' CLK 0.09276f
C569 And_Gate_7.Inverter_0.Vin a_125845_47663# 0.05964f
C570 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout EN 0.07459f
C571 Nand_Gate_5.Vout And_Gate_7.Inverter_0.Vin 0.10129f
C572 D_FlipFlop_6.Inverter_0.Vout a_134897_20636# 0.04995f
C573 a_54085_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.04443f
C574 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.Nand_Gate_1.Vout 0.30154f
C575 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout VDD 1.99837f
C576 D_FlipFlop_1.Q' EN 0.04711f
C577 CDAC8_0.switch_8.Z CDAC8_0.switch_9.Z 7.4006f
C578 a_83875_13083# a_84489_13083# 0.05935f
C579 D_FlipFlop_3.Nand_Gate_1.Vout a_128237_40571# 0.04444f
C580 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_0.Vout 0.0846f
C581 D_FlipFlop_3.3-input-nand_2.C a_132311_40571# 0.05964f
C582 a_87949_13083# VDD 0.02578f
C583 D_FlipFlop_3.3-input-nand_0.Vout a_134897_43285# 0.01335f
C584 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout a_63767_13083# 0.04995f
C585 a_128237_43285# a_128851_43285# 0.05935f
C586 FFCLR D_FlipFlop_1.3-input-nand_2.Vout 0.88667f
C587 Nand_Gate_7.A a_57415_15797# 0.04995f
C588 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout CLK 0.29759f
C589 D_FlipFlop_5.Inverter_0.Vout a_134897_24200# 0.04995f
C590 RingCounter_0.D_FlipFlop_15.Q' a_50755_13083# 0.06113f
C591 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C EN 0.07732f
C592 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.30154f
C593 D_FlipFlop_0.Nand_Gate_0.Vout VDD 1.48313f
C594 RingCounter_0.D_FlipFlop_13.Q' RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout 0.06632f
C595 CDAC8_0.switch_9.Z Q5 0.65428f
C596 Q1 Q0 0.01156f
C597 a_134283_46849# a_134897_46849# 0.05935f
C598 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_106699_49858# 0.01335f
C599 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_0.Vout 0.0846f
C600 FFCLR D_FlipFlop_3.Nand_Gate_1.Vout 0.60828f
C601 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_120325_49858# 0.05964f
C602 RingCounter_0.D_FlipFlop_5.Q' Nand_Gate_2.B 1.10693f
C603 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.48398f
C604 FFCLR a_132925_24200# 0.045f
C605 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_63153_49858# 0.05964f
C606 a_91279_49858# VDD 0.02906f
C607 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.08671f
C608 D_FlipFlop_6.3-input-nand_1.Vout a_134897_20636# 0.01335f
C609 RingCounter_0.D_FlipFlop_4.Q' RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.11654f
C610 a_63153_52572# CLK 0.04619f
C611 D_FlipFlop_1.Q' a_128237_33443# 0.06113f
C612 EN Q1 0.2481f
C613 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout VDD 2.8604f
C614 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout EN 0.60828f
C615 a_132311_23350# a_132925_23350# 0.05935f
C616 D_FlipFlop_2.Inverter_1.Vout VDD 1.73058f
C617 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout a_35335_13083# 0.04995f
C618 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.0857f
C619 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_2.Vout 0.92808f
C620 CDAC8_0.switch_7.Z Nand_Gate_6.B 7.53946f
C621 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.0846f
C622 a_61795_13083# a_62409_13083# 0.05935f
C623 a_100347_52572# RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.05964f
C624 a_41073_52572# CLK 0.04443f
C625 a_117739_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.01335f
C626 D_FlipFlop_1.Inverter_0.Vout a_134283_33443# 0.04443f
C627 a_43789_13083# VDD 0.02578f
C628 D_FlipFlop_5.3-input-nand_1.Vout a_134897_24200# 0.01335f
C629 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C EN 0.07664f
C630 a_95529_15797# VDD 0.01571f
C631 CDAC8_0.switch_6.Z Nand_Gate_4.B 3.52726f
C632 FFCLR D_FlipFlop_0.3-input-nand_0.Vout 0.08617f
C633 a_128237_23350# Q1 0.06113f
C634 RingCounter_0.D_FlipFlop_16.Q' RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.11654f
C635 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.0846f
C636 RingCounter_0.D_FlipFlop_16.Q' RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.06632f
C637 D_FlipFlop_7.3-input-nand_2.C VDD 2.74431f
C638 CLK Q4 0.11898f
C639 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 1.09975f
C640 Nand_Gate_3.B CLK 0.27944f
C641 a_132311_26914# a_132925_26914# 0.05935f
C642 a_132925_27764# VDD 0.01186f
C643 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout EN 0.06649f
C644 Nand_Gate_5.A Q4 0.46277f
C645 D_FlipFlop_6.Q' a_128237_20636# 0.06113f
C646 D_FlipFlop_0.3-input-nand_2.C D_FlipFlop_0.3-input-nand_0.Vout 0.06594f
C647 Nand_Gate_7.B a_67841_15797# 0.04443f
C648 a_68455_15797# VDD 0.06072f
C649 a_97631_52572# EN 0.045f
C650 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_30647_13083# 0.04443f
C651 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_102319_52572# 0.04444f
C652 D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_4.B 0.66417f
C653 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.06465f
C654 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout CLK 0.15609f
C655 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_0.Vout 0.06594f
C656 a_50755_15797# VDD 0.02906f
C657 D_FlipFlop_4.Nand_Gate_1.Vout a_128851_27764# 0.04995f
C658 a_67227_52572# VDD 0.02521f
C659 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.06503f
C660 a_47119_49858# VDD 0.02906f
C661 a_52113_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.05964f
C662 a_81685_47663# CLK 0.07396f
C663 a_110643_13083# VDD 0.05686f
C664 D_FlipFlop_5.Q' a_128237_24200# 0.06113f
C665 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.06445f
C666 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout CLK 0.27229f
C667 Nand_Gate_0.A a_75898_39392# 0.01513f
C668 a_130209_43285# VDD 0.02521f
C669 Comparator_0.Vinm Q4 1.26254f
C670 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_67227_49858# 0.05964f
C671 Nand_Gate_3.B Comparator_0.Vinm 0.03473f
C672 D_FlipFlop_1.3-input-nand_1.Vout a_134283_33443# 0.05964f
C673 a_128237_43285# D_FlipFlop_3.Nand_Gate_0.Vout 0.04444f
C674 FFCLR a_132925_44135# 0.045f
C675 Nand_Gate_5.A RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.08377f
C676 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout VDD 1.86552f
C677 a_134897_26914# VDD 0.01186f
C678 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C CLK 0.30901f
C679 a_95659_49858# EN 0.07058f
C680 a_113359_52572# Nand_Gate_5.A 0.06113f
C681 a_128237_36157# VDD 0.02521f
C682 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 1.09975f
C683 a_69199_52572# VDD 0.02521f
C684 a_39715_13083# a_40329_13083# 0.05935f
C685 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Nand_Gate_1.Vout 0.04109f
C686 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_76909_13083# 0.05964f
C687 D_FlipFlop_0.3-input-nand_2.C a_132925_44135# 0.01335f
C688 a_75898_21528# VDD 1.33597f
C689 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout EN 0.06649f
C690 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_110643_15797# 0.04995f
C691 FFCLR D_FlipFlop_3.Inverter_0.Vout 0.43823f
C692 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_65869_13083# 0.04443f
C693 D_FlipFlop_4.3-input-nand_1.Vout D_FlipFlop_5.3-input-nand_0.Vout 0.01418f
C694 a_117739_49858# VDD 0.01712f
C695 a_46505_52572# FFCLR 0.01335f
C696 a_134897_33443# VDD 0.01186f
C697 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_120325_52572# 0.04444f
C698 Nand_Gate_2.Vout a_103765_47663# 0.04443f
C699 a_55443_15797# EN 0.045f
C700 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_123041_15797# 0.05964f
C701 VDD Q7 3.793f
C702 FFCLR D_FlipFlop_2.3-input-nand_1.Vout 0.95519f
C703 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout EN 0.09127f
C704 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout VDD 2.73618f
C705 a_132311_23350# D_FlipFlop_6.3-input-nand_0.Vout 0.04444f
C706 FFCLR D_FlipFlop_4.3-input-nand_2.C 0.76213f
C707 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout EN 0.06649f
C708 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout VDD 2.41001f
C709 a_66483_13083# VDD 0.05686f
C710 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout EN 0.24889f
C711 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.08671f
C712 Nand_Gate_1.A a_105955_15797# 0.06113f
C713 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.16415f
C714 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 1.09975f
C715 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121683_13083# 0.01335f
C716 a_75551_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.01335f
C717 a_52727_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.04443f
C718 a_132925_19786# VDD 0.01186f
C719 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_112745_52572# 0.04995f
C720 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout EN 0.61894f
C721 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.C 0.06594f
C722 Nand_Gate_5.B a_123655_15797# 0.04995f
C723 a_132311_26914# D_FlipFlop_5.3-input-nand_0.Vout 0.04444f
C724 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout EN 0.08852f
C725 a_95659_52572# VDD 0.0564f
C726 a_128237_20636# VDD 0.02521f
C727 a_51499_49858# EN 0.07058f
C728 D_FlipFlop_0.3-input-nand_0.Vout a_132925_46849# 0.04995f
C729 RingCounter_0.D_FlipFlop_6.Q' VDD 1.93578f
C730 a_128237_46849# a_128851_46849# 0.05935f
C731 a_62539_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.01335f
C732 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_84489_15797# 0.04995f
C733 CDAC8_0.switch_7.Z CDAC8_0.switch_5.Z 3.08191f
C734 a_100347_52572# RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.04443f
C735 D_FlipFlop_2.3-input-nand_0.Vout a_132925_39721# 0.04995f
C736 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_78881_15797# 0.05964f
C737 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout VDD 2.88547f
C738 RingCounter_0.D_FlipFlop_13.Q' RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.11654f
C739 Nand_Gate_1.B Q2 0.05915f
C740 a_73579_49858# VDD 0.01712f
C741 CDAC8_0.switch_9.Z Q1 0.36574f
C742 Nand_Gate_6.B a_95529_15797# 0.01335f
C743 D_FlipFlop_3.Inverter_0.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.0857f
C744 a_112001_15797# a_112615_15797# 0.05935f
C745 a_92725_16975# VDD 0.02521f
C746 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.3-input-nand_2.Vout 0.06445f
C747 Nand_Gate_1.A a_104137_16975# 0.0476f
C748 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.06465f
C749 a_61795_15797# RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.04444f
C750 CDAC8_0.switch_2.Z EN 0.26953f
C751 Nand_Gate_3.B a_63153_52572# 0.04443f
C752 a_118353_49858# EN 0.01149f
C753 CDAC8_0.switch_8.Z CDAC8_0.switch_6.Z 3.59863f
C754 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.25579f
C755 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C CLK 0.30966f
C756 Nand_Gate_7.B Q1 0.35004f
C757 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.06594f
C758 D_FlipFlop_0.3-input-nand_1.Vout a_134897_44135# 0.01335f
C759 a_40459_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.01335f
C760 a_121069_13083# CLK 0.03129f
C761 a_128237_43285# Q5 0.06113f
C762 Nand_Gate_2.A VDD 7.94482f
C763 D_FlipFlop_6.Inverter_0.Vout VDD 1.3737f
C764 D_FlipFlop_7.Q' Q1 0.01194f
C765 a_102319_52572# RingCounter_0.D_FlipFlop_5.Q' 0.04443f
C766 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_34721_15797# 0.05964f
C767 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout CLK 0.06496f
C768 CDAC8_0.switch_6.Z Q5 0.58263f
C769 D_FlipFlop_4.3-input-nand_1.Vout a_132311_27764# 0.04444f
C770 CLK Q2 0.1175f
C771 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_7.3-input-nand_2.Vout 0.01194f
C772 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.C 0.01194f
C773 CDAC8_0.switch_9.Z a_75898_25104# 0.01232f
C774 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.1541f
C775 D_FlipFlop_1.Q' D_FlipFlop_1.Nand_Gate_1.Vout 0.11654f
C776 FFCLR D_FlipFlop_2.Nand_Gate_1.Vout 0.61212f
C777 RingCounter_0.D_FlipFlop_11.Q' a_94915_15797# 0.04443f
C778 a_98245_52572# VDD 0.02521f
C779 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout VDD 2.16362f
C780 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.30154f
C781 D_FlipFlop_3.Nand_Gate_1.Vout a_130209_40571# 0.05964f
C782 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout CLK 0.30735f
C783 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.06503f
C784 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout CLK 0.03436f
C785 a_89921_13083# VDD 0.02865f
C786 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.06594f
C787 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.08671f
C788 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_65125_52572# 0.04444f
C789 a_132311_33443# a_132925_33443# 0.05935f
C790 a_90665_52572# EN 0.04443f
C791 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.06503f
C792 Nand_Gate_6.Vout VDD 1.36733f
C793 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Inverter_1.Vout 0.25963f
C794 CDAC8_0.switch_0.Z VDD 1.38984f
C795 Nand_Gate_7.A RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.08377f
C796 D_FlipFlop_1.Inverter_1.Vout VDD 1.73058f
C797 D_FlipFlop_7.3-input-nand_0.Vout VDD 1.77946f
C798 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.06465f
C799 a_74193_49858# EN 0.01149f
C800 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_108671_49858# 0.04543f
C801 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout CLK 0.23464f
C802 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout VDD 1.76876f
C803 D_FlipFlop_6.3-input-nand_1.Vout VDD 1.78032f
C804 a_76909_13083# CLK 0.03129f
C805 D_FlipFlop_6.Q' D_FlipFlop_6.Nand_Gate_1.Vout 0.11654f
C806 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_88563_15797# 0.01335f
C807 CDAC8_0.switch_7.Z Nand_Gate_4.B 4.09248f
C808 Comparator_0.Vinm Q2 1.64422f
C809 FFCLR D_FlipFlop_6.Inverter_1.Vout 0.56927f
C810 a_75898_46095# CDAC8_0.switch_8.Z 0.33725f
C811 a_128237_46849# D_FlipFlop_0.Nand_Gate_0.Vout 0.04444f
C812 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.08671f
C813 FFCLR a_134897_24200# 0.04005f
C814 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.04109f
C815 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_65125_49858# 0.04444f
C816 a_96273_49858# VDD 0.0325f
C817 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.06445f
C818 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.06445f
C819 a_44403_15797# EN 0.045f
C820 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout CLK 0.20785f
C821 D_FlipFlop_5.Q' D_FlipFlop_5.Nand_Gate_1.Vout 0.11654f
C822 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_65869_15797# 0.05964f
C823 a_110029_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.04444f
C824 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.16429f
C825 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C EN 0.07601f
C826 D_FlipFlop_3.3-input-nand_2.C VDD 2.74431f
C827 a_106569_15797# VDD 0.01571f
C828 a_56801_15797# VDD 0.03119f
C829 a_128851_24200# VDD 0.01186f
C830 FFCLR a_134283_36157# 0.01145f
C831 a_45761_13083# VDD 0.02865f
C832 RingCounter_0.D_FlipFlop_10.Q' RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.11654f
C833 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout CLK 0.71041f
C834 a_128237_30478# Q3 0.06113f
C835 D_FlipFlop_1.3-input-nand_2.Vout a_132311_36157# 0.05964f
C836 a_134897_27764# VDD 0.01186f
C837 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout CLK 0.70923f
C838 a_130209_39721# VDD 0.02521f
C839 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.06594f
C840 a_75898_35820# CDAC8_0.switch_7.Z 0.26998f
C841 FFCLR a_132925_40571# 0.045f
C842 Nand_Gate_2.Vout VDD 1.37836f
C843 Nand_Gate_7.B RingCounter_0.D_FlipFlop_14.Inverter_0.Vout 0.29374f
C844 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C EN 0.07732f
C845 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_33363_13083# 0.01335f
C846 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout VDD 2.04843f
C847 a_128237_30478# VDD 0.02521f
C848 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.3-input-nand_2.Vout 0.16429f
C849 a_90535_13083# EN 0.0452f
C850 a_32749_13083# CLK 0.02953f
C851 D_FlipFlop_2.Q' a_128237_39721# 0.04443f
C852 a_52113_49858# VDD 0.0325f
C853 a_103765_47663# CLK 0.07396f
C854 FFCLR D_FlipFlop_2.Inverter_0.Vout 0.43598f
C855 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_112745_49858# 0.04995f
C856 a_112615_13083# VDD 0.01327f
C857 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_44403_15797# 0.01335f
C858 FFCLR D_FlipFlop_4.3-input-nand_0.Vout 0.12261f
C859 CDAC8_0.switch_9.Z CDAC8_0.switch_2.Z 0.28677f
C860 a_85233_52572# CLK 0.04619f
C861 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C EN 0.09031f
C862 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.08671f
C863 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout VDD 2.8604f
C864 Nand_Gate_0.A D_FlipFlop_2.Q' 0.06938f
C865 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_69199_49858# 0.04444f
C866 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout EN 0.60828f
C867 FFCLR a_134897_44135# 0.04005f
C868 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout a_89921_13083# 0.04443f
C869 a_75551_52572# a_76165_52572# 0.05935f
C870 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_1.Vout 0.08671f
C871 RingCounter_0.D_FlipFlop_6.Q' m3_125329_49141# 0.04886f
C872 And_Gate_0.Inverter_0.Vin EN 0.01805f
C873 a_99603_13083# CLK 0.03129f
C874 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C VDD 3.56545f
C875 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout EN 0.78747f
C876 Nand_Gate_7.B CDAC8_0.switch_2.Z 0.33658f
C877 a_84489_15797# EN 0.04443f
C878 D_FlipFlop_6.Nand_Gate_1.Vout VDD 1.46545f
C879 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_112615_15797# 0.01335f
C880 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout VDD 2.73618f
C881 a_119711_49858# VDD 0.06071f
C882 Nand_Gate_0.B CLK 0.40903f
C883 RingCounter_0.D_FlipFlop_17.Q' FFCLR 1.10693f
C884 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.04109f
C885 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout a_100347_52572# 0.04443f
C886 Nand_Gate_2.A Nand_Gate_2.B 0.07727f
C887 Nand_Gate_0.A Nand_Gate_5.B 0.06463f
C888 a_128851_44135# VDD 0.01186f
C889 Nand_Gate_5.B CDAC8_0.switch_7.Z 0.08438f
C890 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout EN 0.09127f
C891 a_89921_15797# CLK 0.04619f
C892 a_119711_52572# EN 0.045f
C893 a_46375_13083# EN 0.0452f
C894 a_121069_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.04444f
C895 And_Gate_1.Inverter_0.Vin EN 0.01805f
C896 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.25963f
C897 Nand_Gate_6.B Nand_Gate_6.Vout 2.38777f
C898 D_FlipFlop_3.3-input-nand_1.Vout a_132925_40571# 0.04543f
C899 a_123785_52572# Nand_Gate_5.B 0.01335f
C900 a_89307_52572# VDD 0.02521f
C901 a_132925_43285# VDD 0.01186f
C902 a_68455_13083# VDD 0.01327f
C903 CDAC8_0.switch_6.Z Q1 0.74949f
C904 Nand_Gate_2.B RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.08035f
C905 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout CLK 0.29759f
C906 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout VDD 1.56255f
C907 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 1.09975f
C908 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_99603_15797# 0.04995f
C909 a_134283_19786# VDD 0.02521f
C910 D_FlipFlop_0.Inverter_0.Vout a_134897_44135# 0.04995f
C911 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_7.Q' 0.06632f
C912 a_50755_15797# a_51369_15797# 0.05935f
C913 a_85847_15797# VDD 0.02906f
C914 FFCLR D_FlipFlop_5.Q' 0.03748f
C915 Nand_Gate_0.B Comparator_0.Vinm 0.03263f
C916 Nand_Gate_5.B RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.08377f
C917 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout CLK 0.03574f
C918 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout VDD 1.86552f
C919 a_130209_20636# VDD 0.02521f
C920 a_91279_52572# VDD 0.02521f
C921 FFCLR a_132925_17072# 0.045f
C922 Nand_Gate_4.A a_39715_15797# 0.06113f
C923 Nand_Gate_0.A CDAC8_0.switch_8.Z 2.01979f
C924 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C CLK 0.30901f
C925 CDAC8_0.switch_8.Z CDAC8_0.switch_7.Z 1.87529f
C926 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_2.C 0.15106f
C927 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Q' 1.16087f
C928 D_FlipFlop_2.Nand_Gate_1.Vout a_128237_37007# 0.04444f
C929 a_55443_13083# CLK 0.03129f
C930 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout VDD 2.88547f
C931 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_105955_13083# 0.04444f
C932 D_FlipFlop_2.3-input-nand_2.C a_132311_37007# 0.05964f
C933 RingCounter_0.D_FlipFlop_11.Q' a_95529_13083# 0.01335f
C934 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_98989_13083# 0.04444f
C935 D_FlipFlop_2.3-input-nand_0.Vout a_134897_39721# 0.01335f
C936 a_43045_52572# VDD 0.02865f
C937 a_58159_52572# Nand_Gate_3.B 0.06113f
C938 D_FlipFlop_4.Inverter_0.Vout a_134283_27764# 0.04443f
C939 a_75551_49858# VDD 0.06071f
C940 a_76909_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.04444f
C941 a_134897_46849# VDD 0.01186f
C942 a_128237_39721# a_128851_39721# 0.05935f
C943 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Nand_Gate_1.Vout 0.04109f
C944 And_Gate_5.Inverter_0.Vin a_59605_47663# 0.06113f
C945 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout VDD 2.07373f
C946 D_FlipFlop_0.3-input-nand_2.Vout VDD 2.77266f
C947 D_FlipFlop_6.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.06465f
C948 D_FlipFlop_4.3-input-nand_2.Vout a_132311_30478# 0.05964f
C949 D_FlipFlop_4.Q' a_128237_27764# 0.06113f
C950 Nand_Gate_1.B a_116995_15797# 0.06113f
C951 D_FlipFlop_0.Q' a_128237_44135# 0.06113f
C952 Nand_Gate_4.B a_50755_15797# 0.06113f
C953 Nand_Gate_2.A D_FlipFlop_3.Q' 0.06962f
C954 a_114805_16975# VDD 0.02521f
C955 CDAC8_0.switch_7.Z Q5 1.11487f
C956 a_128237_37007# Q6 0.04443f
C957 Nand_Gate_0.A a_128851_39721# 0.04625f
C958 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C CLK 0.30966f
C959 FFCLR EN 2.20871f
C960 a_45761_15797# VDD 0.03119f
C961 Nand_Gate_1.B Q3 0.25213f
C962 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.Nand_Gate_1.Vout 0.1541f
C963 a_123041_13083# CLK 0.04443f
C964 a_73579_52572# a_74193_52572# 0.05935f
C965 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 0.25579f
C966 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.06465f
C967 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.0857f
C968 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout a_118967_15797# 0.04443f
C969 a_59605_47663# VDD 0.02521f
C970 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.1182f
C971 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Nand_Gate_1.Vout 0.04109f
C972 a_130209_19786# D_FlipFlop_7.3-input-nand_2.Vout 0.04443f
C973 Nand_Gate_1.B VDD 7.74643f
C974 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout EN 0.08852f
C975 a_117739_52572# VDD 0.0564f
C976 RingCounter_0.D_FlipFlop_8.Q' RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.11654f
C977 a_32749_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.04444f
C978 D_FlipFlop_4.3-input-nand_1.Vout a_134283_27764# 0.05964f
C979 Nand_Gate_2.B Nand_Gate_2.Vout 2.18021f
C980 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_57545_52572# 0.04995f
C981 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_54829_15797# 0.04443f
C982 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout a_51499_49858# 0.04995f
C983 a_64511_52572# VDD 0.01186f
C984 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_3.Inverter_1.Vout 0.01422f
C985 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_117739_49858# 0.01335f
C986 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Nand_Gate_1.Vout 0.04109f
C987 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout EN 0.78734f
C988 And_Gate_5.Inverter_0.Vin CLK 0.4651f
C989 a_87205_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.05964f
C990 a_94915_13083# VDD 0.02521f
C991 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout Nand_Gate_5.B 0.11443f
C992 a_112745_49858# a_113359_49858# 0.05935f
C993 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout EN 0.13192f
C994 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110029_15797# 0.04443f
C995 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_74193_49858# 0.05964f
C996 D_FlipFlop_3.3-input-nand_0.Vout VDD 1.77946f
C997 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.30154f
C998 a_128237_17072# Q0 0.04443f
C999 CLK Q3 0.1175f
C1000 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C EN 0.76392f
C1001 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout a_74807_15797# 0.04443f
C1002 a_40459_52572# EN 0.04454f
C1003 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_0.Vout 0.06594f
C1004 Nand_Gate_0.A a_74193_52572# 0.04443f
C1005 a_68585_52572# Nand_Gate_0.A 0.01335f
C1006 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout a_74807_13083# 0.04995f
C1007 D_FlipFlop_2.3-input-nand_2.C VDD 2.74431f
C1008 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_43789_15797# 0.05964f
C1009 a_78881_13083# CLK 0.04619f
C1010 CDAC8_0.switch_5.Z CDAC8_0.switch_0.Z 0.09134f
C1011 Nand_Gate_4.B a_132925_19786# 0.04741f
C1012 VDD CLK 82.60049f
C1013 a_98245_49858# VDD 0.0301f
C1014 RingCounter_0.D_FlipFlop_14.Q' a_61795_13083# 0.06113f
C1015 RingCounter_0.D_FlipFlop_2.Q' RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.11654f
C1016 D_FlipFlop_3.Nand_Gate_0.Vout a_130209_43285# 0.05964f
C1017 Nand_Gate_7.B And_Gate_0.Inverter_0.Vin 0.04751f
C1018 Nand_Gate_5.A VDD 7.76004f
C1019 a_99603_15797# VDD 0.03339f
C1020 Nand_Gate_1.A a_100961_15797# 0.04443f
C1021 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.1541f
C1022 a_130209_36157# VDD 0.02521f
C1023 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout CLK 0.30735f
C1024 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_75551_52572# 0.04995f
C1025 And_Gate_5.Inverter_0.Vin Comparator_0.Vinm 0.02725f
C1026 a_128237_39721# D_FlipFlop_2.Nand_Gate_0.Vout 0.04444f
C1027 FFCLR a_132925_37007# 0.045f
C1028 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_52727_15797# 0.05964f
C1029 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout VDD 2.31704f
C1030 D_FlipFlop_6.3-input-nand_0.Vout a_134897_23350# 0.01335f
C1031 a_75898_42964# Comparator_0.Vinm 0.03709f
C1032 Nand_Gate_2.A a_128851_43285# 0.04627f
C1033 And_Gate_3.Inverter_0.Vin a_114805_16975# 0.05964f
C1034 a_75898_35820# Q7 0.4968f
C1035 Comparator_0.Vinm Q3 1.64934f
C1036 Nand_Gate_0.A D_FlipFlop_2.Nand_Gate_0.Vout 0.6452f
C1037 a_120325_52572# VDD 0.02521f
C1038 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout VDD 1.70415f
C1039 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout a_56187_49858# 0.04995f
C1040 a_85233_49858# CLK 0.04619f
C1041 a_50755_13083# VDD 0.02521f
C1042 a_132311_24200# VDD 0.02521f
C1043 a_54829_15797# VDD 0.03178f
C1044 FFCLR D_FlipFlop_1.Inverter_0.Vout 0.44538f
C1045 a_90665_49858# a_91279_49858# 0.05935f
C1046 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.06465f
C1047 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout a_30647_15797# 0.04443f
C1048 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout VDD 1.56255f
C1049 D_FlipFlop_7.3-input-nand_0.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.04107f
C1050 Nand_Gate_4.A VDD 4.19998f
C1051 a_112745_52572# EN 0.04443f
C1052 D_FlipFlop_5.3-input-nand_0.Vout a_134897_26914# 0.01335f
C1053 Comparator_0.Vinm VDD 16.9841f
C1054 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_107927_13083# 0.04443f
C1055 FFCLR a_134897_40571# 0.04005f
C1056 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.08671f
C1057 Nand_Gate_1.B And_Gate_3.Inverter_0.Vin 0.03063f
C1058 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_78267_49858# 0.05964f
C1059 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout VDD 1.76886f
C1060 Comparator_0.Vinm CDAC8_0.switch_1.Z 6.31039f
C1061 a_34721_13083# CLK 0.04619f
C1062 a_132311_46849# VDD 0.02521f
C1063 a_54085_49858# VDD 0.0301f
C1064 a_125845_47663# CLK 0.07396f
C1065 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.16429f
C1066 a_117609_13083# VDD 0.0563f
C1067 Nand_Gate_0.A a_69199_49858# 0.04741f
C1068 Nand_Gate_5.Vout CLK 2.38056f
C1069 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout EN 0.41175f
C1070 a_128851_40571# VDD 0.01186f
C1071 a_123785_52572# a_124399_52572# 0.05935f
C1072 Nand_Gate_5.A Nand_Gate_5.Vout 0.1063f
C1073 RingCounter_0.D_FlipFlop_12.Q' RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.11654f
C1074 FFCLR D_FlipFlop_1.3-input-nand_1.Vout 0.15444f
C1075 RingCounter_0.D_FlipFlop_9.Q' VDD 1.95446f
C1076 FFCLR CDAC8_0.switch_9.Z 2.17565f
C1077 RingCounter_0.D_FlipFlop_15.Q' VDD 1.95446f
C1078 a_76165_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.04443f
C1079 Nand_Gate_5.B Q7 0.06203f
C1080 Nand_Gate_1.B Nand_Gate_6.B 0.05373f
C1081 D_FlipFlop_1.3-input-nand_0.Vout a_132925_36157# 0.04995f
C1082 a_41073_49858# CLK 0.04443f
C1083 D_FlipFlop_1.3-input-nand_2.Vout EN 0.07759f
C1084 a_132925_39721# VDD 0.01186f
C1085 a_68585_49858# a_69199_49858# 0.05935f
C1086 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout Nand_Gate_0.A 0.12214f
C1087 CDAC8_0.switch_7.Z Q1 1.51854f
C1088 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_0.Vout 1.0203f
C1089 a_122427_49858# VDD 0.03726f
C1090 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout CLK 0.30735f
C1091 And_Gate_3.Inverter_0.Vin CLK 0.49672f
C1092 FFCLR Nand_Gate_7.B 0.93907f
C1093 D_FlipFlop_2.Inverter_0.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.0857f
C1094 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout FFCLR 0.12214f
C1095 a_132311_27764# a_132925_27764# 0.05935f
C1096 Nand_Gate_6.B a_94915_13083# 0.04443f
C1097 a_132311_44135# VDD 0.02521f
C1098 Nand_Gate_5.Vout Comparator_0.Vinm 0.02011f
C1099 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C EN 0.07667f
C1100 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout CLK 0.15609f
C1101 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_87949_13083# 0.05964f
C1102 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout VDD 2.04843f
C1103 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout EN 0.97489f
C1104 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_0.Vout 0.06594f
C1105 FFCLR D_FlipFlop_7.Q' 0.03748f
C1106 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_76909_13083# 0.04443f
C1107 D_FlipFlop_4.Q' D_FlipFlop_4.Nand_Gate_1.Vout 0.11654f
C1108 a_67841_15797# a_68455_15797# 0.05935f
C1109 D_FlipFlop_3.3-input-nand_1.Vout a_134897_40571# 0.01335f
C1110 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout CLK 0.03479f
C1111 a_65869_15797# a_66483_15797# 0.05935f
C1112 RingCounter_0.D_FlipFlop_6.Q' Nand_Gate_5.B 1.06171f
C1113 Nand_Gate_2.A D_FlipFlop_3.Nand_Gate_0.Vout 0.64587f
C1114 D_FlipFlop_0.Q' D_FlipFlop_0.Nand_Gate_1.Vout 0.11654f
C1115 Nand_Gate_7.B a_72835_13083# 0.04443f
C1116 a_134897_43285# VDD 0.01186f
C1117 a_108671_49858# CLK 0.03129f
C1118 a_73449_13083# VDD 0.0563f
C1119 CDAC8_0.switch_8.Z Q7 0.29972f
C1120 D_FlipFlop_2.Nand_Gate_1.Vout Q6 0.06503f
C1121 Nand_Gate_1.A Nand_Gate_1.Vout 0.0689f
C1122 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.1541f
C1123 a_107313_52572# CLK 0.04619f
C1124 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_101575_15797# 0.01335f
C1125 D_FlipFlop_7.Inverter_0.Vout VDD 1.3737f
C1126 Nand_Gate_3.B And_Gate_5.Inverter_0.Vin 0.02391f
C1127 And_Gate_2.Inverter_0.Vin Q0 0.05118f
C1128 Nand_Gate_6.B CLK 0.52286f
C1129 Nand_Gate_6.A EN 0.42008f
C1130 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.Inverter_1.Vout 0.25963f
C1131 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout EN 0.60828f
C1132 a_63153_52572# VDD 0.02521f
C1133 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout EN 0.06649f
C1134 a_132925_20636# VDD 0.01186f
C1135 FFCLR a_51499_52572# 0.04995f
C1136 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.0846f
C1137 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_2.C 1.09975f
C1138 a_122427_52572# RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.05964f
C1139 a_46505_49858# a_47119_49858# 0.05935f
C1140 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Inverter_1.Vout 0.25963f
C1141 D_FlipFlop_2.Nand_Gate_1.Vout a_130209_37007# 0.05964f
C1142 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_107927_13083# 0.05964f
C1143 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.3-input-nand_2.Vout 0.06445f
C1144 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout EN 0.78747f
C1145 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_100961_13083# 0.05964f
C1146 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C EN 0.07664f
C1147 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.06465f
C1148 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_95529_13083# 0.04995f
C1149 a_41073_52572# VDD 0.02865f
C1150 a_78267_49858# VDD 0.04111f
C1151 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_88563_13083# 0.04543f
C1152 a_110029_13083# a_110643_13083# 0.05935f
C1153 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_83875_13083# 0.04444f
C1154 And_Gate_2.Inverter_0.Vin EN 0.01805f
C1155 Nand_Gate_2.B CLK 0.40867f
C1156 FFCLR D_FlipFlop_5.3-input-nand_2.Vout 0.06105f
C1157 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_76909_13083# 0.04444f
C1158 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.Inverter_1.Vout 0.25963f
C1159 RingCounter_0.D_FlipFlop_12.Q' CLK 0.09276f
C1160 Nand_Gate_7.A EN 0.42008f
C1161 FFCLR D_FlipFlop_0.Q' 0.03748f
C1162 VDD Q4 3.72275f
C1163 a_134283_23350# a_134897_23350# 0.05935f
C1164 Nand_Gate_3.B VDD 4.34213f
C1165 Nand_Gate_2.A Nand_Gate_5.B 0.06495f
C1166 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.04107f
C1167 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.1182f
C1168 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_124399_52572# 0.04444f
C1169 a_128851_17072# VDD 0.01186f
C1170 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout a_63153_49858# 0.04443f
C1171 Comparator_0.Vinm Nand_Gate_6.B 1.96281f
C1172 D_FlipFlop_7.Inverter_0.Vout a_134283_17072# 0.04443f
C1173 a_117609_15797# EN 0.04443f
C1174 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout a_57415_13083# 0.04995f
C1175 Nand_Gate_7.A a_62409_15797# 0.01335f
C1176 a_64511_49858# CLK 0.03129f
C1177 a_111387_52572# VDD 0.02521f
C1178 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.25963f
C1179 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout VDD 1.70415f
C1180 a_29289_13083# VDD 0.0563f
C1181 Nand_Gate_1.Vout Q0 0.05051f
C1182 a_74193_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.05964f
C1183 D_FlipFlop_7.Q' a_128237_17072# 0.06113f
C1184 FFCLR D_FlipFlop_7.Inverter_1.Vout 0.56927f
C1185 a_134283_26914# a_134897_26914# 0.05935f
C1186 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.06445f
C1187 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.Nand_Gate_1.Vout 0.30154f
C1188 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.06465f
C1189 a_123041_15797# CLK 0.04443f
C1190 D_FlipFlop_2.3-input-nand_0.Vout VDD 1.77946f
C1191 a_81685_47663# VDD 0.02521f
C1192 a_68585_52572# a_69199_52572# 0.05935f
C1193 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout a_65125_49858# 0.04443f
C1194 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.04109f
C1195 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_40329_13083# 0.04995f
C1196 D_FlipFlop_4.3-input-nand_2.Vout VDD 2.77266f
C1197 a_57545_52572# EN 0.04443f
C1198 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_33363_13083# 0.04543f
C1199 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_28675_13083# 0.04444f
C1200 Nand_Gate_2.B Comparator_0.Vinm 0.03245f
C1201 RingCounter_0.D_FlipFlop_14.Q' RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.06632f
C1202 D_FlipFlop_5.3-input-nand_1.Vout D_FlipFlop_6.3-input-nand_0.Vout 0.01418f
C1203 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout VDD 1.86552f
C1204 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C CLK 0.30901f
C1205 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_52727_13083# 0.04443f
C1206 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_1.Q' 0.06632f
C1207 a_113359_52572# VDD 0.02521f
C1208 D_FlipFlop_1.3-input-nand_2.C VDD 2.74431f
C1209 Nand_Gate_1.Vout EN 0.10633f
C1210 a_134283_46849# VDD 0.02521f
C1211 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C VDD 3.61245f
C1212 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_119711_49858# 0.04543f
C1213 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.08671f
C1214 D_FlipFlop_4.3-input-nand_0.Vout a_132925_30478# 0.04995f
C1215 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.1541f
C1216 a_87949_13083# a_88563_13083# 0.05935f
C1217 FFCLR D_FlipFlop_4.Inverter_0.Vout 0.43823f
C1218 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout EN 1.03094f
C1219 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout CLK 0.69703f
C1220 a_96887_13083# VDD 0.02578f
C1221 a_118967_15797# VDD 0.02906f
C1222 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout EN 0.06649f
C1223 FFCLR D_FlipFlop_6.3-input-nand_2.C 0.76213f
C1224 a_29289_15797# EN 0.04443f
C1225 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_76165_49858# 0.04444f
C1226 And_Gate_6.Inverter_0.Vin EN 0.0623f
C1227 a_134283_33443# a_134897_33443# 0.05935f
C1228 And_Gate_1.Inverter_0.Vin a_48565_16975# 0.05964f
C1229 Nand_Gate_4.A a_37897_16975# 0.0476f
C1230 Nand_Gate_2.A Q5 1.05014f
C1231 a_75898_39392# Comparator_0.Vinm 0.0374f
C1232 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.06465f
C1233 D_FlipFlop_6.Q' Q2 0.01194f
C1234 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout EN 0.08653f
C1235 a_34721_15797# CLK 0.04619f
C1236 D_FlipFlop_4.Inverter_1.Vout a_130209_27764# 0.04995f
C1237 RingCounter_0.D_FlipFlop_2.Q' Nand_Gate_0.A 1.10693f
C1238 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_42431_49858# 0.01335f
C1239 D_FlipFlop_1.Q' a_128237_36157# 0.04443f
C1240 a_73449_15797# VDD 0.01571f
C1241 D_FlipFlop_7.3-input-nand_2.Vout a_132925_19786# 0.01335f
C1242 FFCLR RingCounter_0.D_FlipFlop_1.Inverter_0.Vout 0.29368f
C1243 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout 0.0846f
C1244 a_101705_49858# VDD 0.06015f
C1245 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.1541f
C1246 a_97631_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.01335f
C1247 Nand_Gate_1.A RingCounter_0.D_FlipFlop_11.Inverter_0.Vout 0.29374f
C1248 a_101575_15797# VDD 0.06072f
C1249 Nand_Gate_0.B a_80239_49858# 0.04741f
C1250 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.C 0.06594f
C1251 FFCLR a_134897_37007# 0.04055f
C1252 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout EN 0.08852f
C1253 D_FlipFlop_6.3-input-nand_2.C a_132311_20636# 0.05964f
C1254 a_83875_15797# VDD 0.02906f
C1255 RingCounter_0.D_FlipFlop_2.Q' a_68585_49858# 0.01335f
C1256 CDAC8_0.switch_5.Z CLK 0.21166f
C1257 FFCLR D_FlipFlop_4.3-input-nand_1.Vout 0.95389f
C1258 a_30647_15797# VDD 0.02521f
C1259 a_67227_52572# RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.05964f
C1260 D_FlipFlop_1.Q' Q7 1.06172f
C1261 Nand_Gate_4.A a_34721_15797# 0.04443f
C1262 a_84619_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.01335f
C1263 a_122427_52572# RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.04443f
C1264 a_86591_52572# VDD 0.01186f
C1265 a_65869_13083# a_66483_13083# 0.05935f
C1266 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.06465f
C1267 a_87205_49858# CLK 0.03129f
C1268 a_134283_24200# VDD 0.02521f
C1269 a_52727_13083# VDD 0.02578f
C1270 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.Inverter_1.Vout 0.25579f
C1271 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout CLK 0.03574f
C1272 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_123785_49858# 0.04995f
C1273 D_FlipFlop_5.3-input-nand_2.C a_132311_24200# 0.05964f
C1274 a_128851_37007# VDD 0.01186f
C1275 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110643_13083# 0.01335f
C1276 a_52113_52572# CLK 0.04619f
C1277 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_69199_52572# 0.04444f
C1278 FFCLR CDAC8_0.switch_6.Z 6.54715f
C1279 D_FlipFlop_7.3-input-nand_2.C a_132311_19786# 0.04443f
C1280 Nand_Gate_1.B a_112001_15797# 0.04443f
C1281 Nand_Gate_4.B a_45761_15797# 0.04443f
C1282 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 1.09975f
C1283 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout EN 0.60828f
C1284 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_80239_49858# 0.04444f
C1285 D_FlipFlop_2.3-input-nand_1.Vout a_132925_37007# 0.04543f
C1286 Nand_Gate_0.B a_85233_52572# 0.04443f
C1287 RingCounter_0.D_FlipFlop_1.Q' a_58159_49858# 0.06113f
C1288 D_FlipFlop_3.Q' a_128851_40571# 0.01335f
C1289 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_110643_13083# 0.04543f
C1290 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout EN 0.78668f
C1291 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.25579f
C1292 a_75898_21528# Q1 0.49857f
C1293 CDAC8_0.switch_5.Z Comparator_0.Vinm 52.8265f
C1294 a_132925_36157# VDD 0.01186f
C1295 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C VDD 3.56545f
C1296 a_57545_49858# VDD 0.06015f
C1297 Nand_Gate_1.B Nand_Gate_4.B 0.05965f
C1298 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.08671f
C1299 a_121069_13083# VDD 0.02578f
C1300 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_117609_15797# 0.04995f
C1301 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.Nand_Gate_1.Vout 0.04109f
C1302 a_88563_15797# EN 0.045f
C1303 D_FlipFlop_3.Inverter_0.Vout a_134897_40571# 0.04995f
C1304 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 0.25579f
C1305 a_124399_52572# RingCounter_0.D_FlipFlop_6.Q' 0.04443f
C1306 a_132311_40571# VDD 0.02521f
C1307 a_128237_26914# Q2 0.06113f
C1308 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout EN 0.09127f
C1309 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout a_84619_49858# 0.04995f
C1310 Nand_Gate_7.B Nand_Gate_7.A 0.07512f
C1311 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout VDD 1.62198f
C1312 a_43789_13083# a_44403_13083# 0.05935f
C1313 D_FlipFlop_1.3-input-nand_0.Vout a_134897_36157# 0.01335f
C1314 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout EN 0.24889f
C1315 VDD Q2 3.59902f
C1316 a_43045_49858# CLK 0.03129f
C1317 a_96887_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.04443f
C1318 Nand_Gate_4.A a_39715_13083# 0.04443f
C1319 a_134897_39721# VDD 0.01186f
C1320 a_128237_36157# a_128851_36157# 0.05935f
C1321 a_56187_52572# VDD 0.02521f
C1322 EN Q6 0.2481f
C1323 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_43789_13083# 0.04444f
C1324 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout EN 0.61894f
C1325 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_0.Vout 0.0846f
C1326 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout a_100961_13083# 0.04443f
C1327 a_132311_30478# VDD 0.02521f
C1328 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_87205_52572# 0.04444f
C1329 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout VDD 2.31704f
C1330 a_112001_15797# CLK 0.04619f
C1331 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout VDD 1.60037f
C1332 a_124399_49858# VDD 0.02521f
C1333 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout EN 0.80245f
C1334 a_128237_20636# Q1 0.04443f
C1335 a_134283_44135# VDD 0.02521f
C1336 Nand_Gate_4.B CLK 0.53366f
C1337 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout a_74193_49858# 0.04443f
C1338 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout CLK 0.68588f
C1339 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_73449_15797# 0.04995f
C1340 a_58159_52572# VDD 0.02521f
C1341 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C CLK 0.30901f
C1342 FFCLR D_FlipFlop_4.Nand_Gate_1.Vout 0.60828f
C1343 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout a_107927_13083# 0.04995f
C1344 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_67841_15797# 0.05964f
C1345 Nand_Gate_0.B RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.08035f
C1346 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout VDD 2.88547f
C1347 a_128851_36157# Q7 0.01335f
C1348 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_121683_13083# 0.04543f
C1349 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_116995_13083# 0.04444f
C1350 a_76909_13083# VDD 0.02578f
C1351 a_47119_52572# VDD 0.02521f
C1352 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout a_46505_52572# 0.04995f
C1353 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout EN 0.41175f
C1354 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.16429f
C1355 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout a_76165_49858# 0.04443f
C1356 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.06594f
C1357 a_50755_15797# RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.04444f
C1358 D_FlipFlop_3.Q' Q4 0.01194f
C1359 a_134897_20636# VDD 0.01186f
C1360 Nand_Gate_4.B a_50755_13083# 0.04443f
C1361 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout VDD 2.29866f
C1362 FFCLR RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.08377f
C1363 a_132311_19786# a_132925_19786# 0.05935f
C1364 Nand_Gate_6.A a_78881_15797# 0.04443f
C1365 a_67227_52572# RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.04443f
C1366 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_64511_49858# 0.01335f
C1367 Nand_Gate_4.B Nand_Gate_4.A 0.07538f
C1368 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout a_89307_49858# 0.04995f
C1369 Comparator_0.Vinm Nand_Gate_4.B 1.16732f
C1370 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_90535_13083# 0.01335f
C1371 D_FlipFlop_1.3-input-nand_0.Vout VDD 1.77126f
C1372 a_80239_49858# VDD 0.02906f
C1373 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_85847_13083# 0.05964f
C1374 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_78881_13083# 0.05964f
C1375 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_29289_15797# 0.04995f
C1376 D_FlipFlop_5.Inverter_1.Vout VDD 1.73058f
C1377 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_73449_13083# 0.04995f
C1378 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121683_15797# 0.01335f
C1379 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout a_112615_13083# 0.04995f
C1380 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_66483_13083# 0.04543f
C1381 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout VDD 2.73332f
C1382 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_61795_13083# 0.04444f
C1383 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_54829_13083# 0.04444f
C1384 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.0857f
C1385 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout VDD 2.73618f
C1386 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout a_41073_49858# 0.04443f
C1387 RingCounter_0.D_FlipFlop_9.Q' a_106569_13083# 0.01335f
C1388 Nand_Gate_5.B Nand_Gate_1.B 0.06366f
C1389 FFCLR D_FlipFlop_6.3-input-nand_0.Vout 0.1261f
C1390 a_132311_17072# VDD 0.02521f
C1391 D_FlipFlop_0.Nand_Gate_0.Vout a_130209_46849# 0.05964f
C1392 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout EN 0.08852f
C1393 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0846f
C1394 Nand_Gate_6.Vout a_82057_16975# 0.05964f
C1395 a_130209_43285# D_FlipFlop_3.3-input-nand_2.Vout 0.04443f
C1396 FFCLR D_FlipFlop_3.Inverter_1.Vout 0.56927f
C1397 a_128237_46849# Q4 0.06113f
C1398 RingCounter_0.D_FlipFlop_12.Q' a_83875_15797# 0.04443f
C1399 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_54085_49858# 0.05964f
C1400 D_FlipFlop_7.Inverter_0.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.0857f
C1401 a_32749_13083# VDD 0.02578f
C1402 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.06594f
C1403 D_FlipFlop_2.Nand_Gate_0.Vout a_130209_39721# 0.05964f
C1404 CDAC8_0.switch_0.Z Q1 0.0732f
C1405 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.16429f
C1406 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout CLK 0.06496f
C1407 a_103765_47663# VDD 0.02521f
C1408 a_69199_52572# RingCounter_0.D_FlipFlop_2.Q' 0.04443f
C1409 a_128237_36157# D_FlipFlop_1.Nand_Gate_0.Vout 0.04444f
C1410 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Q' 1.05791f
C1411 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Q' 1.05791f
C1412 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_35335_13083# 0.01335f
C1413 D_FlipFlop_6.Inverter_1.Vout a_130209_23350# 0.04443f
C1414 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_85233_49858# 0.05964f
C1415 a_75898_18814# Q0 0.49857f
C1416 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_30647_13083# 0.05964f
C1417 a_75898_35820# Comparator_0.Vinm 0.04018f
C1418 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_2.Vout 0.88855f
C1419 a_85233_52572# VDD 0.02521f
C1420 And_Gate_0.Inverter_0.Vin a_70645_16975# 0.05964f
C1421 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout CLK 0.23464f
C1422 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_5.3-input-nand_2.C 0.01194f
C1423 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_5.3-input-nand_2.Vout 0.01194f
C1424 a_97631_52572# a_98245_52572# 0.05935f
C1425 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_55443_13083# 0.01335f
C1426 RingCounter_0.D_FlipFlop_3.Q' a_79625_49858# 0.01335f
C1427 RingCounter_0.D_FlipFlop_17.Q' EN 0.03751f
C1428 Nand_Gate_1.A EN 0.42008f
C1429 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout a_77523_15797# 0.01335f
C1430 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout 0.06445f
C1431 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout CLK 0.03574f
C1432 a_75898_21528# CDAC8_0.switch_2.Z 0.2969f
C1433 D_FlipFlop_4.3-input-nand_0.Vout a_134283_30478# 0.05964f
C1434 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout EN 0.78747f
C1435 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.08671f
C1436 a_40329_15797# EN 0.04443f
C1437 a_99603_13083# VDD 0.05686f
C1438 Nand_Gate_5.A RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.08024f
C1439 D_FlipFlop_5.Inverter_1.Vout a_130209_26914# 0.04443f
C1440 D_FlipFlop_1.Nand_Gate_0.Vout Q7 0.11443f
C1441 Nand_Gate_6.B Q2 0.34858f
C1442 Nand_Gate_5.B CLK 0.28816f
C1443 a_117739_49858# a_118353_49858# 0.05935f
C1444 Nand_Gate_1.B RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.0839f
C1445 Nand_Gate_4.B RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0839f
C1446 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout a_122427_52572# 0.04443f
C1447 Nand_Gate_0.B VDD 4.34213f
C1448 Nand_Gate_5.A Nand_Gate_5.B 0.13465f
C1449 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.06594f
C1450 Nand_Gate_7.A a_61795_13083# 0.04443f
C1451 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_54829_15797# 0.05964f
C1452 a_89921_15797# VDD 0.03119f
C1453 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout CLK 0.15609f
C1454 a_75898_25104# CDAC8_0.switch_0.Z 0.29588f
C1455 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.16429f
C1456 a_84619_49858# EN 0.07058f
C1457 a_39715_15797# VDD 0.02906f
C1458 CDAC8_0.switch_9.Z Q6 0.24469f
C1459 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110029_13083# 0.04443f
C1460 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_45147_49858# 0.04443f
C1461 RingCounter_0.D_FlipFlop_11.Q' RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.11654f
C1462 a_132311_19786# D_FlipFlop_7.3-input-nand_0.Vout 0.04444f
C1463 RingCounter_0.D_FlipFlop_10.Q' CLK 0.09298f
C1464 Nand_Gate_4.B D_FlipFlop_7.Inverter_0.Vout 0.25902f
C1465 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_40329_15797# 0.04995f
C1466 a_106699_49858# VDD 0.01712f
C1467 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 1.09975f
C1468 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_33363_15797# 0.01335f
C1469 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout VDD 2.04843f
C1470 D_FlipFlop_7.Inverter_1.Vout a_130209_17072# 0.04995f
C1471 FFCLR Nand_Gate_0.A 0.92619f
C1472 a_79625_52572# EN 0.04443f
C1473 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout a_85847_13083# 0.04995f
C1474 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.06445f
C1475 FFCLR CDAC8_0.switch_7.Z 11.2108f
C1476 Nand_Gate_5.B Comparator_0.Vinm 0.11402f
C1477 a_41687_15797# VDD 0.02906f
C1478 CDAC8_0.switch_8.Z CLK 0.35798f
C1479 EN Q0 0.24699f
C1480 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout EN 0.06649f
C1481 And_Gate_4.Inverter_0.Vin CLK 0.50205f
C1482 RingCounter_0.D_FlipFlop_13.Q' a_72835_13083# 0.06113f
C1483 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout VDD 2.16362f
C1484 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout a_95659_49858# 0.04995f
C1485 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_89307_49858# 0.05964f
C1486 Nand_Gate_4.A RingCounter_0.D_FlipFlop_16.Inverter_0.Vout 0.29374f
C1487 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout a_41687_15797# 0.04443f
C1488 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout CLK 0.29759f
C1489 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C VDD 3.61245f
C1490 Nand_Gate_7.B D_FlipFlop_6.Inverter_1.Vout 0.12286f
C1491 a_80239_52572# Nand_Gate_0.B 0.06113f
C1492 D_FlipFlop_6.Q' VDD 1.89809f
C1493 a_55443_13083# VDD 0.05686f
C1494 a_95659_49858# a_96273_49858# 0.05935f
C1495 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout EN 1.03094f
C1496 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.16429f
C1497 CLK Q5 0.1175f
C1498 RingCounter_0.D_FlipFlop_16.Q a_40459_52572# 0.04995f
C1499 a_132311_37007# VDD 0.02521f
C1500 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_2.Vout 0.8898f
C1501 a_40459_49858# EN 0.02716f
C1502 Nand_Gate_1.B RingCounter_0.D_FlipFlop_9.Inverter_0.Vout 0.29374f
C1503 Nand_Gate_4.B RingCounter_0.D_FlipFlop_8.Inverter_0.Vout 0.29374f
C1504 Nand_Gate_6.B D_FlipFlop_5.Inverter_1.Vout 0.12143f
C1505 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.1541f
C1506 D_FlipFlop_2.3-input-nand_1.Vout a_134897_37007# 0.01335f
C1507 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_112615_13083# 0.01335f
C1508 CDAC8_0.switch_8.Z Comparator_0.Vinm 0.10659p
C1509 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.0857f
C1510 D_FlipFlop_6.Nand_Gate_1.Vout Q1 0.06503f
C1511 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C VDD 3.56545f
C1512 a_134897_36157# VDD 0.01186f
C1513 a_62409_15797# EN 0.04443f
C1514 a_43045_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.05964f
C1515 And_Gate_4.Inverter_0.Vin Comparator_0.Vinm 0.02739f
C1516 a_95659_52572# a_96273_52572# 0.05935f
C1517 a_62539_49858# VDD 0.01712f
C1518 a_128237_20636# a_128851_20636# 0.05935f
C1519 RingCounter_0.D_FlipFlop_10.Q' a_117609_13083# 0.01335f
C1520 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.3-input-nand_1.Vout 0.08671f
C1521 a_123041_13083# VDD 0.02865f
C1522 RingCounter_0.D_FlipFlop_16.Q a_28675_13083# 0.04443f
C1523 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.04107f
C1524 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout EN 0.61894f
C1525 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.04109f
C1526 a_67841_15797# CLK 0.04619f
C1527 a_134283_40571# VDD 0.02521f
C1528 D_FlipFlop_7.Nand_Gate_1.Vout a_128851_17072# 0.04995f
C1529 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.06465f
C1530 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.3-input-nand_2.Vout 0.06445f
C1531 Comparator_0.Vinm Q5 0.78239f
C1532 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout a_79625_52572# 0.04995f
C1533 D_FlipFlop_1.3-input-nand_2.C a_132311_33443# 0.05964f
C1534 a_107313_49858# EN 0.01149f
C1535 a_128237_24200# a_128851_24200# 0.05935f
C1536 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.3-input-nand_2.Vout 0.06445f
C1537 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.04107f
C1538 a_108671_52572# VDD 0.01186f
C1539 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_75551_49858# 0.01335f
C1540 a_73579_49858# a_74193_49858# 0.05935f
C1541 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout CLK 0.29759f
C1542 a_110029_13083# CLK 0.03129f
C1543 a_94915_15797# a_95529_15797# 0.05935f
C1544 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout a_100347_49858# 0.04995f
C1545 a_109285_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.05964f
C1546 D_FlipFlop_1.Nand_Gate_0.Vout D_FlipFlop_1.Inverter_1.Vout 0.25963f
C1547 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout EN 0.78734f
C1548 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout CLK 0.70923f
C1549 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_45761_13083# 0.05964f
C1550 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout EN 0.06649f
C1551 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout CLK 0.15614f
C1552 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_88563_15797# 0.04995f
C1553 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout a_67227_52572# 0.04443f
C1554 a_116995_15797# VDD 0.0299f
C1555 And_Gate_5.Inverter_0.Vin VDD 1.43186f
C1556 Nand_Gate_0.A a_71017_47663# 0.04705f
C1557 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.Nand_Gate_1.Vout 0.30154f
C1558 CDAC8_0.switch_0.Z CDAC8_0.switch_2.Z 0.1201f
C1559 a_63767_15797# VDD 0.02906f
C1560 CDAC8_0.switch_5.Z Q2 0.06367f
C1561 a_134283_27764# a_134897_27764# 0.05935f
C1562 a_74193_52572# CLK 0.04619f
C1563 a_75898_42964# VDD 1.30491f
C1564 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout EN 0.60828f
C1565 Nand_Gate_2.A a_96273_52572# 0.04443f
C1566 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_7.Inverter_1.Vout 0.01422f
C1567 VDD Q3 3.60342f
C1568 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.04109f
C1569 a_90665_52572# Nand_Gate_2.A 0.01335f
C1570 a_128237_26914# VDD 0.02521f
C1571 a_65869_15797# RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.04444f
C1572 Nand_Gate_6.B a_89921_15797# 0.04443f
C1573 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_123655_13083# 0.01335f
C1574 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.16429f
C1575 a_78881_13083# VDD 0.02865f
C1576 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_118967_13083# 0.05964f
C1577 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_98989_13083# 0.05964f
C1578 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.C 1.09975f
C1579 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout EN 0.78747f
C1580 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_2.C 1.09975f
C1581 a_128851_23350# VDD 0.01186f
C1582 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Q' 0.06632f
C1583 D_FlipFlop_6.Q' D_FlipFlop_6.Nand_Gate_0.Vout 0.06632f
C1584 Nand_Gate_5.A a_113359_49858# 0.04741f
C1585 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout a_97631_52572# 0.04995f
C1586 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_87949_13083# 0.04443f
C1587 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.06465f
C1588 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C CLK 0.30966f
C1589 Nand_Gate_5.B Q4 0.06203f
C1590 D_FlipFlop_1.Inverter_0.Vout EN 0.39551f
C1591 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout VDD 2.31704f
C1592 CDAC8_0.switch_1.Z VDD 1.11454f
C1593 a_63153_49858# EN 0.01149f
C1594 FFCLR D_FlipFlop_2.Inverter_1.Vout 0.57257f
C1595 a_28675_15797# VDD 0.02521f
C1596 Nand_Gate_6.A RingCounter_0.D_FlipFlop_13.Inverter_0.Vout 0.29374f
C1597 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_67227_49858# 0.04443f
C1598 a_123655_13083# EN 0.0452f
C1599 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.3-input-nand_2.C 0.25579f
C1600 D_FlipFlop_3.Inverter_1.Vout a_130209_40571# 0.04995f
C1601 a_65869_13083# CLK 0.03129f
C1602 a_51499_49858# a_52113_49858# 0.05935f
C1603 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.C 0.25579f
C1604 a_121683_15797# EN 0.045f
C1605 D_FlipFlop_5.Q' D_FlipFlop_5.Nand_Gate_0.Vout 0.06632f
C1606 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout CLK 0.23404f
C1607 a_78267_52572# VDD 0.02521f
C1608 a_112001_13083# a_112615_13083# 0.05935f
C1609 a_85233_49858# VDD 0.0325f
C1610 Nand_Gate_1.B Q1 0.05915f
C1611 FFCLR D_FlipFlop_7.3-input-nand_2.C 0.76213f
C1612 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_98989_15797# 0.04443f
C1613 CDAC8_0.switch_9.Z Q0 0.14628f
C1614 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_68455_13083# 0.01335f
C1615 D_FlipFlop_4.3-input-nand_2.C D_FlipFlop_4.Nand_Gate_1.Vout 0.1541f
C1616 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_63767_13083# 0.05964f
C1617 FFCLR a_132925_27764# 0.045f
C1618 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_56801_13083# 0.05964f
C1619 Nand_Gate_5.A D_FlipFlop_0.Inverter_1.Vout 0.15693f
C1620 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_51369_13083# 0.04995f
C1621 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.3-input-nand_2.C 0.25579f
C1622 a_134283_17072# VDD 0.02521f
C1623 RingCounter_0.D_FlipFlop_4.Q' a_91279_49858# 0.06113f
C1624 D_FlipFlop_4.Q' a_128237_30478# 0.04443f
C1625 CDAC8_0.switch_8.Z Q4 0.55536f
C1626 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C CLK 0.30901f
C1627 a_80239_52572# VDD 0.02521f
C1628 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout EN 0.61894f
C1629 a_105955_15797# a_106569_15797# 0.05935f
C1630 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout EN 0.78734f
C1631 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.06465f
C1632 Nand_Gate_7.A RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout 0.1182f
C1633 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_51499_49858# 0.01335f
C1634 a_34721_13083# VDD 0.02865f
C1635 D_FlipFlop_1.3-input-nand_1.Vout EN 0.97444f
C1636 a_130209_26914# VDD 0.02521f
C1637 CDAC8_0.switch_9.Z EN 5.40382f
C1638 FFCLR a_47119_49858# 0.04741f
C1639 a_125845_47663# VDD 0.02521f
C1640 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout EN 0.41175f
C1641 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout CLK 0.03574f
C1642 Nand_Gate_5.Vout VDD 1.47723f
C1643 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout a_68455_13083# 0.04995f
C1644 a_33363_15797# EN 0.04775f
C1645 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_87205_49858# 0.04444f
C1646 D_FlipFlop_7.Q' Q0 1.09842f
C1647 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout a_63767_15797# 0.04443f
C1648 a_79495_13083# EN 0.0452f
C1649 a_98245_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.04443f
C1650 CDAC8_0.switch_6.Z Q6 0.84618f
C1651 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.1541f
C1652 FFCLR a_134897_26914# 0.08419f
C1653 CLK Q1 0.1175f
C1654 Nand_Gate_7.B EN 1.37686f
C1655 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout CLK 0.03479f
C1656 D_FlipFlop_4.3-input-nand_2.C a_130209_27764# 0.04443f
C1657 And_Gate_4.Inverter_0.Vin a_81685_47663# 0.05964f
C1658 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.04109f
C1659 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout a_96887_15797# 0.05964f
C1660 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_2.A 0.12214f
C1661 a_89921_13083# a_90535_13083# 0.05935f
C1662 a_41073_49858# VDD 0.02521f
C1663 a_77523_15797# VDD 0.03339f
C1664 a_101575_13083# VDD 0.01327f
C1665 Nand_Gate_1.A a_105955_13083# 0.04443f
C1666 D_FlipFlop_7.3-input-nand_1.Vout a_132311_17072# 0.04444f
C1667 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C CLK 0.30966f
C1668 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_63767_13083# 0.04443f
C1669 D_FlipFlop_3.3-input-nand_2.Vout a_132925_43285# 0.01335f
C1670 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout EN 0.64426f
C1671 FFCLR a_134897_33443# 0.0607f
C1672 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout VDD 2.31704f
C1673 RingCounter_0.D_FlipFlop_16.Q' a_29289_13083# 0.01335f
C1674 And_Gate_3.Inverter_0.Vin VDD 1.53086f
C1675 D_FlipFlop_6.Nand_Gate_0.Vout a_128851_23350# 0.04995f
C1676 D_FlipFlop_6.Nand_Gate_0.Vout VDD 1.48313f
C1677 D_FlipFlop_2.Q' a_128851_37007# 0.01335f
C1678 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout CLK 0.71041f
C1679 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout EN 0.08852f
C1680 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout VDD 1.70415f
C1681 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout a_107313_49858# 0.04443f
C1682 a_128237_44135# a_128851_44135# 0.05935f
C1683 a_87949_15797# VDD 0.03178f
C1684 FFCLR Q7 0.77041f
C1685 a_88563_13083# CLK 0.03129f
C1686 a_134897_30478# VDD 0.01186f
C1687 a_53471_52572# VDD 0.01186f
C1688 Nand_Gate_7.B a_72835_15797# 0.06113f
C1689 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout VDD 1.56255f
C1690 Comparator_0.Vinm Q1 1.64919f
C1691 D_FlipFlop_2.Inverter_0.Vout a_134897_37007# 0.04995f
C1692 D_FlipFlop_5.Nand_Gate_0.Vout a_128851_26914# 0.04995f
C1693 a_108671_49858# VDD 0.06071f
C1694 a_45147_52572# VDD 0.02865f
C1695 a_128851_33443# VDD 0.01186f
C1696 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout a_109285_49858# 0.04443f
C1697 Nand_Gate_5.Vout a_125845_47663# 0.04443f
C1698 D_FlipFlop_4.3-input-nand_2.Vout a_132311_27764# 0.04443f
C1699 D_FlipFlop_6.Nand_Gate_1.Vout a_128851_20636# 0.04995f
C1700 a_107313_52572# VDD 0.02521f
C1701 D_FlipFlop_4.3-input-nand_0.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.04107f
C1702 Nand_Gate_6.B VDD 7.84453f
C1703 a_35335_13083# EN 0.0452f
C1704 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.0846f
C1705 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout a_91279_49858# 0.04444f
C1706 a_128237_30478# a_128851_30478# 0.05935f
C1707 a_67841_13083# a_68455_13083# 0.05935f
C1708 RingCounter_0.D_FlipFlop_16.Q a_29289_15797# 0.0156f
C1709 D_FlipFlop_3.3-input-nand_2.C a_132311_43285# 0.04443f
C1710 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout EN 0.13192f
C1711 a_57415_13083# VDD 0.01327f
C1712 a_105955_15797# RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.04444f
C1713 D_FlipFlop_1.Inverter_0.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.0857f
C1714 D_FlipFlop_5.Nand_Gate_1.Vout a_128851_24200# 0.04995f
C1715 D_FlipFlop_1.Nand_Gate_1.Vout EN 0.6398f
C1716 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout CLK 0.71041f
C1717 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.08377f
C1718 a_134283_37007# VDD 0.02521f
C1719 Nand_Gate_2.B VDD 4.34213f
C1720 RingCounter_0.D_FlipFlop_12.Q' VDD 1.95446f
C1721 Comparator_0.Vinm a_75898_25104# 0.03583f
C1722 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_1.Vout 0.07775f
C1723 a_42431_49858# EN 0.04775f
C1724 a_128851_19786# Q0 0.01335f
C1725 D_FlipFlop_6.3-input-nand_2.Vout VDD 2.77266f
C1726 RingCounter_0.D_FlipFlop_8.Q' RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.06632f
C1727 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C a_87205_49858# 0.05964f
C1728 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout a_107927_15797# 0.05964f
C1729 a_44403_13083# CLK 0.03129f
C1730 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.25963f
C1731 a_110643_15797# EN 0.045f
C1732 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout CLK 0.30735f
C1733 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.08671f
C1734 Nand_Gate_5.B Q2 0.06203f
C1735 a_96273_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout 0.05964f
C1736 a_64511_49858# VDD 0.06071f
C1737 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout CLK 0.71041f
C1738 m3_125329_49141# VDD 0.10297f
C1739 a_90665_52572# a_91279_52572# 0.05935f
C1740 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout EN 0.97489f
C1741 a_123041_15797# VDD 0.02734f
C1742 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout CLK 0.15609f
C1743 Nand_Gate_5.B a_124399_49858# 0.04484f
C1744 FFCLR Nand_Gate_2.A 0.93793f
C1745 a_101705_52572# EN 0.04443f
C1746 FFCLR D_FlipFlop_6.Inverter_0.Vout 0.43823f
C1747 a_75898_39392# VDD 1.30474f
C1748 D_FlipFlop_4.Q' Nand_Gate_1.B 0.03509f
C1749 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_3.3-input-nand_0.Vout 0.0846f
C1750 a_37897_16975# VDD 0.02521f
C1751 a_107927_15797# RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.04443f
C1752 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Q' 0.06632f
C1753 RingCounter_0.D_FlipFlop_7.Q' a_112745_49858# 0.01335f
C1754 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout CLK 0.03479f
C1755 a_56801_15797# a_57415_15797# 0.05935f
C1756 D_FlipFlop_1.Nand_Gate_1.Vout a_128237_33443# 0.04444f
C1757 a_54829_15797# a_55443_15797# 0.05935f
C1758 a_42431_52572# a_43045_52572# 0.05935f
C1759 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout CLK 0.03574f
C1760 a_45761_13083# a_46375_13083# 0.05935f
C1761 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout EN 0.58846f
C1762 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout CLK 0.30716f
C1763 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C VDD 3.61245f
C1764 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C a_78267_49858# 0.04443f
C1765 a_112001_13083# CLK 0.04619f
C1766 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.Inverter_1.Vout 0.25963f
C1767 a_128237_19786# VDD 0.02521f
C1768 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_2.3-input-nand_2.Vout 0.01194f
C1769 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout EN 1.03094f
C1770 D_FlipFlop_3.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.C 0.01194f
C1771 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout a_90535_15797# 0.01335f
C1772 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout VDD 1.84669f
C1773 a_130209_46849# D_FlipFlop_0.3-input-nand_2.Vout 0.04443f
C1774 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout EN 0.41172f
C1775 CDAC8_0.switch_9.Z Nand_Gate_7.B 1.10291f
C1776 D_FlipFlop_3.Q' VDD 1.89796f
C1777 RingCounter_0.D_FlipFlop_2.Q' CLK 0.09276f
C1778 a_130209_39721# D_FlipFlop_2.3-input-nand_2.Vout 0.04443f
C1779 FFCLR D_FlipFlop_1.Inverter_1.Vout 0.16183f
C1780 Nand_Gate_3.B RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.08035f
C1781 FFCLR D_FlipFlop_7.3-input-nand_0.Vout 0.1263f
C1782 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C EN 0.07664f
C1783 RingCounter_0.D_FlipFlop_5.Q' a_102319_49858# 0.06113f
C1784 RingCounter_0.D_FlipFlop_4.Q' Nand_Gate_2.A 1.10693f
C1785 a_34721_15797# VDD 0.03119f
C1786 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_41687_13083# 0.04443f
C1787 D_FlipFlop_1.Nand_Gate_0.Vout a_130209_36157# 0.05964f
C1788 CDAC8_0.switch_2.Z CLK 0.08199f
C1789 FFCLR D_FlipFlop_6.3-input-nand_1.Vout 0.95389f
C1790 Nand_Gate_6.B RingCounter_0.D_FlipFlop_12.Inverter_0.Vout 0.29374f
C1791 a_118353_49858# CLK 0.04619f
C1792 a_83875_13083# VDD 0.02521f
C1793 a_132311_43285# a_132925_43285# 0.05935f
C1794 a_128237_30478# D_FlipFlop_4.Nand_Gate_0.Vout 0.04444f
C1795 RingCounter_0.D_FlipFlop_14.Q' CLK 0.09276f
C1796 CDAC8_0.switch_6.Z Q0 0.28955f
C1797 a_119711_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 0.01335f
C1798 CDAC8_0.switch_5.Z Q3 0.5952f
C1799 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout 0.04107f
C1800 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.C 0.06594f
C1801 D_FlipFlop_5.3-input-nand_2.C VDD 2.74431f
C1802 a_128237_46849# VDD 0.02521f
C1803 Nand_Gate_2.A D_FlipFlop_3.3-input-nand_1.Vout 0.07758f
C1804 a_89307_52572# RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout 0.05964f
C1805 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_1.Vout 0.06465f
C1806 D_FlipFlop_7.3-input-nand_0.Vout a_134897_19786# 0.01335f
C1807 CDAC8_0.switch_5.Z VDD 1.3927f
C1808 a_106699_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout 0.01335f
C1809 Nand_Gate_1.B D_FlipFlop_4.Inverter_1.Vout 0.12092f
C1810 Nand_Gate_1.B a_104137_16975# 0.04443f
C1811 D_FlipFlop_7.Nand_Gate_0.Vout Q0 0.1147f
C1812 a_67841_13083# CLK 0.04619f
C1813 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.3-input-nand_2.Vout 0.16429f
C1814 FFCLR D_FlipFlop_3.3-input-nand_2.C 0.76213f
C1815 CDAC8_0.switch_6.Z EN 11.3849f
C1816 FFCLR a_128851_24200# 0.04443f
C1817 a_87205_49858# VDD 0.0301f
C1818 a_128237_39721# Q6 0.06113f
C1819 Comparator_0.Vinm CDAC8_0.switch_2.Z 14.3922f
C1820 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.0857f
C1821 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.04109f
C1822 D_FlipFlop_6.3-input-nand_1.Vout a_132311_20636# 0.04444f
C1823 a_54085_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.05964f
C1824 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout 0.0846f
C1825 RingCounter_0.D_FlipFlop_9.Q' RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.11654f
C1826 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout VDD 2.07373f
C1827 RingCounter_0.D_FlipFlop_15.Q' RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.06632f
C1828 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout CLK 0.03574f
C1829 FFCLR a_134897_27764# 0.04005f
C1830 a_96273_52572# CLK 0.04619f
C1831 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout a_91279_52572# 0.04444f
C1832 Nand_Gate_0.A Q6 1.38518f
C1833 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout EN 0.60828f
C1834 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_96273_49858# 0.05964f
C1835 a_52113_52572# VDD 0.02521f
C1836 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.3-input-nand_2.Vout 0.16429f
C1837 Nand_Gate_2.B a_107313_52572# 0.04443f
C1838 CDAC8_0.switch_7.Z Q6 1.11431f
C1839 a_128851_30478# Nand_Gate_1.B 0.04732f
C1840 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.04107f
C1841 D_FlipFlop_7.3-input-nand_1.Vout VDD 1.78032f
C1842 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.Inverter_1.Vout 0.25579f
C1843 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout a_118353_49858# 0.04443f
C1844 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_9.Inverter_1.Vout 0.25963f
C1845 a_74193_49858# CLK 0.04619f
C1846 a_39715_13083# VDD 0.02521f
C1847 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout a_53471_49858# 0.04543f
C1848 D_FlipFlop_5.3-input-nand_1.Vout a_132311_24200# 0.04444f
C1849 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout a_46505_49858# 0.04995f
C1850 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout EN 0.78747f
C1851 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_41073_49858# 0.05964f
C1852 D_FlipFlop_0.Nand_Gate_1.Vout a_128851_44135# 0.04995f
C1853 a_128851_27764# VDD 0.01186f
C1854 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.06503f
C1855 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout a_120325_49858# 0.04443f
C1856 a_132311_23350# VDD 0.02521f
C1857 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout 0.06445f
C1858 a_128851_43285# VDD 0.01186f
C1859 D_FlipFlop_0.3-input-nand_1.Vout D_FlipFlop_3.3-input-nand_0.Vout 0.01418f
C1860 a_51369_15797# VDD 0.01571f
C1861 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_108671_49858# 0.01335f
C1862 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout 0.0846f
C1863 D_FlipFlop_4.3-input-nand_2.C a_132925_27764# 0.01335f
C1864 Nand_Gate_2.A RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.08024f
C1865 a_43045_49858# VDD 0.02568f
C1866 a_100347_52572# VDD 0.02521f
C1867 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.1541f
C1868 a_79495_15797# VDD 0.06072f
C1869 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C CLK 0.30966f
C1870 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout a_109285_52572# 0.04444f
C1871 a_106569_13083# VDD 0.0563f
C1872 D_FlipFlop_7.3-input-nand_1.Vout a_134283_17072# 0.05964f
C1873 FFCLR D_FlipFlop_6.Nand_Gate_1.Vout 0.60828f
C1874 a_119711_49858# a_120325_49858# 0.05935f
C1875 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.3-input-nand_1.Vout 0.08671f
C1876 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C a_66483_13083# 0.01335f
C1877 a_132311_43285# D_FlipFlop_3.3-input-nand_0.Vout 0.04444f
C1878 a_112001_15797# VDD 0.03119f
C1879 a_61795_15797# VDD 0.02906f
C1880 RingCounter_0.D_FlipFlop_9.Q' a_105955_15797# 0.04443f
C1881 FFCLR a_128851_44135# 0.04443f
C1882 D_FlipFlop_7.3-input-nand_2.C a_130209_17072# 0.04443f
C1883 a_132925_26914# VDD 0.01186f
C1884 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_1.Vout 0.0775f
C1885 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C CLK 0.30901f
C1886 a_102319_52572# VDD 0.02521f
C1887 Nand_Gate_4.B VDD 8.59026f
C1888 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout VDD 2.73618f
C1889 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.06465f
C1890 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C a_98245_49858# 0.05964f
C1891 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_100347_49858# 0.05964f
C1892 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C VDD 3.61242f
C1893 Nand_Gate_0.B And_Gate_4.Inverter_0.Vin 0.02391f
C1894 Nand_Gate_0.A D_FlipFlop_2.Inverter_0.Vout 0.26421f
C1895 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_2.C 0.11436f
C1896 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.0857f
C1897 a_64511_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 0.01335f
C1898 a_111387_49858# VDD 0.04111f
C1899 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout EN 1.03094f
C1900 a_132311_33443# VDD 0.02521f
C1901 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout 0.04107f
C1902 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout 0.25963f
C1903 CDAC8_0.switch_1.Z Nand_Gate_4.B 1.47073f
C1904 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout a_123041_13083# 0.04443f
C1905 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout 0.16429f
C1906 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout 0.0846f
C1907 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout a_57545_49858# 0.04995f
C1908 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.C 1.09975f
C1909 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C CLK 0.19377f
C1910 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.3-input-nand_2.Vout 0.06445f
C1911 a_89307_52572# RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.04443f
C1912 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout CLK 0.03479f
C1913 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_2.C 0.1129f
C1914 RingCounter_0.D_FlipFlop_6.Q' a_123785_49858# 0.01335f
C1915 D_FlipFlop_4.Nand_Gate_0.Vout Nand_Gate_1.B 0.67556f
C1916 Comparator_0.Vinm Vin 0.02469f
C1917 And_Gate_2.Inverter_0.Vin a_92725_16975# 0.05964f
C1918 a_97631_49858# CLK 0.03129f
C1919 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout a_96887_13083# 0.04995f
C1920 D_FlipFlop_7.Nand_Gate_1.Vout VDD 1.46545f
C1921 a_62409_13083# VDD 0.0563f
C1922 And_Gate_0.Inverter_0.Vin CLK 0.63116f
C1923 a_66483_15797# EN 0.045f
C1924 a_97631_49858# a_98245_49858# 0.05935f
C1925 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_2.Nand_Gate_1.Vout 0.30154f
C1926 D_FlipFlop_7.3-input-nand_2.Vout a_132311_17072# 0.04443f
C1927 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout 0.04109f
C1928 FFCLR a_134897_46849# 0.04454f
C1929 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout CLK 0.23464f
C1930 FFCLR D_FlipFlop_0.3-input-nand_2.Vout 0.06105f
C1931 a_75898_35820# VDD 1.30478f
C1932 RingCounter_0.D_FlipFlop_12.Q' a_83875_13083# 0.06113f
C1933 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout EN 0.09127f
C1934 Nand_Gate_1.B a_116995_13083# 0.04443f
C1935 a_134283_19786# a_134897_19786# 0.05935f
C1936 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout EN 0.08852f
C1937 a_128237_44135# Q4 0.04443f
C1938 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.Inverter_1.Vout 0.25579f
C1939 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_2.C 1.09975f
C1940 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout EN 0.24889f
C1941 CDAC8_0.switch_9.Z CDAC8_0.switch_6.Z 10.0827f
C1942 a_85847_15797# RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.04443f
C1943 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout CLK 0.30735f
C1944 D_FlipFlop_3.Nand_Gate_0.Vout VDD 1.48313f
C1945 And_Gate_1.Inverter_0.Vin CLK 0.59514f
C1946 a_75551_52572# VDD 0.01186f
C1947 D_FlipFlop_5.3-input-nand_2.Vout D_FlipFlop_6.3-input-nand_2.C 0.01194f
C1948 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_6.3-input-nand_2.Vout 0.01194f
C1949 Nand_Gate_6.A Nand_Gate_6.Vout 0.0689f
C1950 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_2.C 1.09975f
C1951 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout EN 0.61894f
C1952 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout 0.04107f
C1953 a_67227_49858# VDD 0.04111f
C1954 a_91279_52572# RingCounter_0.D_FlipFlop_4.Q' 0.04443f
C1955 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_44403_15797# 0.04995f
C1956 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout VDD 1.70248f
C1957 CDAC8_0.switch_6.Z Nand_Gate_7.B 3.32256f
C1958 D_FlipFlop_2.Q' VDD 1.89795f
C1959 a_121069_15797# VDD 0.03178f
C1960 D_FlipFlop_3.3-input-nand_2.C D_FlipFlop_3.Nand_Gate_1.Vout 0.1541f
C1961 FFCLR Nand_Gate_1.B 0.91491f
C1962 a_59977_16975# VDD 0.02521f
C1963 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout a_62409_15797# 0.04995f
C1964 a_119711_52572# a_120325_52572# 0.05935f
C1965 D_FlipFlop_2.Inverter_1.Vout a_130209_37007# 0.04995f
C1966 Nand_Gate_6.Vout And_Gate_2.Inverter_0.Vin 0.24808f
C1967 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout a_56801_15797# 0.05964f
C1968 D_FlipFlop_1.Nand_Gate_1.Vout a_130209_33443# 0.05964f
C1969 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout VDD 2.88547f
C1970 Nand_Gate_5.B Q3 0.06203f
C1971 a_43045_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.C 0.04443f
C1972 a_132925_33443# EN 0.05084f
C1973 D_FlipFlop_5.3-input-nand_0.Vout VDD 1.77946f
C1974 a_53471_49858# CLK 0.03129f
C1975 D_FlipFlop_0.3-input-nand_1.Vout a_132311_44135# 0.04444f
C1976 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout 0.0846f
C1977 CDAC8_0.switch_6.Z a_75898_28676# 0.01232f
C1978 RingCounter_0.D_FlipFlop_16.Q EN 0.259f
C1979 a_75551_49858# a_76165_49858# 0.05935f
C1980 a_94915_15797# RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.04444f
C1981 a_75898_25104# Q2 0.49874f
C1982 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout VDD 2.16362f
C1983 Nand_Gate_2.A D_FlipFlop_3.Inverter_0.Vout 0.26407f
C1984 CDAC8_0.switch_7.Z Q0 0.57741f
C1985 RingCounter_0.D_FlipFlop_10.Q' a_116995_15797# 0.04443f
C1986 Nand_Gate_7.B a_132925_23350# 0.0478f
C1987 Nand_Gate_5.B VDD 4.32141f
C1988 FFCLR D_FlipFlop_3.3-input-nand_0.Vout 0.1263f
C1989 a_139696_27690# Comparator_0.Vinm 0.34941f
C1990 D_FlipFlop_7.Q' D_FlipFlop_7.Nand_Gate_0.Vout 0.06632f
C1991 D_FlipFlop_6.Inverter_0.Vout a_134283_20636# 0.04443f
C1992 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_44403_13083# 0.01335f
C1993 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout VDD 1.70415f
C1994 Nand_Gate_0.A EN 0.73819f
C1995 FFCLR D_FlipFlop_2.3-input-nand_2.C 0.76542f
C1996 a_32749_15797# VDD 0.02793f
C1997 CDAC8_0.switch_7.Z EN 21.4209f
C1998 CDAC8_0.switch_8.Z a_75898_42964# 0.01003f
C1999 Nand_Gate_6.B a_132925_26914# 0.04784f
C2000 D_FlipFlop_6.3-input-nand_2.Vout a_132311_23350# 0.05964f
C2001 a_120325_49858# CLK 0.02953f
C2002 D_FlipFlop_3.3-input-nand_2.C a_130209_40571# 0.04443f
C2003 a_85847_13083# VDD 0.02578f
C2004 RingCounter_0.D_FlipFlop_10.Q' VDD 1.96961f
C2005 D_FlipFlop_3.3-input-nand_0.Vout a_134283_43285# 0.05964f
C2006 FFCLR CLK 0.38481f
C2007 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout 0.08671f
C2008 Nand_Gate_6.B Nand_Gate_4.B 0.062f
C2009 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout 1.09975f
C2010 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout 0.04107f
C2011 D_FlipFlop_4.Nand_Gate_1.Vout D_FlipFlop_5.Nand_Gate_0.Vout 0.01681f
C2012 FFCLR Nand_Gate_5.A 0.61625f
C2013 a_123785_52572# EN 0.04443f
C2014 Nand_Gate_3.B a_48937_47663# 0.04443f
C2015 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.Inverter_1.Vout 0.06445f
C2016 Nand_Gate_7.A a_56801_15797# 0.04443f
C2017 D_FlipFlop_5.Inverter_0.Vout a_134283_24200# 0.04443f
C2018 CDAC8_0.switch_8.Z VDD 1.45501f
C2019 a_128237_24200# Q2 0.04443f
C2020 RingCounter_0.D_FlipFlop_13.Q' a_72835_15797# 0.04443f
C2021 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_2.C 0.14342f
C2022 a_45761_15797# a_46375_15797# 0.05935f
C2023 a_75898_42964# Q5 0.4968f
C2024 D_FlipFlop_5.3-input-nand_2.Vout a_132311_26914# 0.05964f
C2025 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout EN 0.06649f
C2026 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_4.3-input-nand_2.Vout 0.06445f
C2027 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout CLK 0.30716f
C2028 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.06594f
C2029 And_Gate_4.Inverter_0.Vin VDD 1.43186f
C2030 D_FlipFlop_0.3-input-nand_2.Vout a_132925_46849# 0.01335f
C2031 a_53471_49858# a_54085_49858# 0.05935f
C2032 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_119711_49858# 0.01335f
C2033 a_102319_52572# Nand_Gate_2.B 0.06113f
C2034 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout EN 0.97427f
C2035 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_98989_13083# 0.04443f
C2036 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout VDD 2.04843f
C2037 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_62539_49858# 0.01335f
C2038 a_90665_49858# VDD 0.06015f
C2039 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.04109f
C2040 a_116995_13083# a_117609_13083# 0.05935f
C2041 D_FlipFlop_2.3-input-nand_2.Vout a_132925_39721# 0.01335f
C2042 Nand_Gate_2.A a_93097_47663# 0.04705f
C2043 D_FlipFlop_6.3-input-nand_1.Vout a_134283_20636# 0.05964f
C2044 D_FlipFlop_4.Inverter_0.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.0857f
C2045 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout CLK 0.23464f
C2046 FFCLR Comparator_0.Vinm 7.20175f
C2047 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout EN 0.41172f
C2048 VDD Q5 3.80025f
C2049 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout CLK 0.70923f
C2050 Nand_Gate_5.B Nand_Gate_5.Vout 2.12832f
C2051 RingCounter_0.D_FlipFlop_4.Q' CLK 0.09276f
C2052 a_128851_39721# VDD 0.01186f
C2053 a_128237_40571# a_128851_40571# 0.05935f
C2054 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout a_98245_49858# 0.04444f
C2055 RingCounter_0.D_FlipFlop_16.Q' VDD 1.93566f
C2056 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout a_34721_13083# 0.04443f
C2057 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout a_66483_15797# 0.01335f
C2058 D_FlipFlop_3.3-input-nand_2.Vout a_132311_40571# 0.04443f
C2059 D_FlipFlop_3.3-input-nand_0.Vout D_FlipFlop_3.3-input-nand_1.Vout 0.04107f
C2060 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.06465f
C2061 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout 0.06445f
C2062 D_FlipFlop_7.Nand_Gate_0.Vout D_FlipFlop_7.Inverter_1.Vout 0.25963f
C2063 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C CLK 0.30862f
C2064 a_117739_52572# a_118353_52572# 0.05935f
C2065 a_76165_49858# CLK 0.03129f
C2066 a_41687_13083# VDD 0.02578f
C2067 D_FlipFlop_5.3-input-nand_1.Vout a_134283_24200# 0.05964f
C2068 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout a_43045_49858# 0.04444f
C2069 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout a_98989_15797# 0.05964f
C2070 Nand_Gate_5.A D_FlipFlop_0.Inverter_0.Vout 0.26399f
C2071 RingCounter_0.D_FlipFlop_16.Q' a_28675_15797# 0.04443f
C2072 Nand_Gate_4.B a_37897_16975# 0.04443f
C2073 a_132311_27764# VDD 0.02521f
C2074 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout a_41687_13083# 0.04995f
C2075 D_FlipFlop_0.3-input-nand_2.C a_132311_46849# 0.04443f
C2076 FFCLR a_128851_40571# 0.04443f
C2077 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_0.Vout 1.02969f
C2078 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.1541f
C2079 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout EN 1.01751f
C2080 a_67841_15797# VDD 0.03119f
C2081 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout 0.16429f
C2082 a_64511_52572# a_65125_52572# 0.05935f
C2083 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout a_101705_52572# 0.04995f
C2084 D_FlipFlop_7.Nand_Gate_0.Vout a_128851_19786# 0.04995f
C2085 D_FlipFlop_2.3-input-nand_2.C a_132311_39721# 0.04443f
C2086 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C a_111387_49858# 0.04443f
C2087 D_FlipFlop_4.Nand_Gate_1.Vout a_128237_27764# 0.04444f
C2088 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout a_79495_13083# 0.04995f
C2089 RingCounter_0.D_FlipFlop_17.Q' a_47119_49858# 0.06113f
C2090 Nand_Gate_2.Vout And_Gate_6.Inverter_0.Vin 0.10129f
C2091 a_46505_49858# VDD 0.01571f
C2092 a_94915_13083# a_95529_13083# 0.05935f
C2093 a_71017_47663# CLK 0.02953f
C2094 a_51499_52572# RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout 0.01335f
C2095 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout VDD 2.04843f
C2096 a_110029_13083# VDD 0.02578f
C2097 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout a_89307_52572# 0.04443f
C2098 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_0.Vout 1.03021f
C2099 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout VDD 2.73618f
C2100 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout VDD 1.70415f
C2101 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.1541f
C2102 a_118353_52572# CLK 0.04619f
C2103 D_FlipFlop_1.3-input-nand_1.Vout a_132925_33443# 0.04543f
C2104 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout EN 0.60828f
C2105 D_FlipFlop_7.3-input-nand_2.C a_132925_17072# 0.01335f
C2106 a_74193_52572# VDD 0.02521f
C2107 Nand_Gate_5.A a_118353_52572# 0.04443f
C2108 a_134283_26914# VDD 0.02521f
C2109 Nand_Gate_5.B Nand_Gate_6.B 0.06371f
C2110 a_112745_52572# Nand_Gate_5.A 0.01335f
C2111 a_68585_52572# VDD 0.01186f
C2112 D_FlipFlop_6.Q' Q1 1.06476f
C2113 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout a_46375_13083# 0.04995f
C2114 D_FlipFlop_7.3-input-nand_2.Vout VDD 2.77266f
C2115 Nand_Gate_5.A a_132925_46849# 0.04685f
C2116 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.06503f
C2117 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_74807_13083# 0.04443f
C2118 D_FlipFlop_0.3-input-nand_2.C a_132311_44135# 0.05964f
C2119 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout a_102319_49858# 0.04444f
C2120 D_FlipFlop_0.3-input-nand_0.Vout a_134897_46849# 0.01335f
C2121 a_43789_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.04444f
C2122 RingCounter_0.D_FlipFlop_8.Q' a_40329_13083# 0.01335f
C2123 D_FlipFlop_0.Nand_Gate_1.Vout Q4 0.06503f
C2124 D_FlipFlop_0.3-input-nand_2.Vout D_FlipFlop_0.3-input-nand_0.Vout 0.0846f
C2125 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout EN 0.78747f
C2126 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout 1.09975f
C2127 a_110029_15797# a_110643_15797# 0.05935f
C2128 FFCLR a_134897_43285# 0.08419f
C2129 a_113359_49858# VDD 0.02906f
C2130 a_134283_33443# VDD 0.02521f
C2131 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout a_119711_52572# 0.04995f
C2132 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_2.3-input-nand_0.Vout 0.0846f
C2133 FFCLR D_FlipFlop_7.Inverter_0.Vout 0.39255f
C2134 Nand_Gate_2.Vout a_93097_47663# 0.05964f
C2135 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_121683_15797# 0.04995f
C2136 Nand_Gate_0.A CDAC8_0.switch_9.Z 0.22762f
C2137 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C VDD 3.56545f
C2138 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout CLK 0.155f
C2139 CDAC8_0.switch_9.Z CDAC8_0.switch_7.Z 3.75058f
C2140 a_95529_15797# EN 0.04443f
C2141 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout CLK 0.03574f
C2142 FFCLR a_132925_20636# 0.045f
C2143 D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.48313f
C2144 Nand_Gate_7.B RingCounter_0.D_FlipFlop_13.Q' 1.05791f
C2145 D_FlipFlop_4.Nand_Gate_0.Vout D_FlipFlop_4.3-input-nand_2.Vout 0.16429f
C2146 a_134283_43285# a_134897_43285# 0.05935f
C2147 a_72835_13083# a_73449_13083# 0.05935f
C2148 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.06503f
C2149 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.06465f
C2150 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_1.3-input-nand_2.Vout 0.01194f
C2151 D_FlipFlop_2.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.C 0.01194f
C2152 RingCounter_0.D_FlipFlop_16.Q RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout 0.14519f
C2153 a_122427_52572# VDD 0.02521f
C2154 a_65869_13083# VDD 0.02578f
C2155 a_100961_15797# CLK 0.04619f
C2156 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout VDD 3.68398f
C2157 D_FlipFlop_3.Q' D_FlipFlop_3.Nand_Gate_0.Vout 0.06632f
C2158 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121069_13083# 0.05964f
C2159 Nand_Gate_5.B m3_125329_49141# 0.18891f
C2160 D_FlipFlop_1.Q' VDD 1.89794f
C2161 CDAC8_0.switch_7.Z Nand_Gate_7.B 7.65138f
C2162 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout CLK 0.03574f
C2163 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout a_54085_52572# 0.04444f
C2164 D_FlipFlop_0.Inverter_1.Vout VDD 1.73058f
C2165 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_1.Vout 0.07411f
C2166 FFCLR Nand_Gate_3.B 0.07771f
C2167 a_130209_36157# D_FlipFlop_1.3-input-nand_2.Vout 0.04443f
C2168 Nand_Gate_5.B a_123041_15797# 0.04443f
C2169 a_132311_46849# a_132925_46849# 0.05935f
C2170 FFCLR a_128851_17072# 0.04443f
C2171 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout 0.1541f
C2172 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C CLK 0.19377f
C2173 a_124399_52572# VDD 0.02521f
C2174 a_62539_52572# a_63153_52572# 0.05935f
C2175 a_83875_15797# a_84489_15797# 0.05935f
C2176 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout CLK 0.29759f
C2177 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C VDD 3.61242f
C2178 a_132311_39721# a_132925_39721# 0.05935f
C2179 a_96887_15797# VDD 0.02906f
C2180 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_77523_15797# 0.04995f
C2181 a_69199_49858# VDD 0.02906f
C2182 a_132311_20636# a_132925_20636# 0.05935f
C2183 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout EN 1.03094f
C2184 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.C 0.25579f
C2185 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout a_43789_13083# 0.04443f
C2186 FFCLR D_FlipFlop_2.3-input-nand_0.Vout 0.1263f
C2187 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout a_46375_15797# 0.01335f
C2188 Nand_Gate_4.B a_51369_15797# 0.01335f
C2189 Nand_Gate_1.B a_117609_15797# 0.01335f
C2190 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_0.Vout 0.06594f
C2191 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout VDD 2.16362f
C2192 FFCLR D_FlipFlop_4.3-input-nand_2.Vout 0.06105f
C2193 Nand_Gate_1.Vout a_114805_16975# 0.04995f
C2194 a_82057_16975# VDD 0.02521f
C2195 D_FlipFlop_7.Inverter_1.Vout a_130209_19786# 0.04443f
C2196 Nand_Gate_6.A CLK 0.38549f
C2197 a_120325_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.04443f
C2198 Nand_Gate_3.B a_62539_52572# 0.04995f
C2199 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout CLK 0.03479f
C2200 a_117739_49858# EN 0.07058f
C2201 a_132311_24200# a_132925_24200# 0.05935f
C2202 FFCLR D_FlipFlop_1.3-input-nand_2.C 0.14795f
C2203 a_50755_13083# a_51369_13083# 0.05935f
C2204 a_54829_15797# RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.04444f
C2205 a_134897_33443# EN 0.04286f
C2206 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout a_43045_52572# 0.04444f
C2207 a_128851_23350# Q1 0.01335f
C2208 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout CLK 0.71041f
C2209 VDD Q1 3.61051f
C2210 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout Nand_Gate_5.A 0.12214f
C2211 a_40459_52572# a_41073_52572# 0.05935f
C2212 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout VDD 1.48392f
C2213 D_FlipFlop_0.3-input-nand_1.Vout a_134283_44135# 0.05964f
C2214 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.04109f
C2215 D_FlipFlop_5.Nand_Gate_1.Vout Q2 0.06503f
C2216 Nand_Gate_5.A D_FlipFlop_0.3-input-nand_0.Vout 1.01439f
C2217 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout a_45147_49858# 0.04995f
C2218 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_0.Vout 0.06594f
C2219 EN Q7 0.26571f
C2220 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout CLK 0.23464f
C2221 a_134897_23350# VDD 0.01186f
C2222 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C CLK 0.30966f
C2223 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout EN 0.13192f
C2224 Nand_Gate_1.B Nand_Gate_1.Vout 2.35665f
C2225 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C VDD 3.56545f
C2226 And_Gate_2.Inverter_0.Vin CLK 0.63116f
C2227 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_33363_15797# 0.04995f
C2228 Nand_Gate_7.A CLK 0.38549f
C2229 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout EN 0.0879f
C2230 D_FlipFlop_4.Inverter_1.Vout D_FlipFlop_5.Inverter_1.Vout 0.01422f
C2231 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout VDD 2.73332f
C2232 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.C 0.25579f
C2233 a_97631_52572# VDD 0.01186f
C2234 a_128237_17072# a_128851_17072# 0.05935f
C2235 D_FlipFlop_3.Nand_Gate_1.Vout a_128851_40571# 0.04995f
C2236 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_2.C 0.11237f
C2237 D_FlipFlop_3.3-input-nand_2.C a_132925_40571# 0.01335f
C2238 a_88563_13083# VDD 0.05686f
C2239 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_87949_15797# 0.04443f
C2240 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout a_64511_52572# 0.04995f
C2241 D_FlipFlop_3.Nand_Gate_0.Vout a_128851_43285# 0.04995f
C2242 a_75898_25104# VDD 1.30969f
C2243 Nand_Gate_7.A RingCounter_0.D_FlipFlop_15.Inverter_0.Vout 0.29374f
C2244 a_128851_36157# VDD 0.01186f
C2245 RingCounter_0.D_FlipFlop_15.Q' a_51369_13083# 0.01335f
C2246 a_132311_19786# VDD 0.02521f
C2247 D_FlipFlop_3.3-input-nand_1.Vout D_FlipFlop_2.3-input-nand_0.Vout 0.01418f
C2248 a_128237_33443# Q7 0.04443f
C2249 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout EN 0.78734f
C2250 a_73579_49858# EN 0.07058f
C2251 a_28675_13083# a_29289_13083# 0.05935f
C2252 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_107313_49858# 0.05964f
C2253 D_FlipFlop_3.Q' Q5 1.06173f
C2254 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.Nand_Gate_1.Vout 0.30154f
C2255 a_132311_46849# D_FlipFlop_0.3-input-nand_0.Vout 0.04444f
C2256 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C a_122427_49858# 0.04443f
C2257 Nand_Gate_1.Vout CLK 2.75415f
C2258 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.0857f
C2259 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout a_64511_49858# 0.04543f
C2260 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.3-input-nand_1.Vout 0.08671f
C2261 a_95659_49858# VDD 0.01712f
C2262 CDAC8_0.switch_8.Z CDAC8_0.switch_5.Z 0.09134f
C2263 a_132311_39721# D_FlipFlop_2.3-input-nand_0.Vout 0.04444f
C2264 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout a_45147_52572# 0.04443f
C2265 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.C 0.25579f
C2266 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout a_52727_15797# 0.04443f
C2267 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout CLK 0.29644f
C2268 D_FlipFlop_1.Q' a_128851_33443# 0.01335f
C2269 FFCLR a_128851_37007# 0.04443f
C2270 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout VDD 2.73332f
C2271 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout CLK 0.68706f
C2272 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.Nand_Gate_1.Vout 0.30154f
C2273 And_Gate_6.Inverter_0.Vin CLK 0.50205f
C2274 D_FlipFlop_6.3-input-nand_0.Vout a_132925_23350# 0.04995f
C2275 a_130209_30478# D_FlipFlop_4.3-input-nand_2.Vout 0.04443f
C2276 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout 0.04107f
C2277 Nand_Gate_2.A EN 0.61039f
C2278 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout a_85847_15797# 0.05964f
C2279 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.25963f
C2280 Nand_Gate_1.A a_106569_15797# 0.01335f
C2281 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout CLK 0.28425f
C2282 Nand_Gate_3.B RingCounter_0.D_FlipFlop_2.Inverter_0.Vout 0.29368f
C2283 a_55443_15797# VDD 0.03339f
C2284 D_FlipFlop_1.Inverter_0.Vout a_134897_33443# 0.04995f
C2285 a_118353_52572# RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout 0.05964f
C2286 FFCLR a_132925_36157# 0.0468f
C2287 a_128237_24200# VDD 0.02521f
C2288 a_44403_13083# VDD 0.05686f
C2289 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout VDD 2.31704f
C2290 D_FlipFlop_6.Nand_Gate_0.Vout Q1 0.11443f
C2291 Nand_Gate_6.Vout Q0 0.05048f
C2292 a_112745_52572# a_113359_52572# 0.05935f
C2293 D_FlipFlop_5.3-input-nand_0.Vout a_132925_26914# 0.04995f
C2294 a_134283_27764# VDD 0.02521f
C2295 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout VDD 2.73332f
C2296 D_FlipFlop_6.Inverter_1.Vout a_130209_20636# 0.04995f
C2297 Nand_Gate_0.A a_134897_37007# 0.04682f
C2298 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C a_43789_15797# 0.04443f
C2299 D_FlipFlop_6.Q' a_128851_20636# 0.01335f
C2300 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout VDD 1.70415f
C2301 Nand_Gate_7.B a_68455_15797# 0.04995f
C2302 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_32749_13083# 0.05964f
C2303 a_65125_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.04443f
C2304 a_65869_15797# VDD 0.03178f
C2305 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout 0.04109f
C2306 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Q' 0.06632f
C2307 D_FlipFlop_7.Nand_Gate_0.Vout a_130209_19786# 0.05964f
C2308 D_FlipFlop_0.Q' D_FlipFlop_0.Nand_Gate_0.Vout 0.06632f
C2309 Nand_Gate_0.A RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.08024f
C2310 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout CLK 0.30716f
C2311 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout VDD 1.56255f
C2312 And_Gate_6.Inverter_0.Vin Comparator_0.Vinm 0.02639f
C2313 D_FlipFlop_4.Nand_Gate_1.Vout a_130209_27764# 0.05964f
C2314 Nand_Gate_6.B a_82057_16975# 0.04443f
C2315 Nand_Gate_6.Vout EN 0.10992f
C2316 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout VDD 2.07373f
C2317 Nand_Gate_5.B Nand_Gate_4.B 0.06408f
C2318 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout VDD 2.46653f
C2319 CDAC8_0.switch_0.Z EN 0.56688f
C2320 a_51499_49858# VDD 0.01712f
C2321 D_FlipFlop_5.Inverter_1.Vout a_130209_24200# 0.04995f
C2322 a_93097_47663# CLK 0.02953f
C2323 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.30154f
C2324 FFCLR a_134897_39721# 0.08419f
C2325 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_111387_49858# 0.05964f
C2326 D_FlipFlop_1.Inverter_1.Vout EN 0.59727f
C2327 a_112001_13083# VDD 0.02865f
C2328 Nand_Gate_1.B a_132925_30478# 0.04789f
C2329 D_FlipFlop_5.Q' a_128851_24200# 0.01335f
C2330 Nand_Gate_6.B Q1 0.06203f
C2331 FFCLR RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.08024f
C2332 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout EN 0.41172f
C2333 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout a_68585_49858# 0.04995f
C2334 Nand_Gate_0.A CDAC8_0.switch_6.Z 9.49208f
C2335 D_FlipFlop_3.3-input-nand_2.Vout VDD 2.77266f
C2336 D_FlipFlop_1.3-input-nand_1.Vout a_134897_33443# 0.01335f
C2337 RingCounter_0.D_FlipFlop_7.Q' CLK 0.09401f
C2338 CDAC8_0.switch_6.Z CDAC8_0.switch_7.Z 14.5275f
C2339 D_FlipFlop_5.Inverter_0.Vout VDD 1.37371f
C2340 a_96273_49858# EN 0.01149f
C2341 RingCounter_0.D_FlipFlop_7.Q' Nand_Gate_5.A 1.10693f
C2342 RingCounter_0.D_FlipFlop_2.Q' VDD 1.96503f
C2343 a_132311_44135# a_132925_44135# 0.05935f
C2344 D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.48313f
C2345 D_FlipFlop_4.Q' Q3 1.06575f
C2346 RingCounter_0.D_FlipFlop_6.Q' RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout 0.11654f
C2347 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_2.C 1.09975f
C2348 a_128851_43285# Q5 0.01335f
C2349 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout CLK 0.03479f
C2350 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_77523_13083# 0.01335f
C2351 CDAC8_0.switch_9.Z Q7 0.29749f
C2352 a_98989_13083# CLK 0.03129f
C2353 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout CLK 0.23464f
C2354 CDAC8_0.switch_2.Z VDD 1.31283f
C2355 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout a_112001_15797# 0.05964f
C2356 a_118353_49858# VDD 0.0325f
C2357 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.06465f
C2358 D_FlipFlop_4.Q' VDD 1.89806f
C2359 a_47119_52572# FFCLR 0.06113f
C2360 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.0857f
C2361 RingCounter_0.D_FlipFlop_14.Q' VDD 1.95446f
C2362 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_6.3-input-nand_2.C 0.06594f
C2363 D_FlipFlop_2.3-input-nand_2.C D_FlipFlop_2.Nand_Gate_1.Vout 0.1541f
C2364 a_128237_44135# VDD 0.02521f
C2365 a_106569_15797# EN 0.04443f
C2366 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout a_123655_15797# 0.01335f
C2367 CDAC8_0.switch_2.Z CDAC8_0.switch_1.Z 0.06088f
C2368 a_111387_52572# RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout 0.05964f
C2369 FFCLR a_134897_20636# 0.04005f
C2370 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout CLK 0.30735f
C2371 D_FlipFlop_3.3-input-nand_1.Vout a_132311_40571# 0.04444f
C2372 D_FlipFlop_7.Inverter_1.Vout D_FlipFlop_7.3-input-nand_2.C 0.25579f
C2373 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.15399f
C2374 a_67841_13083# VDD 0.02865f
C2375 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout CLK 0.15609f
C2376 Nand_Gate_2.Vout EN 0.11847f
C2377 a_105955_15797# VDD 0.02906f
C2378 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout 0.1182f
C2379 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout EN 0.97489f
C2380 D_FlipFlop_5.3-input-nand_1.Vout VDD 1.78032f
C2381 FFCLR D_FlipFlop_1.3-input-nand_0.Vout 1.1762f
C2382 a_100961_15797# a_101575_15797# 0.05935f
C2383 a_76165_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.05964f
C2384 a_98989_15797# a_99603_15797# 0.05935f
C2385 FFCLR D_FlipFlop_5.Inverter_1.Vout 0.56927f
C2386 CLK Q6 0.1175f
C2387 D_FlipFlop_7.3-input-nand_2.Vout D_FlipFlop_7.3-input-nand_1.Vout 0.06465f
C2388 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout CLK 0.03479f
C2389 D_FlipFlop_0.Inverter_0.Vout a_134283_44135# 0.04443f
C2390 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout a_113359_52572# 0.04444f
C2391 Nand_Gate_5.B RingCounter_0.D_FlipFlop_10.Inverter_0.Vout 0.29368f
C2392 Nand_Gate_2.A a_134897_40571# 0.0468f
C2393 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout CLK 0.12047f
C2394 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout VDD 2.07373f
C2395 a_96273_52572# VDD 0.02521f
C2396 a_52113_49858# EN 0.01149f
C2397 a_128851_20636# VDD 0.01186f
C2398 D_FlipFlop_0.3-input-nand_0.Vout a_134283_46849# 0.05964f
C2399 a_90665_52572# VDD 0.01186f
C2400 a_112615_13083# EN 0.0452f
C2401 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout 0.04107f
C2402 a_63153_52572# RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.05964f
C2403 a_54829_13083# CLK 0.03129f
C2404 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout 0.30154f
C2405 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_12.Inverter_1.Vout 0.25963f
C2406 a_107927_15797# VDD 0.02906f
C2407 D_FlipFlop_2.3-input-nand_2.C a_130209_37007# 0.04443f
C2408 RingCounter_0.D_FlipFlop_11.Q' a_94915_13083# 0.06113f
C2409 D_FlipFlop_2.3-input-nand_0.Vout a_134283_39721# 0.05964f
C2410 a_42431_52572# VDD 0.05686f
C2411 a_57545_52572# Nand_Gate_3.B 0.01335f
C2412 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout a_79495_15797# 0.01335f
C2413 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout EN 0.78685f
C2414 a_74193_49858# VDD 0.0325f
C2415 a_130209_46849# VDD 0.02521f
C2416 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_0.Vout 1.03054f
C2417 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout CLK 0.155f
C2418 D_FlipFlop_4.Inverter_1.Vout VDD 1.73058f
C2419 a_104137_16975# VDD 0.02521f
C2420 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C EN 0.07664f
C2421 Comparator_0.Vinm Q6 0.5602f
C2422 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout EN 0.13192f
C2423 Nand_Gate_3.B RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout 0.08377f
C2424 RingCounter_0.D_FlipFlop_11.Q' CLK 0.09276f
C2425 a_44403_15797# VDD 0.03339f
C2426 a_128851_30478# Q3 0.01335f
C2427 a_41073_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout 0.05964f
C2428 D_FlipFlop_1.3-input-nand_2.Vout a_132925_36157# 0.01335f
C2429 a_121683_13083# CLK 0.03129f
C2430 D_FlipFlop_1.Nand_Gate_1.Vout Q7 0.06503f
C2431 D_FlipFlop_3.Nand_Gate_0.Vout Q5 0.11443f
C2432 Nand_Gate_6.A a_83875_15797# 0.06113f
C2433 a_48937_47663# VDD 0.02521f
C2434 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout 0.30154f
C2435 Nand_Gate_7.B D_FlipFlop_6.Inverter_0.Vout 0.25826f
C2436 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C VDD 3.56545f
C2437 a_128237_37007# a_128851_37007# 0.05935f
C2438 a_128851_30478# VDD 0.01186f
C2439 Nand_Gate_1.B Nand_Gate_1.A 0.07512f
C2440 Nand_Gate_4.B D_FlipFlop_7.3-input-nand_2.Vout 0.90723f
C2441 D_FlipFlop_2.3-input-nand_0.Vout D_FlipFlop_2.3-input-nand_1.Vout 0.04107f
C2442 D_FlipFlop_2.3-input-nand_2.Vout a_132311_37007# 0.04443f
C2443 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout a_35335_15797# 0.01335f
C2444 a_68455_13083# EN 0.0452f
C2445 D_FlipFlop_4.3-input-nand_1.Vout a_132925_27764# 0.04543f
C2446 D_FlipFlop_2.Q' Q5 0.01194f
C2447 D_FlipFlop_0.3-input-nand_1.Vout VDD 1.78032f
C2448 CDAC8_0.switch_9.Z CDAC8_0.switch_0.Z 3.66237f
C2449 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout EN 0.61894f
C2450 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout CLK 0.30716f
C2451 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_2.C 1.09975f
C2452 RingCounter_0.D_FlipFlop_11.Q' RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout 0.06632f
C2453 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout a_43045_49858# 0.04443f
C2454 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C VDD 3.61242f
C2455 Nand_Gate_6.B D_FlipFlop_5.Inverter_0.Vout 0.25819f
C2456 a_86591_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 0.01335f
C2457 a_90535_13083# VDD 0.01327f
C2458 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout EN 1.03094f
C2459 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_2.C 0.06594f
C2460 a_132311_43285# VDD 0.02521f
C2461 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_73579_49858# 0.01335f
C2462 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout 0.16429f
C2463 CDAC8_0.switch_0.Z Nand_Gate_7.B 3.36457f
C2464 D_FlipFlop_5.Nand_Gate_1.Vout VDD 1.46545f
C2465 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout EN 0.78734f
C2466 Nand_Gate_5.A a_134897_44135# 0.0468f
C2467 Nand_Gate_5.B Q5 0.06203f
C2468 D_FlipFlop_1.3-input-nand_2.C a_132311_36157# 0.04443f
C2469 RingCounter_0.D_FlipFlop_1.Q' CLK 0.09276f
C2470 Nand_Gate_0.A a_73579_52572# 0.04995f
C2471 a_111387_52572# RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.04443f
C2472 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout a_109285_49858# 0.04444f
C2473 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C VDD 3.54707f
C2474 Nand_Gate_7.B D_FlipFlop_6.3-input-nand_1.Vout 0.07303f
C2475 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.48392f
C2476 a_77523_13083# CLK 0.03129f
C2477 RingCounter_0.D_FlipFlop_17.Q' CLK 0.09276f
C2478 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout 0.04107f
C2479 Nand_Gate_1.A CLK 0.38549f
C2480 FFCLR D_FlipFlop_6.Q' 0.03748f
C2481 a_97631_49858# VDD 0.06071f
C2482 And_Gate_0.Inverter_0.Vin VDD 1.38853f
C2483 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout CLK 0.23464f
C2484 Nand_Gate_1.B Q0 0.06233f
C2485 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout Nand_Gate_3.B 0.12214f
C2486 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout VDD 2.8604f
C2487 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.06465f
C2488 a_84489_15797# VDD 0.01571f
C2489 Nand_Gate_6.B D_FlipFlop_5.3-input-nand_1.Vout 0.07299f
C2490 D_FlipFlop_6.3-input-nand_0.Vout a_134283_23350# 0.05964f
C2491 RingCounter_0.D_FlipFlop_16.Q CDAC8_0.switch_7.Z 0.08064f
C2492 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.Inverter_1.Vout 0.25579f
C2493 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0846f
C2494 CDAC8_0.switch_8.Z Q5 0.32925f
C2495 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout VDD 2.31704f
C2496 a_57415_15797# VDD 0.06072f
C2497 a_119711_52572# VDD 0.01186f
C2498 FFCLR a_134897_36157# 0.04564f
C2499 a_46375_13083# VDD 0.01327f
C2500 a_130209_24200# VDD 0.02521f
C2501 Nand_Gate_1.B EN 1.13628f
C2502 And_Gate_1.Inverter_0.Vin VDD 1.39208f
C2503 a_94915_15797# VDD 0.02906f
C2504 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout a_118967_13083# 0.04995f
C2505 D_FlipFlop_4.Nand_Gate_0.Vout Q3 0.11443f
C2506 a_113359_52572# RingCounter_0.D_FlipFlop_7.Q' 0.04443f
C2507 D_FlipFlop_1.3-input-nand_2.Vout D_FlipFlop_1.3-input-nand_0.Vout 0.0846f
C2508 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout 0.1541f
C2509 D_FlipFlop_5.3-input-nand_0.Vout a_134283_26914# 0.05964f
C2510 Nand_Gate_0.B a_71017_47663# 0.04443f
C2511 Nand_Gate_0.A CDAC8_0.switch_7.Z 7.14466f
C2512 D_FlipFlop_2.3-input-nand_2.Vout VDD 2.77266f
C2513 a_64511_52572# EN 0.045f
C2514 Nand_Gate_4.A a_40329_15797# 0.01335f
C2515 Nand_Gate_7.B RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout 0.0839f
C2516 D_FlipFlop_4.Nand_Gate_0.Vout VDD 1.48313f
C2517 a_134283_39721# a_134897_39721# 0.05935f
C2518 Comparator_0.Vinm a_75898_18814# 0.0277f
C2519 a_33363_13083# CLK 0.02953f
C2520 CDAC8_0.switch_6.Z Q7 0.66797f
C2521 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout CLK 0.69657f
C2522 CLK Q0 1.75855f
C2523 D_FlipFlop_0.Nand_Gate_1.Vout VDD 1.46545f
C2524 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout 0.0846f
C2525 D_FlipFlop_1.Inverter_1.Vout D_FlipFlop_1.Nand_Gate_1.Vout 0.30154f
C2526 D_FlipFlop_2.Q' D_FlipFlop_2.Nand_Gate_0.Vout 0.06632f
C2527 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_2.C 1.09975f
C2528 a_53471_49858# VDD 0.06071f
C2529 a_115177_47663# CLK 0.06925f
C2530 a_118967_15797# RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.04443f
C2531 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout a_113359_49858# 0.04444f
C2532 D_FlipFlop_4.3-input-nand_2.Vout a_132925_30478# 0.01335f
C2533 a_116995_13083# VDD 0.02521f
C2534 a_123785_49858# a_124399_49858# 0.05935f
C2535 Nand_Gate_5.A a_115177_47663# 0.04443f
C2536 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout CLK 0.29644f
C2537 a_128237_40571# VDD 0.02521f
C2538 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout a_90535_13083# 0.04995f
C2539 Nand_Gate_1.A RingCounter_0.D_FlipFlop_9.Q' 1.05791f
C2540 D_FlipFlop_5.Nand_Gate_1.Vout D_FlipFlop_6.Nand_Gate_0.Vout 0.01681f
C2541 EN CLK 8.56602f
C2542 a_99603_15797# EN 0.045f
C2543 a_132311_36157# a_132925_36157# 0.05935f
C2544 Nand_Gate_5.A EN 0.49282f
C2545 Nand_Gate_0.A RingCounter_0.D_FlipFlop_3.Inverter_0.Vout 0.29368f
C2546 a_100961_13083# CLK 0.04619f
C2547 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_2.Inverter_1.Vout 0.01422f
C2548 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout EN 0.09127f
C2549 Comparator_0.Vinm Q0 0.13685f
C2550 a_120325_49858# VDD 0.0301f
C2551 Nand_Gate_3.B a_58159_49858# 0.04741f
C2552 FFCLR VDD 28.0963f
C2553 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_5.Inverter_1.Vout 0.06445f
C2554 a_57545_52572# a_58159_52572# 0.05935f
C2555 a_130209_44135# VDD 0.02521f
C2556 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_85847_13083# 0.04443f
C2557 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout EN 0.24889f
C2558 D_FlipFlop_1.Inverter_1.Vout a_130209_33443# 0.04995f
C2559 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout CLK 0.03479f
C2560 a_43789_15797# VDD 0.03178f
C2561 a_74807_15797# RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.04443f
C2562 D_FlipFlop_0.3-input-nand_2.C VDD 2.74431f
C2563 Nand_Gate_4.A EN 0.42016f
C2564 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout EN 0.61894f
C2565 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.06465f
C2566 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.3-input-nand_1.Vout 0.08671f
C2567 D_FlipFlop_4.3-input-nand_2.C a_132311_30478# 0.04443f
C2568 D_FlipFlop_3.3-input-nand_1.Vout a_134283_40571# 0.05964f
C2569 Comparator_0.Vinm EN 14.0874f
C2570 a_124399_52572# Nand_Gate_5.B 0.06113f
C2571 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout VDD 2.46653f
C2572 a_107313_49858# CLK 0.04619f
C2573 a_72835_13083# VDD 0.02521f
C2574 a_134283_43285# VDD 0.02521f
C2575 a_46505_52572# a_47119_52572# 0.05935f
C2576 a_101705_49858# a_102319_49858# 0.05935f
C2577 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout a_100961_15797# 0.05964f
C2578 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout CLK 0.23464f
C2579 a_134897_19786# VDD 0.01186f
C2580 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout EN 0.41121f
C2581 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout CLK 0.71041f
C2582 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout a_51369_15797# 0.04995f
C2583 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout VDD 2.88547f
C2584 Nand_Gate_2.A CDAC8_0.switch_6.Z 3.68553f
C2585 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.3-input-nand_1.Vout 0.08671f
C2586 a_62539_52572# VDD 0.0564f
C2587 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout 0.1541f
C2588 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout VDD 2.73618f
C2589 a_132311_20636# VDD 0.02521f
C2590 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.1182f
C2591 RingCounter_0.D_FlipFlop_4.Q' VDD 1.96503f
C2592 a_56801_13083# CLK 0.04619f
C2593 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout CLK 0.03479f
C2594 D_FlipFlop_2.Nand_Gate_1.Vout a_128851_37007# 0.04995f
C2595 D_FlipFlop_0.Nand_Gate_0.Vout a_128851_46849# 0.04995f
C2596 D_FlipFlop_2.3-input-nand_2.C a_132925_37007# 0.01335f
C2597 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout a_106569_13083# 0.04995f
C2598 D_FlipFlop_3.Inverter_1.Vout a_130209_43285# 0.04443f
C2599 a_83875_15797# RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.04444f
C2600 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_99603_13083# 0.04543f
C2601 RingCounter_0.D_FlipFlop_1.Q' Nand_Gate_3.B 1.10693f
C2602 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C VDD 2.99599f
C2603 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_94915_13083# 0.04444f
C2604 a_40459_52572# VDD 0.01606f
C2605 Nand_Gate_5.B Q1 0.06203f
C2606 a_134283_20636# a_134897_20636# 0.05935f
C2607 D_FlipFlop_4.Inverter_0.Vout a_134897_27764# 0.04995f
C2608 a_76165_49858# VDD 0.0301f
C2609 a_30647_15797# RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.04443f
C2610 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_87949_13083# 0.04444f
C2611 D_FlipFlop_0.Inverter_0.Vout VDD 1.37367f
C2612 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout a_121069_13083# 0.04443f
C2613 D_FlipFlop_2.Nand_Gate_0.Vout a_128851_39721# 0.04995f
C2614 D_FlipFlop_4.Q' a_128851_27764# 0.01335f
C2615 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.0857f
C2616 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_0.Vout 0.0846f
C2617 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout CLK 0.23464f
C2618 D_FlipFlop_2.3-input-nand_1.Vout D_FlipFlop_1.3-input-nand_0.Vout 0.01418f
C2619 Nand_Gate_6.B a_94915_15797# 0.06113f
C2620 Nand_Gate_4.B RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout 0.1182f
C2621 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout 0.1182f
C2622 D_FlipFlop_0.Q' a_128851_44135# 0.01335f
C2623 a_86591_52572# a_87205_52572# 0.05935f
C2624 a_128237_17072# VDD 0.02521f
C2625 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout a_123785_52572# 0.04995f
C2626 D_FlipFlop_3.3-input-nand_1.Vout VDD 1.78032f
C2627 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout a_62539_49858# 0.04995f
C2628 Nand_Gate_0.A D_FlipFlop_2.Inverter_1.Vout 0.16179f
C2629 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout a_56801_13083# 0.04443f
C2630 a_134283_24200# a_134897_24200# 0.05935f
C2631 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.04109f
C2632 a_63153_49858# CLK 0.04619f
C2633 a_56187_52572# RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout 0.05964f
C2634 a_28675_13083# VDD 0.02521f
C2635 a_46375_15797# VDD 0.06072f
C2636 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout CLK 0.03574f
C2637 a_73579_52572# RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.01335f
C2638 a_79625_49858# a_80239_49858# 0.05935f
C2639 a_132311_36157# D_FlipFlop_1.3-input-nand_0.Vout 0.04444f
C2640 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout 0.04107f
C2641 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout a_111387_52572# 0.04443f
C2642 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout 0.06445f
C2643 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout EN 0.97489f
C2644 a_71017_47663# VDD 0.02521f
C2645 a_132311_39721# VDD 0.02521f
C2646 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_39715_13083# 0.04444f
C2647 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_32749_13083# 0.04444f
C2648 a_130209_30478# VDD 0.02521f
C2649 Nand_Gate_1.B Nand_Gate_7.B 0.0543f
C2650 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout a_30647_13083# 0.04995f
C2651 RingCounter_0.D_FlipFlop_14.Q' a_61795_15797# 0.04443f
C2652 a_118353_52572# VDD 0.02521f
C2653 D_FlipFlop_4.3-input-nand_1.Vout a_134897_27764# 0.01335f
C2654 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout a_58159_52572# 0.04444f
C2655 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout a_52113_49858# 0.04443f
C2656 a_112745_52572# VDD 0.01186f
C2657 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout 0.06594f
C2658 And_Gate_6.Inverter_0.Vin a_103765_47663# 0.05964f
C2659 a_132925_46849# VDD 0.01186f
C2660 a_65125_52572# VDD 0.02521f
C2661 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_118353_49858# 0.05964f
C2662 a_132311_30478# a_132925_30478# 0.05935f
C2663 D_FlipFlop_6.3-input-nand_2.C D_FlipFlop_6.Nand_Gate_1.Vout 0.1541f
C2664 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout 0.04109f
C2665 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout 1.09975f
C2666 FFCLR a_134897_30478# 0.08418f
C2667 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout CLK 0.03479f
C2668 a_95529_13083# VDD 0.0563f
C2669 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout CLK 0.23464f
C2670 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout 0.06594f
C2671 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout a_75551_49858# 0.04543f
C2672 CDAC8_0.switch_9.Z CLK 0.19385f
C2673 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout a_54085_49858# 0.04443f
C2674 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout a_55443_15797# 0.01335f
C2675 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.04107f
C2676 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout CLK 0.155f
C2677 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout 0.06445f
C2678 FFCLR Nand_Gate_6.B 0.93903f
C2679 Nand_Gate_0.A RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout 0.08377f
C2680 D_FlipFlop_5.3-input-nand_2.C D_FlipFlop_5.Nand_Gate_1.Vout 0.1541f
C2681 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout VDD 1.76876f
C2682 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.0857f
C2683 a_69199_52572# Nand_Gate_0.A 0.06113f
C2684 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout VDD 2.16362f
C2685 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout a_67227_49858# 0.04995f
C2686 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout 0.0846f
C2687 a_57545_49858# a_58159_49858# 0.05935f
C2688 EN Q4 0.2481f
C2689 Nand_Gate_3.B EN 0.99738f
C2690 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout a_87949_15797# 0.05964f
C2691 Nand_Gate_7.B CLK 0.58232f
C2692 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110643_15797# 0.01335f
C2693 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout CLK 0.03342f
C2694 a_100347_49858# VDD 0.04111f
C2695 RingCounter_0.D_FlipFlop_14.Q' a_62409_13083# 0.01335f
C2696 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.3-input-nand_2.Vout 0.16429f
C2697 a_121069_13083# a_121683_13083# 0.05935f
C2698 a_100961_15797# VDD 0.03119f
C2699 Nand_Gate_1.A a_101575_15797# 0.04995f
C2700 D_FlipFlop_1.3-input-nand_2.Vout VDD 2.77266f
C2701 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout a_76165_52572# 0.04444f
C2702 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout 0.16429f
C2703 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout EN 0.24889f
C2704 D_FlipFlop_6.3-input-nand_2.C a_130209_20636# 0.04443f
C2705 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout VDD 2.07373f
C2706 a_132311_40571# a_132925_40571# 0.05935f
C2707 CDAC8_0.switch_9.Z Comparator_0.Vinm 0.22008p
C2708 Nand_Gate_2.A D_FlipFlop_3.Inverter_1.Vout 0.16207f
C2709 CDAC8_0.switch_7.Z Q7 1.88874f
C2710 a_84619_52572# a_85233_52572# 0.05935f
C2711 FFCLR D_FlipFlop_6.3-input-nand_2.Vout 0.06105f
C2712 D_FlipFlop_3.Nand_Gate_1.Vout VDD 1.46545f
C2713 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout CLK 0.30716f
C2714 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C VDD 3.59745f
C2715 a_86591_49858# CLK 0.03129f
C2716 a_51369_13083# VDD 0.0563f
C2717 a_132925_24200# VDD 0.01186f
C2718 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout VDD 2.04843f
C2719 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout 0.06445f
C2720 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout EN 1.03094f
C2721 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_122427_49858# 0.05964f
C2722 D_FlipFlop_5.3-input-nand_2.C a_130209_24200# 0.04443f
C2723 a_128237_37007# VDD 0.02521f
C2724 Comparator_0.Vinm Nand_Gate_7.B 2.56398f
C2725 D_FlipFlop_1.3-input-nand_2.C EN 0.79121f
C2726 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C a_110029_13083# 0.05964f
C2727 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C EN 0.07732f
C2728 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout a_68585_52572# 0.04995f
C2729 RingCounter_0.D_FlipFlop_3.Q' CLK 0.09276f
C2730 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout a_79625_49858# 0.04995f
C2731 D_FlipFlop_2.3-input-nand_1.Vout a_132311_37007# 0.04444f
C2732 Nand_Gate_0.B a_84619_52572# 0.04995f
C2733 D_FlipFlop_3.Q' a_128237_40571# 0.06113f
C2734 RingCounter_0.D_FlipFlop_1.Q' a_57545_49858# 0.01335f
C2735 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_110029_13083# 0.04444f
C2736 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.30154f
C2737 Nand_Gate_6.A VDD 4.18085f
C2738 a_75898_28676# Comparator_0.Vinm 0.03583f
C2739 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.0857f
C2740 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout VDD 1.48392f
C2741 D_FlipFlop_6.Nand_Gate_1.Vout D_FlipFlop_7.Nand_Gate_0.Vout 0.01681f
C2742 a_56187_52572# RingCounter_0.D_FlipFlop_1.Inverter_1.Vout 0.04443f
C2743 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_6.Inverter_1.Vout 0.01422f
C2744 D_FlipFlop_0.3-input-nand_0.Vout VDD 1.77946f
C2745 a_56187_49858# VDD 0.04111f
C2746 RingCounter_0.D_FlipFlop_8.Q' CLK 0.09276f
C2747 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout VDD 2.73332f
C2748 a_98989_13083# a_99603_13083# 0.05935f
C2749 D_FlipFlop_6.3-input-nand_0.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.04107f
C2750 a_132311_30478# D_FlipFlop_4.3-input-nand_0.Vout 0.04444f
C2751 D_FlipFlop_6.3-input-nand_2.Vout a_132311_20636# 0.04443f
C2752 a_118967_13083# VDD 0.02578f
C2753 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout CLK 0.70923f
C2754 Nand_Gate_1.B D_FlipFlop_4.Inverter_0.Vout 0.25807f
C2755 a_116995_15797# a_117609_15797# 0.05935f
C2756 D_FlipFlop_3.Inverter_0.Vout a_134283_40571# 0.04443f
C2757 Nand_Gate_5.A D_FlipFlop_0.Q' 0.06453f
C2758 a_130209_40571# VDD 0.02521f
C2759 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout a_32749_13083# 0.04443f
C2760 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout VDD 2.8604f
C2761 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C VDD 3.56545f
C2762 a_73449_15797# EN 0.04443f
C2763 FFCLR D_FlipFlop_3.Q' 0.03748f
C2764 RingCounter_0.D_FlipFlop_5.Q' RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout 0.11654f
C2765 And_Gate_2.Inverter_0.Vin VDD 1.38853f
C2766 Nand_Gate_7.A VDD 4.18085f
C2767 a_139696_27690# a_138318_16817# 0.4942f
C2768 a_134283_44135# a_134897_44135# 0.05935f
C2769 D_FlipFlop_1.3-input-nand_0.Vout a_134283_36157# 0.05964f
C2770 a_42431_49858# CLK 0.03129f
C2771 D_FlipFlop_5.3-input-nand_2.Vout a_132311_24200# 0.04443f
C2772 D_FlipFlop_5.3-input-nand_0.Vout D_FlipFlop_5.3-input-nand_1.Vout 0.04107f
C2773 a_78881_15797# CLK 0.04619f
C2774 a_134283_39721# VDD 0.02521f
C2775 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.0857f
C2776 Nand_Gate_4.A RingCounter_0.D_FlipFlop_8.Q' 1.05791f
C2777 D_FlipFlop_7.3-input-nand_2.Vout a_132311_19786# 0.05964f
C2778 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout a_86591_52572# 0.04995f
C2779 RingCounter_0.D_FlipFlop_17.Q' RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.11654f
C2780 a_117609_15797# VDD 0.01571f
C2781 a_123785_49858# VDD 0.0563f
C2782 D_FlipFlop_3.Inverter_1.Vout D_FlipFlop_3.3-input-nand_2.C 0.25579f
C2783 Nand_Gate_2.A CDAC8_0.switch_7.Z 7.18772f
C2784 a_86591_52572# EN 0.045f
C2785 a_132925_44135# VDD 0.01186f
C2786 a_58159_52572# RingCounter_0.D_FlipFlop_1.Q' 0.04443f
C2787 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C a_88563_13083# 0.01335f
C2788 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout CLK 0.29759f
C2789 FFCLR D_FlipFlop_5.3-input-nand_2.C 0.76213f
C2790 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout 0.30154f
C2791 a_72835_15797# a_73449_15797# 0.05935f
C2792 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout a_73579_49858# 0.04995f
C2793 Nand_Gate_1.B D_FlipFlop_4.3-input-nand_1.Vout 0.07295f
C2794 a_57545_52572# VDD 0.01186f
C2795 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_66483_15797# 0.04995f
C2796 a_74807_15797# VDD 0.02906f
C2797 a_76909_13083# a_77523_13083# 0.05935f
C2798 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_121069_13083# 0.04444f
C2799 a_109285_49858# CLK 0.03129f
C2800 D_FlipFlop_5.Q' Q2 1.06526f
C2801 D_FlipFlop_3.Inverter_0.Vout VDD 1.37367f
C2802 a_74807_13083# VDD 0.02578f
C2803 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.08671f
C2804 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout CLK 0.30606f
C2805 a_47119_52572# RingCounter_0.D_FlipFlop_17.Q' 0.04443f
C2806 a_46505_52572# VDD 0.0563f
C2807 Nand_Gate_1.Vout VDD 1.40515f
C2808 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout CLK 0.29644f
C2809 a_98989_15797# RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.04444f
C2810 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C a_121069_15797# 0.04443f
C2811 D_FlipFlop_2.3-input-nand_1.Vout VDD 1.78032f
C2812 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout VDD 1.86552f
C2813 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout 0.04107f
C2814 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout VDD 2.73332f
C2815 CDAC8_0.switch_9.Z Q4 0.29232f
C2816 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C EN 0.07664f
C2817 a_134283_20636# VDD 0.02521f
C2818 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout CLK 0.155f
C2819 a_29289_15797# VDD 0.01186f
C2820 And_Gate_6.Inverter_0.Vin VDD 1.43186f
C2821 FFCLR a_52113_52572# 0.04443f
C2822 Nand_Gate_4.B And_Gate_1.Inverter_0.Vin 0.06473f
C2823 D_FlipFlop_4.3-input-nand_2.C VDD 2.74431f
C2824 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.25963f
C2825 Nand_Gate_0.B RingCounter_0.D_FlipFlop_4.Inverter_0.Vout 0.29368f
C2826 FFCLR D_FlipFlop_7.3-input-nand_1.Vout 0.95252f
C2827 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout a_101575_13083# 0.01335f
C2828 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C CLK 0.30966f
C2829 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout a_96887_13083# 0.05964f
C2830 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout VDD 2.75373f
C2831 a_79625_49858# VDD 0.06015f
C2832 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout a_89921_13083# 0.05964f
C2833 a_132311_36157# VDD 0.02521f
C2834 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout a_84489_13083# 0.04995f
C2835 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_77523_13083# 0.04543f
C2836 a_28675_15797# a_29289_15797# 0.05935f
C2837 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_72835_13083# 0.04444f
C2838 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout EN 0.48849f
C2839 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout a_112001_13083# 0.04443f
C2840 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_65869_13083# 0.04444f
C2841 FFCLR a_128851_27764# 0.04443f
C2842 EN Q2 0.2481f
C2843 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout CLK 0.03574f
C2844 RingCounter_0.D_FlipFlop_9.Q' a_105955_13083# 0.06113f
C2845 a_87205_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.04443f
C2846 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout a_40459_49858# 0.04995f
C2847 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_6.Q' 0.06632f
C2848 a_130209_17072# VDD 0.02521f
C2849 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_2.C 0.25579f
C2850 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout a_110029_15797# 0.05964f
C2851 D_FlipFlop_7.Inverter_0.Vout a_134897_17072# 0.04995f
C2852 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout EN 0.09065f
C2853 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout EN 0.6089f
C2854 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_53471_49858# 0.01335f
C2855 a_54829_13083# a_55443_13083# 0.05935f
C2856 a_65125_49858# CLK 0.03129f
C2857 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout VDD 2.46653f
C2858 a_30647_13083# VDD 0.02578f
C2859 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout a_78267_49858# 0.04995f
C2860 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C a_76909_15797# 0.04443f
C2861 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout 0.08671f
C2862 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.3-input-nand_1.Vout 0.08671f
C2863 D_FlipFlop_7.Q' a_128851_17072# 0.01335f
C2864 Nand_Gate_6.B Nand_Gate_6.A 0.07512f
C2865 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout a_118967_15797# 0.05964f
C2866 a_93097_47663# VDD 0.02521f
C2867 CDAC8_0.switch_6.Z CLK 0.21538f
C2868 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_8.3-input-nand_2.C 1.09975f
C2869 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout a_41687_13083# 0.05964f
C2870 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout a_34721_13083# 0.05964f
C2871 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_84619_49858# 0.01335f
C2872 a_48565_16975# CLK 0.04479f
C2873 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout a_29289_13083# 0.04995f
C2874 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout EN 0.78734f
C2875 a_84619_52572# VDD 0.0564f
C2876 RingCounter_0.D_FlipFlop_7.Q' VDD 1.96539f
C2877 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C a_54829_13083# 0.05964f
C2878 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout CLK 0.03479f
C2879 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout a_120325_49858# 0.04444f
C2880 FFCLR Nand_Gate_4.B 0.89725f
C2881 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout a_96887_15797# 0.04443f
C2882 Nand_Gate_6.B And_Gate_2.Inverter_0.Vin 0.04751f
C2883 a_132311_17072# a_132925_17072# 0.05935f
C2884 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout VDD 1.48392f
C2885 Nand_Gate_6.A RingCounter_0.D_FlipFlop_12.Q' 1.05791f
C2886 a_98989_13083# VDD 0.02578f
C2887 a_128237_36157# Q7 0.06113f
C2888 a_128851_26914# Q2 0.01335f
C2889 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout VDD 2.88547f
C2890 Nand_Gate_2.A a_91279_49858# 0.04741f
C2891 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout EN 0.10495f
C2892 Nand_Gate_1.Vout And_Gate_3.Inverter_0.Vin 0.2638f
C2893 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout CLK 0.23464f
C2894 D_FlipFlop_0.Q' Q4 1.06174f
C2895 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C a_32749_15797# 0.04443f
C2896 CDAC8_0.switch_6.Z Comparator_0.Vinm 0.45096p
C2897 D_FlipFlop_0.Nand_Gate_1.Vout D_FlipFlop_3.Nand_Gate_0.Vout 0.01681f
C2898 a_134283_36157# a_134897_36157# 0.05935f
C2899 a_88563_15797# VDD 0.03339f
C2900 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout a_74807_15797# 0.05964f
C2901 D_FlipFlop_1.3-input-nand_0.Vout EN 0.08617f
C2902 a_32749_13083# a_33363_13083# 0.05935f
C2903 D_FlipFlop_2.Nand_Gate_1.Vout VDD 1.46545f
C2904 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout 0.04107f
C2905 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C a_43045_49858# 0.05964f
C2906 D_FlipFlop_1.Q' D_FlipFlop_1.Nand_Gate_0.Vout 0.06632f
C2907 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout EN 0.06649f
C2908 Nand_Gate_7.B a_73449_15797# 0.01335f
C2909 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout VDD 2.31704f
C2910 a_132925_30478# VDD 0.01186f
C2911 a_39715_15797# a_40329_15797# 0.05935f
C2912 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout EN 0.13192f
C2913 FFCLR D_FlipFlop_7.Nand_Gate_1.Vout 0.60828f
C2914 D_FlipFlop_3.Q' D_FlipFlop_3.Nand_Gate_1.Vout 0.11654f
C2915 a_102319_49858# VDD 0.02906f
C2916 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout VDD 1.70415f
C2917 a_98245_52572# RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.05964f
C2918 a_98989_15797# VDD 0.03178f
C2919 Nand_Gate_1.A RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout 0.08377f
C2920 Nand_Gate_1.B RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout 0.06503f
C2921 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout a_56187_52572# 0.04443f
C2922 VDD Q6 3.79753f
C2923 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout VDD 1.56255f
C2924 D_FlipFlop_6.3-input-nand_2.C a_132925_20636# 0.01335f
C2925 RingCounter_0.D_FlipFlop_2.Q' a_69199_49858# 0.06113f
C2926 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout VDD 2.86518f
C2927 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout 0.25963f
C2928 Nand_Gate_4.A a_35335_15797# 0.04995f
C2929 a_85233_52572# RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.05964f
C2930 a_87205_52572# VDD 0.02521f
C2931 D_FlipFlop_6.Inverter_1.Vout VDD 1.73058f
C2932 D_FlipFlop_2.Inverter_1.Vout D_FlipFlop_1.Inverter_1.Vout 0.01422f
C2933 a_79625_52572# Nand_Gate_0.B 0.01335f
C2934 a_134897_24200# VDD 0.01186f
C2935 a_54829_13083# VDD 0.02578f
C2936 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout 0.1541f
C2937 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout a_30647_15797# 0.05964f
C2938 D_FlipFlop_1.3-input-nand_2.C D_FlipFlop_1.Nand_Gate_1.Vout 0.1541f
C2939 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout a_124399_49858# 0.04444f
C2940 D_FlipFlop_5.3-input-nand_2.C a_132925_24200# 0.01335f
C2941 a_130209_37007# VDD 0.02521f
C2942 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_2.Q' 0.06632f
C2943 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout CLK 0.29644f
C2944 FFCLR D_FlipFlop_2.Q' 0.03748f
C2945 D_FlipFlop_7.3-input-nand_2.C D_FlipFlop_7.3-input-nand_0.Vout 0.06594f
C2946 Nand_Gate_1.B a_112615_15797# 0.04995f
C2947 Nand_Gate_4.B a_46375_15797# 0.04995f
C2948 D_FlipFlop_2.3-input-nand_1.Vout a_134283_37007# 0.05964f
C2949 Nand_Gate_0.B RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout 0.08377f
C2950 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout a_112001_13083# 0.05964f
C2951 Nand_Gate_6.A a_83875_13083# 0.04443f
C2952 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout VDD 1.76876f
C2953 CDAC8_0.switch_2.Z Q1 0.50779f
C2954 a_75898_46095# Comparator_0.Vinm 0.04537f
C2955 Nand_Gate_2.B And_Gate_6.Inverter_0.Vin 0.02391f
C2956 a_134283_36157# VDD 0.02521f
C2957 FFCLR D_FlipFlop_5.3-input-nand_0.Vout 0.1261f
C2958 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout CLK 0.03574f
C2959 Nand_Gate_0.B EN 0.99738f
C2960 a_42431_52572# RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout 0.01335f
C2961 RingCounter_0.D_FlipFlop_11.Q' VDD 1.95446f
C2962 a_58159_49858# VDD 0.02906f
C2963 RingCounter_0.D_FlipFlop_10.Q' a_116995_13083# 0.06113f
C2964 CDAC8_0.switch_9.Z Q2 0.38677f
C2965 a_121683_13083# VDD 0.05686f
C2966 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_10.Inverter_1.Vout 0.25963f
C2967 D_FlipFlop_5.Nand_Gate_0.Vout Q2 0.11443f
C2968 a_132925_40571# VDD 0.01186f
C2969 D_FlipFlop_7.Nand_Gate_1.Vout a_128237_17072# 0.04444f
C2970 FFCLR Nand_Gate_5.B 0.06347f
C2971 D_FlipFlop_0.Inverter_1.Vout a_130209_46849# 0.04443f
C2972 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout a_85233_49858# 0.04443f
C2973 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout CLK 0.30735f
C2974 a_106699_49858# EN 0.07058f
C2975 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout 0.0857f
C2976 D_FlipFlop_2.Inverter_1.Vout a_130209_39721# 0.04443f
C2977 D_FlipFlop_1.3-input-nand_2.C a_130209_33443# 0.04443f
C2978 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout CLK 0.30716f
C2979 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout EN 0.97489f
C2980 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout CLK 0.15609f
C2981 D_FlipFlop_2.Inverter_0.Vout VDD 1.37367f
C2982 a_108671_52572# RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout 0.01335f
C2983 D_FlipFlop_1.Nand_Gate_0.Vout a_128851_36157# 0.04995f
C2984 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout VDD 2.46653f
C2985 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout a_44403_13083# 0.04543f
C2986 a_89921_15797# a_90535_15797# 0.05935f
C2987 D_FlipFlop_4.3-input-nand_0.Vout VDD 1.77946f
C2988 a_87949_15797# a_88563_15797# 0.05935f
C2989 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_4.3-input-nand_2.C 0.06594f
C2990 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout a_101575_13083# 0.04995f
C2991 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout 0.04109f
C2992 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout CLK 0.03479f
C2993 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout 0.16429f
C2994 a_39715_15797# RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout 0.04444f
C2995 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout a_87205_49858# 0.04443f
C2996 Nand_Gate_2.B a_93097_47663# 0.04443f
C2997 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C EN 0.07732f
C2998 a_134897_44135# VDD 0.01186f
C2999 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout 0.06465f
C3000 CDAC8_0.switch_6.Z Q4 0.65162f
C3001 CDAC8_0.switch_7.Z Nand_Gate_1.B 4.80579f
C3002 a_128237_40571# Q5 0.04443f
C3003 Nand_Gate_2.A a_95659_52572# 0.04995f
C3004 RingCounter_0.D_FlipFlop_5.Q' CLK 0.09276f
C3005 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_13.Inverter_1.Vout 0.25963f
C3006 D_FlipFlop_4.3-input-nand_2.Vout D_FlipFlop_4.3-input-nand_1.Vout 0.06465f
C3007 FFCLR CDAC8_0.switch_8.Z 2.17565f
C3008 RingCounter_0.D_FlipFlop_1.Q' VDD 1.96503f
C3009 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout a_68455_15797# 0.01335f
C3010 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout a_123041_13083# 0.05964f
C3011 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout a_41687_15797# 0.05964f
C3012 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout a_117609_13083# 0.04995f
C3013 a_77523_13083# VDD 0.05686f
C3014 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C a_96887_13083# 0.04443f
C3015 D_FlipFlop_6.Nand_Gate_0.Vout D_FlipFlop_6.Inverter_1.Vout 0.25963f
C3016 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout 0.04107f
C3017 a_106699_49858# a_107313_49858# 0.05935f
C3018 RingCounter_0.D_FlipFlop_17.Q' VDD 1.9286f
C3019 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout Nand_Gate_0.B 0.12214f
C3020 Nand_Gate_1.A VDD 4.18085f
C3021 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout a_47119_52572# 0.04444f
C3022 D_FlipFlop_6.Q' a_128237_23350# 0.04443f
C3023 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout 0.1541f
C3024 RingCounter_0.D_FlipFlop_16.Q CLK 0.06351f
C3025 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout VDD 2.8604f
C3026 D_FlipFlop_1.3-input-nand_2.Vout a_132311_33443# 0.04443f
C3027 D_FlipFlop_1.3-input-nand_0.Vout D_FlipFlop_1.3-input-nand_1.Vout 0.03449f
C3028 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C EN 0.07664f
C3029 a_134897_36157# EN 0.04443f
C3030 a_40329_15797# VDD 0.01571f
C3031 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout CLK 0.03574f
C3032 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C RingCounter_0.D_FlipFlop_7.Inverter_1.Vout 0.25579f
C3033 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout 0.08671f
C3034 a_75898_18814# VDD 1.34284f
C3035 a_62539_49858# EN 0.07058f
C3036 Nand_Gate_7.B a_134897_20636# 0.04548f
C3037 RingCounter_0.D_FlipFlop_13.Q' CLK 0.09276f
C3038 Nand_Gate_6.A a_79495_15797# 0.04995f
C3039 D_FlipFlop_7.3-input-nand_0.Vout a_132925_19786# 0.04995f
C3040 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C a_65125_49858# 0.05964f
C3041 a_41687_15797# RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout 0.04443f
C3042 D_FlipFlop_5.Nand_Gate_0.Vout D_FlipFlop_5.Inverter_1.Vout 0.25963f
C3043 D_FlipFlop_5.Q' Q3 0.01194f
C3044 Nand_Gate_0.A D_FlipFlop_2.3-input-nand_2.C 0.14842f
C3045 D_FlipFlop_5.Q' a_128237_26914# 0.04443f
C3046 Nand_Gate_0.A CLK 0.70112f
C3047 a_84619_49858# VDD 0.01712f
C3048 a_75898_18814# CDAC8_0.switch_1.Z 0.28193f
C3049 CDAC8_0.switch_7.Z CLK 5.70593f
C3050 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout 0.30154f
C3051 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout a_79495_13083# 0.01335f
C3052 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_16.Inverter_1.Vout 0.25963f
C3053 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout a_74807_13083# 0.05964f
C3054 Nand_Gate_2.B a_102319_49858# 0.04741f
C3055 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout a_67841_13083# 0.05964f
C3056 D_FlipFlop_5.Q' VDD 1.89808f
C3057 Nand_Gate_5.A CDAC8_0.switch_7.Z 3.15716f
C3058 Nand_Gate_6.B a_134897_24200# 0.04546f
C3059 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout a_62409_13083# 0.04995f
C3060 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout a_55443_13083# 0.04543f
C3061 a_108671_52572# EN 0.045f
C3062 And_Gate_7.Inverter_0.Vin CLK 0.32457f
C3063 Nand_Gate_5.A a_128851_46849# 0.04628f
C3064 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout a_50755_13083# 0.04444f
C3065 RingCounter_0.D_FlipFlop_16.Q Comparator_0.Vinm 0.02272f
C3066 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout 0.04109f
C3067 a_132925_17072# VDD 0.01186f
C3068 RingCounter_0.D_FlipFlop_4.Q' a_90665_49858# 0.01335f
C3069 D_FlipFlop_0.Nand_Gate_0.Vout D_FlipFlop_0.3-input-nand_2.Vout 0.16429f
C3070 Nand_Gate_6.Vout a_92725_16975# 0.04995f
C3071 a_75898_46095# Q4 0.57423f
C3072 RingCounter_0.D_FlipFlop_12.Q' RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout 0.06632f
C3073 a_79625_52572# VDD 0.01186f
C3074 And_Gate_5.Inverter_0.Vin EN 0.0623f
C3075 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C a_56187_49858# 0.04443f
C3076 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout 0.0846f
C3077 Nand_Gate_7.A a_61795_15797# 0.06113f
C3078 a_33363_13083# VDD 0.05686f
C3079 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout VDD 2.73332f
C3080 D_FlipFlop_2.Nand_Gate_0.Vout D_FlipFlop_2.3-input-nand_2.Vout 0.16429f
C3081 VDD Q0 4.32026f
C3082 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout CLK 0.71041f
C3083 a_84619_49858# a_85233_49858# 0.05935f
C3084 a_115177_47663# VDD 0.03918f
C3085 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout CLK 0.28375f
C3086 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout 0.08671f
C3087 EN Q3 0.2481f
C3088 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout a_67841_13083# 0.04443f
C3089 Nand_Gate_6.B RingCounter_0.D_FlipFlop_11.Q' 1.05791f
C3090 Nand_Gate_0.A Comparator_0.Vinm 4.9842f
C3091 a_70645_16975# CLK 0.04479f
C3092 a_132311_37007# a_132925_37007# 0.05935f
C3093 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout a_86591_49858# 0.04543f
C3094 D_FlipFlop_6.Inverter_1.Vout D_FlipFlop_6.3-input-nand_2.Vout 0.06445f
C3095 CDAC8_0.switch_7.Z Comparator_0.Vinm 0.90965p
C3096 CDAC8_0.switch_1.Z Q0 0.17234f
C3097 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout VDD 1.86552f
C3098 D_FlipFlop_3.Nand_Gate_0.Vout D_FlipFlop_3.Nand_Gate_1.Vout 0.04109f
C3099 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout CLK 0.155f
C3100 RingCounter_0.D_FlipFlop_3.Q' a_80239_49858# 0.06113f
C3101 a_75898_39392# Q6 0.4968f
C3102 VDD EN 0.14532p
C3103 Nand_Gate_2.A RingCounter_0.D_FlipFlop_5.Inverter_0.Vout 0.29368f
C3104 FFCLR D_FlipFlop_7.3-input-nand_2.Vout 0.06105f
C3105 D_FlipFlop_4.3-input-nand_0.Vout a_134897_30478# 0.01335f
C3106 D_FlipFlop_6.Inverter_0.Vout D_FlipFlop_6.3-input-nand_1.Vout 0.0857f
C3107 a_40459_49858# VDD 0.05707f
C3108 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout EN 0.09127f
C3109 D_FlipFlop_0.Inverter_1.Vout D_FlipFlop_0.Nand_Gate_1.Vout 0.30154f
C3110 a_100961_13083# VDD 0.02865f
C3111 D_FlipFlop_5.Inverter_1.Vout D_FlipFlop_5.3-input-nand_2.Vout 0.06445f
C3112 Q0 Vbias 16.49397f
C3113 Q1 Vbias 20.30872f
C3114 Q2 Vbias 20.09656f
C3115 Vin Vbias 1.33035f
C3116 Q3 Vbias 19.86623f
C3117 Q7 Vbias 22.24283f
C3118 Q6 Vbias 22.23229f
C3119 Q5 Vbias 22.23164f
C3120 Q4 Vbias 22.21854f
C3121 CLK Vbias 0.15632p
C3122 EN Vbias 0.19957p
C3123 VDD Vbias 1.9306p
C3124 m3_125329_49141# Vbias 0.68315f $ **FLOATING
C3125 a_123655_13083# Vbias 0.43953f
C3126 a_123041_13083# Vbias 0.3792f
C3127 a_121683_13083# Vbias 0.43856f
C3128 a_121069_13083# Vbias 0.3792f
C3129 a_118967_13083# Vbias 0.43856f
C3130 a_117609_13083# Vbias 0.43856f
C3131 a_116995_13083# Vbias 0.37919f
C3132 a_112615_13083# Vbias 0.43953f
C3133 a_112001_13083# Vbias 0.3792f
C3134 a_110643_13083# Vbias 0.43856f
C3135 a_110029_13083# Vbias 0.3792f
C3136 a_107927_13083# Vbias 0.43856f
C3137 a_106569_13083# Vbias 0.43856f
C3138 a_105955_13083# Vbias 0.37919f
C3139 a_101575_13083# Vbias 0.43953f
C3140 a_100961_13083# Vbias 0.3792f
C3141 a_99603_13083# Vbias 0.43856f
C3142 a_98989_13083# Vbias 0.3792f
C3143 a_96887_13083# Vbias 0.43856f
C3144 a_95529_13083# Vbias 0.43856f
C3145 a_94915_13083# Vbias 0.37919f
C3146 a_90535_13083# Vbias 0.43953f
C3147 a_89921_13083# Vbias 0.3792f
C3148 a_88563_13083# Vbias 0.43856f
C3149 a_87949_13083# Vbias 0.3792f
C3150 a_85847_13083# Vbias 0.43856f
C3151 a_84489_13083# Vbias 0.43856f
C3152 a_83875_13083# Vbias 0.37919f
C3153 a_79495_13083# Vbias 0.43953f
C3154 a_78881_13083# Vbias 0.3792f
C3155 a_77523_13083# Vbias 0.43856f
C3156 a_76909_13083# Vbias 0.3792f
C3157 a_74807_13083# Vbias 0.43856f
C3158 a_73449_13083# Vbias 0.43856f
C3159 a_72835_13083# Vbias 0.37919f
C3160 a_68455_13083# Vbias 0.43953f
C3161 a_67841_13083# Vbias 0.3792f
C3162 a_66483_13083# Vbias 0.43856f
C3163 a_65869_13083# Vbias 0.3792f
C3164 a_63767_13083# Vbias 0.43856f
C3165 a_62409_13083# Vbias 0.43856f
C3166 a_61795_13083# Vbias 0.37919f
C3167 a_57415_13083# Vbias 0.43953f
C3168 a_56801_13083# Vbias 0.3792f
C3169 a_55443_13083# Vbias 0.43856f
C3170 a_54829_13083# Vbias 0.3792f
C3171 a_52727_13083# Vbias 0.43856f
C3172 a_51369_13083# Vbias 0.43856f
C3173 a_50755_13083# Vbias 0.37919f
C3174 a_46375_13083# Vbias 0.43953f
C3175 a_45761_13083# Vbias 0.3792f
C3176 a_44403_13083# Vbias 0.43856f
C3177 a_43789_13083# Vbias 0.3792f
C3178 a_41687_13083# Vbias 0.43856f
C3179 a_40329_13083# Vbias 0.43856f
C3180 a_39715_13083# Vbias 0.37919f
C3181 a_35335_13083# Vbias 0.43953f
C3182 a_34721_13083# Vbias 0.3792f
C3183 a_33363_13083# Vbias 0.43856f
C3184 a_32749_13083# Vbias 0.3792f
C3185 a_30647_13083# Vbias 0.43856f
C3186 a_29289_13083# Vbias 0.43856f
C3187 a_28675_13083# Vbias 0.37919f
C3188 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout Vbias 1.05086f
C3189 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout Vbias 1.23023f
C3190 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout Vbias 1.05086f
C3191 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout Vbias 1.23023f
C3192 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout Vbias 1.05086f
C3193 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout Vbias 1.23023f
C3194 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout Vbias 1.05086f
C3195 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout Vbias 1.23023f
C3196 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout Vbias 1.05086f
C3197 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout Vbias 1.23023f
C3198 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout Vbias 1.05086f
C3199 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout Vbias 1.23023f
C3200 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout Vbias 1.05086f
C3201 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout Vbias 1.23023f
C3202 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout Vbias 1.05086f
C3203 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout Vbias 1.23023f
C3204 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout Vbias 1.05086f
C3205 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout Vbias 1.23023f
C3206 RingCounter_0.D_FlipFlop_10.Inverter_0.Vout Vbias 1.95482f
C3207 a_123655_15797# Vbias 0.43953f
C3208 a_123041_15797# Vbias 0.3792f
C3209 a_121683_15797# Vbias 0.43856f
C3210 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout Vbias 1.14622f
C3211 a_121069_15797# Vbias 0.37919f
C3212 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C Vbias 1.9637f
C3213 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout Vbias 2.17382f
C3214 a_118967_15797# Vbias 0.43856f
C3215 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout Vbias 2.19874f
C3216 a_117609_15797# Vbias 0.43856f
C3217 RingCounter_0.D_FlipFlop_10.Nand_Gate_0.Vout Vbias 1.56071f
C3218 a_116995_15797# Vbias 0.37919f
C3219 RingCounter_0.D_FlipFlop_10.Q' Vbias 1.71102f
C3220 RingCounter_0.D_FlipFlop_9.Inverter_0.Vout Vbias 1.95464f
C3221 a_112615_15797# Vbias 0.43953f
C3222 a_112001_15797# Vbias 0.3792f
C3223 a_110643_15797# Vbias 0.43856f
C3224 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout Vbias 1.11152f
C3225 a_110029_15797# Vbias 0.37919f
C3226 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C Vbias 1.96419f
C3227 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout Vbias 2.17422f
C3228 a_107927_15797# Vbias 0.43856f
C3229 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout Vbias 2.19923f
C3230 a_106569_15797# Vbias 0.43856f
C3231 RingCounter_0.D_FlipFlop_9.Nand_Gate_0.Vout Vbias 1.5612f
C3232 a_105955_15797# Vbias 0.37919f
C3233 RingCounter_0.D_FlipFlop_9.Q' Vbias 1.71151f
C3234 RingCounter_0.D_FlipFlop_11.Inverter_0.Vout Vbias 1.95464f
C3235 a_101575_15797# Vbias 0.43953f
C3236 a_100961_15797# Vbias 0.3792f
C3237 a_99603_15797# Vbias 0.43856f
C3238 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout Vbias 1.11152f
C3239 a_98989_15797# Vbias 0.37919f
C3240 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C Vbias 1.96419f
C3241 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout Vbias 2.17422f
C3242 a_96887_15797# Vbias 0.43856f
C3243 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout Vbias 2.19923f
C3244 a_95529_15797# Vbias 0.43856f
C3245 RingCounter_0.D_FlipFlop_11.Nand_Gate_0.Vout Vbias 1.5612f
C3246 a_94915_15797# Vbias 0.37919f
C3247 RingCounter_0.D_FlipFlop_11.Q' Vbias 1.71151f
C3248 RingCounter_0.D_FlipFlop_12.Inverter_0.Vout Vbias 1.95464f
C3249 a_90535_15797# Vbias 0.43953f
C3250 a_89921_15797# Vbias 0.3792f
C3251 a_88563_15797# Vbias 0.43856f
C3252 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout Vbias 1.11152f
C3253 a_87949_15797# Vbias 0.37919f
C3254 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C Vbias 1.96419f
C3255 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout Vbias 2.17422f
C3256 a_85847_15797# Vbias 0.43856f
C3257 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout Vbias 2.19923f
C3258 a_84489_15797# Vbias 0.43856f
C3259 RingCounter_0.D_FlipFlop_12.Nand_Gate_0.Vout Vbias 1.5612f
C3260 a_83875_15797# Vbias 0.37919f
C3261 RingCounter_0.D_FlipFlop_12.Q' Vbias 1.71151f
C3262 RingCounter_0.D_FlipFlop_13.Inverter_0.Vout Vbias 1.95464f
C3263 a_79495_15797# Vbias 0.43953f
C3264 a_78881_15797# Vbias 0.3792f
C3265 a_77523_15797# Vbias 0.4389f
C3266 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout Vbias 1.11158f
C3267 a_76909_15797# Vbias 0.37919f
C3268 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C Vbias 1.96419f
C3269 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout Vbias 2.17422f
C3270 a_74807_15797# Vbias 0.43856f
C3271 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout Vbias 2.19923f
C3272 a_73449_15797# Vbias 0.43856f
C3273 RingCounter_0.D_FlipFlop_13.Nand_Gate_0.Vout Vbias 1.5612f
C3274 a_72835_15797# Vbias 0.37919f
C3275 RingCounter_0.D_FlipFlop_13.Q' Vbias 1.71151f
C3276 RingCounter_0.D_FlipFlop_14.Inverter_0.Vout Vbias 1.95464f
C3277 a_68455_15797# Vbias 0.43953f
C3278 a_67841_15797# Vbias 0.3792f
C3279 a_66483_15797# Vbias 0.43856f
C3280 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout Vbias 1.11152f
C3281 a_65869_15797# Vbias 0.37919f
C3282 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C Vbias 1.96419f
C3283 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout Vbias 2.17422f
C3284 a_63767_15797# Vbias 0.43856f
C3285 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout Vbias 2.19923f
C3286 a_62409_15797# Vbias 0.43856f
C3287 RingCounter_0.D_FlipFlop_14.Nand_Gate_0.Vout Vbias 1.5612f
C3288 a_61795_15797# Vbias 0.37919f
C3289 RingCounter_0.D_FlipFlop_14.Q' Vbias 1.71151f
C3290 RingCounter_0.D_FlipFlop_15.Inverter_0.Vout Vbias 1.95464f
C3291 a_57415_15797# Vbias 0.43953f
C3292 a_56801_15797# Vbias 0.3792f
C3293 a_55443_15797# Vbias 0.43856f
C3294 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout Vbias 1.11152f
C3295 a_54829_15797# Vbias 0.37919f
C3296 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C Vbias 1.96419f
C3297 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout Vbias 2.17422f
C3298 a_52727_15797# Vbias 0.43856f
C3299 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout Vbias 2.19923f
C3300 a_51369_15797# Vbias 0.43856f
C3301 RingCounter_0.D_FlipFlop_15.Nand_Gate_0.Vout Vbias 1.5612f
C3302 a_50755_15797# Vbias 0.37919f
C3303 RingCounter_0.D_FlipFlop_15.Q' Vbias 1.71151f
C3304 RingCounter_0.D_FlipFlop_8.Inverter_0.Vout Vbias 1.95464f
C3305 a_46375_15797# Vbias 0.43953f
C3306 a_45761_15797# Vbias 0.3792f
C3307 a_44403_15797# Vbias 0.43856f
C3308 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout Vbias 1.11152f
C3309 a_43789_15797# Vbias 0.37919f
C3310 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C Vbias 1.96419f
C3311 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout Vbias 2.17422f
C3312 a_41687_15797# Vbias 0.43856f
C3313 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout Vbias 2.19923f
C3314 a_40329_15797# Vbias 0.43856f
C3315 RingCounter_0.D_FlipFlop_8.Nand_Gate_0.Vout Vbias 1.5612f
C3316 a_39715_15797# Vbias 0.37919f
C3317 RingCounter_0.D_FlipFlop_8.Q' Vbias 1.71151f
C3318 RingCounter_0.D_FlipFlop_16.Inverter_0.Vout Vbias 1.95464f
C3319 a_35335_15797# Vbias 0.43953f
C3320 a_34721_15797# Vbias 0.3792f
C3321 a_33363_15797# Vbias 0.43856f
C3322 RingCounter_0.D_FlipFlop_16.3-input-nand_0.Vout Vbias 1.5861f
C3323 a_32749_15797# Vbias 0.37919f
C3324 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C Vbias 1.98054f
C3325 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout Vbias 2.17384f
C3326 a_30647_15797# Vbias 0.43856f
C3327 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout Vbias 2.19883f
C3328 a_29289_15797# Vbias 0.43856f
C3329 RingCounter_0.D_FlipFlop_16.Nand_Gate_0.Vout Vbias 1.60955f
C3330 a_28675_15797# Vbias 0.37919f
C3331 RingCounter_0.D_FlipFlop_16.Q' Vbias 1.71125f
C3332 a_138318_16817# Vbias 10.4148f
C3333 a_134897_17072# Vbias 0.43953f
C3334 a_134283_17072# Vbias 0.3792f
C3335 a_132925_17072# Vbias 0.43856f
C3336 a_132311_17072# Vbias 0.3792f
C3337 a_130209_17072# Vbias 0.43856f
C3338 a_128851_17072# Vbias 0.43856f
C3339 a_128237_17072# Vbias 0.37919f
C3340 a_114805_16975# Vbias 0.47806f
C3341 a_104137_16975# Vbias 0.43856f
C3342 a_92725_16975# Vbias 0.43856f
C3343 a_82057_16975# Vbias 0.43856f
C3344 a_70645_16975# Vbias 0.43856f
C3345 a_59977_16975# Vbias 0.43856f
C3346 a_48565_16975# Vbias 0.43856f
C3347 a_37897_16975# Vbias 0.43856f
C3348 D_FlipFlop_7.3-input-nand_1.Vout Vbias 1.5225f
C3349 D_FlipFlop_7.Nand_Gate_1.Vout Vbias 1.63772f
C3350 And_Gate_3.Inverter_0.Vin Vbias 1.69781f
C3351 Nand_Gate_1.Vout Vbias 2.308f
C3352 Nand_Gate_1.A Vbias 6.47266f
C3353 And_Gate_2.Inverter_0.Vin Vbias 1.64253f
C3354 Nand_Gate_6.Vout Vbias 2.25417f
C3355 Nand_Gate_6.A Vbias 6.47266f
C3356 And_Gate_0.Inverter_0.Vin Vbias 1.70239f
C3357 Nand_Gate_7.A Vbias 6.5083f
C3358 And_Gate_1.Inverter_0.Vin Vbias 1.70234f
C3359 Nand_Gate_4.A Vbias 6.50322f
C3360 D_FlipFlop_7.Inverter_0.Vout Vbias 1.94621f
C3361 a_134897_19786# Vbias 0.43917f
C3362 a_134283_19786# Vbias 0.3792f
C3363 a_132925_19786# Vbias 0.43856f
C3364 D_FlipFlop_7.3-input-nand_0.Vout Vbias 1.58878f
C3365 a_132311_19786# Vbias 0.37919f
C3366 D_FlipFlop_7.3-input-nand_2.C Vbias 2.14024f
C3367 D_FlipFlop_7.3-input-nand_2.Vout Vbias 2.18913f
C3368 a_130209_19786# Vbias 0.43856f
C3369 D_FlipFlop_7.Inverter_1.Vout Vbias 2.76312f
C3370 Nand_Gate_4.B Vbias 17.14899f
C3371 a_128851_19786# Vbias 0.43856f
C3372 D_FlipFlop_7.Nand_Gate_0.Vout Vbias 1.62586f
C3373 a_128237_19786# Vbias 0.37919f
C3374 D_FlipFlop_7.Q' Vbias 1.69494f
C3375 CDAC8_0.switch_1.Z Vbias 2.69005f
C3376 a_75898_18814# Vbias 2.05996f
C3377 a_134897_20636# Vbias 0.43917f
C3378 a_134283_20636# Vbias 0.3792f
C3379 a_132925_20636# Vbias 0.43856f
C3380 a_132311_20636# Vbias 0.3792f
C3381 a_130209_20636# Vbias 0.43856f
C3382 a_128851_20636# Vbias 0.43856f
C3383 a_128237_20636# Vbias 0.37919f
C3384 D_FlipFlop_6.3-input-nand_1.Vout Vbias 1.513f
C3385 D_FlipFlop_6.Nand_Gate_1.Vout Vbias 1.61501f
C3386 CDAC8_0.switch_2.Z Vbias 4.87994f
C3387 a_75898_21528# Vbias 2.07315f
C3388 D_FlipFlop_6.Inverter_0.Vout Vbias 1.92077f
C3389 a_134897_23350# Vbias 0.43917f
C3390 a_134283_23350# Vbias 0.3792f
C3391 a_132925_23350# Vbias 0.43856f
C3392 D_FlipFlop_6.3-input-nand_0.Vout Vbias 1.58878f
C3393 a_132311_23350# Vbias 0.37919f
C3394 D_FlipFlop_6.3-input-nand_2.C Vbias 2.13068f
C3395 D_FlipFlop_6.3-input-nand_2.Vout Vbias 2.1796f
C3396 a_130209_23350# Vbias 0.43856f
C3397 D_FlipFlop_6.Inverter_1.Vout Vbias 2.74117f
C3398 Nand_Gate_7.B Vbias 15.5696f
C3399 a_128851_23350# Vbias 0.43856f
C3400 D_FlipFlop_6.Nand_Gate_0.Vout Vbias 1.62586f
C3401 a_128237_23350# Vbias 0.37919f
C3402 D_FlipFlop_6.Q' Vbias 1.69798f
C3403 a_134897_24200# Vbias 0.43917f
C3404 a_134283_24200# Vbias 0.3792f
C3405 a_132925_24200# Vbias 0.43856f
C3406 a_132311_24200# Vbias 0.3792f
C3407 a_130209_24200# Vbias 0.43856f
C3408 a_128851_24200# Vbias 0.43856f
C3409 a_128237_24200# Vbias 0.37919f
C3410 D_FlipFlop_5.3-input-nand_1.Vout Vbias 1.513f
C3411 D_FlipFlop_5.Nand_Gate_1.Vout Vbias 1.61501f
C3412 CDAC8_0.switch_0.Z Vbias 8.90899f
C3413 a_75898_25104# Vbias 2.10689f
C3414 D_FlipFlop_5.Inverter_0.Vout Vbias 1.92059f
C3415 a_134897_26914# Vbias 0.43917f
C3416 a_134283_26914# Vbias 0.3792f
C3417 a_132925_26914# Vbias 0.43856f
C3418 D_FlipFlop_5.3-input-nand_0.Vout Vbias 1.58878f
C3419 a_132311_26914# Vbias 0.37919f
C3420 D_FlipFlop_5.3-input-nand_2.C Vbias 2.13068f
C3421 D_FlipFlop_5.3-input-nand_2.Vout Vbias 2.1796f
C3422 a_130209_26914# Vbias 0.43856f
C3423 D_FlipFlop_5.Inverter_1.Vout Vbias 2.74117f
C3424 Nand_Gate_6.B Vbias 16.04721f
C3425 a_128851_26914# Vbias 0.43856f
C3426 D_FlipFlop_5.Nand_Gate_0.Vout Vbias 1.62586f
C3427 a_128237_26914# Vbias 0.37919f
C3428 D_FlipFlop_5.Q' Vbias 1.69798f
C3429 Comparator_0.Vinm Vbias 0.48532p
C3430 a_139696_27690# Vbias 8.75751f
C3431 a_134897_27764# Vbias 0.43917f
C3432 a_134283_27764# Vbias 0.3792f
C3433 a_132925_27764# Vbias 0.43856f
C3434 a_132311_27764# Vbias 0.3792f
C3435 a_130209_27764# Vbias 0.43856f
C3436 a_128851_27764# Vbias 0.43856f
C3437 a_128237_27764# Vbias 0.37919f
C3438 D_FlipFlop_4.3-input-nand_1.Vout Vbias 1.513f
C3439 D_FlipFlop_4.Nand_Gate_1.Vout Vbias 1.61501f
C3440 CDAC8_0.switch_5.Z Vbias 16.42038f
C3441 a_75898_28676# Vbias 2.1069f
C3442 D_FlipFlop_4.Inverter_0.Vout Vbias 1.92082f
C3443 a_134897_30478# Vbias 0.43917f
C3444 a_134283_30478# Vbias 0.3792f
C3445 a_132925_30478# Vbias 0.43856f
C3446 D_FlipFlop_4.3-input-nand_0.Vout Vbias 1.66474f
C3447 a_132311_30478# Vbias 0.37919f
C3448 D_FlipFlop_4.3-input-nand_2.C Vbias 2.14021f
C3449 D_FlipFlop_4.3-input-nand_2.Vout Vbias 2.18874f
C3450 a_130209_30478# Vbias 0.43856f
C3451 D_FlipFlop_4.Inverter_1.Vout Vbias 2.7507f
C3452 Nand_Gate_1.B Vbias 18.0878f
C3453 a_128851_30478# Vbias 0.43856f
C3454 D_FlipFlop_4.Nand_Gate_0.Vout Vbias 1.64856f
C3455 a_128237_30478# Vbias 0.37919f
C3456 D_FlipFlop_4.Q' Vbias 1.70751f
C3457 a_134897_33443# Vbias 0.43917f
C3458 a_134283_33443# Vbias 0.3792f
C3459 a_132925_33443# Vbias 0.43856f
C3460 a_132311_33443# Vbias 0.3792f
C3461 a_130209_33443# Vbias 0.43856f
C3462 a_128851_33443# Vbias 0.43856f
C3463 a_128237_33443# Vbias 0.37919f
C3464 D_FlipFlop_1.3-input-nand_1.Vout Vbias 1.5225f
C3465 D_FlipFlop_1.Nand_Gate_1.Vout Vbias 1.63772f
C3466 D_FlipFlop_1.Inverter_0.Vout Vbias 1.93118f
C3467 a_134897_36157# Vbias 0.43917f
C3468 a_134283_36157# Vbias 0.3792f
C3469 a_132925_36157# Vbias 0.43856f
C3470 D_FlipFlop_1.3-input-nand_0.Vout Vbias 1.59129f
C3471 a_132311_36157# Vbias 0.37919f
C3472 D_FlipFlop_1.3-input-nand_2.C Vbias 2.14024f
C3473 D_FlipFlop_1.3-input-nand_2.Vout Vbias 2.18913f
C3474 a_130209_36157# Vbias 0.43856f
C3475 D_FlipFlop_1.Inverter_1.Vout Vbias 2.76312f
C3476 a_128851_36157# Vbias 0.43856f
C3477 D_FlipFlop_1.Nand_Gate_0.Vout Vbias 1.62586f
C3478 a_128237_36157# Vbias 0.37919f
C3479 D_FlipFlop_1.Q' Vbias 1.7018f
C3480 CDAC8_0.switch_7.Z Vbias 0.26689p
C3481 a_75898_35820# Vbias 2.11281f
C3482 a_134897_37007# Vbias 0.43917f
C3483 a_134283_37007# Vbias 0.3792f
C3484 a_132925_37007# Vbias 0.43856f
C3485 a_132311_37007# Vbias 0.3792f
C3486 a_130209_37007# Vbias 0.43856f
C3487 a_128851_37007# Vbias 0.43856f
C3488 a_128237_37007# Vbias 0.37919f
C3489 D_FlipFlop_2.3-input-nand_1.Vout Vbias 1.513f
C3490 D_FlipFlop_2.Nand_Gate_1.Vout Vbias 1.61501f
C3491 D_FlipFlop_2.Inverter_0.Vout Vbias 1.92088f
C3492 a_134897_39721# Vbias 0.43917f
C3493 a_134283_39721# Vbias 0.3792f
C3494 a_132925_39721# Vbias 0.43856f
C3495 D_FlipFlop_2.3-input-nand_0.Vout Vbias 1.58878f
C3496 a_132311_39721# Vbias 0.37919f
C3497 D_FlipFlop_2.3-input-nand_2.C Vbias 2.13068f
C3498 D_FlipFlop_2.3-input-nand_2.Vout Vbias 2.1796f
C3499 a_130209_39721# Vbias 0.43856f
C3500 D_FlipFlop_2.Inverter_1.Vout Vbias 2.74117f
C3501 a_128851_39721# Vbias 0.43856f
C3502 D_FlipFlop_2.Nand_Gate_0.Vout Vbias 1.62586f
C3503 a_128237_39721# Vbias 0.37919f
C3504 D_FlipFlop_2.Q' Vbias 1.69798f
C3505 CDAC8_0.switch_6.Z Vbias 0.12229p
C3506 a_75898_39392# Vbias 2.11281f
C3507 a_134897_40571# Vbias 0.43917f
C3508 a_134283_40571# Vbias 0.3792f
C3509 a_132925_40571# Vbias 0.43856f
C3510 a_132311_40571# Vbias 0.3792f
C3511 a_130209_40571# Vbias 0.43856f
C3512 a_128851_40571# Vbias 0.43856f
C3513 a_128237_40571# Vbias 0.37919f
C3514 D_FlipFlop_3.3-input-nand_1.Vout Vbias 1.513f
C3515 D_FlipFlop_3.Nand_Gate_1.Vout Vbias 1.61501f
C3516 D_FlipFlop_3.Inverter_0.Vout Vbias 1.92078f
C3517 a_134897_43285# Vbias 0.43917f
C3518 a_134283_43285# Vbias 0.3792f
C3519 a_132925_43285# Vbias 0.43856f
C3520 D_FlipFlop_3.3-input-nand_0.Vout Vbias 1.58878f
C3521 a_132311_43285# Vbias 0.37919f
C3522 D_FlipFlop_3.3-input-nand_2.C Vbias 2.13068f
C3523 D_FlipFlop_3.3-input-nand_2.Vout Vbias 2.1796f
C3524 a_130209_43285# Vbias 0.43856f
C3525 D_FlipFlop_3.Inverter_1.Vout Vbias 2.74117f
C3526 a_128851_43285# Vbias 0.43856f
C3527 D_FlipFlop_3.Nand_Gate_0.Vout Vbias 1.62586f
C3528 a_128237_43285# Vbias 0.37919f
C3529 D_FlipFlop_3.Q' Vbias 1.69798f
C3530 CDAC8_0.switch_9.Z Vbias 56.99755f
C3531 a_75898_42964# Vbias 2.11275f
C3532 a_134897_44135# Vbias 0.43917f
C3533 a_134283_44135# Vbias 0.3792f
C3534 a_132925_44135# Vbias 0.43856f
C3535 a_132311_44135# Vbias 0.3792f
C3536 a_130209_44135# Vbias 0.43856f
C3537 a_128851_44135# Vbias 0.43856f
C3538 a_128237_44135# Vbias 0.37919f
C3539 D_FlipFlop_0.3-input-nand_1.Vout Vbias 1.513f
C3540 D_FlipFlop_0.Nand_Gate_1.Vout Vbias 1.61501f
C3541 D_FlipFlop_0.Inverter_0.Vout Vbias 1.92075f
C3542 a_134897_46849# Vbias 0.43953f
C3543 a_134283_46849# Vbias 0.3792f
C3544 a_132925_46849# Vbias 0.43856f
C3545 D_FlipFlop_0.3-input-nand_0.Vout Vbias 1.66474f
C3546 a_132311_46849# Vbias 0.37919f
C3547 D_FlipFlop_0.3-input-nand_2.C Vbias 2.14021f
C3548 D_FlipFlop_0.3-input-nand_2.Vout Vbias 2.18874f
C3549 a_130209_46849# Vbias 0.43856f
C3550 D_FlipFlop_0.Inverter_1.Vout Vbias 2.7507f
C3551 a_128851_46849# Vbias 0.43856f
C3552 D_FlipFlop_0.Nand_Gate_0.Vout Vbias 1.64856f
C3553 CDAC8_0.switch_8.Z Vbias 30.17742f
C3554 a_75898_46095# Vbias 2.10708f
C3555 a_128237_46849# Vbias 0.37919f
C3556 D_FlipFlop_0.Q' Vbias 1.70751f
C3557 a_125845_47663# Vbias 0.43856f
C3558 a_115177_47663# Vbias 0.44123f
C3559 a_103765_47663# Vbias 0.43856f
C3560 a_93097_47663# Vbias 0.43856f
C3561 a_81685_47663# Vbias 0.43856f
C3562 a_71017_47663# Vbias 0.43856f
C3563 a_59605_47663# Vbias 0.43856f
C3564 a_48937_47663# Vbias 0.43856f
C3565 And_Gate_7.Inverter_0.Vin Vbias 1.72676f
C3566 Nand_Gate_5.Vout Vbias 2.54583f
C3567 And_Gate_6.Inverter_0.Vin Vbias 1.65848f
C3568 Nand_Gate_2.Vout Vbias 2.37367f
C3569 And_Gate_4.Inverter_0.Vin Vbias 1.65848f
C3570 And_Gate_5.Inverter_0.Vin Vbias 1.69344f
C3571 a_124399_49858# Vbias 0.37919f
C3572 a_123785_49858# Vbias 0.43856f
C3573 a_122427_49858# Vbias 0.43856f
C3574 a_120325_49858# Vbias 0.3792f
C3575 a_119711_49858# Vbias 0.43856f
C3576 a_118353_49858# Vbias 0.3792f
C3577 a_117739_49858# Vbias 0.43953f
C3578 a_113359_49858# Vbias 0.37919f
C3579 a_112745_49858# Vbias 0.43856f
C3580 a_111387_49858# Vbias 0.43856f
C3581 a_109285_49858# Vbias 0.3792f
C3582 a_108671_49858# Vbias 0.43856f
C3583 a_107313_49858# Vbias 0.3792f
C3584 a_106699_49858# Vbias 0.43953f
C3585 a_102319_49858# Vbias 0.37919f
C3586 a_101705_49858# Vbias 0.43856f
C3587 a_100347_49858# Vbias 0.43856f
C3588 a_98245_49858# Vbias 0.3792f
C3589 a_97631_49858# Vbias 0.43856f
C3590 a_96273_49858# Vbias 0.3792f
C3591 a_95659_49858# Vbias 0.43953f
C3592 a_91279_49858# Vbias 0.37919f
C3593 a_90665_49858# Vbias 0.43856f
C3594 a_89307_49858# Vbias 0.43856f
C3595 a_87205_49858# Vbias 0.3792f
C3596 a_86591_49858# Vbias 0.43856f
C3597 a_85233_49858# Vbias 0.3792f
C3598 a_84619_49858# Vbias 0.43953f
C3599 a_80239_49858# Vbias 0.37919f
C3600 a_79625_49858# Vbias 0.43856f
C3601 a_78267_49858# Vbias 0.43856f
C3602 a_76165_49858# Vbias 0.3792f
C3603 a_75551_49858# Vbias 0.43856f
C3604 a_74193_49858# Vbias 0.3792f
C3605 a_73579_49858# Vbias 0.43953f
C3606 a_69199_49858# Vbias 0.37919f
C3607 a_68585_49858# Vbias 0.43856f
C3608 a_67227_49858# Vbias 0.43856f
C3609 a_65125_49858# Vbias 0.3792f
C3610 a_64511_49858# Vbias 0.43856f
C3611 a_63153_49858# Vbias 0.3792f
C3612 a_62539_49858# Vbias 0.43953f
C3613 a_58159_49858# Vbias 0.37919f
C3614 a_57545_49858# Vbias 0.43856f
C3615 a_56187_49858# Vbias 0.43856f
C3616 a_54085_49858# Vbias 0.3792f
C3617 a_53471_49858# Vbias 0.43856f
C3618 a_52113_49858# Vbias 0.3792f
C3619 a_51499_49858# Vbias 0.43953f
C3620 a_47119_49858# Vbias 0.37919f
C3621 a_46505_49858# Vbias 0.43856f
C3622 a_45147_49858# Vbias 0.43856f
C3623 a_43045_49858# Vbias 0.3792f
C3624 a_42431_49858# Vbias 0.43856f
C3625 a_41073_49858# Vbias 0.3792f
C3626 a_40459_49858# Vbias 0.43953f
C3627 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout Vbias 1.33211f
C3628 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout Vbias 1.17113f
C3629 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout Vbias 1.23794f
C3630 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout Vbias 1.17113f
C3631 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout Vbias 1.23794f
C3632 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout Vbias 1.17113f
C3633 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout Vbias 1.23794f
C3634 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout Vbias 1.17113f
C3635 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout Vbias 1.23794f
C3636 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout Vbias 1.17113f
C3637 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout Vbias 1.23794f
C3638 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout Vbias 1.17113f
C3639 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout Vbias 1.23794f
C3640 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout Vbias 1.17113f
C3641 RingCounter_0.D_FlipFlop_17.Nand_Gate_1.Vout Vbias 1.55597f
C3642 RingCounter_0.D_FlipFlop_17.3-input-nand_1.Vout Vbias 1.5225f
C3643 Nand_Gate_5.B Vbias 21.21678f
C3644 RingCounter_0.D_FlipFlop_6.Q' Vbias 1.69086f
C3645 a_124399_52572# Vbias 0.37919f
C3646 a_123785_52572# Vbias 0.43856f
C3647 RingCounter_0.D_FlipFlop_6.Nand_Gate_0.Vout Vbias 1.64856f
C3648 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout Vbias 2.22335f
C3649 a_122427_52572# Vbias 0.43856f
C3650 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout Vbias 2.18869f
C3651 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C Vbias 2.10099f
C3652 a_120325_52572# Vbias 0.37919f
C3653 a_119711_52572# Vbias 0.43856f
C3654 RingCounter_0.D_FlipFlop_6.3-input-nand_0.Vout Vbias 1.66474f
C3655 a_118353_52572# Vbias 0.3792f
C3656 a_117739_52572# Vbias 0.43953f
C3657 RingCounter_0.D_FlipFlop_6.Inverter_0.Vout Vbias 1.85585f
C3658 Nand_Gate_5.A Vbias 14.28068f
C3659 RingCounter_0.D_FlipFlop_7.Q' Vbias 1.66178f
C3660 a_113359_52572# Vbias 0.37919f
C3661 a_112745_52572# Vbias 0.43856f
C3662 RingCounter_0.D_FlipFlop_7.Nand_Gate_0.Vout Vbias 1.64393f
C3663 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout Vbias 2.15263f
C3664 a_111387_52572# Vbias 0.43856f
C3665 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout Vbias 2.18869f
C3666 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C Vbias 2.10089f
C3667 a_109285_52572# Vbias 0.37919f
C3668 a_108671_52572# Vbias 0.43856f
C3669 RingCounter_0.D_FlipFlop_7.3-input-nand_0.Vout Vbias 1.66474f
C3670 a_107313_52572# Vbias 0.3792f
C3671 a_106699_52572# Vbias 0.43953f
C3672 RingCounter_0.D_FlipFlop_7.Inverter_0.Vout Vbias 1.85585f
C3673 Nand_Gate_2.B Vbias 8.32586f
C3674 RingCounter_0.D_FlipFlop_5.Q' Vbias 1.66178f
C3675 a_102319_52572# Vbias 0.37919f
C3676 a_101705_52572# Vbias 0.43856f
C3677 RingCounter_0.D_FlipFlop_5.Nand_Gate_0.Vout Vbias 1.64393f
C3678 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout Vbias 2.15263f
C3679 a_100347_52572# Vbias 0.43856f
C3680 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout Vbias 2.18869f
C3681 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C Vbias 2.10089f
C3682 a_98245_52572# Vbias 0.37919f
C3683 a_97631_52572# Vbias 0.43856f
C3684 RingCounter_0.D_FlipFlop_5.3-input-nand_0.Vout Vbias 1.66474f
C3685 a_96273_52572# Vbias 0.3792f
C3686 a_95659_52572# Vbias 0.43953f
C3687 RingCounter_0.D_FlipFlop_5.Inverter_0.Vout Vbias 1.85585f
C3688 Nand_Gate_2.A Vbias 14.65982f
C3689 RingCounter_0.D_FlipFlop_4.Q' Vbias 1.66178f
C3690 a_91279_52572# Vbias 0.37919f
C3691 a_90665_52572# Vbias 0.43856f
C3692 RingCounter_0.D_FlipFlop_4.Nand_Gate_0.Vout Vbias 1.64393f
C3693 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout Vbias 2.15263f
C3694 a_89307_52572# Vbias 0.43856f
C3695 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout Vbias 2.18869f
C3696 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C Vbias 2.10089f
C3697 a_87205_52572# Vbias 0.37919f
C3698 a_86591_52572# Vbias 0.43856f
C3699 RingCounter_0.D_FlipFlop_4.3-input-nand_0.Vout Vbias 1.66474f
C3700 a_85233_52572# Vbias 0.3792f
C3701 a_84619_52572# Vbias 0.43953f
C3702 RingCounter_0.D_FlipFlop_4.Inverter_0.Vout Vbias 1.85585f
C3703 Nand_Gate_0.B Vbias 8.32586f
C3704 RingCounter_0.D_FlipFlop_3.Q' Vbias 1.66178f
C3705 a_80239_52572# Vbias 0.37919f
C3706 a_79625_52572# Vbias 0.43856f
C3707 RingCounter_0.D_FlipFlop_3.Nand_Gate_0.Vout Vbias 1.64393f
C3708 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout Vbias 2.15263f
C3709 a_78267_52572# Vbias 0.43856f
C3710 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout Vbias 2.18869f
C3711 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C Vbias 2.10089f
C3712 a_76165_52572# Vbias 0.37919f
C3713 a_75551_52572# Vbias 0.43856f
C3714 RingCounter_0.D_FlipFlop_3.3-input-nand_0.Vout Vbias 1.66474f
C3715 a_74193_52572# Vbias 0.3792f
C3716 a_73579_52572# Vbias 0.43953f
C3717 RingCounter_0.D_FlipFlop_3.Inverter_0.Vout Vbias 1.85585f
C3718 Nand_Gate_0.A Vbias 16.40797f
C3719 RingCounter_0.D_FlipFlop_2.Q' Vbias 1.66178f
C3720 a_69199_52572# Vbias 0.37919f
C3721 a_68585_52572# Vbias 0.43856f
C3722 RingCounter_0.D_FlipFlop_2.Nand_Gate_0.Vout Vbias 1.64393f
C3723 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout Vbias 2.15263f
C3724 a_67227_52572# Vbias 0.43856f
C3725 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout Vbias 2.18869f
C3726 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C Vbias 2.10089f
C3727 a_65125_52572# Vbias 0.37919f
C3728 a_64511_52572# Vbias 0.43856f
C3729 RingCounter_0.D_FlipFlop_2.3-input-nand_0.Vout Vbias 1.66474f
C3730 a_63153_52572# Vbias 0.3792f
C3731 a_62539_52572# Vbias 0.43953f
C3732 RingCounter_0.D_FlipFlop_2.Inverter_0.Vout Vbias 1.85585f
C3733 Nand_Gate_3.B Vbias 8.33895f
C3734 RingCounter_0.D_FlipFlop_1.Q' Vbias 1.66178f
C3735 a_58159_52572# Vbias 0.37919f
C3736 a_57545_52572# Vbias 0.43856f
C3737 RingCounter_0.D_FlipFlop_1.Nand_Gate_0.Vout Vbias 1.64393f
C3738 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout Vbias 2.15263f
C3739 a_56187_52572# Vbias 0.43856f
C3740 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout Vbias 2.18869f
C3741 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C Vbias 2.10089f
C3742 a_54085_52572# Vbias 0.37919f
C3743 a_53471_52572# Vbias 0.43856f
C3744 RingCounter_0.D_FlipFlop_1.3-input-nand_0.Vout Vbias 1.66474f
C3745 a_52113_52572# Vbias 0.3792f
C3746 a_51499_52572# Vbias 0.43953f
C3747 RingCounter_0.D_FlipFlop_1.Inverter_0.Vout Vbias 1.85585f
C3748 FFCLR Vbias 34.75264f
C3749 RingCounter_0.D_FlipFlop_17.Q' Vbias 1.66178f
C3750 a_47119_52572# Vbias 0.37919f
C3751 a_46505_52572# Vbias 0.43856f
C3752 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout Vbias 1.10101f
C3753 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout Vbias 2.22697f
C3754 a_45147_52572# Vbias 0.43856f
C3755 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout Vbias 2.02639f
C3756 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C Vbias 2.17854f
C3757 a_43045_52572# Vbias 0.37919f
C3758 a_42431_52572# Vbias 0.43856f
C3759 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout Vbias 1.01307f
C3760 a_41073_52572# Vbias 0.3792f
C3761 a_40459_52572# Vbias 0.43953f
C3762 RingCounter_0.D_FlipFlop_17.Inverter_0.Vout Vbias 1.93442f
C3763 RingCounter_0.D_FlipFlop_16.Q Vbias 24.46742f
C3764 dw_138090_16601# Vbias 0.32071p $ **FLOATING
C3765 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t1 Vbias 0.05958f
C3766 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n0 Vbias 0.0577f
C3767 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n1 Vbias 0.12257f
C3768 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t6 Vbias 0.23742f
C3769 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t4 Vbias 0.45664f
C3770 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n2 Vbias 0.1334f
C3771 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n3 Vbias 0.05705f
C3772 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n4 Vbias 0.10533f
C3773 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n5 Vbias 0.18236f
C3774 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n6 Vbias 0.13574f
C3775 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n7 Vbias 0.06431f
C3776 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t5 Vbias 0.45666f
C3777 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n8 Vbias 0.47347f
C3778 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n9 Vbias 0.05122f
C3779 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n10 Vbias 0.06839f
C3780 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t7 Vbias 0.22727f
C3781 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t0 Vbias 0.06194f
C3782 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n11 Vbias 0.39067f
C3783 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t3 Vbias 0.06323f
C3784 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.t2 Vbias 0.06194f
C3785 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n12 Vbias 0.35224f
C3786 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n13 Vbias 0.11629f
C3787 RingCounter_0.D_FlipFlop_2.3-input-nand_2.C.n14 Vbias 0.16533f
C3788 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t1 Vbias 0.06358f
C3789 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n0 Vbias 0.03611f
C3790 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n1 Vbias 0.06992f
C3791 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t3 Vbias 0.25335f
C3792 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n2 Vbias 0.24817f
C3793 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n3 Vbias 0.05234f
C3794 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t4 Vbias 0.48726f
C3795 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n4 Vbias 0.14234f
C3796 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n5 Vbias 0.03542f
C3797 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n6 Vbias 0.05152f
C3798 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n7 Vbias 0.13202f
C3799 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C3800 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n9 Vbias 0.06862f
C3801 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t0 Vbias 0.06624f
C3802 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.t2 Vbias 0.07883f
C3803 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n10 Vbias 0.39844f
C3804 RingCounter_0.D_FlipFlop_3.Nand_Gate_1.Vout.n11 Vbias 0.20187f
C3805 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t4 Vbias 0.45666f
C3806 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n0 Vbias 0.47347f
C3807 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n1 Vbias 0.05122f
C3808 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n2 Vbias 0.06839f
C3809 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t6 Vbias 0.22727f
C3810 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t1 Vbias 0.06194f
C3811 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n3 Vbias 0.39067f
C3812 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t3 Vbias 0.06323f
C3813 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t2 Vbias 0.06194f
C3814 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n4 Vbias 0.35224f
C3815 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n5 Vbias 0.11629f
C3816 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n6 Vbias 0.16533f
C3817 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n7 Vbias 0.06431f
C3818 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t7 Vbias 0.23742f
C3819 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t5 Vbias 0.45664f
C3820 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n8 Vbias 0.1334f
C3821 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n9 Vbias 0.05705f
C3822 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n10 Vbias 0.10533f
C3823 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n11 Vbias 0.18236f
C3824 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n12 Vbias 0.13574f
C3825 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n13 Vbias 0.12257f
C3826 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.n14 Vbias 0.0577f
C3827 RingCounter_0.D_FlipFlop_5.3-input-nand_2.C.t0 Vbias 0.05958f
C3828 And_Gate_0.B.t1 Vbias 0.07874f
C3829 Nand_Gate_7.Vout Vbias -0.158f
C3830 And_Gate_0.B.n0 Vbias 0.04472f
C3831 And_Gate_0.B.n1 Vbias 0.0866f
C3832 And_Gate_0.B.t3 Vbias 0.31378f
C3833 And_Gate_0.Nand_Gate_0.B Vbias -0.2359f
C3834 And_Gate_0.B.n2 Vbias 0.30737f
C3835 And_Gate_0.B.n3 Vbias 0.06483f
C3836 And_Gate_0.B.t4 Vbias 0.60348f
C3837 And_Gate_0.B.n4 Vbias 0.17629f
C3838 And_Gate_0.B.n5 Vbias 0.04387f
C3839 And_Gate_0.B.n6 Vbias 0.06381f
C3840 And_Gate_0.B.n7 Vbias 1.30112f
C3841 And_Gate_0.B.n8 Vbias 1.30112f
C3842 And_Gate_0.B.n9 Vbias 0.08499f
C3843 And_Gate_0.B.t2 Vbias 0.08204f
C3844 And_Gate_0.B.t0 Vbias 0.09763f
C3845 And_Gate_0.B.n10 Vbias 0.49348f
C3846 And_Gate_0.B.n11 Vbias 0.25003f
C3847 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t3 Vbias 0.05201f
C3848 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n0 Vbias 0.22649f
C3849 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n1 Vbias 0.05616f
C3850 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t4 Vbias 0.39877f
C3851 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n2 Vbias 0.39189f
C3852 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n3 Vbias 0.04283f
C3853 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t5 Vbias 0.20732f
C3854 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n4 Vbias 0.05972f
C3855 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n5 Vbias 0.02559f
C3856 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n6 Vbias 0.04796f
C3857 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n7 Vbias 0.10804f
C3858 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n8 Vbias 0.10804f
C3859 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n9 Vbias 0.06475f
C3860 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t2 Vbias 0.05421f
C3861 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t0 Vbias 0.05522f
C3862 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.t1 Vbias 0.05409f
C3863 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n10 Vbias 0.30759f
C3864 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n11 Vbias 0.17406f
C3865 RingCounter_0.D_FlipFlop_14.3-input-nand_0.Vout.n12 Vbias 0.03715f
C3866 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t2 Vbias 0.07037f
C3867 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n0 Vbias 0.16004f
C3868 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n1 Vbias 0.07725f
C3869 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t5 Vbias 0.2799f
C3870 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n2 Vbias 0.27418f
C3871 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n3 Vbias 0.05783f
C3872 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t4 Vbias 0.53832f
C3873 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n4 Vbias 0.15726f
C3874 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n5 Vbias 0.03913f
C3875 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n6 Vbias 0.05692f
C3876 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n7 Vbias 0.14585f
C3877 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n8 Vbias 0.14585f
C3878 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n9 Vbias 0.07581f
C3879 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t3 Vbias 0.07318f
C3880 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t0 Vbias 0.07454f
C3881 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.t1 Vbias 0.07302f
C3882 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n10 Vbias 0.41525f
C3883 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n11 Vbias 0.23391f
C3884 RingCounter_0.D_FlipFlop_9.3-input-nand_1.Vout.n12 Vbias 0.22303f
C3885 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t2 Vbias 0.05201f
C3886 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n0 Vbias 0.22649f
C3887 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n1 Vbias 0.05616f
C3888 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t4 Vbias 0.39877f
C3889 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n2 Vbias 0.39189f
C3890 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n3 Vbias 0.04283f
C3891 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t5 Vbias 0.20732f
C3892 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n4 Vbias 0.05972f
C3893 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n5 Vbias 0.02559f
C3894 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n6 Vbias 0.04796f
C3895 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n7 Vbias 0.10804f
C3896 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n8 Vbias 0.10804f
C3897 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n9 Vbias 0.06475f
C3898 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t3 Vbias 0.05421f
C3899 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t1 Vbias 0.05522f
C3900 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.t0 Vbias 0.05409f
C3901 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n10 Vbias 0.30759f
C3902 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n11 Vbias 0.17406f
C3903 RingCounter_0.D_FlipFlop_10.3-input-nand_0.Vout.n12 Vbias 0.03715f
C3904 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t2 Vbias 0.07037f
C3905 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n0 Vbias 0.16004f
C3906 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n1 Vbias 0.07725f
C3907 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t5 Vbias 0.2799f
C3908 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n2 Vbias 0.27418f
C3909 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n3 Vbias 0.05783f
C3910 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t4 Vbias 0.53832f
C3911 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n4 Vbias 0.15726f
C3912 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n5 Vbias 0.03913f
C3913 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n6 Vbias 0.05692f
C3914 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n7 Vbias 0.14585f
C3915 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n8 Vbias 0.14585f
C3916 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n9 Vbias 0.07581f
C3917 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t3 Vbias 0.07318f
C3918 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t0 Vbias 0.07454f
C3919 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.t1 Vbias 0.07302f
C3920 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n10 Vbias 0.41525f
C3921 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n11 Vbias 0.23391f
C3922 RingCounter_0.D_FlipFlop_15.3-input-nand_1.Vout.n12 Vbias 0.22303f
C3923 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t2 Vbias 0.07024f
C3924 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n0 Vbias 0.03989f
C3925 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n1 Vbias 0.07725f
C3926 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t5 Vbias 0.2799f
C3927 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n2 Vbias 0.27418f
C3928 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n3 Vbias 0.05783f
C3929 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t4 Vbias 0.53832f
C3930 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n4 Vbias 0.15726f
C3931 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n5 Vbias 0.03913f
C3932 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n6 Vbias 0.05692f
C3933 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n7 Vbias 0.14585f
C3934 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n8 Vbias 0.14585f
C3935 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n9 Vbias 0.07581f
C3936 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t3 Vbias 0.07318f
C3937 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t0 Vbias 0.07454f
C3938 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.t1 Vbias 0.07302f
C3939 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n10 Vbias 0.41525f
C3940 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n11 Vbias 0.23391f
C3941 RingCounter_0.D_FlipFlop_7.3-input-nand_1.Vout.n12 Vbias 0.22303f
C3942 Nand_Gate_0.B.t11 Vbias 0.33127f
C3943 Nand_Gate_0.B.n0 Vbias 0.09677f
C3944 Nand_Gate_0.B.n1 Vbias 0.04199f
C3945 Nand_Gate_0.B.n2 Vbias 0.18462f
C3946 Nand_Gate_0.B.t5 Vbias 0.15408f
C3947 Nand_Gate_0.B.n3 Vbias 0.04834f
C3948 Nand_Gate_0.B.t3 Vbias 0.04321f
C3949 Nand_Gate_0.B.n4 Vbias 0.18816f
C3950 Nand_Gate_0.B.n5 Vbias 0.04665f
C3951 Nand_Gate_0.B.t9 Vbias 0.33129f
C3952 Nand_Gate_0.B.n6 Vbias 0.32557f
C3953 Nand_Gate_0.B.n7 Vbias 0.03558f
C3954 Nand_Gate_0.B.t10 Vbias 0.17224f
C3955 Nand_Gate_0.B.n8 Vbias 0.04961f
C3956 Nand_Gate_0.B.n9 Vbias 0.02126f
C3957 Nand_Gate_0.B.n10 Vbias 0.03984f
C3958 Nand_Gate_0.B.n11 Vbias 0.05014f
C3959 Nand_Gate_0.B.t6 Vbias 0.33129f
C3960 Nand_Gate_0.B.n12 Vbias 0.32557f
C3961 Nand_Gate_0.B.n13 Vbias 0.03558f
C3962 Nand_Gate_0.B.t7 Vbias 0.17224f
C3963 Nand_Gate_0.B.n14 Vbias 0.04961f
C3964 Nand_Gate_0.B.n15 Vbias 0.02126f
C3965 Nand_Gate_0.B.n16 Vbias 0.03984f
C3966 Nand_Gate_0.B.n18 Vbias 0.15033f
C3967 Nand_Gate_0.B.n19 Vbias 0.41862f
C3968 Nand_Gate_0.B.n20 Vbias 0.18785f
C3969 Nand_Gate_0.B.t4 Vbias 0.17224f
C3970 Nand_Gate_0.B.t8 Vbias 0.33127f
C3971 Nand_Gate_0.B.n21 Vbias 0.09677f
C3972 Nand_Gate_0.B.n22 Vbias 0.04139f
C3973 Nand_Gate_0.B.n23 Vbias 0.07641f
C3974 Nand_Gate_0.B.n24 Vbias 0.87221f
C3975 Nand_Gate_0.B.n25 Vbias 1.18609f
C3976 Nand_Gate_0.B.n26 Vbias 0.05328f
C3977 Nand_Gate_0.B.n27 Vbias 0.01961f
C3978 Nand_Gate_0.B.n29 Vbias 0.05379f
C3979 Nand_Gate_0.B.n30 Vbias 0.02717f
C3980 Nand_Gate_0.B.t0 Vbias 0.04587f
C3981 Nand_Gate_0.B.t1 Vbias 0.04493f
C3982 Nand_Gate_0.B.n31 Vbias 0.25554f
C3983 Nand_Gate_0.B.n32 Vbias 0.08338f
C3984 Nand_Gate_0.B.t2 Vbias 0.04493f
C3985 Nand_Gate_0.B.n33 Vbias 0.06922f
C3986 Nand_Gate_0.B.n34 Vbias 0.12256f
C3987 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t1 Vbias 0.0608f
C3988 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C3989 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C3990 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C3991 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C3992 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C3993 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C3994 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C3995 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C3996 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C3997 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C3998 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C3999 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C4000 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t2 Vbias 0.06323f
C4001 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C4002 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C4003 RingCounter_0.D_FlipFlop_12.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C4004 Q0.t6 Vbias 0.14104f
C4005 Q0.n0 Vbias 0.0412f
C4006 Q0.n1 Vbias 0.01788f
C4007 Q0.n2 Vbias 0.0786f
C4008 Q0.t9 Vbias 0.0656f
C4009 Q0.n3 Vbias 0.0176f
C4010 Q0.n4 Vbias 0.04807f
C4011 Q0.t3 Vbias 0.0184f
C4012 Q0.n5 Vbias 0.09022f
C4013 Q0.n6 Vbias 0.02214f
C4014 Q0.t1 Vbias 0.01953f
C4015 Q0.t0 Vbias 0.01913f
C4016 Q0.n7 Vbias 0.10879f
C4017 Q0.n8 Vbias 0.0362f
C4018 Q0.t2 Vbias 0.01913f
C4019 Q0.n9 Vbias 0.02645f
C4020 Q0.n10 Vbias 0.01124f
C4021 Q0.n11 Vbias 6.2933f
C4022 Q0.t7 Vbias 0.07345f
C4023 Q0.t8 Vbias 0.07345f
C4024 Q0.t5 Vbias 0.14141f
C4025 Q0.n12 Vbias 0.11441f
C4026 Q0.n13 Vbias 0.11507f
C4027 Q0.t4 Vbias 0.12571f
C4028 Q0.n14 Vbias 1.44692f
C4029 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t1 Vbias 0.04607f
C4030 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n0 Vbias 0.10477f
C4031 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n1 Vbias 0.05057f
C4032 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t3 Vbias 0.35243f
C4033 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n2 Vbias 0.3654f
C4034 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n3 Vbias 0.03953f
C4035 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n4 Vbias 0.05278f
C4036 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t2 Vbias 0.27708f
C4037 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t5 Vbias 0.27709f
C4038 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n5 Vbias 0.17949f
C4039 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n6 Vbias 0.03786f
C4040 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t4 Vbias 0.35241f
C4041 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n7 Vbias 0.10295f
C4042 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n8 Vbias 0.02562f
C4043 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n9 Vbias 0.03726f
C4044 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n10 Vbias 0.09548f
C4045 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n11 Vbias 0.09548f
C4046 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n12 Vbias 0.04963f
C4047 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.t0 Vbias 0.04792f
C4048 RingCounter_0.D_FlipFlop_11.Inverter_1.Vout.n13 Vbias 0.28399f
C4049 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t1 Vbias 0.04998f
C4050 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n0 Vbias 0.02839f
C4051 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n1 Vbias 0.05497f
C4052 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t3 Vbias 0.38308f
C4053 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n2 Vbias 0.39717f
C4054 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n3 Vbias 0.04297f
C4055 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n4 Vbias 0.05737f
C4056 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t4 Vbias 0.30118f
C4057 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t2 Vbias 0.30119f
C4058 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n5 Vbias 0.1951f
C4059 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n6 Vbias 0.04115f
C4060 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t5 Vbias 0.38306f
C4061 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n7 Vbias 0.1119f
C4062 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n8 Vbias 0.02784f
C4063 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n9 Vbias 0.0405f
C4064 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n10 Vbias 0.10379f
C4065 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n11 Vbias 0.10379f
C4066 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n12 Vbias 0.05395f
C4067 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.t0 Vbias 0.05208f
C4068 RingCounter_0.D_FlipFlop_4.Inverter_1.Vout.n13 Vbias 0.30868f
C4069 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t6 Vbias 0.36784f
C4070 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n0 Vbias 0.10746f
C4071 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n1 Vbias 0.04662f
C4072 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t3 Vbias 0.04798f
C4073 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n2 Vbias 0.22815f
C4074 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n3 Vbias 0.0518f
C4075 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t5 Vbias 0.36785f
C4076 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n4 Vbias 0.38072f
C4077 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t4 Vbias 0.19125f
C4078 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n5 Vbias 0.18752f
C4079 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n6 Vbias 0.10934f
C4080 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n7 Vbias 0.01378f
C4081 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n8 Vbias 0.01095f
C4082 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t0 Vbias 0.05094f
C4083 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t1 Vbias 0.04989f
C4084 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n9 Vbias 0.28374f
C4085 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n10 Vbias 0.09258f
C4086 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t2 Vbias 0.04989f
C4087 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n11 Vbias 0.31407f
C4088 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.t7 Vbias 0.1838f
C4089 RingCounter_0.D_FlipFlop_1.3-input-nand_2.Vout.n12 Vbias 0.205f
C4090 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t5 Vbias 0.36784f
C4091 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n0 Vbias 0.10746f
C4092 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n1 Vbias 0.04662f
C4093 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t3 Vbias 0.04798f
C4094 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n2 Vbias 0.22815f
C4095 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n3 Vbias 0.0518f
C4096 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t6 Vbias 0.36785f
C4097 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n4 Vbias 0.38072f
C4098 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t7 Vbias 0.19125f
C4099 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n5 Vbias 0.18752f
C4100 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n6 Vbias 0.10934f
C4101 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n7 Vbias 0.01378f
C4102 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n8 Vbias 0.01506f
C4103 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t0 Vbias 0.05094f
C4104 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t1 Vbias 0.04989f
C4105 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n9 Vbias 0.28374f
C4106 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n10 Vbias 0.09441f
C4107 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t2 Vbias 0.04989f
C4108 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n11 Vbias 0.31407f
C4109 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.t4 Vbias 0.1838f
C4110 RingCounter_0.D_FlipFlop_10.3-input-nand_2.Vout.n12 Vbias 0.205f
C4111 Nand_Gate_6.Vout.t1 Vbias 0.08204f
C4112 Nand_Gate_6.Vout.t2 Vbias 0.09763f
C4113 Nand_Gate_6.Vout.n0 Vbias 0.49348f
C4114 Nand_Gate_6.Vout.n1 Vbias 0.25003f
C4115 Nand_Gate_6.Vout.n2 Vbias 0.08499f
C4116 Nand_Gate_6.Vout.t3 Vbias 0.31378f
C4117 Nand_Gate_6.Vout.n3 Vbias 0.30737f
C4118 Nand_Gate_6.Vout.n4 Vbias 0.06483f
C4119 Nand_Gate_6.Vout.t4 Vbias 0.60348f
C4120 Nand_Gate_6.Vout.n5 Vbias 0.17629f
C4121 Nand_Gate_6.Vout.n6 Vbias 0.04387f
C4122 Nand_Gate_6.Vout.n7 Vbias 0.06381f
C4123 Nand_Gate_6.Vout.n8 Vbias 1.30112f
C4124 Nand_Gate_6.Vout.n9 Vbias 1.30112f
C4125 Nand_Gate_6.Vout.n10 Vbias 0.0866f
C4126 Nand_Gate_6.Vout.n11 Vbias 0.04472f
C4127 Nand_Gate_6.Vout.t0 Vbias 0.07874f
C4128 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t7 Vbias 0.36784f
C4129 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n0 Vbias 0.10746f
C4130 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n1 Vbias 0.04662f
C4131 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t2 Vbias 0.04798f
C4132 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n2 Vbias 0.22815f
C4133 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n3 Vbias 0.0518f
C4134 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t4 Vbias 0.36785f
C4135 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n4 Vbias 0.38072f
C4136 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t6 Vbias 0.19125f
C4137 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n5 Vbias 0.18752f
C4138 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n6 Vbias 0.10934f
C4139 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n7 Vbias 0.01378f
C4140 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n8 Vbias 0.01506f
C4141 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t0 Vbias 0.05094f
C4142 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t1 Vbias 0.04989f
C4143 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n9 Vbias 0.28374f
C4144 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n10 Vbias 0.09441f
C4145 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t3 Vbias 0.04989f
C4146 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n11 Vbias 0.31407f
C4147 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.t5 Vbias 0.1838f
C4148 RingCounter_0.D_FlipFlop_16.3-input-nand_2.Vout.n12 Vbias 0.205f
C4149 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t7 Vbias 0.36784f
C4150 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n0 Vbias 0.10746f
C4151 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n1 Vbias 0.04662f
C4152 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t2 Vbias 0.04798f
C4153 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n2 Vbias 0.22815f
C4154 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n3 Vbias 0.0518f
C4155 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t6 Vbias 0.36785f
C4156 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n4 Vbias 0.38072f
C4157 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t5 Vbias 0.19125f
C4158 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n5 Vbias 0.18752f
C4159 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n6 Vbias 0.10934f
C4160 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n7 Vbias 0.01378f
C4161 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n8 Vbias 0.01506f
C4162 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t0 Vbias 0.05094f
C4163 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t1 Vbias 0.04989f
C4164 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n9 Vbias 0.28374f
C4165 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n10 Vbias 0.09441f
C4166 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t3 Vbias 0.04989f
C4167 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n11 Vbias 0.31407f
C4168 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.t4 Vbias 0.1838f
C4169 RingCounter_0.D_FlipFlop_11.3-input-nand_2.Vout.n12 Vbias 0.205f
C4170 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t1 Vbias 0.04607f
C4171 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n0 Vbias 0.10477f
C4172 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n1 Vbias 0.05057f
C4173 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t3 Vbias 0.35243f
C4174 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n2 Vbias 0.3654f
C4175 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n3 Vbias 0.03953f
C4176 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n4 Vbias 0.05278f
C4177 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t2 Vbias 0.27708f
C4178 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t5 Vbias 0.27709f
C4179 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n5 Vbias 0.17949f
C4180 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n6 Vbias 0.03786f
C4181 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t4 Vbias 0.35241f
C4182 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n7 Vbias 0.10295f
C4183 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n8 Vbias 0.02562f
C4184 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n9 Vbias 0.03726f
C4185 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n10 Vbias 0.09548f
C4186 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n11 Vbias 0.09548f
C4187 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n12 Vbias 0.04963f
C4188 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.t0 Vbias 0.04792f
C4189 RingCounter_0.D_FlipFlop_15.Inverter_1.Vout.n13 Vbias 0.28399f
C4190 D_FlipFlop_6.3-input-nand_2.Vout.t5 Vbias 0.35515f
C4191 D_FlipFlop_6.3-input-nand_2.Vout.n0 Vbias 0.10375f
C4192 D_FlipFlop_6.3-input-nand_2.Vout.n1 Vbias 0.04502f
C4193 D_FlipFlop_6.3-input-nand_2.Vout.n2 Vbias 0.19793f
C4194 D_FlipFlop_6.3-input-nand_2.Vout.t7 Vbias 0.17747f
C4195 D_FlipFlop_6.3-input-nand_2.Vout.t1 Vbias 0.04817f
C4196 D_FlipFlop_6.3-input-nand_2.Vout.n3 Vbias 0.30324f
C4197 D_FlipFlop_6.3-input-nand_2.Vout.t3 Vbias 0.04918f
C4198 D_FlipFlop_6.3-input-nand_2.Vout.t2 Vbias 0.04817f
C4199 D_FlipFlop_6.3-input-nand_2.Vout.n4 Vbias 0.27396f
C4200 D_FlipFlop_6.3-input-nand_2.Vout.n5 Vbias 0.09115f
C4201 D_FlipFlop_6.3-input-nand_2.Vout.n6 Vbias 0.01454f
C4202 D_FlipFlop_6.3-input-nand_2.Vout.n7 Vbias 0.01331f
C4203 D_FlipFlop_6.3-input-nand_2.Vout.t4 Vbias 0.35517f
C4204 D_FlipFlop_6.3-input-nand_2.Vout.n8 Vbias 0.36759f
C4205 D_FlipFlop_6.3-input-nand_2.Vout.t6 Vbias 0.18465f
C4206 D_FlipFlop_6.3-input-nand_2.Vout.n9 Vbias 0.18106f
C4207 D_FlipFlop_6.3-input-nand_2.Vout.n10 Vbias 0.10557f
C4208 D_FlipFlop_6.3-input-nand_2.Vout.n11 Vbias 0.05002f
C4209 D_FlipFlop_6.3-input-nand_2.Vout.t0 Vbias 0.04632f
C4210 D_FlipFlop_6.3-input-nand_2.Vout.n12 Vbias 0.22028f
C4211 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t1 Vbias 0.06069f
C4212 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n0 Vbias 0.03447f
C4213 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C4214 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C4215 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C4216 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C4217 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C4218 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C4219 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C4220 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C4221 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C4222 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C4223 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C4224 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t0 Vbias 0.06323f
C4225 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.t2 Vbias 0.07525f
C4226 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C4227 RingCounter_0.D_FlipFlop_6.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C4228 D_FlipFlop_2.3-input-nand_2.Vout.t5 Vbias 0.35515f
C4229 D_FlipFlop_2.3-input-nand_2.Vout.n0 Vbias 0.10375f
C4230 D_FlipFlop_2.3-input-nand_2.Vout.n1 Vbias 0.04502f
C4231 D_FlipFlop_2.3-input-nand_2.Vout.t2 Vbias 0.04632f
C4232 D_FlipFlop_2.3-input-nand_2.Vout.n2 Vbias 0.22028f
C4233 D_FlipFlop_2.3-input-nand_2.Vout.n3 Vbias 0.05002f
C4234 D_FlipFlop_2.3-input-nand_2.Vout.t4 Vbias 0.35517f
C4235 D_FlipFlop_2.3-input-nand_2.Vout.n4 Vbias 0.36759f
C4236 D_FlipFlop_2.3-input-nand_2.Vout.t6 Vbias 0.18465f
C4237 D_FlipFlop_2.3-input-nand_2.Vout.n5 Vbias 0.18106f
C4238 D_FlipFlop_2.3-input-nand_2.Vout.n6 Vbias 0.10557f
C4239 D_FlipFlop_2.3-input-nand_2.Vout.n7 Vbias 0.01331f
C4240 D_FlipFlop_2.3-input-nand_2.Vout.n8 Vbias 0.01454f
C4241 D_FlipFlop_2.3-input-nand_2.Vout.t3 Vbias 0.04918f
C4242 D_FlipFlop_2.3-input-nand_2.Vout.t0 Vbias 0.04817f
C4243 D_FlipFlop_2.3-input-nand_2.Vout.n9 Vbias 0.27396f
C4244 D_FlipFlop_2.3-input-nand_2.Vout.n10 Vbias 0.09115f
C4245 D_FlipFlop_2.3-input-nand_2.Vout.t1 Vbias 0.04817f
C4246 D_FlipFlop_2.3-input-nand_2.Vout.n11 Vbias 0.30324f
C4247 D_FlipFlop_2.3-input-nand_2.Vout.t7 Vbias 0.17747f
C4248 D_FlipFlop_2.3-input-nand_2.Vout.n12 Vbias 0.19793f
C4249 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t1 Vbias 0.06624f
C4250 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t2 Vbias 0.07883f
C4251 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n0 Vbias 0.39844f
C4252 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n1 Vbias 0.20187f
C4253 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n2 Vbias 0.06862f
C4254 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t4 Vbias 0.25335f
C4255 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n3 Vbias 0.24817f
C4256 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n4 Vbias 0.05234f
C4257 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t3 Vbias 0.48726f
C4258 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n5 Vbias 0.14234f
C4259 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n6 Vbias 0.03542f
C4260 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n7 Vbias 0.05152f
C4261 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C4262 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n9 Vbias 0.13202f
C4263 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n10 Vbias 0.06992f
C4264 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.n11 Vbias 0.03611f
C4265 RingCounter_0.D_FlipFlop_2.Nand_Gate_1.Vout.t0 Vbias 0.06358f
C4266 And_Gate_1.B.t1 Vbias 0.0378f
C4267 Nand_Gate_4.Vout Vbias -0.07584f
C4268 And_Gate_1.B.n0 Vbias 0.02147f
C4269 And_Gate_1.B.n1 Vbias 0.04157f
C4270 And_Gate_1.B.t3 Vbias 0.15061f
C4271 And_Gate_1.Nand_Gate_0.B Vbias -0.11323f
C4272 And_Gate_1.B.n2 Vbias 0.14754f
C4273 And_Gate_1.B.n3 Vbias 0.03112f
C4274 And_Gate_1.B.t4 Vbias 0.28967f
C4275 And_Gate_1.B.n4 Vbias 0.08462f
C4276 And_Gate_1.B.n5 Vbias 0.02106f
C4277 And_Gate_1.B.n6 Vbias 0.03063f
C4278 And_Gate_1.B.n7 Vbias 0.62454f
C4279 And_Gate_1.B.n8 Vbias 0.62454f
C4280 And_Gate_1.B.n9 Vbias 0.04079f
C4281 And_Gate_1.B.t2 Vbias 0.03938f
C4282 And_Gate_1.B.t0 Vbias 0.04686f
C4283 And_Gate_1.B.n10 Vbias 0.23687f
C4284 And_Gate_1.B.n11 Vbias 0.12001f
C4285 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t1 Vbias 0.05803f
C4286 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n0 Vbias 0.15518f
C4287 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n1 Vbias 0.11917f
C4288 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t7 Vbias 0.23082f
C4289 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t4 Vbias 0.44396f
C4290 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n2 Vbias 0.12969f
C4291 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n3 Vbias 0.05546f
C4292 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n4 Vbias 0.1024f
C4293 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n5 Vbias 0.1773f
C4294 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n6 Vbias 0.13197f
C4295 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n7 Vbias 0.06252f
C4296 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t5 Vbias 0.44398f
C4297 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n8 Vbias 0.46032f
C4298 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n9 Vbias 0.0498f
C4299 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n10 Vbias 0.06649f
C4300 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t6 Vbias 0.22095f
C4301 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t0 Vbias 0.06022f
C4302 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n11 Vbias 0.37982f
C4303 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t3 Vbias 0.06148f
C4304 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.t2 Vbias 0.06022f
C4305 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n12 Vbias 0.34246f
C4306 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n13 Vbias 0.11306f
C4307 RingCounter_0.D_FlipFlop_16.3-input-nand_2.C.n14 Vbias 0.16074f
C4308 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t6 Vbias 0.36784f
C4309 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n0 Vbias 0.10746f
C4310 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n1 Vbias 0.04662f
C4311 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t2 Vbias 0.04798f
C4312 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n2 Vbias 0.22815f
C4313 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n3 Vbias 0.0518f
C4314 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t7 Vbias 0.36785f
C4315 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n4 Vbias 0.38072f
C4316 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t5 Vbias 0.19125f
C4317 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n5 Vbias 0.18752f
C4318 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n6 Vbias 0.10934f
C4319 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n7 Vbias 0.01378f
C4320 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n8 Vbias 0.01095f
C4321 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t0 Vbias 0.05094f
C4322 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t1 Vbias 0.04989f
C4323 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n9 Vbias 0.28374f
C4324 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n10 Vbias 0.09258f
C4325 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t3 Vbias 0.04989f
C4326 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n11 Vbias 0.31407f
C4327 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.t4 Vbias 0.1838f
C4328 RingCounter_0.D_FlipFlop_4.3-input-nand_2.Vout.n12 Vbias 0.205f
C4329 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t1 Vbias 0.04607f
C4330 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n0 Vbias 0.10477f
C4331 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n1 Vbias 0.05057f
C4332 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t3 Vbias 0.35243f
C4333 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n2 Vbias 0.3654f
C4334 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n3 Vbias 0.03953f
C4335 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n4 Vbias 0.05278f
C4336 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t2 Vbias 0.27708f
C4337 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t5 Vbias 0.27709f
C4338 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n5 Vbias 0.17949f
C4339 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n6 Vbias 0.03786f
C4340 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t4 Vbias 0.35241f
C4341 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n7 Vbias 0.10295f
C4342 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n8 Vbias 0.02562f
C4343 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n9 Vbias 0.03726f
C4344 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n10 Vbias 0.09548f
C4345 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n11 Vbias 0.09548f
C4346 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n12 Vbias 0.04963f
C4347 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.t0 Vbias 0.04792f
C4348 RingCounter_0.D_FlipFlop_12.Inverter_1.Vout.n13 Vbias 0.28399f
C4349 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t2 Vbias 0.0608f
C4350 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C4351 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C4352 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t3 Vbias 0.24183f
C4353 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C4354 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C4355 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t4 Vbias 0.46511f
C4356 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C4357 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C4358 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C4359 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C4360 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C4361 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C4362 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t1 Vbias 0.06323f
C4363 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C4364 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C4365 RingCounter_0.D_FlipFlop_13.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C4366 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t4 Vbias 0.45666f
C4367 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n0 Vbias 0.47347f
C4368 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n1 Vbias 0.05122f
C4369 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t2 Vbias 0.05969f
C4370 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n2 Vbias 0.15961f
C4371 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n3 Vbias 0.12257f
C4372 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t5 Vbias 0.23742f
C4373 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t7 Vbias 0.45664f
C4374 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n4 Vbias 0.1334f
C4375 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n5 Vbias 0.05705f
C4376 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n6 Vbias 0.10533f
C4377 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n7 Vbias 0.18236f
C4378 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n8 Vbias 0.13574f
C4379 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n9 Vbias 0.06431f
C4380 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n10 Vbias 0.16533f
C4381 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t3 Vbias 0.06323f
C4382 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t0 Vbias 0.06194f
C4383 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n11 Vbias 0.35224f
C4384 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n12 Vbias 0.11629f
C4385 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t1 Vbias 0.06194f
C4386 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n13 Vbias 0.39067f
C4387 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.t6 Vbias 0.22727f
C4388 RingCounter_0.D_FlipFlop_10.3-input-nand_2.C.n14 Vbias 0.06839f
C4389 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t2 Vbias 0.07037f
C4390 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n0 Vbias 0.16004f
C4391 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n1 Vbias 0.07725f
C4392 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t4 Vbias 0.2799f
C4393 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n2 Vbias 0.27418f
C4394 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n3 Vbias 0.05783f
C4395 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t5 Vbias 0.53832f
C4396 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n4 Vbias 0.15726f
C4397 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n5 Vbias 0.03913f
C4398 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n6 Vbias 0.05692f
C4399 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n7 Vbias 0.14585f
C4400 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n8 Vbias 0.14585f
C4401 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n9 Vbias 0.07581f
C4402 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t3 Vbias 0.07318f
C4403 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t0 Vbias 0.07454f
C4404 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.t1 Vbias 0.07302f
C4405 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n10 Vbias 0.41525f
C4406 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n11 Vbias 0.23391f
C4407 RingCounter_0.D_FlipFlop_10.3-input-nand_1.Vout.n12 Vbias 0.22303f
C4408 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t2 Vbias 0.07024f
C4409 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n0 Vbias 0.03989f
C4410 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n1 Vbias 0.07725f
C4411 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t5 Vbias 0.2799f
C4412 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n2 Vbias 0.27418f
C4413 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n3 Vbias 0.05783f
C4414 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t4 Vbias 0.53832f
C4415 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n4 Vbias 0.15726f
C4416 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n5 Vbias 0.03913f
C4417 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n6 Vbias 0.05692f
C4418 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n7 Vbias 0.14585f
C4419 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n8 Vbias 0.14585f
C4420 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n9 Vbias 0.07581f
C4421 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t3 Vbias 0.07318f
C4422 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t0 Vbias 0.07454f
C4423 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.t1 Vbias 0.07302f
C4424 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n10 Vbias 0.41525f
C4425 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n11 Vbias 0.23391f
C4426 RingCounter_0.D_FlipFlop_6.3-input-nand_1.Vout.n12 Vbias 0.22303f
C4427 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t5 Vbias 0.45666f
C4428 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n0 Vbias 0.47347f
C4429 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n1 Vbias 0.05122f
C4430 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t1 Vbias 0.05969f
C4431 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n2 Vbias 0.15961f
C4432 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n3 Vbias 0.12257f
C4433 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t7 Vbias 0.23742f
C4434 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t4 Vbias 0.45664f
C4435 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n4 Vbias 0.1334f
C4436 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n5 Vbias 0.05705f
C4437 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n6 Vbias 0.10533f
C4438 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n7 Vbias 0.18236f
C4439 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n8 Vbias 0.13574f
C4440 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n9 Vbias 0.06431f
C4441 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n10 Vbias 0.16533f
C4442 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t3 Vbias 0.06323f
C4443 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t0 Vbias 0.06194f
C4444 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n11 Vbias 0.35224f
C4445 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n12 Vbias 0.11629f
C4446 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t2 Vbias 0.06194f
C4447 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n13 Vbias 0.39067f
C4448 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.t6 Vbias 0.22727f
C4449 RingCounter_0.D_FlipFlop_14.3-input-nand_2.C.n14 Vbias 0.06839f
C4450 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t1 Vbias 0.04998f
C4451 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n0 Vbias 0.02839f
C4452 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n1 Vbias 0.05497f
C4453 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t2 Vbias 0.38308f
C4454 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n2 Vbias 0.39717f
C4455 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n3 Vbias 0.04297f
C4456 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n4 Vbias 0.05737f
C4457 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t3 Vbias 0.30118f
C4458 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t5 Vbias 0.30119f
C4459 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n5 Vbias 0.1951f
C4460 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n6 Vbias 0.04115f
C4461 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t4 Vbias 0.38306f
C4462 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n7 Vbias 0.1119f
C4463 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n8 Vbias 0.02784f
C4464 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n9 Vbias 0.0405f
C4465 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n10 Vbias 0.10379f
C4466 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n11 Vbias 0.10379f
C4467 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n12 Vbias 0.05395f
C4468 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.t0 Vbias 0.05208f
C4469 RingCounter_0.D_FlipFlop_5.Inverter_1.Vout.n13 Vbias 0.30868f
C4470 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t1 Vbias 0.06067f
C4471 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n0 Vbias 0.26418f
C4472 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n1 Vbias 0.0655f
C4473 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t3 Vbias 0.46513f
C4474 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n2 Vbias 0.4571f
C4475 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n3 Vbias 0.04996f
C4476 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t4 Vbias 0.24182f
C4477 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n4 Vbias 0.06966f
C4478 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n5 Vbias 0.02985f
C4479 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n6 Vbias 0.05594f
C4480 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n7 Vbias 0.12602f
C4481 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n8 Vbias 0.12602f
C4482 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n9 Vbias 0.07553f
C4483 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n10 Vbias 0.03814f
C4484 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t0 Vbias 0.06323f
C4485 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.t2 Vbias 0.07525f
C4486 RingCounter_0.D_FlipFlop_17.Nand_Gate_0.Vout.n11 Vbias 0.37895f
C4487 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t1 Vbias 0.03999f
C4488 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n0 Vbias 0.02271f
C4489 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n1 Vbias 0.04398f
C4490 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t2 Vbias 0.30646f
C4491 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n2 Vbias 0.31774f
C4492 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n3 Vbias 0.03438f
C4493 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n4 Vbias 0.0459f
C4494 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t3 Vbias 0.24094f
C4495 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t5 Vbias 0.24095f
C4496 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n5 Vbias 0.15608f
C4497 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n6 Vbias 0.03292f
C4498 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t4 Vbias 0.30645f
C4499 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n7 Vbias 0.08952f
C4500 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n8 Vbias 0.02228f
C4501 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n9 Vbias 0.0324f
C4502 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n10 Vbias 0.08303f
C4503 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n11 Vbias 0.08303f
C4504 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n12 Vbias 0.04316f
C4505 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.t0 Vbias 0.04167f
C4506 RingCounter_0.D_FlipFlop_17.Inverter_1.Vout.n13 Vbias 0.24695f
C4507 RingCounter_0.D_FlipFlop_16.Q.t5 Vbias 0.09863f
C4508 RingCounter_0.D_FlipFlop_16.Q.n0 Vbias 0.02881f
C4509 RingCounter_0.D_FlipFlop_16.Q.n1 Vbias 0.0125f
C4510 RingCounter_0.D_FlipFlop_16.Q.n2 Vbias 0.05497f
C4511 RingCounter_0.D_FlipFlop_16.Q.t8 Vbias 0.04587f
C4512 RingCounter_0.D_FlipFlop_16.Q.n3 Vbias 0.01439f
C4513 RingCounter_0.D_FlipFlop_16.Q.t4 Vbias 0.09863f
C4514 RingCounter_0.D_FlipFlop_16.Q.n4 Vbias 0.09693f
C4515 RingCounter_0.D_FlipFlop_16.Q.n5 Vbias 0.01059f
C4516 RingCounter_0.D_FlipFlop_16.Q.t6 Vbias 0.05128f
C4517 RingCounter_0.D_FlipFlop_16.Q.n6 Vbias 0.01477f
C4518 RingCounter_0.D_FlipFlop_16.Q.n8 Vbias 0.01186f
C4519 RingCounter_0.D_FlipFlop_16.Q.n9 Vbias 0.01493f
C4520 RingCounter_0.D_FlipFlop_16.Q.t9 Vbias 0.09863f
C4521 RingCounter_0.D_FlipFlop_16.Q.n10 Vbias 0.09693f
C4522 RingCounter_0.D_FlipFlop_16.Q.n11 Vbias 0.01059f
C4523 RingCounter_0.D_FlipFlop_16.Q.t7 Vbias 0.05128f
C4524 RingCounter_0.D_FlipFlop_16.Q.n12 Vbias 0.01477f
C4525 RingCounter_0.D_FlipFlop_16.Q.n14 Vbias 0.01186f
C4526 RingCounter_0.D_FlipFlop_16.Q.n16 Vbias 0.83774f
C4527 RingCounter_0.D_FlipFlop_16.Q.t1 Vbias 0.01286f
C4528 RingCounter_0.D_FlipFlop_16.Q.n17 Vbias 0.06309f
C4529 RingCounter_0.D_FlipFlop_16.Q.n18 Vbias 0.01548f
C4530 RingCounter_0.D_FlipFlop_16.Q.t0 Vbias 0.01366f
C4531 RingCounter_0.D_FlipFlop_16.Q.t3 Vbias 0.01338f
C4532 RingCounter_0.D_FlipFlop_16.Q.n19 Vbias 0.07608f
C4533 RingCounter_0.D_FlipFlop_16.Q.n20 Vbias 0.02531f
C4534 RingCounter_0.D_FlipFlop_16.Q.t2 Vbias 0.01338f
C4535 RingCounter_0.D_FlipFlop_16.Q.n21 Vbias 0.02059f
C4536 RingCounter_0.D_FlipFlop_16.Q.n22 Vbias 1.6069f
C4537 RingCounter_0.D_FlipFlop_16.Q.n23 Vbias 0.03074f
C4538 CDAC8_0.switch_0.Z.t1 Vbias 0.03482f
C4539 CDAC8_0.switch_0.Z.t5 Vbias 5.94383f
C4540 CDAC8_0.switch_0.Z.n0 Vbias 2.04684f
C4541 CDAC8_0.switch_0.Z.t7 Vbias 5.94383f
C4542 CDAC8_0.switch_0.Z.t6 Vbias 5.85885f
C4543 CDAC8_0.switch_0.Z.n1 Vbias 2.17361f
C4544 CDAC8_0.switch_0.Z.t4 Vbias 5.85885f
C4545 CDAC8_0.switch_0.Z.n2 Vbias 2.17361f
C4546 CDAC8_0.switch_0.Z.n3 Vbias 2.00334f
C4547 CDAC8_0.switch_0.Z.n4 Vbias 0.50573f
C4548 CDAC8_0.switch_0.Z.t2 Vbias 0.0348f
C4549 CDAC8_0.switch_0.Z.n5 Vbias 0.11883f
C4550 CDAC8_0.switch_0.Z.t3 Vbias 0.03316f
C4551 CDAC8_0.switch_0.Z.t0 Vbias 0.03316f
C4552 CDAC8_0.switch_0.Z.n6 Vbias 0.11982f
C4553 CDAC8_0.switch_0.Z.n7 Vbias 0.27578f
C4554 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t1 Vbias 0.06323f
C4555 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t2 Vbias 0.07525f
C4556 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n0 Vbias 0.38033f
C4557 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n1 Vbias 0.1927f
C4558 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n2 Vbias 0.0655f
C4559 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t3 Vbias 0.24183f
C4560 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n3 Vbias 0.23689f
C4561 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n4 Vbias 0.04996f
C4562 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t4 Vbias 0.46511f
C4563 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n5 Vbias 0.13587f
C4564 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n6 Vbias 0.03381f
C4565 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n7 Vbias 0.04918f
C4566 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C4567 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n9 Vbias 0.12602f
C4568 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n10 Vbias 0.06674f
C4569 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.t0 Vbias 0.0608f
C4570 RingCounter_0.D_FlipFlop_8.Nand_Gate_1.Vout.n11 Vbias 0.13827f
C4571 D_FlipFlop_4.3-input-nand_2.C.t5 Vbias 0.3425f
C4572 D_FlipFlop_4.3-input-nand_2.C.n0 Vbias 0.3551f
C4573 D_FlipFlop_4.3-input-nand_2.C.n1 Vbias 0.03842f
C4574 D_FlipFlop_4.3-input-nand_2.C.n2 Vbias 0.05129f
C4575 D_FlipFlop_4.3-input-nand_2.C.t4 Vbias 0.17045f
C4576 D_FlipFlop_4.3-input-nand_2.C.t1 Vbias 0.04645f
C4577 D_FlipFlop_4.3-input-nand_2.C.n3 Vbias 0.293f
C4578 D_FlipFlop_4.3-input-nand_2.C.t3 Vbias 0.04742f
C4579 D_FlipFlop_4.3-input-nand_2.C.t2 Vbias 0.04645f
C4580 D_FlipFlop_4.3-input-nand_2.C.n4 Vbias 0.26418f
C4581 D_FlipFlop_4.3-input-nand_2.C.n5 Vbias 0.08722f
C4582 D_FlipFlop_4.3-input-nand_2.C.n6 Vbias 0.124f
C4583 D_FlipFlop_4.3-input-nand_2.C.n7 Vbias 0.04823f
C4584 D_FlipFlop_4.3-input-nand_2.C.t6 Vbias 0.17806f
C4585 D_FlipFlop_4.3-input-nand_2.C.t7 Vbias 0.34248f
C4586 D_FlipFlop_4.3-input-nand_2.C.n8 Vbias 0.10005f
C4587 D_FlipFlop_4.3-input-nand_2.C.n9 Vbias 0.04279f
C4588 D_FlipFlop_4.3-input-nand_2.C.n10 Vbias 0.079f
C4589 D_FlipFlop_4.3-input-nand_2.C.n11 Vbias 0.13677f
C4590 D_FlipFlop_4.3-input-nand_2.C.n12 Vbias 0.10181f
C4591 D_FlipFlop_4.3-input-nand_2.C.n13 Vbias 0.09193f
C4592 D_FlipFlop_4.3-input-nand_2.C.t0 Vbias 0.04477f
C4593 D_FlipFlop_4.3-input-nand_2.C.n14 Vbias 0.11971f
C4594 D_FlipFlop_4.3-input-nand_2.Vout.t4 Vbias 0.35515f
C4595 D_FlipFlop_4.3-input-nand_2.Vout.n0 Vbias 0.10375f
C4596 D_FlipFlop_4.3-input-nand_2.Vout.n1 Vbias 0.04502f
C4597 D_FlipFlop_4.3-input-nand_2.Vout.t3 Vbias 0.04632f
C4598 D_FlipFlop_4.3-input-nand_2.Vout.n2 Vbias 0.22028f
C4599 D_FlipFlop_4.3-input-nand_2.Vout.n3 Vbias 0.05002f
C4600 D_FlipFlop_4.3-input-nand_2.Vout.t6 Vbias 0.35517f
C4601 D_FlipFlop_4.3-input-nand_2.Vout.n4 Vbias 0.36759f
C4602 D_FlipFlop_4.3-input-nand_2.Vout.t5 Vbias 0.18465f
C4603 D_FlipFlop_4.3-input-nand_2.Vout.n5 Vbias 0.18106f
C4604 D_FlipFlop_4.3-input-nand_2.Vout.n6 Vbias 0.10557f
C4605 D_FlipFlop_4.3-input-nand_2.Vout.n7 Vbias 0.01331f
C4606 D_FlipFlop_4.3-input-nand_2.Vout.n8 Vbias 0.01454f
C4607 D_FlipFlop_4.3-input-nand_2.Vout.t0 Vbias 0.04918f
C4608 D_FlipFlop_4.3-input-nand_2.Vout.t1 Vbias 0.04817f
C4609 D_FlipFlop_4.3-input-nand_2.Vout.n9 Vbias 0.27396f
C4610 D_FlipFlop_4.3-input-nand_2.Vout.n10 Vbias 0.09115f
C4611 D_FlipFlop_4.3-input-nand_2.Vout.t2 Vbias 0.04817f
C4612 D_FlipFlop_4.3-input-nand_2.Vout.n11 Vbias 0.30324f
C4613 D_FlipFlop_4.3-input-nand_2.Vout.t7 Vbias 0.17747f
C4614 D_FlipFlop_4.3-input-nand_2.Vout.n12 Vbias 0.19793f
C4615 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t2 Vbias 0.07024f
C4616 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n0 Vbias 0.03989f
C4617 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n1 Vbias 0.07725f
C4618 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t4 Vbias 0.2799f
C4619 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n2 Vbias 0.27418f
C4620 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n3 Vbias 0.05783f
C4621 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t5 Vbias 0.53832f
C4622 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n4 Vbias 0.15726f
C4623 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n5 Vbias 0.03913f
C4624 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n6 Vbias 0.05692f
C4625 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n7 Vbias 0.14585f
C4626 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n8 Vbias 0.14585f
C4627 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n9 Vbias 0.07581f
C4628 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t3 Vbias 0.07318f
C4629 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t0 Vbias 0.07454f
C4630 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.t1 Vbias 0.07302f
C4631 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n10 Vbias 0.41525f
C4632 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n11 Vbias 0.23391f
C4633 RingCounter_0.D_FlipFlop_1.3-input-nand_1.Vout.n12 Vbias 0.22303f
C4634 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t2 Vbias 0.05201f
C4635 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n0 Vbias 0.22649f
C4636 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n1 Vbias 0.05616f
C4637 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t4 Vbias 0.39877f
C4638 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n2 Vbias 0.39189f
C4639 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n3 Vbias 0.04283f
C4640 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t5 Vbias 0.20732f
C4641 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n4 Vbias 0.05972f
C4642 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n5 Vbias 0.02559f
C4643 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n6 Vbias 0.04796f
C4644 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n7 Vbias 0.10804f
C4645 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n8 Vbias 0.10804f
C4646 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n9 Vbias 0.06475f
C4647 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t3 Vbias 0.05421f
C4648 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t1 Vbias 0.05522f
C4649 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.t0 Vbias 0.05409f
C4650 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n10 Vbias 0.30759f
C4651 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n11 Vbias 0.17406f
C4652 RingCounter_0.D_FlipFlop_15.3-input-nand_0.Vout.n12 Vbias 0.03715f
C4653 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t2 Vbias 0.05201f
C4654 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n0 Vbias 0.22649f
C4655 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n1 Vbias 0.05616f
C4656 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t4 Vbias 0.39877f
C4657 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n2 Vbias 0.39189f
C4658 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n3 Vbias 0.04283f
C4659 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t5 Vbias 0.20732f
C4660 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n4 Vbias 0.05972f
C4661 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n5 Vbias 0.02559f
C4662 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n6 Vbias 0.04796f
C4663 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n7 Vbias 0.10804f
C4664 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n8 Vbias 0.10804f
C4665 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n9 Vbias 0.06475f
C4666 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t3 Vbias 0.05421f
C4667 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t1 Vbias 0.05522f
C4668 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.t0 Vbias 0.05409f
C4669 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n10 Vbias 0.30759f
C4670 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n11 Vbias 0.17406f
C4671 RingCounter_0.D_FlipFlop_9.3-input-nand_0.Vout.n12 Vbias 0.03715f
C4672 And_Gate_5.A.t1 Vbias 0.03721f
C4673 And_Gate_5.A.t2 Vbias 0.04429f
C4674 And_Gate_5.A.n0 Vbias 0.22385f
C4675 Nand_Gate_3.Vout Vbias -0.07167f
C4676 And_Gate_5.A.n1 Vbias 0.11341f
C4677 And_Gate_5.A.n2 Vbias 0.03855f
C4678 And_Gate_5.A.t4 Vbias 0.14233f
C4679 And_Gate_5.Nand_Gate_0.A Vbias -0.10701f
C4680 And_Gate_5.A.n3 Vbias 0.13943f
C4681 And_Gate_5.A.n4 Vbias 0.02941f
C4682 And_Gate_5.A.t3 Vbias 0.27375f
C4683 And_Gate_5.A.n5 Vbias 0.07997f
C4684 And_Gate_5.A.n6 Vbias 0.0199f
C4685 And_Gate_5.A.n7 Vbias 0.02895f
C4686 And_Gate_5.A.n8 Vbias 0.55617f
C4687 And_Gate_5.A.n9 Vbias 0.55617f
C4688 And_Gate_5.A.n10 Vbias 0.03928f
C4689 And_Gate_5.A.n11 Vbias 0.02029f
C4690 And_Gate_5.A.t0 Vbias 0.03572f
C4691 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t6 Vbias 0.45666f
C4692 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n0 Vbias 0.47347f
C4693 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n1 Vbias 0.05122f
C4694 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n2 Vbias 0.06839f
C4695 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t5 Vbias 0.22727f
C4696 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t2 Vbias 0.06194f
C4697 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n3 Vbias 0.39067f
C4698 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t3 Vbias 0.06323f
C4699 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t1 Vbias 0.06194f
C4700 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n4 Vbias 0.35224f
C4701 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n5 Vbias 0.11629f
C4702 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n6 Vbias 0.16533f
C4703 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n7 Vbias 0.06431f
C4704 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t7 Vbias 0.23742f
C4705 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t4 Vbias 0.45664f
C4706 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n8 Vbias 0.1334f
C4707 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n9 Vbias 0.05705f
C4708 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n10 Vbias 0.10533f
C4709 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n11 Vbias 0.18236f
C4710 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n12 Vbias 0.13574f
C4711 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n13 Vbias 0.12257f
C4712 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.t0 Vbias 0.05969f
C4713 RingCounter_0.D_FlipFlop_11.3-input-nand_2.C.n14 Vbias 0.15961f
C4714 And_Gate_0.Vout.t1 Vbias 0.12492f
C4715 And_Gate_0.Inverter_0.Vout Vbias 0.03629f
C4716 And_Gate_0.Vout.n0 Vbias 0.13783f
C4717 And_Gate_0.Vout.t4 Vbias 0.95742f
C4718 D_FlipFlop_6.3-input-nand_0.C Vbias -0.56919f
C4719 And_Gate_0.Vout.n1 Vbias 0.99266f
C4720 And_Gate_0.Vout.n2 Vbias 0.10739f
C4721 And_Gate_0.Vout.n3 Vbias 0.14338f
C4722 And_Gate_0.Vout.t5 Vbias 0.44073f
C4723 D_FlipFlop_6.CLK Vbias -0.01479f
C4724 And_Gate_0.Vout.n4 Vbias 0.35269f
C4725 And_Gate_0.Vout.t3 Vbias 0.95737f
C4726 D_FlipFlop_6.3-input-nand_1.C Vbias -0.32001f
C4727 And_Gate_0.Vout.t6 Vbias 0.49778f
C4728 D_FlipFlop_6.Inverter_1.Vin Vbias -0.3108f
C4729 And_Gate_0.Vout.n5 Vbias 0.52493f
C4730 And_Gate_0.Vout.t2 Vbias 0.95737f
C4731 And_Gate_0.Vout.n6 Vbias 0.84748f
C4732 And_Gate_0.Vout.n7 Vbias 0.84981f
C4733 And_Gate_0.Vout.n8 Vbias 0.53181f
C4734 And_Gate_0.Vout.t7 Vbias 0.44069f
C4735 And_Gate_0.Vout.n9 Vbias 0.0818f
C4736 And_Gate_0.Vout.n10 Vbias 0.19316f
C4737 And_Gate_0.Vout.n11 Vbias 18.7304f
C4738 And_Gate_0.Vout.t0 Vbias 0.13044f
C4739 And_Gate_0.Vout.n12 Vbias 15.2812f
C4740 And_Gate_0.Vout.n13 Vbias 0.29731f
C4741 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t2 Vbias 0.05201f
C4742 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n0 Vbias 0.22649f
C4743 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n1 Vbias 0.05616f
C4744 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t4 Vbias 0.39877f
C4745 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n2 Vbias 0.39189f
C4746 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n3 Vbias 0.04283f
C4747 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t5 Vbias 0.20732f
C4748 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n4 Vbias 0.05972f
C4749 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n5 Vbias 0.02559f
C4750 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n6 Vbias 0.04796f
C4751 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n7 Vbias 0.10804f
C4752 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n8 Vbias 0.10804f
C4753 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n9 Vbias 0.06475f
C4754 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t3 Vbias 0.05421f
C4755 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t1 Vbias 0.05522f
C4756 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.t0 Vbias 0.05409f
C4757 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n10 Vbias 0.30759f
C4758 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n11 Vbias 0.17406f
C4759 RingCounter_0.D_FlipFlop_12.3-input-nand_0.Vout.n12 Vbias 0.03715f
C4760 And_Gate_6.Vout.t1 Vbias 0.09234f
C4761 And_Gate_6.Inverter_0.Vout Vbias -0.29682f
C4762 And_Gate_6.Vout.n0 Vbias 0.05245f
C4763 And_Gate_6.Vout.n1 Vbias 0.10156f
C4764 And_Gate_6.Vout.t5 Vbias 0.70775f
C4765 D_FlipFlop_3.3-input-nand_0.C Vbias -0.42076f
C4766 And_Gate_6.Vout.n2 Vbias 0.7338f
C4767 And_Gate_6.Vout.n3 Vbias 0.07939f
C4768 And_Gate_6.Vout.n4 Vbias 0.10599f
C4769 And_Gate_6.Vout.t2 Vbias 0.32576f
C4770 D_FlipFlop_3.CLK Vbias 0.04733f
C4771 And_Gate_6.Vout.n5 Vbias 0.31014f
C4772 And_Gate_6.Vout.n6 Vbias 0.09329f
C4773 And_Gate_6.Vout.t7 Vbias 0.70772f
C4774 D_FlipFlop_3.3-input-nand_1.C Vbias -0.23656f
C4775 And_Gate_6.Vout.t3 Vbias 0.36798f
C4776 D_FlipFlop_3.Inverter_1.Vin Vbias -0.22976f
C4777 And_Gate_6.Vout.n7 Vbias 0.38805f
C4778 And_Gate_6.Vout.t6 Vbias 0.70772f
C4779 And_Gate_6.Vout.n8 Vbias 0.62648f
C4780 And_Gate_6.Vout.n9 Vbias 0.6282f
C4781 And_Gate_6.Vout.n10 Vbias 0.39313f
C4782 And_Gate_6.Vout.t4 Vbias 0.32577f
C4783 And_Gate_6.Vout.n11 Vbias 7.68586f
C4784 And_Gate_6.Vout.n12 Vbias 5.63698f
C4785 And_Gate_6.Vout.n13 Vbias 0.09967f
C4786 And_Gate_6.Vout.t0 Vbias 0.09623f
C4787 And_Gate_6.Vout.n14 Vbias 0.57031f
C4788 Q4.t1 Vbias 0.01589f
C4789 Q4.n0 Vbias 0.07793f
C4790 Q4.n1 Vbias 0.01912f
C4791 Q4.t3 Vbias 0.01687f
C4792 Q4.t0 Vbias 0.01653f
C4793 Q4.n2 Vbias 0.09398f
C4794 Q4.n3 Vbias 0.03127f
C4795 Q4.t2 Vbias 0.01653f
C4796 Q4.n4 Vbias 0.02546f
C4797 Q4.n5 Vbias 0.03664f
C4798 Q4.n6 Vbias 0.01877f
C4799 Q4.t5 Vbias 0.12183f
C4800 Q4.n7 Vbias 0.03559f
C4801 Q4.n8 Vbias 0.01544f
C4802 Q4.n9 Vbias 0.0679f
C4803 Q4.t9 Vbias 0.05667f
C4804 Q4.n11 Vbias 0.01459f
C4805 Q4.n13 Vbias 3.26567f
C4806 Q4.n14 Vbias 1.24988f
C4807 Q4.t4 Vbias 0.12215f
C4808 Q4.t6 Vbias 0.12215f
C4809 Q4.t8 Vbias 0.06345f
C4810 Q4.n15 Vbias 0.09883f
C4811 Q4.n16 Vbias 0.07245f
C4812 Q4.t7 Vbias 0.06334f
C4813 Q4.n17 Vbias 0.02077f
C4814 Nand_Gate_1.A.t10 Vbias 0.27993f
C4815 Nand_Gate_1.A.n0 Vbias 0.08177f
C4816 Nand_Gate_1.A.n1 Vbias 0.03548f
C4817 Nand_Gate_1.A.n2 Vbias 0.15601f
C4818 Nand_Gate_1.A.t6 Vbias 0.1302f
C4819 Nand_Gate_1.A.n3 Vbias 0.04085f
C4820 Nand_Gate_1.A.t2 Vbias 0.03651f
C4821 Nand_Gate_1.A.n4 Vbias 0.159f
C4822 Nand_Gate_1.A.n5 Vbias 0.03942f
C4823 Nand_Gate_1.A.t7 Vbias 0.27994f
C4824 Nand_Gate_1.A.n6 Vbias 0.27511f
C4825 Nand_Gate_1.A.n7 Vbias 0.03007f
C4826 Nand_Gate_1.A.t11 Vbias 0.14554f
C4827 Nand_Gate_1.A.n8 Vbias 0.04192f
C4828 Nand_Gate_1.A.n9 Vbias 0.01797f
C4829 Nand_Gate_1.A.n10 Vbias 0.03367f
C4830 Nand_Gate_1.A.n11 Vbias 0.04236f
C4831 Nand_Gate_1.A.t9 Vbias 0.27994f
C4832 Nand_Gate_1.A.n12 Vbias 0.27511f
C4833 Nand_Gate_1.A.n13 Vbias 0.03007f
C4834 Nand_Gate_1.A.t4 Vbias 0.14554f
C4835 Nand_Gate_1.A.n14 Vbias 0.04192f
C4836 Nand_Gate_1.A.n15 Vbias 0.01797f
C4837 Nand_Gate_1.A.n16 Vbias 0.03367f
C4838 Nand_Gate_1.A.n18 Vbias 0.12656f
C4839 Nand_Gate_1.A.n19 Vbias 0.03459f
C4840 Nand_Gate_1.A.n20 Vbias 0.09204f
C4841 Nand_Gate_1.A.t5 Vbias 0.14555f
C4842 Nand_Gate_1.A.n21 Vbias 0.14257f
C4843 Nand_Gate_1.A.n22 Vbias 0.03007f
C4844 Nand_Gate_1.A.t8 Vbias 0.27993f
C4845 Nand_Gate_1.A.n23 Vbias 0.08177f
C4846 Nand_Gate_1.A.n24 Vbias 0.02035f
C4847 Nand_Gate_1.A.n25 Vbias 0.0296f
C4848 Nand_Gate_1.A.n26 Vbias 0.14551f
C4849 Nand_Gate_1.A.n27 Vbias 0.25531f
C4850 Nand_Gate_1.A.n28 Vbias 0.15873f
C4851 Nand_Gate_1.A.n29 Vbias 0.34318f
C4852 Nand_Gate_1.A.n31 Vbias 0.04546f
C4853 Nand_Gate_1.A.n32 Vbias 0.02608f
C4854 Nand_Gate_1.A.t0 Vbias 0.03876f
C4855 Nand_Gate_1.A.t1 Vbias 0.03797f
C4856 Nand_Gate_1.A.n33 Vbias 0.21593f
C4857 Nand_Gate_1.A.n34 Vbias 0.07184f
C4858 Nand_Gate_1.A.t3 Vbias 0.03797f
C4859 Nand_Gate_1.A.n35 Vbias 0.05849f
C4860 Nand_Gate_1.A.n36 Vbias 0.10356f
C4861 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t1 Vbias 0.0608f
C4862 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C4863 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C4864 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t3 Vbias 0.24183f
C4865 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C4866 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C4867 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t4 Vbias 0.46511f
C4868 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C4869 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C4870 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C4871 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C4872 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C4873 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C4874 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t2 Vbias 0.06323f
C4875 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C4876 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C4877 RingCounter_0.D_FlipFlop_11.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C4878 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t1 Vbias 0.0608f
C4879 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C4880 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C4881 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C4882 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C4883 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C4884 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C4885 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C4886 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C4887 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C4888 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C4889 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C4890 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C4891 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t2 Vbias 0.06323f
C4892 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C4893 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C4894 RingCounter_0.D_FlipFlop_10.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C4895 Q2.t9 Vbias 0.11806f
C4896 Q2.n0 Vbias 0.03449f
C4897 Q2.n1 Vbias 0.01496f
C4898 Q2.n2 Vbias 0.06579f
C4899 Q2.t8 Vbias 0.05415f
C4900 Q2.t1 Vbias 0.0154f
C4901 Q2.n3 Vbias 0.07552f
C4902 Q2.n4 Vbias 0.01853f
C4903 Q2.t0 Vbias 0.01635f
C4904 Q2.t3 Vbias 0.01601f
C4905 Q2.n5 Vbias 0.09106f
C4906 Q2.n6 Vbias 0.0303f
C4907 Q2.t2 Vbias 0.01601f
C4908 Q2.n7 Vbias 0.02467f
C4909 Q2.n8 Vbias 0.0409f
C4910 Q2.n9 Vbias 0.01975f
C4911 Q2.n11 Vbias 0.03836f
C4912 Q2.n12 Vbias 5.50481f
C4913 Q2.t4 Vbias 0.06148f
C4914 Q2.t7 Vbias 0.11836f
C4915 Q2.t5 Vbias 0.06148f
C4916 Q2.n13 Vbias 0.09576f
C4917 Q2.n14 Vbias 0.09631f
C4918 Q2.t6 Vbias 0.10522f
C4919 Q2.n15 Vbias 1.21113f
C4920 And_Gate_4.A.t2 Vbias 0.07612f
C4921 And_Gate_4.A.t1 Vbias 0.09059f
C4922 And_Gate_4.A.n0 Vbias 0.45787f
C4923 Nand_Gate_0.Vout Vbias -0.1466f
C4924 And_Gate_4.A.n1 Vbias 0.23199f
C4925 And_Gate_4.A.n2 Vbias 0.07886f
C4926 And_Gate_4.A.t3 Vbias 0.29114f
C4927 And_Gate_4.Nand_Gate_0.A Vbias -0.21888f
C4928 And_Gate_4.A.n3 Vbias 0.28519f
C4929 And_Gate_4.A.n4 Vbias 0.06015f
C4930 And_Gate_4.A.t4 Vbias 0.55994f
C4931 And_Gate_4.A.n5 Vbias 0.16357f
C4932 And_Gate_4.A.n6 Vbias 0.0407f
C4933 And_Gate_4.A.n7 Vbias 0.05921f
C4934 And_Gate_4.A.n8 Vbias 1.13762f
C4935 And_Gate_4.A.n9 Vbias 1.13762f
C4936 And_Gate_4.A.n10 Vbias 0.08035f
C4937 And_Gate_4.A.n11 Vbias 0.0415f
C4938 And_Gate_4.A.t0 Vbias 0.07306f
C4939 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t2 Vbias 0.06358f
C4940 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n0 Vbias 0.03611f
C4941 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n1 Vbias 0.06992f
C4942 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t4 Vbias 0.25335f
C4943 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n2 Vbias 0.24817f
C4944 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n3 Vbias 0.05234f
C4945 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t3 Vbias 0.48726f
C4946 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n4 Vbias 0.14234f
C4947 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n5 Vbias 0.03542f
C4948 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n6 Vbias 0.05152f
C4949 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n7 Vbias 0.13202f
C4950 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C4951 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n9 Vbias 0.06862f
C4952 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t0 Vbias 0.06624f
C4953 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.t1 Vbias 0.07883f
C4954 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n10 Vbias 0.39844f
C4955 RingCounter_0.D_FlipFlop_4.Nand_Gate_1.Vout.n11 Vbias 0.20187f
C4956 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t6 Vbias 0.45666f
C4957 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n0 Vbias 0.47347f
C4958 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n1 Vbias 0.05122f
C4959 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n2 Vbias 0.06839f
C4960 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t7 Vbias 0.22727f
C4961 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t2 Vbias 0.06194f
C4962 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n3 Vbias 0.39067f
C4963 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t3 Vbias 0.06323f
C4964 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t1 Vbias 0.06194f
C4965 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n4 Vbias 0.35224f
C4966 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n5 Vbias 0.11629f
C4967 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n6 Vbias 0.16533f
C4968 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n7 Vbias 0.06431f
C4969 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t4 Vbias 0.23742f
C4970 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t5 Vbias 0.45664f
C4971 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n8 Vbias 0.1334f
C4972 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n9 Vbias 0.05705f
C4973 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n10 Vbias 0.10533f
C4974 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n11 Vbias 0.18236f
C4975 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n12 Vbias 0.13574f
C4976 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n13 Vbias 0.12257f
C4977 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.n14 Vbias 0.0577f
C4978 RingCounter_0.D_FlipFlop_4.3-input-nand_2.C.t0 Vbias 0.05958f
C4979 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t2 Vbias 0.07037f
C4980 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n0 Vbias 0.16004f
C4981 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n1 Vbias 0.07725f
C4982 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t5 Vbias 0.2799f
C4983 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n2 Vbias 0.27418f
C4984 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n3 Vbias 0.05783f
C4985 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t4 Vbias 0.53832f
C4986 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n4 Vbias 0.15726f
C4987 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n5 Vbias 0.03913f
C4988 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n6 Vbias 0.05692f
C4989 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n7 Vbias 0.14585f
C4990 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n8 Vbias 0.14585f
C4991 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n9 Vbias 0.07581f
C4992 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t3 Vbias 0.07318f
C4993 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t0 Vbias 0.07454f
C4994 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.t1 Vbias 0.07302f
C4995 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n10 Vbias 0.41525f
C4996 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n11 Vbias 0.23391f
C4997 RingCounter_0.D_FlipFlop_12.3-input-nand_1.Vout.n12 Vbias 0.22303f
C4998 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t2 Vbias 0.07024f
C4999 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n0 Vbias 0.03989f
C5000 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n1 Vbias 0.07725f
C5001 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t5 Vbias 0.2799f
C5002 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n2 Vbias 0.27418f
C5003 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n3 Vbias 0.05783f
C5004 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t4 Vbias 0.53832f
C5005 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n4 Vbias 0.15726f
C5006 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n5 Vbias 0.03913f
C5007 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n6 Vbias 0.05692f
C5008 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n7 Vbias 0.14585f
C5009 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n8 Vbias 0.14585f
C5010 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n9 Vbias 0.07581f
C5011 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t3 Vbias 0.07318f
C5012 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t0 Vbias 0.07454f
C5013 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.t1 Vbias 0.07302f
C5014 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n10 Vbias 0.41525f
C5015 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n11 Vbias 0.23391f
C5016 RingCounter_0.D_FlipFlop_2.3-input-nand_1.Vout.n12 Vbias 0.22303f
C5017 And_Gate_2.Vout.t1 Vbias 0.10621f
C5018 And_Gate_2.Inverter_0.Vout Vbias 0.03085f
C5019 And_Gate_2.Vout.n0 Vbias 0.11719f
C5020 And_Gate_2.Vout.t7 Vbias 0.81407f
C5021 D_FlipFlop_5.3-input-nand_0.C Vbias -0.48397f
C5022 And_Gate_2.Vout.n1 Vbias 0.84403f
C5023 And_Gate_2.Vout.n2 Vbias 0.09131f
C5024 And_Gate_2.Vout.n3 Vbias 0.12192f
C5025 And_Gate_2.Vout.t4 Vbias 0.37472f
C5026 D_FlipFlop_5.CLK Vbias -0.0253f
C5027 And_Gate_2.Vout.n4 Vbias 0.294f
C5028 And_Gate_2.Vout.t3 Vbias 0.81403f
C5029 D_FlipFlop_5.3-input-nand_1.C Vbias -0.2721f
C5030 And_Gate_2.Vout.t5 Vbias 0.42325f
C5031 D_FlipFlop_5.Inverter_1.Vin Vbias -0.26427f
C5032 And_Gate_2.Vout.n5 Vbias 0.44634f
C5033 And_Gate_2.Vout.t2 Vbias 0.81403f
C5034 And_Gate_2.Vout.n6 Vbias 0.72059f
C5035 And_Gate_2.Vout.n7 Vbias 0.72257f
C5036 And_Gate_2.Vout.n8 Vbias 0.45218f
C5037 And_Gate_2.Vout.t6 Vbias 0.37471f
C5038 And_Gate_2.Vout.n9 Vbias 0.07492f
C5039 And_Gate_2.Vout.n10 Vbias 0.17642f
C5040 And_Gate_2.Vout.n11 Vbias 11.6967f
C5041 And_Gate_2.Vout.t0 Vbias 0.11091f
C5042 And_Gate_2.Vout.n12 Vbias 9.27182f
C5043 And_Gate_2.Vout.n13 Vbias 0.2528f
C5044 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t7 Vbias 0.36784f
C5045 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n0 Vbias 0.10746f
C5046 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n1 Vbias 0.04662f
C5047 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t2 Vbias 0.04798f
C5048 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n2 Vbias 0.22815f
C5049 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n3 Vbias 0.0518f
C5050 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t4 Vbias 0.36785f
C5051 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n4 Vbias 0.38072f
C5052 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t6 Vbias 0.19125f
C5053 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n5 Vbias 0.18752f
C5054 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n6 Vbias 0.10934f
C5055 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n7 Vbias 0.01378f
C5056 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n8 Vbias 0.01506f
C5057 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t0 Vbias 0.05094f
C5058 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t3 Vbias 0.04989f
C5059 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n9 Vbias 0.28374f
C5060 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n10 Vbias 0.09441f
C5061 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t1 Vbias 0.04989f
C5062 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n11 Vbias 0.31407f
C5063 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.t5 Vbias 0.1838f
C5064 RingCounter_0.D_FlipFlop_14.3-input-nand_2.Vout.n12 Vbias 0.205f
C5065 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t3 Vbias 0.07037f
C5066 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n0 Vbias 0.16004f
C5067 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n1 Vbias 0.07725f
C5068 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t5 Vbias 0.2799f
C5069 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n2 Vbias 0.27418f
C5070 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n3 Vbias 0.05783f
C5071 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t4 Vbias 0.53832f
C5072 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n4 Vbias 0.15726f
C5073 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n5 Vbias 0.03913f
C5074 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n6 Vbias 0.05692f
C5075 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n7 Vbias 0.14585f
C5076 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n8 Vbias 0.14585f
C5077 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n9 Vbias 0.07581f
C5078 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t2 Vbias 0.07318f
C5079 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t0 Vbias 0.07454f
C5080 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.t1 Vbias 0.07302f
C5081 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n10 Vbias 0.41525f
C5082 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n11 Vbias 0.23391f
C5083 RingCounter_0.D_FlipFlop_13.3-input-nand_1.Vout.n12 Vbias 0.22303f
C5084 D_FlipFlop_5.3-input-nand_2.Vout.t4 Vbias 0.35515f
C5085 D_FlipFlop_5.3-input-nand_2.Vout.n0 Vbias 0.10375f
C5086 D_FlipFlop_5.3-input-nand_2.Vout.n1 Vbias 0.04502f
C5087 D_FlipFlop_5.3-input-nand_2.Vout.t1 Vbias 0.04632f
C5088 D_FlipFlop_5.3-input-nand_2.Vout.n2 Vbias 0.22028f
C5089 D_FlipFlop_5.3-input-nand_2.Vout.n3 Vbias 0.05002f
C5090 D_FlipFlop_5.3-input-nand_2.Vout.t7 Vbias 0.35517f
C5091 D_FlipFlop_5.3-input-nand_2.Vout.n4 Vbias 0.36759f
C5092 D_FlipFlop_5.3-input-nand_2.Vout.t5 Vbias 0.18465f
C5093 D_FlipFlop_5.3-input-nand_2.Vout.n5 Vbias 0.18106f
C5094 D_FlipFlop_5.3-input-nand_2.Vout.n6 Vbias 0.10557f
C5095 D_FlipFlop_5.3-input-nand_2.Vout.n7 Vbias 0.01331f
C5096 D_FlipFlop_5.3-input-nand_2.Vout.n8 Vbias 0.01454f
C5097 D_FlipFlop_5.3-input-nand_2.Vout.t0 Vbias 0.04918f
C5098 D_FlipFlop_5.3-input-nand_2.Vout.t3 Vbias 0.04817f
C5099 D_FlipFlop_5.3-input-nand_2.Vout.n9 Vbias 0.27396f
C5100 D_FlipFlop_5.3-input-nand_2.Vout.n10 Vbias 0.09115f
C5101 D_FlipFlop_5.3-input-nand_2.Vout.t2 Vbias 0.04817f
C5102 D_FlipFlop_5.3-input-nand_2.Vout.n11 Vbias 0.30324f
C5103 D_FlipFlop_5.3-input-nand_2.Vout.t6 Vbias 0.17747f
C5104 D_FlipFlop_5.3-input-nand_2.Vout.n12 Vbias 0.19793f
C5105 Nand_Gate_7.A.t10 Vbias 0.27993f
C5106 Nand_Gate_7.A.n0 Vbias 0.08177f
C5107 Nand_Gate_7.A.n1 Vbias 0.03548f
C5108 Nand_Gate_7.A.n2 Vbias 0.15601f
C5109 Nand_Gate_7.A.t6 Vbias 0.1302f
C5110 Nand_Gate_7.A.n3 Vbias 0.04085f
C5111 Nand_Gate_7.A.t2 Vbias 0.03651f
C5112 Nand_Gate_7.A.n4 Vbias 0.159f
C5113 Nand_Gate_7.A.n5 Vbias 0.03942f
C5114 Nand_Gate_7.A.t7 Vbias 0.27994f
C5115 Nand_Gate_7.A.n6 Vbias 0.27511f
C5116 Nand_Gate_7.A.n7 Vbias 0.03007f
C5117 Nand_Gate_7.A.t5 Vbias 0.14554f
C5118 Nand_Gate_7.A.n8 Vbias 0.04192f
C5119 Nand_Gate_7.A.n9 Vbias 0.01797f
C5120 Nand_Gate_7.A.n10 Vbias 0.03367f
C5121 Nand_Gate_7.A.n11 Vbias 0.04236f
C5122 Nand_Gate_7.A.t4 Vbias 0.27994f
C5123 Nand_Gate_7.A.n12 Vbias 0.27511f
C5124 Nand_Gate_7.A.n13 Vbias 0.03007f
C5125 Nand_Gate_7.A.t8 Vbias 0.14554f
C5126 Nand_Gate_7.A.n14 Vbias 0.04192f
C5127 Nand_Gate_7.A.n15 Vbias 0.01797f
C5128 Nand_Gate_7.A.n16 Vbias 0.03367f
C5129 Nand_Gate_7.A.n18 Vbias 0.12703f
C5130 Nand_Gate_7.A.n19 Vbias 0.0915f
C5131 Nand_Gate_7.A.t9 Vbias 0.14555f
C5132 Nand_Gate_7.A.n20 Vbias 0.14257f
C5133 Nand_Gate_7.A.n21 Vbias 0.03007f
C5134 Nand_Gate_7.A.t11 Vbias 0.27993f
C5135 Nand_Gate_7.A.n22 Vbias 0.08177f
C5136 Nand_Gate_7.A.n23 Vbias 0.02035f
C5137 Nand_Gate_7.A.n24 Vbias 0.0296f
C5138 Nand_Gate_7.A.n25 Vbias 0.14551f
C5139 Nand_Gate_7.A.n26 Vbias 0.25531f
C5140 Nand_Gate_7.A.n27 Vbias 0.15839f
C5141 Nand_Gate_7.A.n28 Vbias 0.34271f
C5142 Nand_Gate_7.A.n30 Vbias 0.04546f
C5143 Nand_Gate_7.A.n31 Vbias 0.02608f
C5144 Nand_Gate_7.A.t0 Vbias 0.03876f
C5145 Nand_Gate_7.A.t3 Vbias 0.03797f
C5146 Nand_Gate_7.A.n32 Vbias 0.21593f
C5147 Nand_Gate_7.A.n33 Vbias 0.07184f
C5148 Nand_Gate_7.A.t1 Vbias 0.03797f
C5149 Nand_Gate_7.A.n34 Vbias 0.05849f
C5150 Nand_Gate_7.A.n35 Vbias 0.10356f
C5151 Nand_Gate_1.Vout.t1 Vbias 0.08532f
C5152 Nand_Gate_1.Vout.t2 Vbias 0.10154f
C5153 Nand_Gate_1.Vout.n0 Vbias 0.51322f
C5154 Nand_Gate_1.Vout.n1 Vbias 0.26003f
C5155 Nand_Gate_1.Vout.n2 Vbias 0.08839f
C5156 Nand_Gate_1.Vout.t4 Vbias 0.32633f
C5157 Nand_Gate_1.Vout.n3 Vbias 0.31966f
C5158 Nand_Gate_1.Vout.n4 Vbias 0.06742f
C5159 Nand_Gate_1.Vout.t3 Vbias 0.62762f
C5160 Nand_Gate_1.Vout.n5 Vbias 0.18335f
C5161 Nand_Gate_1.Vout.n6 Vbias 0.04562f
C5162 Nand_Gate_1.Vout.n7 Vbias 0.06636f
C5163 Nand_Gate_1.Vout.n8 Vbias 1.35316f
C5164 Nand_Gate_1.Vout.n9 Vbias 1.35316f
C5165 Nand_Gate_1.Vout.n10 Vbias 0.09007f
C5166 Nand_Gate_1.Vout.n11 Vbias 0.04651f
C5167 Nand_Gate_1.Vout.t0 Vbias 0.08189f
C5168 D_FlipFlop_7.3-input-nand_2.Vout.t4 Vbias 0.35515f
C5169 D_FlipFlop_7.3-input-nand_2.Vout.n0 Vbias 0.10375f
C5170 D_FlipFlop_7.3-input-nand_2.Vout.n1 Vbias 0.04502f
C5171 D_FlipFlop_7.3-input-nand_2.Vout.t2 Vbias 0.04632f
C5172 D_FlipFlop_7.3-input-nand_2.Vout.n2 Vbias 0.22028f
C5173 D_FlipFlop_7.3-input-nand_2.Vout.n3 Vbias 0.05002f
C5174 D_FlipFlop_7.3-input-nand_2.Vout.t7 Vbias 0.35517f
C5175 D_FlipFlop_7.3-input-nand_2.Vout.n4 Vbias 0.36759f
C5176 D_FlipFlop_7.3-input-nand_2.Vout.t5 Vbias 0.18465f
C5177 D_FlipFlop_7.3-input-nand_2.Vout.n5 Vbias 0.18106f
C5178 D_FlipFlop_7.3-input-nand_2.Vout.n6 Vbias 0.10557f
C5179 D_FlipFlop_7.3-input-nand_2.Vout.n7 Vbias 0.01331f
C5180 D_FlipFlop_7.3-input-nand_2.Vout.n8 Vbias 0.01454f
C5181 D_FlipFlop_7.3-input-nand_2.Vout.t1 Vbias 0.04918f
C5182 D_FlipFlop_7.3-input-nand_2.Vout.t0 Vbias 0.04817f
C5183 D_FlipFlop_7.3-input-nand_2.Vout.n9 Vbias 0.27396f
C5184 D_FlipFlop_7.3-input-nand_2.Vout.n10 Vbias 0.09115f
C5185 D_FlipFlop_7.3-input-nand_2.Vout.t3 Vbias 0.04817f
C5186 D_FlipFlop_7.3-input-nand_2.Vout.n11 Vbias 0.30324f
C5187 D_FlipFlop_7.3-input-nand_2.Vout.t6 Vbias 0.17747f
C5188 D_FlipFlop_7.3-input-nand_2.Vout.n12 Vbias 0.19793f
C5189 D_FlipFlop_7.3-input-nand_2.C.t7 Vbias 0.3425f
C5190 D_FlipFlop_7.3-input-nand_2.C.n0 Vbias 0.3551f
C5191 D_FlipFlop_7.3-input-nand_2.C.n1 Vbias 0.03842f
C5192 D_FlipFlop_7.3-input-nand_2.C.t1 Vbias 0.04477f
C5193 D_FlipFlop_7.3-input-nand_2.C.n2 Vbias 0.11971f
C5194 D_FlipFlop_7.3-input-nand_2.C.n3 Vbias 0.09193f
C5195 D_FlipFlop_7.3-input-nand_2.C.t5 Vbias 0.17806f
C5196 D_FlipFlop_7.3-input-nand_2.C.t6 Vbias 0.34248f
C5197 D_FlipFlop_7.3-input-nand_2.C.n4 Vbias 0.10005f
C5198 D_FlipFlop_7.3-input-nand_2.C.n5 Vbias 0.04279f
C5199 D_FlipFlop_7.3-input-nand_2.C.n6 Vbias 0.079f
C5200 D_FlipFlop_7.3-input-nand_2.C.n7 Vbias 0.13677f
C5201 D_FlipFlop_7.3-input-nand_2.C.n8 Vbias 0.10181f
C5202 D_FlipFlop_7.3-input-nand_2.C.n9 Vbias 0.04823f
C5203 D_FlipFlop_7.3-input-nand_2.C.n10 Vbias 0.124f
C5204 D_FlipFlop_7.3-input-nand_2.C.t3 Vbias 0.04742f
C5205 D_FlipFlop_7.3-input-nand_2.C.t0 Vbias 0.04645f
C5206 D_FlipFlop_7.3-input-nand_2.C.n11 Vbias 0.26418f
C5207 D_FlipFlop_7.3-input-nand_2.C.n12 Vbias 0.08722f
C5208 D_FlipFlop_7.3-input-nand_2.C.t2 Vbias 0.04645f
C5209 D_FlipFlop_7.3-input-nand_2.C.n13 Vbias 0.293f
C5210 D_FlipFlop_7.3-input-nand_2.C.t4 Vbias 0.17045f
C5211 D_FlipFlop_7.3-input-nand_2.C.n14 Vbias 0.05129f
C5212 Q5.t0 Vbias 0.01626f
C5213 Q5.n0 Vbias 0.07974f
C5214 Q5.n1 Vbias 0.01957f
C5215 Q5.t3 Vbias 0.01726f
C5216 Q5.t2 Vbias 0.01691f
C5217 Q5.n2 Vbias 0.09616f
C5218 Q5.n3 Vbias 0.03199f
C5219 Q5.t1 Vbias 0.01691f
C5220 Q5.n4 Vbias 0.02605f
C5221 Q5.n5 Vbias 0.03693f
C5222 Q5.n6 Vbias 0.0192f
C5223 Q5.t8 Vbias 0.12466f
C5224 Q5.n7 Vbias 0.03642f
C5225 Q5.n8 Vbias 0.0158f
C5226 Q5.n9 Vbias 0.06947f
C5227 Q5.t9 Vbias 0.05798f
C5228 Q5.n11 Vbias 0.0161f
C5229 Q5.n13 Vbias 3.34141f
C5230 Q5.t6 Vbias 0.12498f
C5231 Q5.t7 Vbias 0.12498f
C5232 Q5.t5 Vbias 0.06492f
C5233 Q5.n14 Vbias 0.10112f
C5234 Q5.n15 Vbias 0.1017f
C5235 Q5.t4 Vbias 0.05702f
C5236 Q5.n16 Vbias 1.27887f
C5237 And_Gate_5.Vout.t1 Vbias 0.12948f
C5238 And_Gate_5.Inverter_0.Vout Vbias -0.41618f
C5239 And_Gate_5.Vout.n0 Vbias 0.07354f
C5240 And_Gate_5.Vout.n1 Vbias 0.1424f
C5241 And_Gate_5.Vout.t3 Vbias 0.99235f
C5242 D_FlipFlop_1.3-input-nand_0.C Vbias -0.58996f
C5243 And_Gate_5.Vout.n2 Vbias 1.02888f
C5244 And_Gate_5.Vout.n3 Vbias 0.11131f
C5245 And_Gate_5.Vout.n4 Vbias 0.14862f
C5246 And_Gate_5.Vout.t6 Vbias 0.45675f
C5247 D_FlipFlop_1.CLK Vbias 0.04947f
C5248 And_Gate_5.Vout.n5 Vbias 0.43118f
C5249 And_Gate_5.Vout.n6 Vbias 0.13081f
C5250 And_Gate_5.Vout.t5 Vbias 0.99231f
C5251 D_FlipFlop_1.3-input-nand_1.C Vbias -0.33169f
C5252 And_Gate_5.Vout.t7 Vbias 0.51595f
C5253 D_FlipFlop_1.Inverter_1.Vin Vbias -0.32215f
C5254 And_Gate_5.Vout.n7 Vbias 0.54409f
C5255 And_Gate_5.Vout.t4 Vbias 0.99231f
C5256 And_Gate_5.Vout.n8 Vbias 0.87841f
C5257 And_Gate_5.Vout.n9 Vbias 0.88082f
C5258 And_Gate_5.Vout.n10 Vbias 0.55121f
C5259 And_Gate_5.Vout.t2 Vbias 0.45677f
C5260 And_Gate_5.Vout.n11 Vbias 0.0213f
C5261 And_Gate_5.Vout.n12 Vbias 24.0152f
C5262 And_Gate_5.Vout.n13 Vbias 21.6425f
C5263 And_Gate_5.Vout.n14 Vbias 0.13974f
C5264 And_Gate_5.Vout.t0 Vbias 0.13492f
C5265 And_Gate_5.Vout.n15 Vbias 0.79964f
C5266 Q7.t0 Vbias 0.01626f
C5267 Q7.n0 Vbias 0.07974f
C5268 Q7.n1 Vbias 0.01957f
C5269 Q7.t3 Vbias 0.01726f
C5270 Q7.t2 Vbias 0.01691f
C5271 Q7.n2 Vbias 0.09616f
C5272 Q7.n3 Vbias 0.03199f
C5273 Q7.t1 Vbias 0.01691f
C5274 Q7.n4 Vbias 0.02605f
C5275 Q7.n5 Vbias 0.03769f
C5276 Q7.n6 Vbias 0.0192f
C5277 Q7.t5 Vbias 0.12466f
C5278 Q7.n7 Vbias 0.03642f
C5279 Q7.n8 Vbias 0.0158f
C5280 Q7.n9 Vbias 0.06947f
C5281 Q7.t6 Vbias 0.05798f
C5282 Q7.n11 Vbias 0.01451f
C5283 Q7.n13 Vbias 3.34141f
C5284 Q7.t7 Vbias 0.12498f
C5285 Q7.t8 Vbias 0.12498f
C5286 Q7.t4 Vbias 0.06492f
C5287 Q7.n14 Vbias 0.10112f
C5288 Q7.n15 Vbias 0.1017f
C5289 Q7.t9 Vbias 0.05702f
C5290 Q7.n16 Vbias 1.27887f
C5291 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t1 Vbias 0.07024f
C5292 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n0 Vbias 0.03989f
C5293 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n1 Vbias 0.07725f
C5294 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t5 Vbias 0.2799f
C5295 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n2 Vbias 0.27418f
C5296 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n3 Vbias 0.05783f
C5297 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t4 Vbias 0.53832f
C5298 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n4 Vbias 0.15726f
C5299 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n5 Vbias 0.03913f
C5300 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n6 Vbias 0.05692f
C5301 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n7 Vbias 0.14585f
C5302 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n8 Vbias 0.14585f
C5303 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n9 Vbias 0.07581f
C5304 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t2 Vbias 0.07318f
C5305 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t0 Vbias 0.07454f
C5306 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.t3 Vbias 0.07302f
C5307 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n10 Vbias 0.41525f
C5308 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n11 Vbias 0.23391f
C5309 RingCounter_0.D_FlipFlop_5.3-input-nand_1.Vout.n12 Vbias 0.22303f
C5310 Nand_Gate_1.B.t13 Vbias 0.47211f
C5311 Nand_Gate_1.B.n0 Vbias 0.13792f
C5312 Nand_Gate_1.B.n1 Vbias 0.05984f
C5313 Nand_Gate_1.B.n2 Vbias 0.26311f
C5314 Nand_Gate_1.B.t16 Vbias 0.21959f
C5315 Nand_Gate_1.B.n3 Vbias 0.06889f
C5316 Nand_Gate_1.B.t1 Vbias 0.06158f
C5317 Nand_Gate_1.B.n4 Vbias 0.26816f
C5318 Nand_Gate_1.B.n5 Vbias 0.06649f
C5319 Nand_Gate_1.B.t10 Vbias 0.47213f
C5320 Nand_Gate_1.B.n6 Vbias 0.46399f
C5321 Nand_Gate_1.B.n7 Vbias 0.05071f
C5322 Nand_Gate_1.B.t6 Vbias 0.24546f
C5323 Nand_Gate_1.B.n8 Vbias 0.07071f
C5324 Nand_Gate_1.B.n9 Vbias 0.0303f
C5325 Nand_Gate_1.B.n10 Vbias 0.05678f
C5326 Nand_Gate_1.B.n11 Vbias 0.07145f
C5327 Nand_Gate_1.B.t5 Vbias 0.47213f
C5328 Nand_Gate_1.B.n12 Vbias 0.46399f
C5329 Nand_Gate_1.B.n13 Vbias 0.05071f
C5330 Nand_Gate_1.B.t11 Vbias 0.24546f
C5331 Nand_Gate_1.B.n14 Vbias 0.07071f
C5332 Nand_Gate_1.B.n15 Vbias 0.0303f
C5333 Nand_Gate_1.B.n16 Vbias 0.05678f
C5334 Nand_Gate_1.B.n18 Vbias 0.21345f
C5335 Nand_Gate_1.B.n19 Vbias 0.05834f
C5336 Nand_Gate_1.B.n20 Vbias 0.15524f
C5337 Nand_Gate_1.B.t15 Vbias 0.47213f
C5338 Nand_Gate_1.B.n21 Vbias 0.47546f
C5339 Nand_Gate_1.B.n22 Vbias 0.05071f
C5340 Nand_Gate_1.B.t14 Vbias 0.24546f
C5341 Nand_Gate_1.B.n23 Vbias 0.07071f
C5342 Nand_Gate_1.B.n24 Vbias 0.01883f
C5343 Nand_Gate_1.B.n25 Vbias 0.02935f
C5344 Nand_Gate_1.B.n26 Vbias 0.29279f
C5345 Nand_Gate_1.B.t8 Vbias 0.47213f
C5346 Nand_Gate_1.B.n27 Vbias 0.47546f
C5347 Nand_Gate_1.B.n28 Vbias 0.05071f
C5348 Nand_Gate_1.B.t7 Vbias 0.24546f
C5349 Nand_Gate_1.B.n29 Vbias 0.07071f
C5350 Nand_Gate_1.B.n30 Vbias 0.01883f
C5351 Nand_Gate_1.B.n31 Vbias 0.02935f
C5352 Nand_Gate_1.B.n33 Vbias 0.76027f
C5353 Nand_Gate_1.B.n34 Vbias 0.31374f
C5354 Nand_Gate_1.B.n35 Vbias 0.13131f
C5355 Nand_Gate_1.B.t17 Vbias 0.47211f
C5356 Nand_Gate_1.B.n36 Vbias 0.13792f
C5357 Nand_Gate_1.B.n37 Vbias 0.05984f
C5358 Nand_Gate_1.B.n38 Vbias 0.26311f
C5359 Nand_Gate_1.B.t9 Vbias 0.21957f
C5360 Nand_Gate_1.B.n39 Vbias 0.06876f
C5361 Nand_Gate_1.B.n40 Vbias 0.15969f
C5362 Nand_Gate_1.B.n41 Vbias 3.82373f
C5363 Nand_Gate_1.B.t4 Vbias 0.24547f
C5364 Nand_Gate_1.B.n42 Vbias 0.26225f
C5365 Nand_Gate_1.B.t12 Vbias 0.47211f
C5366 Nand_Gate_1.B.n43 Vbias 1.07465f
C5367 Nand_Gate_1.B.n44 Vbias 5.83655f
C5368 Nand_Gate_1.B.n45 Vbias 0.08001f
C5369 Nand_Gate_1.B.n46 Vbias 0.26771f
C5370 Nand_Gate_1.B.n47 Vbias 0.5788f
C5371 Nand_Gate_1.B.n49 Vbias 0.07667f
C5372 Nand_Gate_1.B.n50 Vbias 0.04399f
C5373 Nand_Gate_1.B.t0 Vbias 0.06538f
C5374 Nand_Gate_1.B.t3 Vbias 0.06404f
C5375 Nand_Gate_1.B.n51 Vbias 0.36418f
C5376 Nand_Gate_1.B.n52 Vbias 0.12117f
C5377 Nand_Gate_1.B.t2 Vbias 0.06404f
C5378 Nand_Gate_1.B.n53 Vbias 0.09864f
C5379 Nand_Gate_1.B.n54 Vbias 0.17466f
C5380 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t1 Vbias 0.04998f
C5381 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n0 Vbias 0.02839f
C5382 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n1 Vbias 0.05497f
C5383 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t2 Vbias 0.38308f
C5384 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n2 Vbias 0.39717f
C5385 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n3 Vbias 0.04297f
C5386 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n4 Vbias 0.05737f
C5387 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t3 Vbias 0.30118f
C5388 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t5 Vbias 0.30119f
C5389 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n5 Vbias 0.1951f
C5390 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n6 Vbias 0.04115f
C5391 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t4 Vbias 0.38306f
C5392 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n7 Vbias 0.1119f
C5393 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n8 Vbias 0.02784f
C5394 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n9 Vbias 0.0405f
C5395 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n10 Vbias 0.10379f
C5396 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n11 Vbias 0.10379f
C5397 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n12 Vbias 0.05395f
C5398 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.t0 Vbias 0.05208f
C5399 RingCounter_0.D_FlipFlop_3.Inverter_1.Vout.n13 Vbias 0.30868f
C5400 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t7 Vbias 0.36784f
C5401 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n0 Vbias 0.10746f
C5402 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n1 Vbias 0.04662f
C5403 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t2 Vbias 0.04798f
C5404 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n2 Vbias 0.22815f
C5405 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n3 Vbias 0.0518f
C5406 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t5 Vbias 0.36785f
C5407 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n4 Vbias 0.38072f
C5408 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t4 Vbias 0.19125f
C5409 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n5 Vbias 0.18752f
C5410 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n6 Vbias 0.10934f
C5411 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n7 Vbias 0.01378f
C5412 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n8 Vbias 0.01095f
C5413 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t0 Vbias 0.05094f
C5414 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t3 Vbias 0.04989f
C5415 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n9 Vbias 0.28374f
C5416 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n10 Vbias 0.09258f
C5417 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t1 Vbias 0.04989f
C5418 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n11 Vbias 0.31407f
C5419 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.t6 Vbias 0.1838f
C5420 RingCounter_0.D_FlipFlop_2.3-input-nand_2.Vout.n12 Vbias 0.205f
C5421 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t1 Vbias 0.04607f
C5422 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n0 Vbias 0.10477f
C5423 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n1 Vbias 0.05057f
C5424 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t4 Vbias 0.35243f
C5425 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n2 Vbias 0.3654f
C5426 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n3 Vbias 0.03953f
C5427 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n4 Vbias 0.05278f
C5428 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t3 Vbias 0.27708f
C5429 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t2 Vbias 0.27709f
C5430 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n5 Vbias 0.17949f
C5431 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n6 Vbias 0.03786f
C5432 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t5 Vbias 0.35241f
C5433 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n7 Vbias 0.10295f
C5434 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n8 Vbias 0.02562f
C5435 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n9 Vbias 0.03726f
C5436 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n10 Vbias 0.09548f
C5437 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n11 Vbias 0.09548f
C5438 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n12 Vbias 0.04963f
C5439 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.t0 Vbias 0.04792f
C5440 RingCounter_0.D_FlipFlop_8.Inverter_1.Vout.n13 Vbias 0.28399f
C5441 Nand_Gate_3.B.t9 Vbias 0.33127f
C5442 Nand_Gate_3.B.n0 Vbias 0.09677f
C5443 Nand_Gate_3.B.n1 Vbias 0.04199f
C5444 Nand_Gate_3.B.n2 Vbias 0.18462f
C5445 Nand_Gate_3.B.t7 Vbias 0.15408f
C5446 Nand_Gate_3.B.n3 Vbias 0.04834f
C5447 Nand_Gate_3.B.t2 Vbias 0.04321f
C5448 Nand_Gate_3.B.n4 Vbias 0.18816f
C5449 Nand_Gate_3.B.n5 Vbias 0.04665f
C5450 Nand_Gate_3.B.t11 Vbias 0.33129f
C5451 Nand_Gate_3.B.n6 Vbias 0.32557f
C5452 Nand_Gate_3.B.n7 Vbias 0.03558f
C5453 Nand_Gate_3.B.t5 Vbias 0.17224f
C5454 Nand_Gate_3.B.n8 Vbias 0.04961f
C5455 Nand_Gate_3.B.n9 Vbias 0.02126f
C5456 Nand_Gate_3.B.n10 Vbias 0.03984f
C5457 Nand_Gate_3.B.n11 Vbias 0.05014f
C5458 Nand_Gate_3.B.t4 Vbias 0.33129f
C5459 Nand_Gate_3.B.n12 Vbias 0.32557f
C5460 Nand_Gate_3.B.n13 Vbias 0.03558f
C5461 Nand_Gate_3.B.t10 Vbias 0.17224f
C5462 Nand_Gate_3.B.n14 Vbias 0.04961f
C5463 Nand_Gate_3.B.n15 Vbias 0.02126f
C5464 Nand_Gate_3.B.n16 Vbias 0.03984f
C5465 Nand_Gate_3.B.n18 Vbias 0.15033f
C5466 Nand_Gate_3.B.n19 Vbias 0.41862f
C5467 Nand_Gate_3.B.n20 Vbias 0.18785f
C5468 Nand_Gate_3.B.t6 Vbias 0.17224f
C5469 Nand_Gate_3.B.t8 Vbias 0.33127f
C5470 Nand_Gate_3.B.n21 Vbias 0.09677f
C5471 Nand_Gate_3.B.n22 Vbias 0.04139f
C5472 Nand_Gate_3.B.n23 Vbias 0.07641f
C5473 Nand_Gate_3.B.n24 Vbias 0.87221f
C5474 Nand_Gate_3.B.n25 Vbias 1.18609f
C5475 Nand_Gate_3.B.n26 Vbias 0.05328f
C5476 Nand_Gate_3.B.n27 Vbias 0.01961f
C5477 Nand_Gate_3.B.n29 Vbias 0.05379f
C5478 Nand_Gate_3.B.n30 Vbias 0.02717f
C5479 Nand_Gate_3.B.t0 Vbias 0.04587f
C5480 Nand_Gate_3.B.t1 Vbias 0.04493f
C5481 Nand_Gate_3.B.n31 Vbias 0.25554f
C5482 Nand_Gate_3.B.n32 Vbias 0.08338f
C5483 Nand_Gate_3.B.t3 Vbias 0.04493f
C5484 Nand_Gate_3.B.n33 Vbias 0.06922f
C5485 Nand_Gate_3.B.n34 Vbias 0.12256f
C5486 Nand_Gate_2.Vout.t2 Vbias 0.07306f
C5487 Nand_Gate_2.Vout.n0 Vbias 0.0415f
C5488 Nand_Gate_2.Vout.n1 Vbias 0.08035f
C5489 Nand_Gate_2.Vout.t4 Vbias 0.29114f
C5490 Nand_Gate_2.Vout.n2 Vbias 0.28519f
C5491 Nand_Gate_2.Vout.n3 Vbias 0.06015f
C5492 Nand_Gate_2.Vout.t3 Vbias 0.55994f
C5493 Nand_Gate_2.Vout.n4 Vbias 0.16357f
C5494 Nand_Gate_2.Vout.n5 Vbias 0.0407f
C5495 Nand_Gate_2.Vout.n6 Vbias 0.05921f
C5496 Nand_Gate_2.Vout.n7 Vbias 1.13762f
C5497 Nand_Gate_2.Vout.n8 Vbias 1.13762f
C5498 Nand_Gate_2.Vout.n9 Vbias 0.07886f
C5499 Nand_Gate_2.Vout.t1 Vbias 0.07612f
C5500 Nand_Gate_2.Vout.t0 Vbias 0.09059f
C5501 Nand_Gate_2.Vout.n10 Vbias 0.45787f
C5502 Nand_Gate_2.Vout.n11 Vbias 0.23199f
C5503 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t7 Vbias 0.36784f
C5504 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n0 Vbias 0.10746f
C5505 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n1 Vbias 0.04662f
C5506 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t2 Vbias 0.04798f
C5507 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n2 Vbias 0.22815f
C5508 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n3 Vbias 0.0518f
C5509 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t5 Vbias 0.36785f
C5510 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n4 Vbias 0.38072f
C5511 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t4 Vbias 0.19125f
C5512 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n5 Vbias 0.18752f
C5513 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n6 Vbias 0.10934f
C5514 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n7 Vbias 0.01378f
C5515 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n8 Vbias 0.01095f
C5516 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t0 Vbias 0.05094f
C5517 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t1 Vbias 0.04989f
C5518 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n9 Vbias 0.28374f
C5519 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n10 Vbias 0.09258f
C5520 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t3 Vbias 0.04989f
C5521 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n11 Vbias 0.31407f
C5522 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.t6 Vbias 0.1838f
C5523 RingCounter_0.D_FlipFlop_6.3-input-nand_2.Vout.n12 Vbias 0.205f
C5524 CDAC8_0.switch_1.Z.t2 Vbias 0.0253f
C5525 CDAC8_0.switch_1.Z.t1 Vbias 0.02525f
C5526 CDAC8_0.switch_1.Z.n0 Vbias 0.05629f
C5527 CDAC8_0.switch_1.Z.n1 Vbias 0.01036f
C5528 CDAC8_0.switch_1.Z.t4 Vbias 5.82511f
C5529 CDAC8_0.switch_1.Z.n2 Vbias 0.11275f
C5530 CDAC8_0.switch_1.Z.n3 Vbias 0.02706f
C5531 CDAC8_0.switch_1.Z.t3 Vbias 0.02612f
C5532 CDAC8_0.switch_1.Z.t0 Vbias 0.02612f
C5533 CDAC8_0.switch_1.Z.n4 Vbias 0.09382f
C5534 CDAC8_0.switch_1.Z.n5 Vbias 0.28853f
C5535 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t4 Vbias 0.46931f
C5536 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n0 Vbias 0.1371f
C5537 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n1 Vbias 0.05949f
C5538 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t2 Vbias 0.06121f
C5539 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n2 Vbias 0.29108f
C5540 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n3 Vbias 0.06609f
C5541 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t6 Vbias 0.46933f
C5542 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n4 Vbias 0.48575f
C5543 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t5 Vbias 0.244f
C5544 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n5 Vbias 0.23925f
C5545 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n6 Vbias 0.13951f
C5546 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n7 Vbias 0.01758f
C5547 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n8 Vbias 0.01397f
C5548 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t0 Vbias 0.06499f
C5549 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t1 Vbias 0.06366f
C5550 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n9 Vbias 0.36201f
C5551 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n10 Vbias 0.11813f
C5552 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t3 Vbias 0.06366f
C5553 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n11 Vbias 0.40071f
C5554 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.t7 Vbias 0.23451f
C5555 RingCounter_0.D_FlipFlop_17.3-input-nand_2.Vout.n12 Vbias 0.26155f
C5556 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t1 Vbias 0.05969f
C5557 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n0 Vbias 0.15961f
C5558 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n1 Vbias 0.12257f
C5559 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t7 Vbias 0.23742f
C5560 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t4 Vbias 0.45664f
C5561 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n2 Vbias 0.1334f
C5562 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n3 Vbias 0.05705f
C5563 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n4 Vbias 0.10533f
C5564 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n5 Vbias 0.18236f
C5565 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n6 Vbias 0.13574f
C5566 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n7 Vbias 0.06431f
C5567 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t5 Vbias 0.45666f
C5568 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n8 Vbias 0.47347f
C5569 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n9 Vbias 0.05122f
C5570 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n10 Vbias 0.06839f
C5571 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t6 Vbias 0.22727f
C5572 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t0 Vbias 0.06194f
C5573 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n11 Vbias 0.39067f
C5574 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t2 Vbias 0.06323f
C5575 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.t3 Vbias 0.06194f
C5576 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n12 Vbias 0.35224f
C5577 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n13 Vbias 0.11629f
C5578 RingCounter_0.D_FlipFlop_15.3-input-nand_2.C.n14 Vbias 0.16533f
C5579 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t6 Vbias 0.36784f
C5580 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n0 Vbias 0.10746f
C5581 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n1 Vbias 0.04662f
C5582 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t1 Vbias 0.04798f
C5583 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n2 Vbias 0.22815f
C5584 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n3 Vbias 0.0518f
C5585 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t7 Vbias 0.36785f
C5586 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n4 Vbias 0.38072f
C5587 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t5 Vbias 0.19125f
C5588 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n5 Vbias 0.18752f
C5589 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n6 Vbias 0.10934f
C5590 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n7 Vbias 0.01378f
C5591 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n8 Vbias 0.01506f
C5592 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t0 Vbias 0.05094f
C5593 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t3 Vbias 0.04989f
C5594 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n9 Vbias 0.28374f
C5595 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n10 Vbias 0.09441f
C5596 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t2 Vbias 0.04989f
C5597 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n11 Vbias 0.31407f
C5598 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.t4 Vbias 0.1838f
C5599 RingCounter_0.D_FlipFlop_15.3-input-nand_2.Vout.n12 Vbias 0.205f
C5600 a_138366_35417.t1 Vbias 0.70679f
C5601 a_138366_35417.t2 Vbias 2.14691f
C5602 a_138366_35417.t3 Vbias 3.57208f
C5603 a_138366_35417.n0 Vbias 1.57769f
C5604 a_138366_35417.n1 Vbias 1.3122f
C5605 a_138366_35417.t0 Vbias 2.28434f
C5606 Q1.t8 Vbias 0.11808f
C5607 Q1.n0 Vbias 0.03449f
C5608 Q1.n1 Vbias 0.01497f
C5609 Q1.n2 Vbias 0.06581f
C5610 Q1.t4 Vbias 0.05417f
C5611 Q1.t3 Vbias 0.0154f
C5612 Q1.n3 Vbias 0.07553f
C5613 Q1.n4 Vbias 0.01853f
C5614 Q1.t1 Vbias 0.01635f
C5615 Q1.t0 Vbias 0.01602f
C5616 Q1.n5 Vbias 0.09108f
C5617 Q1.n6 Vbias 0.03031f
C5618 Q1.t2 Vbias 0.01602f
C5619 Q1.n7 Vbias 0.02467f
C5620 Q1.n8 Vbias 0.04119f
C5621 Q1.n9 Vbias 0.01949f
C5622 Q1.n11 Vbias 0.03785f
C5623 Q1.n12 Vbias 5.26881f
C5624 Q1.t7 Vbias 0.06149f
C5625 Q1.t6 Vbias 0.11839f
C5626 Q1.t9 Vbias 0.06149f
C5627 Q1.n13 Vbias 0.09578f
C5628 Q1.n14 Vbias 0.09633f
C5629 Q1.t5 Vbias 0.10524f
C5630 Q1.n15 Vbias 1.21138f
C5631 Nand_Gate_7.B.t5 Vbias 0.74786f
C5632 Nand_Gate_7.B.n0 Vbias 0.21847f
C5633 Nand_Gate_7.B.n1 Vbias 0.09479f
C5634 Nand_Gate_7.B.n2 Vbias 0.41679f
C5635 Nand_Gate_7.B.t15 Vbias 0.34785f
C5636 Nand_Gate_7.B.n3 Vbias 0.10913f
C5637 Nand_Gate_7.B.t2 Vbias 0.09755f
C5638 Nand_Gate_7.B.n4 Vbias 0.42479f
C5639 Nand_Gate_7.B.n5 Vbias 0.10532f
C5640 Nand_Gate_7.B.t10 Vbias 0.7479f
C5641 Nand_Gate_7.B.n6 Vbias 0.735f
C5642 Nand_Gate_7.B.n7 Vbias 0.08033f
C5643 Nand_Gate_7.B.t14 Vbias 0.38883f
C5644 Nand_Gate_7.B.n8 Vbias 0.11201f
C5645 Nand_Gate_7.B.n9 Vbias 0.048f
C5646 Nand_Gate_7.B.n10 Vbias 0.08994f
C5647 Nand_Gate_7.B.n11 Vbias 0.11318f
C5648 Nand_Gate_7.B.t13 Vbias 0.7479f
C5649 Nand_Gate_7.B.n12 Vbias 0.735f
C5650 Nand_Gate_7.B.n13 Vbias 0.08033f
C5651 Nand_Gate_7.B.t11 Vbias 0.38883f
C5652 Nand_Gate_7.B.n14 Vbias 0.11201f
C5653 Nand_Gate_7.B.n15 Vbias 0.048f
C5654 Nand_Gate_7.B.n16 Vbias 0.08994f
C5655 Nand_Gate_7.B.n17 Vbias 0.01348f
C5656 Nand_Gate_7.B.n18 Vbias 0.33812f
C5657 Nand_Gate_7.B.n19 Vbias 0.09242f
C5658 Nand_Gate_7.B.n20 Vbias 0.24591f
C5659 Nand_Gate_7.B.t12 Vbias 0.7479f
C5660 Nand_Gate_7.B.n21 Vbias 0.75317f
C5661 Nand_Gate_7.B.n22 Vbias 0.08033f
C5662 Nand_Gate_7.B.t17 Vbias 0.38883f
C5663 Nand_Gate_7.B.n23 Vbias 0.11201f
C5664 Nand_Gate_7.B.n24 Vbias 0.02983f
C5665 Nand_Gate_7.B.n25 Vbias 0.04649f
C5666 Nand_Gate_7.B.n26 Vbias 0.46381f
C5667 Nand_Gate_7.B.t6 Vbias 0.7479f
C5668 Nand_Gate_7.B.n27 Vbias 0.75317f
C5669 Nand_Gate_7.B.n28 Vbias 0.08033f
C5670 Nand_Gate_7.B.t7 Vbias 0.38883f
C5671 Nand_Gate_7.B.n29 Vbias 0.11201f
C5672 Nand_Gate_7.B.n30 Vbias 0.02983f
C5673 Nand_Gate_7.B.n31 Vbias 0.04649f
C5674 Nand_Gate_7.B.n32 Vbias 0.01348f
C5675 Nand_Gate_7.B.n33 Vbias 1.20433f
C5676 Nand_Gate_7.B.n34 Vbias 0.49857f
C5677 Nand_Gate_7.B.n35 Vbias 0.20801f
C5678 Nand_Gate_7.B.t4 Vbias 0.74786f
C5679 Nand_Gate_7.B.n36 Vbias 0.21847f
C5680 Nand_Gate_7.B.n37 Vbias 0.09479f
C5681 Nand_Gate_7.B.n38 Vbias 0.41679f
C5682 Nand_Gate_7.B.t8 Vbias 0.34781f
C5683 Nand_Gate_7.B.n39 Vbias 0.10735f
C5684 Nand_Gate_7.B.n40 Vbias 0.24938f
C5685 Nand_Gate_7.B.n41 Vbias 13.7543f
C5686 Nand_Gate_7.B.t16 Vbias 0.38885f
C5687 Nand_Gate_7.B.n42 Vbias 0.41543f
C5688 Nand_Gate_7.B.t9 Vbias 0.74786f
C5689 Nand_Gate_7.B.n43 Vbias 1.70233f
C5690 Nand_Gate_7.B.n44 Vbias 16.1738f
C5691 Nand_Gate_7.B.n45 Vbias 0.12675f
C5692 Nand_Gate_7.B.n46 Vbias 0.42407f
C5693 Nand_Gate_7.B.n47 Vbias 0.91686f
C5694 Nand_Gate_7.B.n48 Vbias 0.01376f
C5695 Nand_Gate_7.B.n49 Vbias 0.12144f
C5696 Nand_Gate_7.B.n50 Vbias 0.06968f
C5697 Nand_Gate_7.B.t0 Vbias 0.10356f
C5698 Nand_Gate_7.B.t1 Vbias 0.10144f
C5699 Nand_Gate_7.B.n51 Vbias 0.57688f
C5700 Nand_Gate_7.B.n52 Vbias 0.19194f
C5701 Nand_Gate_7.B.t3 Vbias 0.10144f
C5702 Nand_Gate_7.B.n53 Vbias 0.15626f
C5703 Nand_Gate_7.B.n54 Vbias 0.27668f
C5704 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t4 Vbias 0.36784f
C5705 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n0 Vbias 0.10746f
C5706 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n1 Vbias 0.04662f
C5707 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t3 Vbias 0.04798f
C5708 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n2 Vbias 0.22815f
C5709 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n3 Vbias 0.0518f
C5710 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t7 Vbias 0.36785f
C5711 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n4 Vbias 0.38072f
C5712 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t6 Vbias 0.19125f
C5713 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n5 Vbias 0.18752f
C5714 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n6 Vbias 0.10934f
C5715 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n7 Vbias 0.01378f
C5716 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n8 Vbias 0.01506f
C5717 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t0 Vbias 0.05094f
C5718 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t1 Vbias 0.04989f
C5719 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n9 Vbias 0.28374f
C5720 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n10 Vbias 0.09441f
C5721 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t2 Vbias 0.04989f
C5722 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n11 Vbias 0.31407f
C5723 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.t5 Vbias 0.1838f
C5724 RingCounter_0.D_FlipFlop_8.3-input-nand_2.Vout.n12 Vbias 0.205f
C5725 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t4 Vbias 0.45666f
C5726 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n0 Vbias 0.47347f
C5727 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n1 Vbias 0.05122f
C5728 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n2 Vbias 0.06839f
C5729 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t7 Vbias 0.22727f
C5730 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t1 Vbias 0.06194f
C5731 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n3 Vbias 0.39067f
C5732 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t2 Vbias 0.06323f
C5733 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t3 Vbias 0.06194f
C5734 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n4 Vbias 0.35224f
C5735 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n5 Vbias 0.11629f
C5736 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n6 Vbias 0.16533f
C5737 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n7 Vbias 0.06431f
C5738 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t5 Vbias 0.23742f
C5739 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t6 Vbias 0.45664f
C5740 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n8 Vbias 0.1334f
C5741 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n9 Vbias 0.05705f
C5742 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n10 Vbias 0.10533f
C5743 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n11 Vbias 0.18236f
C5744 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n12 Vbias 0.13574f
C5745 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n13 Vbias 0.12257f
C5746 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.t0 Vbias 0.05969f
C5747 RingCounter_0.D_FlipFlop_8.3-input-nand_2.C.n14 Vbias 0.15961f
C5748 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t2 Vbias 0.07282f
C5749 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n0 Vbias 0.31709f
C5750 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n1 Vbias 0.07862f
C5751 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t4 Vbias 0.55828f
C5752 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n2 Vbias 0.54865f
C5753 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n3 Vbias 0.05997f
C5754 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t5 Vbias 0.29025f
C5755 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n4 Vbias 0.08361f
C5756 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n5 Vbias 0.03583f
C5757 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n6 Vbias 0.06714f
C5758 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n7 Vbias 0.15126f
C5759 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n8 Vbias 0.15126f
C5760 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n9 Vbias 0.09065f
C5761 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n10 Vbias 0.04578f
C5762 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t3 Vbias 0.07589f
C5763 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t0 Vbias 0.0773f
C5764 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.t1 Vbias 0.07572f
C5765 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n11 Vbias 0.43063f
C5766 RingCounter_0.D_FlipFlop_17.3-input-nand_0.Vout.n12 Vbias 0.24092f
C5767 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t2 Vbias 0.07037f
C5768 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n0 Vbias 0.16004f
C5769 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n1 Vbias 0.07725f
C5770 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t4 Vbias 0.2799f
C5771 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n2 Vbias 0.27418f
C5772 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n3 Vbias 0.05783f
C5773 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t5 Vbias 0.53832f
C5774 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n4 Vbias 0.15726f
C5775 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n5 Vbias 0.03913f
C5776 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n6 Vbias 0.05692f
C5777 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n7 Vbias 0.14585f
C5778 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n8 Vbias 0.14585f
C5779 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n9 Vbias 0.07581f
C5780 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t3 Vbias 0.07318f
C5781 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t0 Vbias 0.07454f
C5782 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.t1 Vbias 0.07302f
C5783 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n10 Vbias 0.41525f
C5784 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n11 Vbias 0.23391f
C5785 RingCounter_0.D_FlipFlop_16.3-input-nand_1.Vout.n12 Vbias 0.22303f
C5786 a_139496_37417.t3 Vbias 2.18377f
C5787 a_139496_37417.t0 Vbias 2.18303f
C5788 a_139496_37417.n0 Vbias 1.40282f
C5789 a_139496_37417.t2 Vbias 0.59708f
C5790 a_139496_37417.n1 Vbias 0.93584f
C5791 a_139496_37417.t1 Vbias 1.59747f
C5792 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t2 Vbias 0.07024f
C5793 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n0 Vbias 0.03989f
C5794 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n1 Vbias 0.07725f
C5795 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t5 Vbias 0.2799f
C5796 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n2 Vbias 0.27418f
C5797 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n3 Vbias 0.05783f
C5798 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t4 Vbias 0.53832f
C5799 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n4 Vbias 0.15726f
C5800 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n5 Vbias 0.03913f
C5801 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n6 Vbias 0.05692f
C5802 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n7 Vbias 0.14585f
C5803 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n8 Vbias 0.14585f
C5804 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n9 Vbias 0.07581f
C5805 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t3 Vbias 0.07318f
C5806 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t0 Vbias 0.07454f
C5807 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.t1 Vbias 0.07302f
C5808 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n10 Vbias 0.41525f
C5809 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n11 Vbias 0.23391f
C5810 RingCounter_0.D_FlipFlop_4.3-input-nand_1.Vout.n12 Vbias 0.22303f
C5811 D_FlipFlop_0.3-input-nand_2.C.t6 Vbias 0.3425f
C5812 D_FlipFlop_0.3-input-nand_2.C.n0 Vbias 0.3551f
C5813 D_FlipFlop_0.3-input-nand_2.C.n1 Vbias 0.03842f
C5814 D_FlipFlop_0.3-input-nand_2.C.n2 Vbias 0.05129f
C5815 D_FlipFlop_0.3-input-nand_2.C.t7 Vbias 0.17045f
C5816 D_FlipFlop_0.3-input-nand_2.C.t1 Vbias 0.04645f
C5817 D_FlipFlop_0.3-input-nand_2.C.n3 Vbias 0.293f
C5818 D_FlipFlop_0.3-input-nand_2.C.t3 Vbias 0.04742f
C5819 D_FlipFlop_0.3-input-nand_2.C.t2 Vbias 0.04645f
C5820 D_FlipFlop_0.3-input-nand_2.C.n4 Vbias 0.26418f
C5821 D_FlipFlop_0.3-input-nand_2.C.n5 Vbias 0.08722f
C5822 D_FlipFlop_0.3-input-nand_2.C.n6 Vbias 0.124f
C5823 D_FlipFlop_0.3-input-nand_2.C.n7 Vbias 0.04823f
C5824 D_FlipFlop_0.3-input-nand_2.C.t4 Vbias 0.17806f
C5825 D_FlipFlop_0.3-input-nand_2.C.t5 Vbias 0.34248f
C5826 D_FlipFlop_0.3-input-nand_2.C.n8 Vbias 0.10005f
C5827 D_FlipFlop_0.3-input-nand_2.C.n9 Vbias 0.04279f
C5828 D_FlipFlop_0.3-input-nand_2.C.n10 Vbias 0.079f
C5829 D_FlipFlop_0.3-input-nand_2.C.n11 Vbias 0.13677f
C5830 D_FlipFlop_0.3-input-nand_2.C.n12 Vbias 0.10181f
C5831 D_FlipFlop_0.3-input-nand_2.C.n13 Vbias 0.09193f
C5832 D_FlipFlop_0.3-input-nand_2.C.t0 Vbias 0.04477f
C5833 D_FlipFlop_0.3-input-nand_2.C.n14 Vbias 0.11971f
C5834 D_FlipFlop_3.3-input-nand_2.C.t7 Vbias 0.3425f
C5835 D_FlipFlop_3.3-input-nand_2.C.n0 Vbias 0.3551f
C5836 D_FlipFlop_3.3-input-nand_2.C.n1 Vbias 0.03842f
C5837 D_FlipFlop_3.3-input-nand_2.C.t2 Vbias 0.04477f
C5838 D_FlipFlop_3.3-input-nand_2.C.n2 Vbias 0.11971f
C5839 D_FlipFlop_3.3-input-nand_2.C.n3 Vbias 0.09193f
C5840 D_FlipFlop_3.3-input-nand_2.C.t5 Vbias 0.17806f
C5841 D_FlipFlop_3.3-input-nand_2.C.t6 Vbias 0.34248f
C5842 D_FlipFlop_3.3-input-nand_2.C.n4 Vbias 0.10005f
C5843 D_FlipFlop_3.3-input-nand_2.C.n5 Vbias 0.04279f
C5844 D_FlipFlop_3.3-input-nand_2.C.n6 Vbias 0.079f
C5845 D_FlipFlop_3.3-input-nand_2.C.n7 Vbias 0.13677f
C5846 D_FlipFlop_3.3-input-nand_2.C.n8 Vbias 0.10181f
C5847 D_FlipFlop_3.3-input-nand_2.C.n9 Vbias 0.04823f
C5848 D_FlipFlop_3.3-input-nand_2.C.n10 Vbias 0.124f
C5849 D_FlipFlop_3.3-input-nand_2.C.t3 Vbias 0.04742f
C5850 D_FlipFlop_3.3-input-nand_2.C.t0 Vbias 0.04645f
C5851 D_FlipFlop_3.3-input-nand_2.C.n11 Vbias 0.26418f
C5852 D_FlipFlop_3.3-input-nand_2.C.n12 Vbias 0.08722f
C5853 D_FlipFlop_3.3-input-nand_2.C.t1 Vbias 0.04645f
C5854 D_FlipFlop_3.3-input-nand_2.C.n13 Vbias 0.293f
C5855 D_FlipFlop_3.3-input-nand_2.C.t4 Vbias 0.17045f
C5856 D_FlipFlop_3.3-input-nand_2.C.n14 Vbias 0.05129f
C5857 D_FlipFlop_3.3-input-nand_2.Vout.t4 Vbias 0.35515f
C5858 D_FlipFlop_3.3-input-nand_2.Vout.n0 Vbias 0.10375f
C5859 D_FlipFlop_3.3-input-nand_2.Vout.n1 Vbias 0.04502f
C5860 D_FlipFlop_3.3-input-nand_2.Vout.t1 Vbias 0.04632f
C5861 D_FlipFlop_3.3-input-nand_2.Vout.n2 Vbias 0.22028f
C5862 D_FlipFlop_3.3-input-nand_2.Vout.n3 Vbias 0.05002f
C5863 D_FlipFlop_3.3-input-nand_2.Vout.t7 Vbias 0.35517f
C5864 D_FlipFlop_3.3-input-nand_2.Vout.n4 Vbias 0.36759f
C5865 D_FlipFlop_3.3-input-nand_2.Vout.t5 Vbias 0.18465f
C5866 D_FlipFlop_3.3-input-nand_2.Vout.n5 Vbias 0.18106f
C5867 D_FlipFlop_3.3-input-nand_2.Vout.n6 Vbias 0.10557f
C5868 D_FlipFlop_3.3-input-nand_2.Vout.n7 Vbias 0.01331f
C5869 D_FlipFlop_3.3-input-nand_2.Vout.n8 Vbias 0.01454f
C5870 D_FlipFlop_3.3-input-nand_2.Vout.t2 Vbias 0.04918f
C5871 D_FlipFlop_3.3-input-nand_2.Vout.t3 Vbias 0.04817f
C5872 D_FlipFlop_3.3-input-nand_2.Vout.n9 Vbias 0.27396f
C5873 D_FlipFlop_3.3-input-nand_2.Vout.n10 Vbias 0.09115f
C5874 D_FlipFlop_3.3-input-nand_2.Vout.t0 Vbias 0.04817f
C5875 D_FlipFlop_3.3-input-nand_2.Vout.n11 Vbias 0.30324f
C5876 D_FlipFlop_3.3-input-nand_2.Vout.t6 Vbias 0.17747f
C5877 D_FlipFlop_3.3-input-nand_2.Vout.n12 Vbias 0.19793f
C5878 Nand_Gate_4.B.t9 Vbias 0.65284f
C5879 Nand_Gate_4.B.n0 Vbias 0.19071f
C5880 Nand_Gate_4.B.n1 Vbias 0.08275f
C5881 Nand_Gate_4.B.n2 Vbias 0.36383f
C5882 Nand_Gate_4.B.t17 Vbias 0.30365f
C5883 Nand_Gate_4.B.n3 Vbias 0.09526f
C5884 Nand_Gate_4.B.t2 Vbias 0.08515f
C5885 Nand_Gate_4.B.n4 Vbias 0.37081f
C5886 Nand_Gate_4.B.n5 Vbias 0.09194f
C5887 Nand_Gate_4.B.t13 Vbias 0.65287f
C5888 Nand_Gate_4.B.n6 Vbias 0.6416f
C5889 Nand_Gate_4.B.n7 Vbias 0.07013f
C5890 Nand_Gate_4.B.t16 Vbias 0.33943f
C5891 Nand_Gate_4.B.n8 Vbias 0.09778f
C5892 Nand_Gate_4.B.n9 Vbias 0.0419f
C5893 Nand_Gate_4.B.n10 Vbias 0.07851f
C5894 Nand_Gate_4.B.n11 Vbias 0.0988f
C5895 Nand_Gate_4.B.t14 Vbias 0.65287f
C5896 Nand_Gate_4.B.n12 Vbias 0.6416f
C5897 Nand_Gate_4.B.n13 Vbias 0.07013f
C5898 Nand_Gate_4.B.t6 Vbias 0.33943f
C5899 Nand_Gate_4.B.n14 Vbias 0.09778f
C5900 Nand_Gate_4.B.n15 Vbias 0.0419f
C5901 Nand_Gate_4.B.n16 Vbias 0.07851f
C5902 Nand_Gate_4.B.n17 Vbias 0.01177f
C5903 Nand_Gate_4.B.n18 Vbias 0.29516f
C5904 Nand_Gate_4.B.n19 Vbias 0.08068f
C5905 Nand_Gate_4.B.n20 Vbias 0.21466f
C5906 Nand_Gate_4.B.t5 Vbias 0.65287f
C5907 Nand_Gate_4.B.n21 Vbias 0.65747f
C5908 Nand_Gate_4.B.n22 Vbias 0.07013f
C5909 Nand_Gate_4.B.t11 Vbias 0.33943f
C5910 Nand_Gate_4.B.n23 Vbias 0.09778f
C5911 Nand_Gate_4.B.n24 Vbias 0.02604f
C5912 Nand_Gate_4.B.n25 Vbias 0.04058f
C5913 Nand_Gate_4.B.n26 Vbias 0.40488f
C5914 Nand_Gate_4.B.t12 Vbias 0.65287f
C5915 Nand_Gate_4.B.n27 Vbias 0.65747f
C5916 Nand_Gate_4.B.n28 Vbias 0.07013f
C5917 Nand_Gate_4.B.t4 Vbias 0.33943f
C5918 Nand_Gate_4.B.n29 Vbias 0.09778f
C5919 Nand_Gate_4.B.n30 Vbias 0.02604f
C5920 Nand_Gate_4.B.n31 Vbias 0.04058f
C5921 Nand_Gate_4.B.n32 Vbias 0.01177f
C5922 Nand_Gate_4.B.n33 Vbias 1.0513f
C5923 Nand_Gate_4.B.n34 Vbias 0.45039f
C5924 Nand_Gate_4.B.n35 Vbias 0.18158f
C5925 Nand_Gate_4.B.t15 Vbias 0.65284f
C5926 Nand_Gate_4.B.n36 Vbias 0.19071f
C5927 Nand_Gate_4.B.n37 Vbias 0.08275f
C5928 Nand_Gate_4.B.n38 Vbias 0.36383f
C5929 Nand_Gate_4.B.t7 Vbias 0.30362f
C5930 Nand_Gate_4.B.n39 Vbias 0.07854f
C5931 Nand_Gate_4.B.n40 Vbias 0.1833f
C5932 Nand_Gate_4.B.n41 Vbias 15.2571f
C5933 Nand_Gate_4.B.t10 Vbias 0.33944f
C5934 Nand_Gate_4.B.n42 Vbias 0.36264f
C5935 Nand_Gate_4.B.t8 Vbias 0.65284f
C5936 Nand_Gate_4.B.n43 Vbias 1.46118f
C5937 Nand_Gate_4.B.n44 Vbias 17.2191f
C5938 Nand_Gate_4.B.n45 Vbias 0.11064f
C5939 Nand_Gate_4.B.n46 Vbias 0.37019f
C5940 Nand_Gate_4.B.n47 Vbias 0.80036f
C5941 Nand_Gate_4.B.n48 Vbias 0.01201f
C5942 Nand_Gate_4.B.n49 Vbias 0.10601f
C5943 Nand_Gate_4.B.n50 Vbias 0.06083f
C5944 Nand_Gate_4.B.t1 Vbias 0.0904f
C5945 Nand_Gate_4.B.t0 Vbias 0.08855f
C5946 Nand_Gate_4.B.n51 Vbias 0.50358f
C5947 Nand_Gate_4.B.n52 Vbias 0.16755f
C5948 Nand_Gate_4.B.t3 Vbias 0.08855f
C5949 Nand_Gate_4.B.n53 Vbias 0.1364f
C5950 Nand_Gate_4.B.n54 Vbias 0.24153f
C5951 Nand_Gate_5.A.t16 Vbias 0.37936f
C5952 Nand_Gate_5.A.n0 Vbias 0.11082f
C5953 Nand_Gate_5.A.n1 Vbias 0.04808f
C5954 Nand_Gate_5.A.n2 Vbias 0.21142f
C5955 Nand_Gate_5.A.t7 Vbias 0.17645f
C5956 Nand_Gate_5.A.n3 Vbias 0.05535f
C5957 Nand_Gate_5.A.t3 Vbias 0.04948f
C5958 Nand_Gate_5.A.n4 Vbias 0.21548f
C5959 Nand_Gate_5.A.n5 Vbias 0.05342f
C5960 Nand_Gate_5.A.t8 Vbias 0.37938f
C5961 Nand_Gate_5.A.n6 Vbias 0.37283f
C5962 Nand_Gate_5.A.n7 Vbias 0.04075f
C5963 Nand_Gate_5.A.t12 Vbias 0.19724f
C5964 Nand_Gate_5.A.n8 Vbias 0.05682f
C5965 Nand_Gate_5.A.n9 Vbias 0.02435f
C5966 Nand_Gate_5.A.n10 Vbias 0.04562f
C5967 Nand_Gate_5.A.n11 Vbias 0.05741f
C5968 Nand_Gate_5.A.t13 Vbias 0.37938f
C5969 Nand_Gate_5.A.n12 Vbias 0.37283f
C5970 Nand_Gate_5.A.n13 Vbias 0.04075f
C5971 Nand_Gate_5.A.t11 Vbias 0.19724f
C5972 Nand_Gate_5.A.n14 Vbias 0.05682f
C5973 Nand_Gate_5.A.n15 Vbias 0.02435f
C5974 Nand_Gate_5.A.n16 Vbias 0.04562f
C5975 Nand_Gate_5.A.n18 Vbias 0.17215f
C5976 Nand_Gate_5.A.n19 Vbias 0.47939f
C5977 Nand_Gate_5.A.n20 Vbias 0.21511f
C5978 Nand_Gate_5.A.t15 Vbias 0.37938f
C5979 Nand_Gate_5.A.n21 Vbias 0.38205f
C5980 Nand_Gate_5.A.n22 Vbias 0.04075f
C5981 Nand_Gate_5.A.t5 Vbias 0.19724f
C5982 Nand_Gate_5.A.n23 Vbias 0.05682f
C5983 Nand_Gate_5.A.n24 Vbias 0.01513f
C5984 Nand_Gate_5.A.n25 Vbias 0.02358f
C5985 Nand_Gate_5.A.n26 Vbias 0.23527f
C5986 Nand_Gate_5.A.t6 Vbias 0.37938f
C5987 Nand_Gate_5.A.n27 Vbias 0.38205f
C5988 Nand_Gate_5.A.n28 Vbias 0.04075f
C5989 Nand_Gate_5.A.t14 Vbias 0.19724f
C5990 Nand_Gate_5.A.n29 Vbias 0.05682f
C5991 Nand_Gate_5.A.n30 Vbias 0.01513f
C5992 Nand_Gate_5.A.n31 Vbias 0.02358f
C5993 Nand_Gate_5.A.n33 Vbias 0.6109f
C5994 Nand_Gate_5.A.n34 Vbias 0.28356f
C5995 Nand_Gate_5.A.n35 Vbias 0.10551f
C5996 Nand_Gate_5.A.t10 Vbias 0.37936f
C5997 Nand_Gate_5.A.n36 Vbias 0.11082f
C5998 Nand_Gate_5.A.n37 Vbias 0.04808f
C5999 Nand_Gate_5.A.n38 Vbias 0.21142f
C6000 Nand_Gate_5.A.t17 Vbias 0.17643f
C6001 Nand_Gate_5.A.n39 Vbias 0.0238f
C6002 Nand_Gate_5.A.n40 Vbias 0.05701f
C6003 Nand_Gate_5.A.n41 Vbias 2.28866f
C6004 Nand_Gate_5.A.t9 Vbias 0.19725f
C6005 Nand_Gate_5.A.n42 Vbias 0.19322f
C6006 Nand_Gate_5.A.n43 Vbias 0.04075f
C6007 Nand_Gate_5.A.t4 Vbias 0.37936f
C6008 Nand_Gate_5.A.n44 Vbias 0.11082f
C6009 Nand_Gate_5.A.n45 Vbias 0.02758f
C6010 Nand_Gate_5.A.n46 Vbias 0.04011f
C6011 Nand_Gate_5.A.n47 Vbias 0.05907f
C6012 Nand_Gate_5.A.n48 Vbias 3.11672f
C6013 Nand_Gate_5.A.n49 Vbias 0.20875f
C6014 Nand_Gate_5.A.n50 Vbias 0.06102f
C6015 Nand_Gate_5.A.n51 Vbias 0.02246f
C6016 Nand_Gate_5.A.n53 Vbias 0.0616f
C6017 Nand_Gate_5.A.n54 Vbias 0.03111f
C6018 Nand_Gate_5.A.t0 Vbias 0.05253f
C6019 Nand_Gate_5.A.t1 Vbias 0.05146f
C6020 Nand_Gate_5.A.n55 Vbias 0.29263f
C6021 Nand_Gate_5.A.n56 Vbias 0.09549f
C6022 Nand_Gate_5.A.t2 Vbias 0.05146f
C6023 Nand_Gate_5.A.n57 Vbias 0.07926f
C6024 Nand_Gate_5.A.n58 Vbias 0.14035f
C6025 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t2 Vbias 0.05201f
C6026 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n0 Vbias 0.22649f
C6027 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n1 Vbias 0.05616f
C6028 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t5 Vbias 0.39877f
C6029 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n2 Vbias 0.39189f
C6030 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n3 Vbias 0.04283f
C6031 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t4 Vbias 0.20732f
C6032 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n4 Vbias 0.05972f
C6033 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n5 Vbias 0.02559f
C6034 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n6 Vbias 0.04796f
C6035 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n7 Vbias 0.10804f
C6036 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n8 Vbias 0.10804f
C6037 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n9 Vbias 0.06475f
C6038 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t3 Vbias 0.05421f
C6039 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t0 Vbias 0.05522f
C6040 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.t1 Vbias 0.05409f
C6041 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n10 Vbias 0.30759f
C6042 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n11 Vbias 0.17406f
C6043 RingCounter_0.D_FlipFlop_11.3-input-nand_0.Vout.n12 Vbias 0.03715f
C6044 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t1 Vbias 0.0608f
C6045 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C6046 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C6047 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C6048 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C6049 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C6050 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C6051 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C6052 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C6053 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C6054 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C6055 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C6056 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C6057 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t0 Vbias 0.06323f
C6058 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.t2 Vbias 0.07525f
C6059 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C6060 RingCounter_0.D_FlipFlop_16.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C6061 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t1 Vbias 0.04607f
C6062 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n0 Vbias 0.10477f
C6063 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n1 Vbias 0.05057f
C6064 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t4 Vbias 0.35243f
C6065 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n2 Vbias 0.3654f
C6066 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n3 Vbias 0.03953f
C6067 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n4 Vbias 0.05278f
C6068 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t3 Vbias 0.27708f
C6069 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t2 Vbias 0.27709f
C6070 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n5 Vbias 0.17949f
C6071 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n6 Vbias 0.03786f
C6072 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t5 Vbias 0.35241f
C6073 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n7 Vbias 0.10295f
C6074 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n8 Vbias 0.02562f
C6075 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n9 Vbias 0.03726f
C6076 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n10 Vbias 0.09548f
C6077 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n11 Vbias 0.09548f
C6078 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n12 Vbias 0.04963f
C6079 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.t0 Vbias 0.04792f
C6080 RingCounter_0.D_FlipFlop_16.Inverter_1.Vout.n13 Vbias 0.28399f
C6081 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t1 Vbias 0.04798f
C6082 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n0 Vbias 0.02725f
C6083 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n1 Vbias 0.05277f
C6084 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t5 Vbias 0.36775f
C6085 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n2 Vbias 0.38129f
C6086 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n3 Vbias 0.04125f
C6087 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n4 Vbias 0.05508f
C6088 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t2 Vbias 0.28913f
C6089 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t4 Vbias 0.28914f
C6090 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n5 Vbias 0.1873f
C6091 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n6 Vbias 0.0395f
C6092 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t3 Vbias 0.36774f
C6093 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n7 Vbias 0.10743f
C6094 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n8 Vbias 0.02673f
C6095 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n9 Vbias 0.03888f
C6096 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n10 Vbias 0.09964f
C6097 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n11 Vbias 0.09964f
C6098 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n12 Vbias 0.05179f
C6099 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.t0 Vbias 0.05f
C6100 RingCounter_0.D_FlipFlop_6.Inverter_1.Vout.n13 Vbias 0.29633f
C6101 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t1 Vbias 0.06624f
C6102 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t2 Vbias 0.07883f
C6103 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n0 Vbias 0.39844f
C6104 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n1 Vbias 0.20187f
C6105 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n2 Vbias 0.06862f
C6106 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t3 Vbias 0.25335f
C6107 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n3 Vbias 0.24817f
C6108 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n4 Vbias 0.05234f
C6109 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t4 Vbias 0.48726f
C6110 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n5 Vbias 0.14234f
C6111 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n6 Vbias 0.03542f
C6112 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n7 Vbias 0.05152f
C6113 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C6114 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n9 Vbias 0.13202f
C6115 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n10 Vbias 0.06992f
C6116 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.n11 Vbias 0.03611f
C6117 RingCounter_0.D_FlipFlop_5.Nand_Gate_1.Vout.t0 Vbias 0.06358f
C6118 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t2 Vbias 0.05201f
C6119 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n0 Vbias 0.22649f
C6120 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n1 Vbias 0.05616f
C6121 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t5 Vbias 0.39877f
C6122 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n2 Vbias 0.39189f
C6123 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n3 Vbias 0.04283f
C6124 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t4 Vbias 0.20732f
C6125 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n4 Vbias 0.05972f
C6126 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n5 Vbias 0.02559f
C6127 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n6 Vbias 0.04796f
C6128 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n7 Vbias 0.10804f
C6129 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n8 Vbias 0.10804f
C6130 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n9 Vbias 0.06475f
C6131 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t3 Vbias 0.05421f
C6132 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t1 Vbias 0.05522f
C6133 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.t0 Vbias 0.05409f
C6134 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n10 Vbias 0.30759f
C6135 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n11 Vbias 0.17406f
C6136 RingCounter_0.D_FlipFlop_8.3-input-nand_0.Vout.n12 Vbias 0.03715f
C6137 Nand_Gate_6.B.t16 Vbias 0.66019f
C6138 Nand_Gate_6.B.n0 Vbias 0.19286f
C6139 Nand_Gate_6.B.n1 Vbias 0.08368f
C6140 Nand_Gate_6.B.n2 Vbias 0.36793f
C6141 Nand_Gate_6.B.t5 Vbias 0.30707f
C6142 Nand_Gate_6.B.n3 Vbias 0.09633f
C6143 Nand_Gate_6.B.t2 Vbias 0.08611f
C6144 Nand_Gate_6.B.n4 Vbias 0.37499f
C6145 Nand_Gate_6.B.n5 Vbias 0.09297f
C6146 Nand_Gate_6.B.t10 Vbias 0.66022f
C6147 Nand_Gate_6.B.n6 Vbias 0.64883f
C6148 Nand_Gate_6.B.n7 Vbias 0.07092f
C6149 Nand_Gate_6.B.t17 Vbias 0.34325f
C6150 Nand_Gate_6.B.n8 Vbias 0.09888f
C6151 Nand_Gate_6.B.n9 Vbias 0.04237f
C6152 Nand_Gate_6.B.n10 Vbias 0.0794f
C6153 Nand_Gate_6.B.n11 Vbias 0.09991f
C6154 Nand_Gate_6.B.t15 Vbias 0.66022f
C6155 Nand_Gate_6.B.n12 Vbias 0.64883f
C6156 Nand_Gate_6.B.n13 Vbias 0.07092f
C6157 Nand_Gate_6.B.t11 Vbias 0.34325f
C6158 Nand_Gate_6.B.n14 Vbias 0.09888f
C6159 Nand_Gate_6.B.n15 Vbias 0.04237f
C6160 Nand_Gate_6.B.n16 Vbias 0.0794f
C6161 Nand_Gate_6.B.n17 Vbias 0.0119f
C6162 Nand_Gate_6.B.n18 Vbias 0.29848f
C6163 Nand_Gate_6.B.n19 Vbias 0.08159f
C6164 Nand_Gate_6.B.n20 Vbias 0.21708f
C6165 Nand_Gate_6.B.t6 Vbias 0.66022f
C6166 Nand_Gate_6.B.n21 Vbias 0.66487f
C6167 Nand_Gate_6.B.n22 Vbias 0.07092f
C6168 Nand_Gate_6.B.t12 Vbias 0.34325f
C6169 Nand_Gate_6.B.n23 Vbias 0.09888f
C6170 Nand_Gate_6.B.n24 Vbias 0.02633f
C6171 Nand_Gate_6.B.n25 Vbias 0.04104f
C6172 Nand_Gate_6.B.n26 Vbias 0.40943f
C6173 Nand_Gate_6.B.t13 Vbias 0.66022f
C6174 Nand_Gate_6.B.n27 Vbias 0.66487f
C6175 Nand_Gate_6.B.n28 Vbias 0.07092f
C6176 Nand_Gate_6.B.t7 Vbias 0.34325f
C6177 Nand_Gate_6.B.n29 Vbias 0.09888f
C6178 Nand_Gate_6.B.n30 Vbias 0.02633f
C6179 Nand_Gate_6.B.n31 Vbias 0.04104f
C6180 Nand_Gate_6.B.n32 Vbias 0.0119f
C6181 Nand_Gate_6.B.n33 Vbias 1.06314f
C6182 Nand_Gate_6.B.n34 Vbias 0.43942f
C6183 Nand_Gate_6.B.n35 Vbias 0.18362f
C6184 Nand_Gate_6.B.t4 Vbias 0.66019f
C6185 Nand_Gate_6.B.n36 Vbias 0.19286f
C6186 Nand_Gate_6.B.n37 Vbias 0.08368f
C6187 Nand_Gate_6.B.n38 Vbias 0.36793f
C6188 Nand_Gate_6.B.t9 Vbias 0.30704f
C6189 Nand_Gate_6.B.n39 Vbias 0.09546f
C6190 Nand_Gate_6.B.n40 Vbias 0.22172f
C6191 Nand_Gate_6.B.n41 Vbias 8.79656f
C6192 Nand_Gate_6.B.t8 Vbias 0.34326f
C6193 Nand_Gate_6.B.n42 Vbias 0.36672f
C6194 Nand_Gate_6.B.t14 Vbias 0.66019f
C6195 Nand_Gate_6.B.n43 Vbias 1.50275f
C6196 Nand_Gate_6.B.n44 Vbias 11.1675f
C6197 Nand_Gate_6.B.n45 Vbias 0.11189f
C6198 Nand_Gate_6.B.n46 Vbias 0.37436f
C6199 Nand_Gate_6.B.n47 Vbias 0.80937f
C6200 Nand_Gate_6.B.n48 Vbias 0.01215f
C6201 Nand_Gate_6.B.n49 Vbias 0.10721f
C6202 Nand_Gate_6.B.n50 Vbias 0.06151f
C6203 Nand_Gate_6.B.t0 Vbias 0.09142f
C6204 Nand_Gate_6.B.t1 Vbias 0.08955f
C6205 Nand_Gate_6.B.n51 Vbias 0.50925f
C6206 Nand_Gate_6.B.n52 Vbias 0.16944f
C6207 Nand_Gate_6.B.t3 Vbias 0.08955f
C6208 Nand_Gate_6.B.n53 Vbias 0.13794f
C6209 Nand_Gate_6.B.n54 Vbias 0.24424f
C6210 Nand_Gate_5.Vout.t2 Vbias 0.07306f
C6211 Nand_Gate_5.Vout.n0 Vbias 0.0415f
C6212 Nand_Gate_5.Vout.n1 Vbias 0.08035f
C6213 Nand_Gate_5.Vout.t3 Vbias 0.29114f
C6214 Nand_Gate_5.Vout.n2 Vbias 0.28519f
C6215 Nand_Gate_5.Vout.n3 Vbias 0.06015f
C6216 Nand_Gate_5.Vout.t4 Vbias 0.55994f
C6217 Nand_Gate_5.Vout.n4 Vbias 0.16357f
C6218 Nand_Gate_5.Vout.n5 Vbias 0.0407f
C6219 Nand_Gate_5.Vout.n6 Vbias 0.05921f
C6220 Nand_Gate_5.Vout.n7 Vbias 1.13762f
C6221 Nand_Gate_5.Vout.n8 Vbias 1.13762f
C6222 Nand_Gate_5.Vout.n9 Vbias 0.07886f
C6223 Nand_Gate_5.Vout.t1 Vbias 0.07612f
C6224 Nand_Gate_5.Vout.t0 Vbias 0.09059f
C6225 Nand_Gate_5.Vout.n10 Vbias 0.45787f
C6226 Nand_Gate_5.Vout.n11 Vbias 0.23199f
C6227 CDAC8_0.switch_5.Z.t2 Vbias 0.03054f
C6228 CDAC8_0.switch_5.Z.t1 Vbias 0.03054f
C6229 CDAC8_0.switch_5.Z.n0 Vbias 0.11035f
C6230 CDAC8_0.switch_5.Z.n1 Vbias 0.254f
C6231 CDAC8_0.switch_5.Z.t3 Vbias 0.03207f
C6232 CDAC8_0.switch_5.Z.t6 Vbias 5.60901f
C6233 CDAC8_0.switch_5.Z.n2 Vbias 1.99837f
C6234 CDAC8_0.switch_5.Z.t5 Vbias 5.4744f
C6235 CDAC8_0.switch_5.Z.t9 Vbias 5.4744f
C6236 CDAC8_0.switch_5.Z.t7 Vbias 5.39614f
C6237 CDAC8_0.switch_5.Z.n3 Vbias 1.42238f
C6238 CDAC8_0.switch_5.Z.t4 Vbias 5.39614f
C6239 CDAC8_0.switch_5.Z.n4 Vbias 1.67019f
C6240 CDAC8_0.switch_5.Z.n5 Vbias 2.09417f
C6241 CDAC8_0.switch_5.Z.n6 Vbias 2.09417f
C6242 CDAC8_0.switch_5.Z.t8 Vbias 5.39614f
C6243 CDAC8_0.switch_5.Z.n7 Vbias 1.67019f
C6244 CDAC8_0.switch_5.Z.t11 Vbias 5.39614f
C6245 CDAC8_0.switch_5.Z.n8 Vbias 1.42238f
C6246 CDAC8_0.switch_5.Z.t10 Vbias 5.60901f
C6247 CDAC8_0.switch_5.Z.n9 Vbias 1.95831f
C6248 CDAC8_0.switch_5.Z.n10 Vbias 0.46579f
C6249 CDAC8_0.switch_5.Z.n11 Vbias 0.10945f
C6250 CDAC8_0.switch_5.Z.t0 Vbias 0.03205f
C6251 Q3.t8 Vbias 0.11803f
C6252 Q3.n0 Vbias 0.03448f
C6253 Q3.n1 Vbias 0.01496f
C6254 Q3.n2 Vbias 0.06578f
C6255 Q3.t5 Vbias 0.05414f
C6256 Q3.t1 Vbias 0.0154f
C6257 Q3.n3 Vbias 0.0755f
C6258 Q3.n4 Vbias 0.01853f
C6259 Q3.t0 Vbias 0.01634f
C6260 Q3.t3 Vbias 0.01601f
C6261 Q3.n5 Vbias 0.09105f
C6262 Q3.n6 Vbias 0.03029f
C6263 Q3.t2 Vbias 0.01601f
C6264 Q3.n7 Vbias 0.02466f
C6265 Q3.n8 Vbias 0.04061f
C6266 Q3.n9 Vbias 0.02001f
C6267 Q3.n11 Vbias 0.03887f
C6268 Q3.n12 Vbias 5.74071f
C6269 Q3.t6 Vbias 0.06147f
C6270 Q3.t4 Vbias 0.11834f
C6271 Q3.t7 Vbias 0.06147f
C6272 Q3.n13 Vbias 0.09574f
C6273 Q3.n14 Vbias 0.09629f
C6274 Q3.t9 Vbias 0.1052f
C6275 Q3.n15 Vbias 1.21087f
C6276 CDAC8_0.switch_2.Z.t2 Vbias 0.03087f
C6277 CDAC8_0.switch_2.Z.t1 Vbias 0.03087f
C6278 CDAC8_0.switch_2.Z.n0 Vbias 0.12722f
C6279 CDAC8_0.switch_2.Z.t5 Vbias 6.50564f
C6280 CDAC8_0.switch_2.Z.t4 Vbias 6.4338f
C6281 CDAC8_0.switch_2.Z.n1 Vbias 1.02469f
C6282 CDAC8_0.switch_2.Z.n2 Vbias 0.01025f
C6283 CDAC8_0.switch_2.Z.n3 Vbias 0.03182f
C6284 CDAC8_0.switch_2.Z.t3 Vbias 0.02943f
C6285 CDAC8_0.switch_2.Z.t0 Vbias 0.02943f
C6286 CDAC8_0.switch_2.Z.n4 Vbias 0.10631f
C6287 CDAC8_0.switch_2.Z.n5 Vbias 0.24452f
C6288 Q6.t3 Vbias 0.01626f
C6289 Q6.n0 Vbias 0.07974f
C6290 Q6.n1 Vbias 0.01957f
C6291 Q6.t1 Vbias 0.01726f
C6292 Q6.t0 Vbias 0.01691f
C6293 Q6.n2 Vbias 0.09616f
C6294 Q6.n3 Vbias 0.03199f
C6295 Q6.t2 Vbias 0.01691f
C6296 Q6.n4 Vbias 0.02605f
C6297 Q6.n5 Vbias 0.0372f
C6298 Q6.n6 Vbias 0.0192f
C6299 Q6.t8 Vbias 0.12466f
C6300 Q6.n7 Vbias 0.03642f
C6301 Q6.n8 Vbias 0.0158f
C6302 Q6.n9 Vbias 0.06947f
C6303 Q6.t6 Vbias 0.05798f
C6304 Q6.n11 Vbias 0.01555f
C6305 Q6.n13 Vbias 3.34141f
C6306 Q6.t4 Vbias 0.12498f
C6307 Q6.t5 Vbias 0.12498f
C6308 Q6.t9 Vbias 0.06492f
C6309 Q6.n14 Vbias 0.10112f
C6310 Q6.n15 Vbias 0.1017f
C6311 Q6.t7 Vbias 0.05702f
C6312 Q6.n16 Vbias 1.27887f
C6313 D_FlipFlop_5.3-input-nand_2.C.t5 Vbias 0.3425f
C6314 D_FlipFlop_5.3-input-nand_2.C.n0 Vbias 0.3551f
C6315 D_FlipFlop_5.3-input-nand_2.C.n1 Vbias 0.03842f
C6316 D_FlipFlop_5.3-input-nand_2.C.n2 Vbias 0.05129f
C6317 D_FlipFlop_5.3-input-nand_2.C.t6 Vbias 0.17045f
C6318 D_FlipFlop_5.3-input-nand_2.C.t1 Vbias 0.04645f
C6319 D_FlipFlop_5.3-input-nand_2.C.n3 Vbias 0.293f
C6320 D_FlipFlop_5.3-input-nand_2.C.t3 Vbias 0.04742f
C6321 D_FlipFlop_5.3-input-nand_2.C.t2 Vbias 0.04645f
C6322 D_FlipFlop_5.3-input-nand_2.C.n4 Vbias 0.26418f
C6323 D_FlipFlop_5.3-input-nand_2.C.n5 Vbias 0.08722f
C6324 D_FlipFlop_5.3-input-nand_2.C.n6 Vbias 0.124f
C6325 D_FlipFlop_5.3-input-nand_2.C.n7 Vbias 0.04823f
C6326 D_FlipFlop_5.3-input-nand_2.C.t7 Vbias 0.17806f
C6327 D_FlipFlop_5.3-input-nand_2.C.t4 Vbias 0.34248f
C6328 D_FlipFlop_5.3-input-nand_2.C.n8 Vbias 0.10005f
C6329 D_FlipFlop_5.3-input-nand_2.C.n9 Vbias 0.04279f
C6330 D_FlipFlop_5.3-input-nand_2.C.n10 Vbias 0.079f
C6331 D_FlipFlop_5.3-input-nand_2.C.n11 Vbias 0.13677f
C6332 D_FlipFlop_5.3-input-nand_2.C.n12 Vbias 0.10181f
C6333 D_FlipFlop_5.3-input-nand_2.C.n13 Vbias 0.09193f
C6334 D_FlipFlop_5.3-input-nand_2.C.t0 Vbias 0.04477f
C6335 D_FlipFlop_5.3-input-nand_2.C.n14 Vbias 0.11971f
C6336 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t4 Vbias 0.36784f
C6337 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6338 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6339 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t1 Vbias 0.04798f
C6340 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6341 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6342 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t6 Vbias 0.36785f
C6343 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6344 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t5 Vbias 0.19125f
C6345 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6346 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6347 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6348 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n8 Vbias 0.01095f
C6349 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t0 Vbias 0.05094f
C6350 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t3 Vbias 0.04989f
C6351 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6352 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n10 Vbias 0.09258f
C6353 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t2 Vbias 0.04989f
C6354 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6355 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.t7 Vbias 0.1838f
C6356 RingCounter_0.D_FlipFlop_3.3-input-nand_2.Vout.n12 Vbias 0.205f
C6357 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t1 Vbias 0.04998f
C6358 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n0 Vbias 0.02839f
C6359 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n1 Vbias 0.05497f
C6360 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t5 Vbias 0.38308f
C6361 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n2 Vbias 0.39717f
C6362 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n3 Vbias 0.04297f
C6363 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n4 Vbias 0.05737f
C6364 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t2 Vbias 0.30118f
C6365 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t4 Vbias 0.30119f
C6366 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n5 Vbias 0.1951f
C6367 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n6 Vbias 0.04115f
C6368 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t3 Vbias 0.38306f
C6369 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n7 Vbias 0.1119f
C6370 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n8 Vbias 0.02784f
C6371 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n9 Vbias 0.0405f
C6372 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n10 Vbias 0.10379f
C6373 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n11 Vbias 0.10379f
C6374 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n12 Vbias 0.05395f
C6375 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.t0 Vbias 0.05208f
C6376 RingCounter_0.D_FlipFlop_2.Inverter_1.Vout.n13 Vbias 0.30868f
C6377 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t5 Vbias 0.45666f
C6378 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n0 Vbias 0.47347f
C6379 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n1 Vbias 0.05122f
C6380 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n2 Vbias 0.06839f
C6381 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t6 Vbias 0.22727f
C6382 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t1 Vbias 0.06194f
C6383 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n3 Vbias 0.39067f
C6384 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t3 Vbias 0.06323f
C6385 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t2 Vbias 0.06194f
C6386 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n4 Vbias 0.35224f
C6387 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n5 Vbias 0.11629f
C6388 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n6 Vbias 0.16533f
C6389 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n7 Vbias 0.06431f
C6390 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t7 Vbias 0.23742f
C6391 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t4 Vbias 0.45664f
C6392 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n8 Vbias 0.1334f
C6393 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n9 Vbias 0.05705f
C6394 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n10 Vbias 0.10533f
C6395 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n11 Vbias 0.18236f
C6396 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n12 Vbias 0.13574f
C6397 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n13 Vbias 0.12257f
C6398 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.t0 Vbias 0.05969f
C6399 RingCounter_0.D_FlipFlop_12.3-input-nand_2.C.n14 Vbias 0.15961f
C6400 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t6 Vbias 0.36784f
C6401 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6402 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6403 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t2 Vbias 0.04798f
C6404 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6405 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6406 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t7 Vbias 0.36785f
C6407 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6408 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t5 Vbias 0.19125f
C6409 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6410 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6411 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6412 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n8 Vbias 0.01506f
C6413 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t0 Vbias 0.05094f
C6414 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t1 Vbias 0.04989f
C6415 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6416 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n10 Vbias 0.09441f
C6417 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t3 Vbias 0.04989f
C6418 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6419 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.t4 Vbias 0.1838f
C6420 RingCounter_0.D_FlipFlop_12.3-input-nand_2.Vout.n12 Vbias 0.205f
C6421 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t7 Vbias 0.45666f
C6422 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n0 Vbias 0.47347f
C6423 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n1 Vbias 0.05122f
C6424 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n2 Vbias 0.06839f
C6425 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t4 Vbias 0.22727f
C6426 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t1 Vbias 0.06194f
C6427 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n3 Vbias 0.39067f
C6428 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t2 Vbias 0.06323f
C6429 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t3 Vbias 0.06194f
C6430 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n4 Vbias 0.35224f
C6431 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n5 Vbias 0.11629f
C6432 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n6 Vbias 0.16533f
C6433 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n7 Vbias 0.06431f
C6434 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t5 Vbias 0.23742f
C6435 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t6 Vbias 0.45664f
C6436 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n8 Vbias 0.1334f
C6437 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n9 Vbias 0.05705f
C6438 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n10 Vbias 0.10533f
C6439 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n11 Vbias 0.18236f
C6440 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n12 Vbias 0.13574f
C6441 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n13 Vbias 0.12257f
C6442 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.t0 Vbias 0.05969f
C6443 RingCounter_0.D_FlipFlop_9.3-input-nand_2.C.n14 Vbias 0.15961f
C6444 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t4 Vbias 0.36784f
C6445 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6446 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6447 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t3 Vbias 0.04798f
C6448 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6449 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6450 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t5 Vbias 0.36785f
C6451 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6452 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t7 Vbias 0.19125f
C6453 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6454 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6455 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6456 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n8 Vbias 0.01506f
C6457 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t1 Vbias 0.05094f
C6458 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t2 Vbias 0.04989f
C6459 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6460 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n10 Vbias 0.09441f
C6461 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t0 Vbias 0.04989f
C6462 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6463 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.t6 Vbias 0.1838f
C6464 RingCounter_0.D_FlipFlop_9.3-input-nand_2.Vout.n12 Vbias 0.205f
C6465 D_FlipFlop_0.3-input-nand_2.Vout.t6 Vbias 0.35515f
C6466 D_FlipFlop_0.3-input-nand_2.Vout.n0 Vbias 0.10375f
C6467 D_FlipFlop_0.3-input-nand_2.Vout.n1 Vbias 0.04502f
C6468 D_FlipFlop_0.3-input-nand_2.Vout.t1 Vbias 0.04632f
C6469 D_FlipFlop_0.3-input-nand_2.Vout.n2 Vbias 0.22028f
C6470 D_FlipFlop_0.3-input-nand_2.Vout.n3 Vbias 0.05002f
C6471 D_FlipFlop_0.3-input-nand_2.Vout.t5 Vbias 0.35517f
C6472 D_FlipFlop_0.3-input-nand_2.Vout.n4 Vbias 0.36759f
C6473 D_FlipFlop_0.3-input-nand_2.Vout.t7 Vbias 0.18465f
C6474 D_FlipFlop_0.3-input-nand_2.Vout.n5 Vbias 0.18106f
C6475 D_FlipFlop_0.3-input-nand_2.Vout.n6 Vbias 0.10557f
C6476 D_FlipFlop_0.3-input-nand_2.Vout.n7 Vbias 0.01331f
C6477 D_FlipFlop_0.3-input-nand_2.Vout.n8 Vbias 0.01454f
C6478 D_FlipFlop_0.3-input-nand_2.Vout.t3 Vbias 0.04918f
C6479 D_FlipFlop_0.3-input-nand_2.Vout.t2 Vbias 0.04817f
C6480 D_FlipFlop_0.3-input-nand_2.Vout.n9 Vbias 0.27396f
C6481 D_FlipFlop_0.3-input-nand_2.Vout.n10 Vbias 0.09115f
C6482 D_FlipFlop_0.3-input-nand_2.Vout.t0 Vbias 0.04817f
C6483 D_FlipFlop_0.3-input-nand_2.Vout.n11 Vbias 0.30324f
C6484 D_FlipFlop_0.3-input-nand_2.Vout.t4 Vbias 0.17747f
C6485 D_FlipFlop_0.3-input-nand_2.Vout.n12 Vbias 0.19793f
C6486 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t4 Vbias 0.36784f
C6487 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6488 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6489 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t1 Vbias 0.04798f
C6490 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6491 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6492 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t6 Vbias 0.36785f
C6493 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6494 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t7 Vbias 0.19125f
C6495 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6496 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6497 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6498 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n8 Vbias 0.01506f
C6499 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t0 Vbias 0.05094f
C6500 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t3 Vbias 0.04989f
C6501 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6502 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n10 Vbias 0.09441f
C6503 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t2 Vbias 0.04989f
C6504 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6505 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.t5 Vbias 0.1838f
C6506 RingCounter_0.D_FlipFlop_13.3-input-nand_2.Vout.n12 Vbias 0.205f
C6507 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t4 Vbias 0.45666f
C6508 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n0 Vbias 0.47347f
C6509 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n1 Vbias 0.05122f
C6510 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n2 Vbias 0.06839f
C6511 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t7 Vbias 0.22727f
C6512 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t1 Vbias 0.06194f
C6513 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n3 Vbias 0.39067f
C6514 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t3 Vbias 0.06323f
C6515 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t2 Vbias 0.06194f
C6516 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n4 Vbias 0.35224f
C6517 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n5 Vbias 0.11629f
C6518 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n6 Vbias 0.16533f
C6519 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n7 Vbias 0.06431f
C6520 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t5 Vbias 0.23742f
C6521 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t6 Vbias 0.45664f
C6522 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n8 Vbias 0.1334f
C6523 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n9 Vbias 0.05705f
C6524 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n10 Vbias 0.10533f
C6525 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n11 Vbias 0.18236f
C6526 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n12 Vbias 0.13574f
C6527 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n13 Vbias 0.12257f
C6528 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.t0 Vbias 0.05969f
C6529 RingCounter_0.D_FlipFlop_13.3-input-nand_2.C.n14 Vbias 0.15961f
C6530 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t7 Vbias 0.36784f
C6531 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6532 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6533 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t3 Vbias 0.04798f
C6534 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6535 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6536 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t5 Vbias 0.36785f
C6537 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6538 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t4 Vbias 0.19125f
C6539 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6540 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6541 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6542 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n8 Vbias 0.01095f
C6543 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t0 Vbias 0.05094f
C6544 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t1 Vbias 0.04989f
C6545 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6546 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n10 Vbias 0.09258f
C6547 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t2 Vbias 0.04989f
C6548 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6549 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.t6 Vbias 0.1838f
C6550 RingCounter_0.D_FlipFlop_5.3-input-nand_2.Vout.n12 Vbias 0.205f
C6551 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t7 Vbias 0.38055f
C6552 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n0 Vbias 0.39456f
C6553 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n1 Vbias 0.04269f
C6554 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t2 Vbias 0.04965f
C6555 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n2 Vbias 0.04808f
C6556 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n3 Vbias 0.10214f
C6557 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t4 Vbias 0.19785f
C6558 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t6 Vbias 0.38054f
C6559 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n4 Vbias 0.11117f
C6560 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n5 Vbias 0.04754f
C6561 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n6 Vbias 0.08777f
C6562 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n7 Vbias 0.15197f
C6563 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n8 Vbias 0.11312f
C6564 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n9 Vbias 0.05359f
C6565 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n10 Vbias 0.13778f
C6566 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t0 Vbias 0.05269f
C6567 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t3 Vbias 0.05162f
C6568 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n11 Vbias 0.29353f
C6569 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n12 Vbias 0.09691f
C6570 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t1 Vbias 0.05162f
C6571 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n13 Vbias 0.32556f
C6572 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.t5 Vbias 0.18939f
C6573 RingCounter_0.D_FlipFlop_17.3-input-nand_2.C.n14 Vbias 0.05699f
C6574 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t5 Vbias 0.45666f
C6575 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n0 Vbias 0.47347f
C6576 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n1 Vbias 0.05122f
C6577 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n2 Vbias 0.06839f
C6578 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t7 Vbias 0.22727f
C6579 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t1 Vbias 0.06194f
C6580 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n3 Vbias 0.39067f
C6581 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t2 Vbias 0.06323f
C6582 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t3 Vbias 0.06194f
C6583 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n4 Vbias 0.35224f
C6584 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n5 Vbias 0.11629f
C6585 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n6 Vbias 0.16533f
C6586 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n7 Vbias 0.06431f
C6587 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t6 Vbias 0.23742f
C6588 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t4 Vbias 0.45664f
C6589 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n8 Vbias 0.1334f
C6590 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n9 Vbias 0.05705f
C6591 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n10 Vbias 0.10533f
C6592 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n11 Vbias 0.18236f
C6593 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n12 Vbias 0.13574f
C6594 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n13 Vbias 0.12257f
C6595 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.n14 Vbias 0.0577f
C6596 RingCounter_0.D_FlipFlop_6.3-input-nand_2.C.t0 Vbias 0.05958f
C6597 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t4 Vbias 0.36784f
C6598 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n0 Vbias 0.10746f
C6599 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n1 Vbias 0.04662f
C6600 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t1 Vbias 0.04798f
C6601 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n2 Vbias 0.22815f
C6602 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n3 Vbias 0.0518f
C6603 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t7 Vbias 0.36785f
C6604 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n4 Vbias 0.38072f
C6605 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t6 Vbias 0.19125f
C6606 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n5 Vbias 0.18752f
C6607 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n6 Vbias 0.10934f
C6608 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n7 Vbias 0.01378f
C6609 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n8 Vbias 0.01095f
C6610 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t0 Vbias 0.05094f
C6611 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t3 Vbias 0.04989f
C6612 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n9 Vbias 0.28374f
C6613 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n10 Vbias 0.09258f
C6614 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t2 Vbias 0.04989f
C6615 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n11 Vbias 0.31407f
C6616 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.t5 Vbias 0.1838f
C6617 RingCounter_0.D_FlipFlop_7.3-input-nand_2.Vout.n12 Vbias 0.205f
C6618 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t4 Vbias 0.45666f
C6619 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n0 Vbias 0.47347f
C6620 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n1 Vbias 0.05122f
C6621 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n2 Vbias 0.06839f
C6622 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t6 Vbias 0.22727f
C6623 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t1 Vbias 0.06194f
C6624 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n3 Vbias 0.39067f
C6625 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t2 Vbias 0.06323f
C6626 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t3 Vbias 0.06194f
C6627 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n4 Vbias 0.35224f
C6628 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n5 Vbias 0.11629f
C6629 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n6 Vbias 0.16533f
C6630 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n7 Vbias 0.06431f
C6631 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t5 Vbias 0.23742f
C6632 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t7 Vbias 0.45664f
C6633 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n8 Vbias 0.1334f
C6634 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n9 Vbias 0.05705f
C6635 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n10 Vbias 0.10533f
C6636 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n11 Vbias 0.18236f
C6637 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n12 Vbias 0.13574f
C6638 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n13 Vbias 0.12257f
C6639 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.n14 Vbias 0.0577f
C6640 RingCounter_0.D_FlipFlop_7.3-input-nand_2.C.t0 Vbias 0.05958f
C6641 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t2 Vbias 0.07037f
C6642 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n0 Vbias 0.16004f
C6643 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n1 Vbias 0.07725f
C6644 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t4 Vbias 0.2799f
C6645 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n2 Vbias 0.27418f
C6646 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n3 Vbias 0.05783f
C6647 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t5 Vbias 0.53832f
C6648 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n4 Vbias 0.15726f
C6649 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n5 Vbias 0.03913f
C6650 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n6 Vbias 0.05692f
C6651 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n7 Vbias 0.14585f
C6652 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n8 Vbias 0.14585f
C6653 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n9 Vbias 0.07581f
C6654 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t3 Vbias 0.07318f
C6655 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t0 Vbias 0.07454f
C6656 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.t1 Vbias 0.07302f
C6657 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n10 Vbias 0.41525f
C6658 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n11 Vbias 0.23391f
C6659 RingCounter_0.D_FlipFlop_14.3-input-nand_1.Vout.n12 Vbias 0.22303f
C6660 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t1 Vbias 0.04607f
C6661 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n0 Vbias 0.10477f
C6662 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n1 Vbias 0.05057f
C6663 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t3 Vbias 0.35243f
C6664 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n2 Vbias 0.3654f
C6665 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n3 Vbias 0.03953f
C6666 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n4 Vbias 0.05278f
C6667 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t2 Vbias 0.27708f
C6668 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t5 Vbias 0.27709f
C6669 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n5 Vbias 0.17949f
C6670 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n6 Vbias 0.03786f
C6671 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t4 Vbias 0.35241f
C6672 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n7 Vbias 0.10295f
C6673 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n8 Vbias 0.02562f
C6674 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n9 Vbias 0.03726f
C6675 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n10 Vbias 0.09548f
C6676 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n11 Vbias 0.09548f
C6677 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n12 Vbias 0.04963f
C6678 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.t0 Vbias 0.04792f
C6679 RingCounter_0.D_FlipFlop_10.Inverter_1.Vout.n13 Vbias 0.28399f
C6680 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t7 Vbias 0.45666f
C6681 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n0 Vbias 0.47347f
C6682 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n1 Vbias 0.05122f
C6683 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t2 Vbias 0.05958f
C6684 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n2 Vbias 0.0577f
C6685 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n3 Vbias 0.12257f
C6686 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t5 Vbias 0.23742f
C6687 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t4 Vbias 0.45664f
C6688 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n4 Vbias 0.1334f
C6689 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n5 Vbias 0.05705f
C6690 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n6 Vbias 0.10533f
C6691 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n7 Vbias 0.18236f
C6692 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n8 Vbias 0.13574f
C6693 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n9 Vbias 0.06431f
C6694 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n10 Vbias 0.16533f
C6695 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t1 Vbias 0.06323f
C6696 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t0 Vbias 0.06194f
C6697 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n11 Vbias 0.35224f
C6698 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n12 Vbias 0.11629f
C6699 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t3 Vbias 0.06194f
C6700 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n13 Vbias 0.39067f
C6701 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.t6 Vbias 0.22727f
C6702 RingCounter_0.D_FlipFlop_1.3-input-nand_2.C.n14 Vbias 0.06839f
C6703 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t2 Vbias 0.0608f
C6704 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C6705 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C6706 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t3 Vbias 0.24183f
C6707 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C6708 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C6709 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t4 Vbias 0.46511f
C6710 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C6711 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C6712 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C6713 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C6714 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C6715 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C6716 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t1 Vbias 0.06323f
C6717 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C6718 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C6719 RingCounter_0.D_FlipFlop_9.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C6720 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t1 Vbias 0.04607f
C6721 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n0 Vbias 0.10477f
C6722 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n1 Vbias 0.05057f
C6723 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t5 Vbias 0.35243f
C6724 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n2 Vbias 0.3654f
C6725 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n3 Vbias 0.03953f
C6726 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n4 Vbias 0.05278f
C6727 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t4 Vbias 0.27708f
C6728 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t3 Vbias 0.27709f
C6729 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n5 Vbias 0.17949f
C6730 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n6 Vbias 0.03786f
C6731 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t2 Vbias 0.35241f
C6732 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n7 Vbias 0.10295f
C6733 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n8 Vbias 0.02562f
C6734 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n9 Vbias 0.03726f
C6735 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n10 Vbias 0.09548f
C6736 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n11 Vbias 0.09548f
C6737 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n12 Vbias 0.04963f
C6738 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.t0 Vbias 0.04792f
C6739 RingCounter_0.D_FlipFlop_9.Inverter_1.Vout.n13 Vbias 0.28399f
C6740 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t1 Vbias 0.06358f
C6741 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n0 Vbias 0.03611f
C6742 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n1 Vbias 0.06992f
C6743 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t3 Vbias 0.25335f
C6744 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n2 Vbias 0.24817f
C6745 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n3 Vbias 0.05234f
C6746 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t4 Vbias 0.48726f
C6747 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n4 Vbias 0.14234f
C6748 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n5 Vbias 0.03542f
C6749 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n6 Vbias 0.05152f
C6750 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n7 Vbias 0.13202f
C6751 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C6752 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n9 Vbias 0.06862f
C6753 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t2 Vbias 0.06624f
C6754 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.t0 Vbias 0.07883f
C6755 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n10 Vbias 0.39844f
C6756 RingCounter_0.D_FlipFlop_7.Nand_Gate_1.Vout.n11 Vbias 0.20187f
C6757 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t1 Vbias 0.04998f
C6758 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n0 Vbias 0.02839f
C6759 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n1 Vbias 0.05497f
C6760 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t5 Vbias 0.38308f
C6761 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n2 Vbias 0.39717f
C6762 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n3 Vbias 0.04297f
C6763 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n4 Vbias 0.05737f
C6764 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t4 Vbias 0.30118f
C6765 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t3 Vbias 0.30119f
C6766 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n5 Vbias 0.1951f
C6767 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n6 Vbias 0.04115f
C6768 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t2 Vbias 0.38306f
C6769 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n7 Vbias 0.1119f
C6770 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n8 Vbias 0.02784f
C6771 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n9 Vbias 0.0405f
C6772 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n10 Vbias 0.10379f
C6773 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n11 Vbias 0.10379f
C6774 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n12 Vbias 0.05395f
C6775 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.t0 Vbias 0.05208f
C6776 RingCounter_0.D_FlipFlop_7.Inverter_1.Vout.n13 Vbias 0.30868f
C6777 FFCLR.t35 Vbias 0.56738f
C6778 FFCLR.n0 Vbias 0.16575f
C6779 FFCLR.n1 Vbias 0.07192f
C6780 FFCLR.n2 Vbias 0.3162f
C6781 FFCLR.t6 Vbias 0.2639f
C6782 FFCLR.n3 Vbias 0.08279f
C6783 FFCLR.t2 Vbias 0.07401f
C6784 FFCLR.n4 Vbias 0.32227f
C6785 FFCLR.n5 Vbias 0.0799f
C6786 FFCLR.t41 Vbias 0.5674f
C6787 FFCLR.n6 Vbias 0.55761f
C6788 FFCLR.n7 Vbias 0.06095f
C6789 FFCLR.t34 Vbias 0.29499f
C6790 FFCLR.n8 Vbias 0.08498f
C6791 FFCLR.n9 Vbias 0.03642f
C6792 FFCLR.n10 Vbias 0.06823f
C6793 FFCLR.n11 Vbias 0.08587f
C6794 FFCLR.t32 Vbias 0.5674f
C6795 FFCLR.n12 Vbias 0.55761f
C6796 FFCLR.n13 Vbias 0.06095f
C6797 FFCLR.t40 Vbias 0.29499f
C6798 FFCLR.n14 Vbias 0.08498f
C6799 FFCLR.n15 Vbias 0.03642f
C6800 FFCLR.n16 Vbias 0.06823f
C6801 FFCLR.n17 Vbias 0.01023f
C6802 FFCLR.n18 Vbias 0.25748f
C6803 FFCLR.n19 Vbias 0.71698f
C6804 FFCLR.n20 Vbias 0.32173f
C6805 FFCLR.t39 Vbias 0.5674f
C6806 FFCLR.n21 Vbias 0.5714f
C6807 FFCLR.n22 Vbias 0.06095f
C6808 FFCLR.t11 Vbias 0.29499f
C6809 FFCLR.n23 Vbias 0.08498f
C6810 FFCLR.n24 Vbias 0.02263f
C6811 FFCLR.n25 Vbias 0.03527f
C6812 FFCLR.n26 Vbias 0.35187f
C6813 FFCLR.t13 Vbias 0.5674f
C6814 FFCLR.n27 Vbias 0.5714f
C6815 FFCLR.n28 Vbias 0.06095f
C6816 FFCLR.t38 Vbias 0.29499f
C6817 FFCLR.n29 Vbias 0.08498f
C6818 FFCLR.n30 Vbias 0.02263f
C6819 FFCLR.n31 Vbias 0.03527f
C6820 FFCLR.n32 Vbias 0.01023f
C6821 FFCLR.n33 Vbias 0.91367f
C6822 FFCLR.n34 Vbias 0.42769f
C6823 FFCLR.n35 Vbias 0.15781f
C6824 FFCLR.t26 Vbias 0.56738f
C6825 FFCLR.n36 Vbias 0.16575f
C6826 FFCLR.n37 Vbias 0.07192f
C6827 FFCLR.n38 Vbias 0.3162f
C6828 FFCLR.t44 Vbias 0.26387f
C6829 FFCLR.n39 Vbias 0.03199f
C6830 FFCLR.n40 Vbias 0.07711f
C6831 FFCLR.n41 Vbias 0.02079f
C6832 FFCLR.t19 Vbias 0.5674f
C6833 FFCLR.n42 Vbias 0.58828f
C6834 FFCLR.n43 Vbias 0.06364f
C6835 FFCLR.n44 Vbias 0.08498f
C6836 FFCLR.t27 Vbias 0.26502f
C6837 FFCLR.n45 Vbias 0.53269f
C6838 FFCLR.n46 Vbias 0.15142f
C6839 FFCLR.t33 Vbias 0.295f
C6840 FFCLR.n47 Vbias 0.27519f
C6841 FFCLR.n48 Vbias 0.06095f
C6842 FFCLR.t53 Vbias 0.56738f
C6843 FFCLR.n49 Vbias 0.16575f
C6844 FFCLR.n50 Vbias 0.05503f
C6845 FFCLR.n51 Vbias 0.09296f
C6846 FFCLR.n52 Vbias 0.35187f
C6847 FFCLR.t8 Vbias 0.295f
C6848 FFCLR.n53 Vbias 0.27519f
C6849 FFCLR.n54 Vbias 0.06095f
C6850 FFCLR.t23 Vbias 0.56738f
C6851 FFCLR.n55 Vbias 0.16575f
C6852 FFCLR.n56 Vbias 0.05503f
C6853 FFCLR.n57 Vbias 0.09296f
C6854 FFCLR.n58 Vbias 0.01023f
C6855 FFCLR.n59 Vbias 0.89353f
C6856 FFCLR.n60 Vbias 0.49808f
C6857 FFCLR.t37 Vbias 0.5674f
C6858 FFCLR.n61 Vbias 0.58828f
C6859 FFCLR.n62 Vbias 0.06364f
C6860 FFCLR.n63 Vbias 0.08498f
C6861 FFCLR.t45 Vbias 0.26498f
C6862 FFCLR.n64 Vbias 0.57621f
C6863 FFCLR.n65 Vbias 0.32094f
C6864 FFCLR.n66 Vbias 0.15142f
C6865 FFCLR.t50 Vbias 0.295f
C6866 FFCLR.n67 Vbias 0.27519f
C6867 FFCLR.n68 Vbias 0.06095f
C6868 FFCLR.t12 Vbias 0.56738f
C6869 FFCLR.n69 Vbias 0.16575f
C6870 FFCLR.n70 Vbias 0.05503f
C6871 FFCLR.n71 Vbias 0.09296f
C6872 FFCLR.n72 Vbias 0.35187f
C6873 FFCLR.t22 Vbias 0.295f
C6874 FFCLR.n73 Vbias 0.27519f
C6875 FFCLR.n74 Vbias 0.06095f
C6876 FFCLR.t42 Vbias 0.56738f
C6877 FFCLR.n75 Vbias 0.16575f
C6878 FFCLR.n76 Vbias 0.05503f
C6879 FFCLR.n77 Vbias 0.09296f
C6880 FFCLR.n78 Vbias 0.01023f
C6881 FFCLR.n79 Vbias 0.89353f
C6882 FFCLR.n80 Vbias 0.49808f
C6883 FFCLR.t14 Vbias 0.5674f
C6884 FFCLR.n81 Vbias 0.58828f
C6885 FFCLR.n82 Vbias 0.06364f
C6886 FFCLR.n83 Vbias 0.08498f
C6887 FFCLR.t7 Vbias 0.26498f
C6888 FFCLR.n84 Vbias 0.57621f
C6889 FFCLR.n85 Vbias 0.32094f
C6890 FFCLR.n86 Vbias 0.15142f
C6891 FFCLR.t24 Vbias 0.295f
C6892 FFCLR.n87 Vbias 0.27519f
C6893 FFCLR.n88 Vbias 0.06095f
C6894 FFCLR.t31 Vbias 0.56738f
C6895 FFCLR.n89 Vbias 0.16575f
C6896 FFCLR.n90 Vbias 0.05503f
C6897 FFCLR.n91 Vbias 0.09296f
C6898 FFCLR.n92 Vbias 0.35187f
C6899 FFCLR.t56 Vbias 0.295f
C6900 FFCLR.n93 Vbias 0.27519f
C6901 FFCLR.n94 Vbias 0.06095f
C6902 FFCLR.t4 Vbias 0.56738f
C6903 FFCLR.n95 Vbias 0.16575f
C6904 FFCLR.n96 Vbias 0.05503f
C6905 FFCLR.n97 Vbias 0.09296f
C6906 FFCLR.n98 Vbias 0.01023f
C6907 FFCLR.n99 Vbias 0.89353f
C6908 FFCLR.n100 Vbias 0.80291f
C6909 FFCLR.n101 Vbias 0.10865f
C6910 FFCLR.t54 Vbias 0.295f
C6911 FFCLR.n102 Vbias 0.27519f
C6912 FFCLR.n103 Vbias 0.06095f
C6913 FFCLR.t17 Vbias 0.56738f
C6914 FFCLR.n104 Vbias 0.16575f
C6915 FFCLR.n105 Vbias 0.05503f
C6916 FFCLR.n106 Vbias 0.09296f
C6917 FFCLR.n107 Vbias 0.35187f
C6918 FFCLR.t28 Vbias 0.295f
C6919 FFCLR.n108 Vbias 0.27519f
C6920 FFCLR.n109 Vbias 0.06095f
C6921 FFCLR.t46 Vbias 0.56738f
C6922 FFCLR.n110 Vbias 0.16575f
C6923 FFCLR.n111 Vbias 0.05503f
C6924 FFCLR.n112 Vbias 0.09296f
C6925 FFCLR.n113 Vbias 0.01023f
C6926 FFCLR.n114 Vbias 0.89353f
C6927 FFCLR.n115 Vbias 0.12822f
C6928 FFCLR.n116 Vbias 0.15142f
C6929 FFCLR.n117 Vbias 0.32094f
C6930 FFCLR.t43 Vbias 0.5674f
C6931 FFCLR.n118 Vbias 0.58828f
C6932 FFCLR.n119 Vbias 0.06364f
C6933 FFCLR.n120 Vbias 0.08498f
C6934 FFCLR.t49 Vbias 0.26498f
C6935 FFCLR.n121 Vbias 0.20635f
C6936 FFCLR.n122 Vbias 0.58864f
C6937 FFCLR.n123 Vbias 1.01138f
C6938 FFCLR.t10 Vbias 0.295f
C6939 FFCLR.n124 Vbias 0.27519f
C6940 FFCLR.n125 Vbias 0.06095f
C6941 FFCLR.t29 Vbias 0.56738f
C6942 FFCLR.n126 Vbias 0.16575f
C6943 FFCLR.n127 Vbias 0.05503f
C6944 FFCLR.n128 Vbias 0.09296f
C6945 FFCLR.n129 Vbias 0.35187f
C6946 FFCLR.t36 Vbias 0.295f
C6947 FFCLR.n130 Vbias 0.27519f
C6948 FFCLR.n131 Vbias 0.06095f
C6949 FFCLR.t59 Vbias 0.56738f
C6950 FFCLR.n132 Vbias 0.16575f
C6951 FFCLR.n133 Vbias 0.05503f
C6952 FFCLR.n134 Vbias 0.09296f
C6953 FFCLR.n135 Vbias 0.01023f
C6954 FFCLR.n136 Vbias 0.89353f
C6955 FFCLR.n137 Vbias 0.12822f
C6956 FFCLR.n138 Vbias 0.15142f
C6957 FFCLR.n139 Vbias 0.32094f
C6958 FFCLR.t15 Vbias 0.5674f
C6959 FFCLR.n140 Vbias 0.58828f
C6960 FFCLR.n141 Vbias 0.06364f
C6961 FFCLR.n142 Vbias 0.08498f
C6962 FFCLR.t9 Vbias 0.26498f
C6963 FFCLR.n143 Vbias 0.20635f
C6964 FFCLR.n144 Vbias 1.12268f
C6965 FFCLR.n145 Vbias 1.59883f
C6966 FFCLR.t21 Vbias 0.295f
C6967 FFCLR.n146 Vbias 0.27519f
C6968 FFCLR.n147 Vbias 0.06095f
C6969 FFCLR.t25 Vbias 0.56738f
C6970 FFCLR.n148 Vbias 0.16575f
C6971 FFCLR.n149 Vbias 0.05503f
C6972 FFCLR.n150 Vbias 0.09296f
C6973 FFCLR.n151 Vbias 0.35187f
C6974 FFCLR.t51 Vbias 0.295f
C6975 FFCLR.n152 Vbias 0.27519f
C6976 FFCLR.n153 Vbias 0.06095f
C6977 FFCLR.t57 Vbias 0.56738f
C6978 FFCLR.n154 Vbias 0.16575f
C6979 FFCLR.n155 Vbias 0.05503f
C6980 FFCLR.n156 Vbias 0.09296f
C6981 FFCLR.n157 Vbias 0.01023f
C6982 FFCLR.n158 Vbias 0.89353f
C6983 FFCLR.n159 Vbias 0.12822f
C6984 FFCLR.n160 Vbias 0.15142f
C6985 FFCLR.n161 Vbias 0.32094f
C6986 FFCLR.t52 Vbias 0.5674f
C6987 FFCLR.n162 Vbias 0.58828f
C6988 FFCLR.n163 Vbias 0.06364f
C6989 FFCLR.n164 Vbias 0.08498f
C6990 FFCLR.t5 Vbias 0.26498f
C6991 FFCLR.n165 Vbias 0.20635f
C6992 FFCLR.n166 Vbias 1.65673f
C6993 FFCLR.n167 Vbias 2.18628f
C6994 FFCLR.t58 Vbias 0.295f
C6995 FFCLR.n168 Vbias 0.27519f
C6996 FFCLR.n169 Vbias 0.06095f
C6997 FFCLR.t18 Vbias 0.56738f
C6998 FFCLR.n170 Vbias 0.16575f
C6999 FFCLR.n171 Vbias 0.05503f
C7000 FFCLR.n172 Vbias 0.09296f
C7001 FFCLR.n173 Vbias 0.35187f
C7002 FFCLR.t30 Vbias 0.295f
C7003 FFCLR.n174 Vbias 0.27519f
C7004 FFCLR.n175 Vbias 0.06095f
C7005 FFCLR.t47 Vbias 0.56738f
C7006 FFCLR.n176 Vbias 0.16575f
C7007 FFCLR.n177 Vbias 0.05503f
C7008 FFCLR.n178 Vbias 0.09296f
C7009 FFCLR.n179 Vbias 0.01023f
C7010 FFCLR.n180 Vbias 0.89353f
C7011 FFCLR.n181 Vbias 0.12822f
C7012 FFCLR.n182 Vbias 0.15142f
C7013 FFCLR.n183 Vbias 0.32094f
C7014 FFCLR.t20 Vbias 0.5674f
C7015 FFCLR.n184 Vbias 0.58828f
C7016 FFCLR.n185 Vbias 0.06364f
C7017 FFCLR.n186 Vbias 0.08498f
C7018 FFCLR.t55 Vbias 0.26498f
C7019 FFCLR.n187 Vbias 0.20635f
C7020 FFCLR.n188 Vbias 2.25881f
C7021 FFCLR.n189 Vbias 3.07138f
C7022 FFCLR.n190 Vbias 0.98757f
C7023 FFCLR.n191 Vbias 15.1698f
C7024 FFCLR.t16 Vbias 0.295f
C7025 FFCLR.n192 Vbias 0.28898f
C7026 FFCLR.n193 Vbias 0.06095f
C7027 FFCLR.t48 Vbias 0.56738f
C7028 FFCLR.n194 Vbias 0.16575f
C7029 FFCLR.n195 Vbias 0.04124f
C7030 FFCLR.n196 Vbias 0.05999f
C7031 FFCLR.n197 Vbias 0.08834f
C7032 FFCLR.n198 Vbias 16.0173f
C7033 FFCLR.n199 Vbias 0.31221f
C7034 FFCLR.n200 Vbias 0.09126f
C7035 FFCLR.n201 Vbias 0.03359f
C7036 FFCLR.n202 Vbias 0.01039f
C7037 FFCLR.n203 Vbias 0.09213f
C7038 FFCLR.n204 Vbias 0.04653f
C7039 FFCLR.t1 Vbias 0.07857f
C7040 FFCLR.t0 Vbias 0.07696f
C7041 FFCLR.n205 Vbias 0.43766f
C7042 FFCLR.n206 Vbias 0.14281f
C7043 FFCLR.t3 Vbias 0.07696f
C7044 FFCLR.n207 Vbias 0.11855f
C7045 FFCLR.n208 Vbias 0.20991f
C7046 Nand_Gate_6.A.t7 Vbias 0.27993f
C7047 Nand_Gate_6.A.n0 Vbias 0.08177f
C7048 Nand_Gate_6.A.n1 Vbias 0.03548f
C7049 Nand_Gate_6.A.n2 Vbias 0.15601f
C7050 Nand_Gate_6.A.t11 Vbias 0.1302f
C7051 Nand_Gate_6.A.n3 Vbias 0.04085f
C7052 Nand_Gate_6.A.t1 Vbias 0.03651f
C7053 Nand_Gate_6.A.n4 Vbias 0.159f
C7054 Nand_Gate_6.A.n5 Vbias 0.03942f
C7055 Nand_Gate_6.A.t4 Vbias 0.27994f
C7056 Nand_Gate_6.A.n6 Vbias 0.27511f
C7057 Nand_Gate_6.A.n7 Vbias 0.03007f
C7058 Nand_Gate_6.A.t10 Vbias 0.14554f
C7059 Nand_Gate_6.A.n8 Vbias 0.04192f
C7060 Nand_Gate_6.A.n9 Vbias 0.01797f
C7061 Nand_Gate_6.A.n10 Vbias 0.03367f
C7062 Nand_Gate_6.A.n11 Vbias 0.04236f
C7063 Nand_Gate_6.A.t6 Vbias 0.27994f
C7064 Nand_Gate_6.A.n12 Vbias 0.27511f
C7065 Nand_Gate_6.A.n13 Vbias 0.03007f
C7066 Nand_Gate_6.A.t8 Vbias 0.14554f
C7067 Nand_Gate_6.A.n14 Vbias 0.04192f
C7068 Nand_Gate_6.A.n15 Vbias 0.01797f
C7069 Nand_Gate_6.A.n16 Vbias 0.03367f
C7070 Nand_Gate_6.A.n18 Vbias 0.12656f
C7071 Nand_Gate_6.A.n19 Vbias 0.03459f
C7072 Nand_Gate_6.A.n20 Vbias 0.09204f
C7073 Nand_Gate_6.A.t9 Vbias 0.14555f
C7074 Nand_Gate_6.A.n21 Vbias 0.14257f
C7075 Nand_Gate_6.A.n22 Vbias 0.03007f
C7076 Nand_Gate_6.A.t5 Vbias 0.27993f
C7077 Nand_Gate_6.A.n23 Vbias 0.08177f
C7078 Nand_Gate_6.A.n24 Vbias 0.02035f
C7079 Nand_Gate_6.A.n25 Vbias 0.0296f
C7080 Nand_Gate_6.A.n26 Vbias 0.14551f
C7081 Nand_Gate_6.A.n27 Vbias 0.25531f
C7082 Nand_Gate_6.A.n28 Vbias 0.15873f
C7083 Nand_Gate_6.A.n29 Vbias 0.34318f
C7084 Nand_Gate_6.A.n31 Vbias 0.04546f
C7085 Nand_Gate_6.A.n32 Vbias 0.02608f
C7086 Nand_Gate_6.A.t0 Vbias 0.03876f
C7087 Nand_Gate_6.A.t3 Vbias 0.03797f
C7088 Nand_Gate_6.A.n33 Vbias 0.21593f
C7089 Nand_Gate_6.A.n34 Vbias 0.07184f
C7090 Nand_Gate_6.A.t2 Vbias 0.03797f
C7091 Nand_Gate_6.A.n35 Vbias 0.05849f
C7092 Nand_Gate_6.A.n36 Vbias 0.10356f
C7093 Nand_Gate_5.B.t9 Vbias 0.09725f
C7094 Nand_Gate_5.B.n0 Vbias 0.02801f
C7095 Nand_Gate_5.B.n1 Vbias 0.01201f
C7096 Nand_Gate_5.B.n2 Vbias 0.02249f
C7097 Nand_Gate_5.B.t8 Vbias 0.18705f
C7098 Nand_Gate_5.B.n3 Vbias 0.18382f
C7099 Nand_Gate_5.B.n4 Vbias 0.02009f
C7100 Nand_Gate_5.B.t11 Vbias 0.09725f
C7101 Nand_Gate_5.B.n5 Vbias 0.02801f
C7102 Nand_Gate_5.B.n6 Vbias 0.01201f
C7103 Nand_Gate_5.B.n7 Vbias 0.02249f
C7104 Nand_Gate_5.B.n8 Vbias 0.05912f
C7105 Nand_Gate_5.B.n9 Vbias 0.05912f
C7106 Nand_Gate_5.B.n10 Vbias 0.02009f
C7107 Nand_Gate_5.B.n11 Vbias 0.18382f
C7108 Nand_Gate_5.B.t10 Vbias 0.16795f
C7109 Nand_Gate_5.B.n12 Vbias 1.59684f
C7110 Nand_Gate_5.B.t6 Vbias 0.09725f
C7111 Nand_Gate_5.B.t4 Vbias 0.18704f
C7112 Nand_Gate_5.B.n13 Vbias 0.05464f
C7113 Nand_Gate_5.B.n14 Vbias 0.02337f
C7114 Nand_Gate_5.B.n15 Vbias 0.04314f
C7115 Nand_Gate_5.B.n16 Vbias 0.36438f
C7116 Nand_Gate_5.B.n17 Vbias 2.13619f
C7117 Nand_Gate_5.B.t5 Vbias 0.16927f
C7118 Nand_Gate_5.B.n18 Vbias 0.05464f
C7119 Nand_Gate_5.B.n19 Vbias 0.02371f
C7120 Nand_Gate_5.B.n20 Vbias 0.10424f
C7121 Nand_Gate_5.B.t7 Vbias 0.087f
C7122 Nand_Gate_5.B.n21 Vbias 0.02729f
C7123 Nand_Gate_5.B.t3 Vbias 0.0244f
C7124 Nand_Gate_5.B.n22 Vbias 0.11964f
C7125 Nand_Gate_5.B.n23 Vbias 0.02727f
C7126 Nand_Gate_5.B.t0 Vbias 0.0259f
C7127 Nand_Gate_5.B.t1 Vbias 0.02537f
C7128 Nand_Gate_5.B.n24 Vbias 0.14428f
C7129 Nand_Gate_5.B.n25 Vbias 0.04708f
C7130 Nand_Gate_5.B.t2 Vbias 0.02537f
C7131 Nand_Gate_5.B.n26 Vbias 0.03908f
C7132 Nand_Gate_5.B.n27 Vbias 0.0692f
C7133 CDAC8_0.switch_9.Z.t2 Vbias 0.03608f
C7134 CDAC8_0.switch_9.Z.t3 Vbias 0.0344f
C7135 CDAC8_0.switch_9.Z.t1 Vbias 0.0344f
C7136 CDAC8_0.switch_9.Z.n0 Vbias 0.12427f
C7137 CDAC8_0.switch_9.Z.n1 Vbias 0.28559f
C7138 CDAC8_0.switch_9.Z.n2 Vbias 0.0372f
C7139 CDAC8_0.switch_9.Z.t25 Vbias 6.43398f
C7140 CDAC8_0.switch_9.Z.t23 Vbias 6.07647f
C7141 CDAC8_0.switch_9.Z.n3 Vbias 3.42262f
C7142 CDAC8_0.switch_9.Z.t32 Vbias 6.07647f
C7143 CDAC8_0.switch_9.Z.n4 Vbias 1.60172f
C7144 CDAC8_0.switch_9.Z.n5 Vbias 1.3726f
C7145 CDAC8_0.switch_9.Z.t28 Vbias 6.43398f
C7146 CDAC8_0.switch_9.Z.t27 Vbias 6.07647f
C7147 CDAC8_0.switch_9.Z.n6 Vbias 3.42262f
C7148 CDAC8_0.switch_9.Z.t35 Vbias 6.07647f
C7149 CDAC8_0.switch_9.Z.n7 Vbias 1.60172f
C7150 CDAC8_0.switch_9.Z.t31 Vbias 6.44737f
C7151 CDAC8_0.switch_9.Z.t24 Vbias 6.07647f
C7152 CDAC8_0.switch_9.Z.n8 Vbias 3.47318f
C7153 CDAC8_0.switch_9.Z.t26 Vbias 6.07647f
C7154 CDAC8_0.switch_9.Z.n9 Vbias 1.75389f
C7155 CDAC8_0.switch_9.Z.t30 Vbias 6.07647f
C7156 CDAC8_0.switch_9.Z.n10 Vbias 1.88076f
C7157 CDAC8_0.switch_9.Z.t10 Vbias 6.07647f
C7158 CDAC8_0.switch_9.Z.n11 Vbias 2.07349f
C7159 CDAC8_0.switch_9.Z.t14 Vbias 6.07647f
C7160 CDAC8_0.switch_9.Z.n12 Vbias 2.07349f
C7161 CDAC8_0.switch_9.Z.t13 Vbias 6.07647f
C7162 CDAC8_0.switch_9.Z.n13 Vbias 2.07349f
C7163 CDAC8_0.switch_9.Z.t18 Vbias 6.07647f
C7164 CDAC8_0.switch_9.Z.n14 Vbias 2.07349f
C7165 CDAC8_0.switch_9.Z.t17 Vbias 6.07647f
C7166 CDAC8_0.switch_9.Z.n15 Vbias 2.07349f
C7167 CDAC8_0.switch_9.Z.t34 Vbias 6.07647f
C7168 CDAC8_0.switch_9.Z.n16 Vbias 2.07349f
C7169 CDAC8_0.switch_9.Z.t6 Vbias 6.07647f
C7170 CDAC8_0.switch_9.Z.n17 Vbias 2.07349f
C7171 CDAC8_0.switch_9.Z.t5 Vbias 6.07647f
C7172 CDAC8_0.switch_9.Z.n18 Vbias 2.07349f
C7173 CDAC8_0.switch_9.Z.t9 Vbias 6.07647f
C7174 CDAC8_0.switch_9.Z.n19 Vbias 1.72859f
C7175 CDAC8_0.switch_9.Z.t29 Vbias 6.44737f
C7176 CDAC8_0.switch_9.Z.t20 Vbias 6.07647f
C7177 CDAC8_0.switch_9.Z.n20 Vbias 3.47318f
C7178 CDAC8_0.switch_9.Z.t22 Vbias 6.07647f
C7179 CDAC8_0.switch_9.Z.n21 Vbias 1.75389f
C7180 CDAC8_0.switch_9.Z.n22 Vbias 1.99f
C7181 CDAC8_0.switch_9.Z.n23 Vbias 1.99f
C7182 CDAC8_0.switch_9.Z.t11 Vbias 6.07647f
C7183 CDAC8_0.switch_9.Z.n24 Vbias 1.72859f
C7184 CDAC8_0.switch_9.Z.t7 Vbias 6.07647f
C7185 CDAC8_0.switch_9.Z.n25 Vbias 2.07349f
C7186 CDAC8_0.switch_9.Z.t8 Vbias 6.07647f
C7187 CDAC8_0.switch_9.Z.n26 Vbias 2.07349f
C7188 CDAC8_0.switch_9.Z.t4 Vbias 6.07647f
C7189 CDAC8_0.switch_9.Z.n27 Vbias 2.07349f
C7190 CDAC8_0.switch_9.Z.t19 Vbias 6.07647f
C7191 CDAC8_0.switch_9.Z.n28 Vbias 2.07349f
C7192 CDAC8_0.switch_9.Z.t21 Vbias 6.07647f
C7193 CDAC8_0.switch_9.Z.n29 Vbias 2.07349f
C7194 CDAC8_0.switch_9.Z.t15 Vbias 6.07647f
C7195 CDAC8_0.switch_9.Z.n30 Vbias 2.07349f
C7196 CDAC8_0.switch_9.Z.t16 Vbias 6.07647f
C7197 CDAC8_0.switch_9.Z.n31 Vbias 2.07349f
C7198 CDAC8_0.switch_9.Z.t12 Vbias 6.07647f
C7199 CDAC8_0.switch_9.Z.n32 Vbias 2.07349f
C7200 CDAC8_0.switch_9.Z.t33 Vbias 6.07647f
C7201 CDAC8_0.switch_9.Z.n33 Vbias 1.88076f
C7202 CDAC8_0.switch_9.Z.n34 Vbias 1.32914f
C7203 CDAC8_0.switch_9.Z.n35 Vbias 1.3012f
C7204 CDAC8_0.switch_9.Z.n36 Vbias 0.01846f
C7205 CDAC8_0.switch_9.Z.t0 Vbias 0.03608f
C7206 CDAC8_0.switch_9.Z.n37 Vbias 0.149f
C7207 D_FlipFlop_2.3-input-nand_2.C.t7 Vbias 0.3425f
C7208 D_FlipFlop_2.3-input-nand_2.C.n0 Vbias 0.3551f
C7209 D_FlipFlop_2.3-input-nand_2.C.n1 Vbias 0.03842f
C7210 D_FlipFlop_2.3-input-nand_2.C.t1 Vbias 0.04477f
C7211 D_FlipFlop_2.3-input-nand_2.C.n2 Vbias 0.11971f
C7212 D_FlipFlop_2.3-input-nand_2.C.n3 Vbias 0.09193f
C7213 D_FlipFlop_2.3-input-nand_2.C.t4 Vbias 0.17806f
C7214 D_FlipFlop_2.3-input-nand_2.C.t5 Vbias 0.34248f
C7215 D_FlipFlop_2.3-input-nand_2.C.n4 Vbias 0.10005f
C7216 D_FlipFlop_2.3-input-nand_2.C.n5 Vbias 0.04279f
C7217 D_FlipFlop_2.3-input-nand_2.C.n6 Vbias 0.079f
C7218 D_FlipFlop_2.3-input-nand_2.C.n7 Vbias 0.13677f
C7219 D_FlipFlop_2.3-input-nand_2.C.n8 Vbias 0.10181f
C7220 D_FlipFlop_2.3-input-nand_2.C.n9 Vbias 0.04823f
C7221 D_FlipFlop_2.3-input-nand_2.C.n10 Vbias 0.124f
C7222 D_FlipFlop_2.3-input-nand_2.C.t0 Vbias 0.04742f
C7223 D_FlipFlop_2.3-input-nand_2.C.t2 Vbias 0.04645f
C7224 D_FlipFlop_2.3-input-nand_2.C.n11 Vbias 0.26418f
C7225 D_FlipFlop_2.3-input-nand_2.C.n12 Vbias 0.08722f
C7226 D_FlipFlop_2.3-input-nand_2.C.t3 Vbias 0.04645f
C7227 D_FlipFlop_2.3-input-nand_2.C.n13 Vbias 0.293f
C7228 D_FlipFlop_2.3-input-nand_2.C.t6 Vbias 0.17045f
C7229 D_FlipFlop_2.3-input-nand_2.C.n14 Vbias 0.05129f
C7230 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t1 Vbias 0.04607f
C7231 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n0 Vbias 0.10477f
C7232 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n1 Vbias 0.05057f
C7233 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t2 Vbias 0.35243f
C7234 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n2 Vbias 0.3654f
C7235 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n3 Vbias 0.03953f
C7236 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n4 Vbias 0.05278f
C7237 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t5 Vbias 0.27708f
C7238 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t4 Vbias 0.27709f
C7239 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n5 Vbias 0.17949f
C7240 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n6 Vbias 0.03786f
C7241 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t3 Vbias 0.35241f
C7242 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n7 Vbias 0.10295f
C7243 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n8 Vbias 0.02562f
C7244 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n9 Vbias 0.03726f
C7245 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n10 Vbias 0.09548f
C7246 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n11 Vbias 0.09548f
C7247 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n12 Vbias 0.04963f
C7248 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.t0 Vbias 0.04792f
C7249 RingCounter_0.D_FlipFlop_13.Inverter_1.Vout.n13 Vbias 0.28399f
C7250 And_Gate_3.Vout.t1 Vbias 0.08912f
C7251 And_Gate_3.Inverter_0.Vout Vbias 0.02589f
C7252 And_Gate_3.Vout.n0 Vbias 0.09833f
C7253 And_Gate_3.Vout.t5 Vbias 0.68307f
C7254 D_FlipFlop_4.3-input-nand_0.C Vbias -0.40609f
C7255 And_Gate_3.Vout.n1 Vbias 0.70821f
C7256 And_Gate_3.Vout.n2 Vbias 0.07662f
C7257 And_Gate_3.Vout.n3 Vbias 0.1023f
C7258 And_Gate_3.Vout.t3 Vbias 0.31442f
C7259 D_FlipFlop_4.CLK Vbias -0.02336f
C7260 And_Gate_3.Vout.n4 Vbias 0.2457f
C7261 And_Gate_3.Vout.t2 Vbias 0.68304f
C7262 D_FlipFlop_4.3-input-nand_1.C Vbias -0.22831f
C7263 And_Gate_3.Vout.t4 Vbias 0.35514f
C7264 D_FlipFlop_4.Inverter_1.Vin Vbias -0.22174f
C7265 And_Gate_3.Vout.n5 Vbias 0.37451f
C7266 And_Gate_3.Vout.t7 Vbias 0.68304f
C7267 And_Gate_3.Vout.n6 Vbias 0.60464f
C7268 And_Gate_3.Vout.n7 Vbias 0.6063f
C7269 And_Gate_3.Vout.n8 Vbias 0.37942f
C7270 And_Gate_3.Vout.t6 Vbias 0.31441f
C7271 And_Gate_3.Vout.n9 Vbias 0.06377f
C7272 And_Gate_3.Vout.n10 Vbias 0.15007f
C7273 And_Gate_3.Vout.n11 Vbias 6.09909f
C7274 And_Gate_3.Vout.t0 Vbias 0.09306f
C7275 And_Gate_3.Vout.n12 Vbias 4.81721f
C7276 And_Gate_3.Vout.n13 Vbias 0.21212f
C7277 And_Gate_7.Vout.t1 Vbias 0.0601f
C7278 And_Gate_7.Inverter_0.Vout Vbias -0.13238f
C7279 And_Gate_7.Vout.t3 Vbias 0.46171f
C7280 D_FlipFlop_0.3-input-nand_0.C Vbias -0.27449f
C7281 And_Gate_7.Vout.n0 Vbias 0.47871f
C7282 And_Gate_7.Vout.n1 Vbias 0.05179f
C7283 And_Gate_7.Vout.n2 Vbias 0.06915f
C7284 And_Gate_7.Vout.t6 Vbias 0.21251f
C7285 And_Gate_7.Vout.n3 Vbias 0.19074f
C7286 And_Gate_7.Vout.n4 Vbias 0.06086f
C7287 And_Gate_7.Vout.t5 Vbias 0.46169f
C7288 D_FlipFlop_0.3-input-nand_1.C Vbias -0.15432f
C7289 And_Gate_7.Vout.t7 Vbias 0.24006f
C7290 D_FlipFlop_0.Inverter_1.Vin Vbias -0.14989f
C7291 And_Gate_7.Vout.n5 Vbias 0.25315f
C7292 And_Gate_7.Vout.t4 Vbias 0.46169f
C7293 And_Gate_7.Vout.n6 Vbias 0.4087f
C7294 And_Gate_7.Vout.n7 Vbias 0.40982f
C7295 And_Gate_7.Vout.n8 Vbias 0.25646f
C7296 And_Gate_7.Vout.t2 Vbias 0.21252f
C7297 And_Gate_7.Vout.n9 Vbias 0.01225f
C7298 And_Gate_7.Vout.n10 Vbias 0.03152f
C7299 And_Gate_7.Vout.n11 Vbias 1.48264f
C7300 And_Gate_7.Vout.n12 Vbias 0.85866f
C7301 And_Gate_7.Vout.n13 Vbias 0.01206f
C7302 And_Gate_7.Vout.n14 Vbias 0.06203f
C7303 And_Gate_7.Vout.t0 Vbias 0.06278f
C7304 And_Gate_7.Vout.n15 Vbias 0.40066f
C7305 And_Gate_4.Vout.t1 Vbias 0.1132f
C7306 And_Gate_4.Inverter_0.Vout Vbias -0.36385f
C7307 And_Gate_4.Vout.n0 Vbias 0.06429f
C7308 And_Gate_4.Vout.n1 Vbias 0.12449f
C7309 And_Gate_4.Vout.t5 Vbias 0.86757f
C7310 D_FlipFlop_2.3-input-nand_0.C Vbias -0.51578f
C7311 And_Gate_4.Vout.n2 Vbias 0.89951f
C7312 And_Gate_4.Vout.n3 Vbias 0.09731f
C7313 And_Gate_4.Vout.n4 Vbias 0.12993f
C7314 And_Gate_4.Vout.t6 Vbias 0.39932f
C7315 D_FlipFlop_2.CLK Vbias 0.05804f
C7316 And_Gate_4.Vout.n5 Vbias 0.3804f
C7317 And_Gate_4.Vout.n6 Vbias 0.11436f
C7318 And_Gate_4.Vout.t4 Vbias 0.86753f
C7319 D_FlipFlop_2.3-input-nand_1.C Vbias -0.28998f
C7320 And_Gate_4.Vout.t7 Vbias 0.45107f
C7321 D_FlipFlop_2.Inverter_1.Vin Vbias -0.28164f
C7322 And_Gate_4.Vout.n7 Vbias 0.47567f
C7323 And_Gate_4.Vout.t3 Vbias 0.86753f
C7324 And_Gate_4.Vout.n8 Vbias 0.76796f
C7325 And_Gate_4.Vout.n9 Vbias 0.77006f
C7326 And_Gate_4.Vout.n10 Vbias 0.4819f
C7327 And_Gate_4.Vout.t2 Vbias 0.39933f
C7328 And_Gate_4.Vout.n11 Vbias 15.5365f
C7329 And_Gate_4.Vout.n12 Vbias 12.546f
C7330 And_Gate_4.Vout.n13 Vbias 0.12217f
C7331 And_Gate_4.Vout.t0 Vbias 0.11796f
C7332 And_Gate_4.Vout.n14 Vbias 0.69909f
C7333 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t2 Vbias 0.0608f
C7334 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C7335 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C7336 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C7337 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C7338 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C7339 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C7340 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C7341 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C7342 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C7343 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C7344 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C7345 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C7346 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t1 Vbias 0.06323f
C7347 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C7348 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C7349 RingCounter_0.D_FlipFlop_14.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C7350 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t1 Vbias 0.04607f
C7351 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n0 Vbias 0.10477f
C7352 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n1 Vbias 0.05057f
C7353 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t4 Vbias 0.35243f
C7354 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n2 Vbias 0.3654f
C7355 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n3 Vbias 0.03953f
C7356 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n4 Vbias 0.05278f
C7357 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t3 Vbias 0.27708f
C7358 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t2 Vbias 0.27709f
C7359 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n5 Vbias 0.17949f
C7360 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n6 Vbias 0.03786f
C7361 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t5 Vbias 0.35241f
C7362 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n7 Vbias 0.10295f
C7363 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n8 Vbias 0.02562f
C7364 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n9 Vbias 0.03726f
C7365 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n10 Vbias 0.09548f
C7366 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n11 Vbias 0.09548f
C7367 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n12 Vbias 0.04963f
C7368 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.t0 Vbias 0.04792f
C7369 RingCounter_0.D_FlipFlop_14.Inverter_1.Vout.n13 Vbias 0.28399f
C7370 Nand_Gate_2.B.t10 Vbias 0.33127f
C7371 Nand_Gate_2.B.n0 Vbias 0.09677f
C7372 Nand_Gate_2.B.n1 Vbias 0.04199f
C7373 Nand_Gate_2.B.n2 Vbias 0.18462f
C7374 Nand_Gate_2.B.t5 Vbias 0.15408f
C7375 Nand_Gate_2.B.n3 Vbias 0.04834f
C7376 Nand_Gate_2.B.t2 Vbias 0.04321f
C7377 Nand_Gate_2.B.n4 Vbias 0.18816f
C7378 Nand_Gate_2.B.n5 Vbias 0.04665f
C7379 Nand_Gate_2.B.t7 Vbias 0.33129f
C7380 Nand_Gate_2.B.n6 Vbias 0.32557f
C7381 Nand_Gate_2.B.n7 Vbias 0.03558f
C7382 Nand_Gate_2.B.t4 Vbias 0.17224f
C7383 Nand_Gate_2.B.n8 Vbias 0.04961f
C7384 Nand_Gate_2.B.n9 Vbias 0.02126f
C7385 Nand_Gate_2.B.n10 Vbias 0.03984f
C7386 Nand_Gate_2.B.n11 Vbias 0.05014f
C7387 Nand_Gate_2.B.t6 Vbias 0.33129f
C7388 Nand_Gate_2.B.n12 Vbias 0.32557f
C7389 Nand_Gate_2.B.n13 Vbias 0.03558f
C7390 Nand_Gate_2.B.t8 Vbias 0.17224f
C7391 Nand_Gate_2.B.n14 Vbias 0.04961f
C7392 Nand_Gate_2.B.n15 Vbias 0.02126f
C7393 Nand_Gate_2.B.n16 Vbias 0.03984f
C7394 Nand_Gate_2.B.n18 Vbias 0.15033f
C7395 Nand_Gate_2.B.n19 Vbias 0.41862f
C7396 Nand_Gate_2.B.n20 Vbias 0.18785f
C7397 Nand_Gate_2.B.t11 Vbias 0.17224f
C7398 Nand_Gate_2.B.t9 Vbias 0.33127f
C7399 Nand_Gate_2.B.n21 Vbias 0.09677f
C7400 Nand_Gate_2.B.n22 Vbias 0.04139f
C7401 Nand_Gate_2.B.n23 Vbias 0.07641f
C7402 Nand_Gate_2.B.n24 Vbias 0.87221f
C7403 Nand_Gate_2.B.n25 Vbias 1.18609f
C7404 Nand_Gate_2.B.n26 Vbias 0.05328f
C7405 Nand_Gate_2.B.n27 Vbias 0.01961f
C7406 Nand_Gate_2.B.n29 Vbias 0.05379f
C7407 Nand_Gate_2.B.n30 Vbias 0.02717f
C7408 Nand_Gate_2.B.t0 Vbias 0.04587f
C7409 Nand_Gate_2.B.t1 Vbias 0.04493f
C7410 Nand_Gate_2.B.n31 Vbias 0.25554f
C7411 Nand_Gate_2.B.n32 Vbias 0.08338f
C7412 Nand_Gate_2.B.t3 Vbias 0.04493f
C7413 Nand_Gate_2.B.n33 Vbias 0.06922f
C7414 Nand_Gate_2.B.n34 Vbias 0.12256f
C7415 And_Gate_1.Vout.t1 Vbias 0.08622f
C7416 And_Gate_1.Inverter_0.Vout Vbias 0.02505f
C7417 And_Gate_1.Vout.n0 Vbias 0.09513f
C7418 And_Gate_1.Vout.t6 Vbias 0.66083f
C7419 D_FlipFlop_7.3-input-nand_0.C Vbias -0.39286f
C7420 And_Gate_1.Vout.n1 Vbias 0.68515f
C7421 And_Gate_1.Vout.n2 Vbias 0.07412f
C7422 And_Gate_1.Vout.n3 Vbias 0.09897f
C7423 And_Gate_1.Vout.t3 Vbias 0.30416f
C7424 D_FlipFlop_7.CLK Vbias -0.06024f
C7425 And_Gate_1.Vout.n4 Vbias 0.24717f
C7426 And_Gate_1.Vout.n5 Vbias 0.08711f
C7427 And_Gate_1.Vout.t2 Vbias 0.6608f
C7428 D_FlipFlop_7.3-input-nand_1.C Vbias -0.22088f
C7429 And_Gate_1.Vout.t4 Vbias 0.34358f
C7430 D_FlipFlop_7.Inverter_1.Vin Vbias -0.21452f
C7431 And_Gate_1.Vout.n6 Vbias 0.36232f
C7432 And_Gate_1.Vout.t7 Vbias 0.6608f
C7433 And_Gate_1.Vout.n7 Vbias 0.58495f
C7434 And_Gate_1.Vout.n8 Vbias 0.58655f
C7435 And_Gate_1.Vout.n9 Vbias 0.36707f
C7436 And_Gate_1.Vout.t5 Vbias 0.30417f
C7437 And_Gate_1.Vout.n10 Vbias 0.04337f
C7438 And_Gate_1.Vout.n11 Vbias 0.10365f
C7439 And_Gate_1.Vout.n12 Vbias 16.2797f
C7440 And_Gate_1.Vout.t0 Vbias 0.09003f
C7441 And_Gate_1.Vout.n13 Vbias 13.6324f
C7442 And_Gate_1.Vout.n14 Vbias 0.20521f
C7443 Nand_Gate_2.A.t8 Vbias 0.62844f
C7444 Nand_Gate_2.A.n0 Vbias 0.18359f
C7445 Nand_Gate_2.A.n1 Vbias 0.07966f
C7446 Nand_Gate_2.A.n2 Vbias 0.35024f
C7447 Nand_Gate_2.A.t11 Vbias 0.2923f
C7448 Nand_Gate_2.A.n3 Vbias 0.0917f
C7449 Nand_Gate_2.A.t2 Vbias 0.08197f
C7450 Nand_Gate_2.A.n4 Vbias 0.35696f
C7451 Nand_Gate_2.A.n5 Vbias 0.0885f
C7452 Nand_Gate_2.A.t16 Vbias 0.62847f
C7453 Nand_Gate_2.A.n6 Vbias 0.61763f
C7454 Nand_Gate_2.A.n7 Vbias 0.06751f
C7455 Nand_Gate_2.A.t17 Vbias 0.32674f
C7456 Nand_Gate_2.A.n8 Vbias 0.09412f
C7457 Nand_Gate_2.A.n9 Vbias 0.04034f
C7458 Nand_Gate_2.A.n10 Vbias 0.07558f
C7459 Nand_Gate_2.A.n11 Vbias 0.09511f
C7460 Nand_Gate_2.A.t4 Vbias 0.62847f
C7461 Nand_Gate_2.A.n12 Vbias 0.61763f
C7462 Nand_Gate_2.A.n13 Vbias 0.06751f
C7463 Nand_Gate_2.A.t15 Vbias 0.32674f
C7464 Nand_Gate_2.A.n14 Vbias 0.09412f
C7465 Nand_Gate_2.A.n15 Vbias 0.04034f
C7466 Nand_Gate_2.A.n16 Vbias 0.07558f
C7467 Nand_Gate_2.A.n17 Vbias 0.01133f
C7468 Nand_Gate_2.A.n18 Vbias 0.28519f
C7469 Nand_Gate_2.A.n19 Vbias 0.79416f
C7470 Nand_Gate_2.A.n20 Vbias 0.35636f
C7471 Nand_Gate_2.A.t6 Vbias 0.62847f
C7472 Nand_Gate_2.A.n21 Vbias 0.6329f
C7473 Nand_Gate_2.A.n22 Vbias 0.06751f
C7474 Nand_Gate_2.A.t9 Vbias 0.32674f
C7475 Nand_Gate_2.A.n23 Vbias 0.09412f
C7476 Nand_Gate_2.A.n24 Vbias 0.02507f
C7477 Nand_Gate_2.A.n25 Vbias 0.03906f
C7478 Nand_Gate_2.A.n26 Vbias 0.38975f
C7479 Nand_Gate_2.A.t10 Vbias 0.62847f
C7480 Nand_Gate_2.A.n27 Vbias 0.6329f
C7481 Nand_Gate_2.A.n28 Vbias 0.06751f
C7482 Nand_Gate_2.A.t5 Vbias 0.32674f
C7483 Nand_Gate_2.A.n29 Vbias 0.09412f
C7484 Nand_Gate_2.A.n30 Vbias 0.02507f
C7485 Nand_Gate_2.A.n31 Vbias 0.03906f
C7486 Nand_Gate_2.A.n32 Vbias 0.01133f
C7487 Nand_Gate_2.A.n33 Vbias 1.01202f
C7488 Nand_Gate_2.A.n34 Vbias 0.47041f
C7489 Nand_Gate_2.A.n35 Vbias 0.17479f
C7490 Nand_Gate_2.A.t13 Vbias 0.62844f
C7491 Nand_Gate_2.A.n36 Vbias 0.18359f
C7492 Nand_Gate_2.A.n37 Vbias 0.07966f
C7493 Nand_Gate_2.A.n38 Vbias 0.35024f
C7494 Nand_Gate_2.A.t7 Vbias 0.29227f
C7495 Nand_Gate_2.A.n39 Vbias 0.03875f
C7496 Nand_Gate_2.A.n40 Vbias 0.09293f
C7497 Nand_Gate_2.A.n41 Vbias 8.01087f
C7498 Nand_Gate_2.A.t14 Vbias 0.32676f
C7499 Nand_Gate_2.A.n42 Vbias 0.32008f
C7500 Nand_Gate_2.A.n43 Vbias 0.06751f
C7501 Nand_Gate_2.A.t12 Vbias 0.62844f
C7502 Nand_Gate_2.A.n44 Vbias 0.18359f
C7503 Nand_Gate_2.A.n45 Vbias 0.04568f
C7504 Nand_Gate_2.A.n46 Vbias 0.06645f
C7505 Nand_Gate_2.A.n47 Vbias 0.09785f
C7506 Nand_Gate_2.A.n48 Vbias 9.45741f
C7507 Nand_Gate_2.A.n49 Vbias 0.34581f
C7508 Nand_Gate_2.A.n50 Vbias 0.10108f
C7509 Nand_Gate_2.A.n51 Vbias 0.0372f
C7510 Nand_Gate_2.A.n52 Vbias 0.01151f
C7511 Nand_Gate_2.A.n53 Vbias 0.10205f
C7512 Nand_Gate_2.A.n54 Vbias 0.05153f
C7513 Nand_Gate_2.A.t0 Vbias 0.08702f
C7514 Nand_Gate_2.A.t3 Vbias 0.08524f
C7515 Nand_Gate_2.A.n55 Vbias 0.48477f
C7516 Nand_Gate_2.A.n56 Vbias 0.15818f
C7517 Nand_Gate_2.A.t1 Vbias 0.08524f
C7518 Nand_Gate_2.A.n57 Vbias 0.13131f
C7519 Nand_Gate_2.A.n58 Vbias 0.2325f
C7520 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t2 Vbias 0.07024f
C7521 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n0 Vbias 0.03989f
C7522 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n1 Vbias 0.07725f
C7523 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t4 Vbias 0.2799f
C7524 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n2 Vbias 0.27418f
C7525 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n3 Vbias 0.05783f
C7526 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t5 Vbias 0.53832f
C7527 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n4 Vbias 0.15726f
C7528 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n5 Vbias 0.03913f
C7529 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n6 Vbias 0.05692f
C7530 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n7 Vbias 0.14585f
C7531 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n8 Vbias 0.14585f
C7532 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n9 Vbias 0.07581f
C7533 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t3 Vbias 0.07318f
C7534 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t0 Vbias 0.07454f
C7535 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.t1 Vbias 0.07302f
C7536 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n10 Vbias 0.41525f
C7537 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n11 Vbias 0.23391f
C7538 RingCounter_0.D_FlipFlop_3.3-input-nand_1.Vout.n12 Vbias 0.22303f
C7539 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t1 Vbias 0.06624f
C7540 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t2 Vbias 0.07883f
C7541 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n0 Vbias 0.39844f
C7542 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n1 Vbias 0.20187f
C7543 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n2 Vbias 0.06862f
C7544 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t3 Vbias 0.25335f
C7545 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n3 Vbias 0.24817f
C7546 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n4 Vbias 0.05234f
C7547 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t4 Vbias 0.48726f
C7548 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n5 Vbias 0.14234f
C7549 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n6 Vbias 0.03542f
C7550 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n7 Vbias 0.05152f
C7551 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n8 Vbias 0.13202f
C7552 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n9 Vbias 0.13202f
C7553 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n10 Vbias 0.06992f
C7554 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.n11 Vbias 0.03611f
C7555 RingCounter_0.D_FlipFlop_1.Nand_Gate_1.Vout.t0 Vbias 0.06358f
C7556 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t1 Vbias 0.04998f
C7557 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n0 Vbias 0.02839f
C7558 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n1 Vbias 0.05497f
C7559 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t5 Vbias 0.38308f
C7560 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n2 Vbias 0.39717f
C7561 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n3 Vbias 0.04297f
C7562 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n4 Vbias 0.05737f
C7563 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t4 Vbias 0.30118f
C7564 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t3 Vbias 0.30119f
C7565 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n5 Vbias 0.1951f
C7566 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n6 Vbias 0.04115f
C7567 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t2 Vbias 0.38306f
C7568 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n7 Vbias 0.1119f
C7569 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n8 Vbias 0.02784f
C7570 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n9 Vbias 0.0405f
C7571 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n10 Vbias 0.10379f
C7572 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n11 Vbias 0.10379f
C7573 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n12 Vbias 0.05395f
C7574 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.t0 Vbias 0.05208f
C7575 RingCounter_0.D_FlipFlop_1.Inverter_1.Vout.n13 Vbias 0.30868f
C7576 Nand_Gate_0.A.t9 Vbias 0.75629f
C7577 Nand_Gate_0.A.n0 Vbias 0.22093f
C7578 Nand_Gate_0.A.n1 Vbias 0.09586f
C7579 Nand_Gate_0.A.n2 Vbias 0.42149f
C7580 Nand_Gate_0.A.t13 Vbias 0.35177f
C7581 Nand_Gate_0.A.n3 Vbias 0.11036f
C7582 Nand_Gate_0.A.t2 Vbias 0.09865f
C7583 Nand_Gate_0.A.n4 Vbias 0.42957f
C7584 Nand_Gate_0.A.n5 Vbias 0.10651f
C7585 Nand_Gate_0.A.t14 Vbias 0.75632f
C7586 Nand_Gate_0.A.n6 Vbias 0.74327f
C7587 Nand_Gate_0.A.n7 Vbias 0.08124f
C7588 Nand_Gate_0.A.t8 Vbias 0.39321f
C7589 Nand_Gate_0.A.n8 Vbias 0.11327f
C7590 Nand_Gate_0.A.n9 Vbias 0.04854f
C7591 Nand_Gate_0.A.n10 Vbias 0.09095f
C7592 Nand_Gate_0.A.n11 Vbias 0.11446f
C7593 Nand_Gate_0.A.t7 Vbias 0.75632f
C7594 Nand_Gate_0.A.n12 Vbias 0.74327f
C7595 Nand_Gate_0.A.n13 Vbias 0.08124f
C7596 Nand_Gate_0.A.t12 Vbias 0.39321f
C7597 Nand_Gate_0.A.n14 Vbias 0.11327f
C7598 Nand_Gate_0.A.n15 Vbias 0.04854f
C7599 Nand_Gate_0.A.n16 Vbias 0.09095f
C7600 Nand_Gate_0.A.n17 Vbias 0.01364f
C7601 Nand_Gate_0.A.n18 Vbias 0.34321f
C7602 Nand_Gate_0.A.n19 Vbias 0.95571f
C7603 Nand_Gate_0.A.n20 Vbias 0.42885f
C7604 Nand_Gate_0.A.t15 Vbias 0.75632f
C7605 Nand_Gate_0.A.n21 Vbias 0.76165f
C7606 Nand_Gate_0.A.n22 Vbias 0.08124f
C7607 Nand_Gate_0.A.t17 Vbias 0.39321f
C7608 Nand_Gate_0.A.n23 Vbias 0.11327f
C7609 Nand_Gate_0.A.n24 Vbias 0.03017f
C7610 Nand_Gate_0.A.n25 Vbias 0.04701f
C7611 Nand_Gate_0.A.n26 Vbias 0.46904f
C7612 Nand_Gate_0.A.t6 Vbias 0.75632f
C7613 Nand_Gate_0.A.n27 Vbias 0.76165f
C7614 Nand_Gate_0.A.n28 Vbias 0.08124f
C7615 Nand_Gate_0.A.t10 Vbias 0.39321f
C7616 Nand_Gate_0.A.n29 Vbias 0.11327f
C7617 Nand_Gate_0.A.n30 Vbias 0.03017f
C7618 Nand_Gate_0.A.n31 Vbias 0.04701f
C7619 Nand_Gate_0.A.n32 Vbias 0.01364f
C7620 Nand_Gate_0.A.n33 Vbias 1.2179f
C7621 Nand_Gate_0.A.n34 Vbias 0.5679f
C7622 Nand_Gate_0.A.n35 Vbias 0.21035f
C7623 Nand_Gate_0.A.t5 Vbias 0.75629f
C7624 Nand_Gate_0.A.n36 Vbias 0.22093f
C7625 Nand_Gate_0.A.n37 Vbias 0.09586f
C7626 Nand_Gate_0.A.n38 Vbias 0.42149f
C7627 Nand_Gate_0.A.t16 Vbias 0.35173f
C7628 Nand_Gate_0.A.n39 Vbias 0.04484f
C7629 Nand_Gate_0.A.n40 Vbias 0.10776f
C7630 Nand_Gate_0.A.n41 Vbias 14.747f
C7631 Nand_Gate_0.A.t11 Vbias 0.39323f
C7632 Nand_Gate_0.A.n42 Vbias 0.38519f
C7633 Nand_Gate_0.A.n43 Vbias 0.08124f
C7634 Nand_Gate_0.A.t4 Vbias 0.75629f
C7635 Nand_Gate_0.A.n44 Vbias 0.22093f
C7636 Nand_Gate_0.A.n45 Vbias 0.05497f
C7637 Nand_Gate_0.A.n46 Vbias 0.07997f
C7638 Nand_Gate_0.A.n47 Vbias 0.11775f
C7639 Nand_Gate_0.A.n48 Vbias 16.5226f
C7640 Nand_Gate_0.A.n49 Vbias 0.41616f
C7641 Nand_Gate_0.A.n50 Vbias 0.12165f
C7642 Nand_Gate_0.A.n51 Vbias 0.04477f
C7643 Nand_Gate_0.A.n52 Vbias 0.01385f
C7644 Nand_Gate_0.A.n53 Vbias 0.12281f
C7645 Nand_Gate_0.A.n54 Vbias 0.06202f
C7646 Nand_Gate_0.A.t0 Vbias 0.10473f
C7647 Nand_Gate_0.A.t1 Vbias 0.10258f
C7648 Nand_Gate_0.A.n55 Vbias 0.58338f
C7649 Nand_Gate_0.A.n56 Vbias 0.19036f
C7650 Nand_Gate_0.A.t3 Vbias 0.10258f
C7651 Nand_Gate_0.A.n57 Vbias 0.15802f
C7652 Nand_Gate_0.A.n58 Vbias 0.2798f
C7653 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t2 Vbias 0.05201f
C7654 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n0 Vbias 0.22649f
C7655 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n1 Vbias 0.05616f
C7656 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t5 Vbias 0.39877f
C7657 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n2 Vbias 0.39189f
C7658 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n3 Vbias 0.04283f
C7659 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t4 Vbias 0.20732f
C7660 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n4 Vbias 0.05972f
C7661 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n5 Vbias 0.02559f
C7662 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n6 Vbias 0.04796f
C7663 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n7 Vbias 0.10804f
C7664 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n8 Vbias 0.10804f
C7665 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n9 Vbias 0.06475f
C7666 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t3 Vbias 0.05421f
C7667 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t0 Vbias 0.05522f
C7668 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.t1 Vbias 0.05409f
C7669 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n10 Vbias 0.30759f
C7670 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n11 Vbias 0.17406f
C7671 RingCounter_0.D_FlipFlop_13.3-input-nand_0.Vout.n12 Vbias 0.03715f
C7672 Comparator_0.Vout Vbias 0.06753f
C7673 D_FlipFlop_0.D.t35 Vbias 0.54627f
C7674 D_FlipFlop_0.D.n0 Vbias 0.15946f
C7675 D_FlipFlop_0.D.t2 Vbias 1.91888f
C7676 D_FlipFlop_0.D.t1 Vbias 0.42801f
C7677 D_FlipFlop_0.D.n1 Vbias 1.48735f
C7678 D_FlipFlop_0.D.t0 Vbias 0.80231f
C7679 D_FlipFlop_0.D.n2 Vbias -3.54159f
C7680 D_FlipFlop_0.D.n3 Vbias 4.00296f
C7681 D_FlipFlop_0.D.n4 Vbias 1.19852f
C7682 D_FlipFlop_0.D.t20 Vbias 0.14499f
C7683 D_FlipFlop_0.Inverter_0.Vin Vbias -0.10555f
C7684 D_FlipFlop_0.D.n5 Vbias 0.14249f
C7685 D_FlipFlop_0.D.n6 Vbias 0.01557f
C7686 D_FlipFlop_0.D.t30 Vbias 0.07538f
C7687 D_FlipFlop_0.D.n7 Vbias 0.02171f
C7688 D_FlipFlop_0.D.n9 Vbias 0.01744f
C7689 D_FlipFlop_0.D.t27 Vbias 0.14499f
C7690 D_FlipFlop_0.3-input-nand_0.B Vbias -0.10555f
C7691 D_FlipFlop_0.D.n11 Vbias 0.14249f
C7692 D_FlipFlop_0.D.n12 Vbias 0.01557f
C7693 D_FlipFlop_0.D.t23 Vbias 0.07538f
C7694 D_FlipFlop_0.D.n13 Vbias 0.02171f
C7695 D_FlipFlop_0.D.n15 Vbias 0.01744f
C7696 D_FlipFlop_0.D.n16 Vbias 0.02184f
C7697 D_FlipFlop_0.D.n17 Vbias 0.10923f
C7698 D_FlipFlop_0.D.t31 Vbias 0.14499f
C7699 D_FlipFlop_3.Inverter_0.Vin Vbias -0.10555f
C7700 D_FlipFlop_0.D.n18 Vbias 0.14249f
C7701 D_FlipFlop_0.D.n19 Vbias 0.01557f
C7702 D_FlipFlop_0.D.t11 Vbias 0.07538f
C7703 D_FlipFlop_0.D.n20 Vbias 0.02171f
C7704 D_FlipFlop_0.D.n22 Vbias 0.01744f
C7705 D_FlipFlop_0.D.t4 Vbias 0.14499f
C7706 D_FlipFlop_3.3-input-nand_0.B Vbias -0.10555f
C7707 D_FlipFlop_0.D.n24 Vbias 0.14249f
C7708 D_FlipFlop_0.D.n25 Vbias 0.01557f
C7709 D_FlipFlop_0.D.t32 Vbias 0.07538f
C7710 D_FlipFlop_0.D.n26 Vbias 0.02171f
C7711 D_FlipFlop_0.D.n28 Vbias 0.01744f
C7712 D_FlipFlop_0.D.n29 Vbias 0.02184f
C7713 D_FlipFlop_0.D.n30 Vbias 0.0728f
C7714 D_FlipFlop_0.D.n31 Vbias 2.33998f
C7715 D_FlipFlop_0.D.t14 Vbias 0.14499f
C7716 D_FlipFlop_2.Inverter_0.Vin Vbias -0.10555f
C7717 D_FlipFlop_0.D.n32 Vbias 0.14249f
C7718 D_FlipFlop_0.D.n33 Vbias 0.01557f
C7719 D_FlipFlop_0.D.t17 Vbias 0.07538f
C7720 D_FlipFlop_0.D.n34 Vbias 0.02171f
C7721 D_FlipFlop_0.D.n36 Vbias 0.01744f
C7722 D_FlipFlop_0.D.t24 Vbias 0.14499f
C7723 D_FlipFlop_2.3-input-nand_0.B Vbias -0.10555f
C7724 D_FlipFlop_0.D.n38 Vbias 0.14249f
C7725 D_FlipFlop_0.D.n39 Vbias 0.01557f
C7726 D_FlipFlop_0.D.t8 Vbias 0.07538f
C7727 D_FlipFlop_0.D.n40 Vbias 0.02171f
C7728 D_FlipFlop_0.D.n42 Vbias 0.01744f
C7729 D_FlipFlop_0.D.n43 Vbias 0.02184f
C7730 D_FlipFlop_0.D.n44 Vbias 0.07368f
C7731 D_FlipFlop_0.D.n45 Vbias 1.52411f
C7732 D_FlipFlop_0.D.t19 Vbias 0.14499f
C7733 D_FlipFlop_1.Inverter_0.Vin Vbias -0.10555f
C7734 D_FlipFlop_0.D.n46 Vbias 0.14249f
C7735 D_FlipFlop_0.D.n47 Vbias 0.01557f
C7736 D_FlipFlop_0.D.t29 Vbias 0.07538f
C7737 D_FlipFlop_0.D.n48 Vbias 0.02171f
C7738 D_FlipFlop_0.D.n50 Vbias 0.01744f
C7739 D_FlipFlop_0.D.t26 Vbias 0.14499f
C7740 D_FlipFlop_1.3-input-nand_0.B Vbias -0.10555f
C7741 D_FlipFlop_0.D.n52 Vbias 0.14249f
C7742 D_FlipFlop_0.D.n53 Vbias 0.01557f
C7743 D_FlipFlop_0.D.t22 Vbias 0.07538f
C7744 D_FlipFlop_0.D.n54 Vbias 0.02171f
C7745 D_FlipFlop_0.D.n56 Vbias 0.01744f
C7746 D_FlipFlop_0.D.n57 Vbias 0.02184f
C7747 D_FlipFlop_0.D.n58 Vbias 0.07308f
C7748 D_FlipFlop_0.D.n59 Vbias 1.95548f
C7749 D_FlipFlop_0.D.t21 Vbias 0.14499f
C7750 D_FlipFlop_4.Inverter_0.Vin Vbias -0.10555f
C7751 D_FlipFlop_0.D.n60 Vbias 0.14249f
C7752 D_FlipFlop_0.D.n61 Vbias 0.01557f
C7753 D_FlipFlop_0.D.t13 Vbias 0.07538f
C7754 D_FlipFlop_0.D.n62 Vbias 0.02171f
C7755 D_FlipFlop_0.D.n64 Vbias 0.01744f
C7756 D_FlipFlop_0.D.t28 Vbias 0.14499f
C7757 D_FlipFlop_4.3-input-nand_0.B Vbias -0.10555f
C7758 D_FlipFlop_0.D.n66 Vbias 0.14249f
C7759 D_FlipFlop_0.D.n67 Vbias 0.01557f
C7760 D_FlipFlop_0.D.t3 Vbias 0.07538f
C7761 D_FlipFlop_0.D.n68 Vbias 0.02171f
C7762 D_FlipFlop_0.D.n70 Vbias 0.01744f
C7763 D_FlipFlop_0.D.n71 Vbias 0.02184f
C7764 D_FlipFlop_0.D.n72 Vbias 0.07316f
C7765 D_FlipFlop_0.D.n73 Vbias 1.95555f
C7766 D_FlipFlop_0.D.t33 Vbias 0.14499f
C7767 D_FlipFlop_7.Inverter_0.Vin Vbias -0.10555f
C7768 D_FlipFlop_0.D.n74 Vbias 0.14249f
C7769 D_FlipFlop_0.D.n75 Vbias 0.01557f
C7770 D_FlipFlop_0.D.t12 Vbias 0.07538f
C7771 D_FlipFlop_0.D.n76 Vbias 0.02171f
C7772 D_FlipFlop_0.D.n78 Vbias 0.01744f
C7773 D_FlipFlop_0.D.t6 Vbias 0.14499f
C7774 D_FlipFlop_7.3-input-nand_0.B Vbias -0.10555f
C7775 D_FlipFlop_0.D.n80 Vbias 0.14249f
C7776 D_FlipFlop_0.D.n81 Vbias 0.01557f
C7777 D_FlipFlop_0.D.t34 Vbias 0.07538f
C7778 D_FlipFlop_0.D.n82 Vbias 0.02171f
C7779 D_FlipFlop_0.D.n84 Vbias 0.01744f
C7780 D_FlipFlop_0.D.n85 Vbias 0.02184f
C7781 D_FlipFlop_0.D.n86 Vbias 0.11007f
C7782 D_FlipFlop_0.D.t15 Vbias 0.14499f
C7783 D_FlipFlop_6.Inverter_0.Vin Vbias -0.10555f
C7784 D_FlipFlop_0.D.n87 Vbias 0.14249f
C7785 D_FlipFlop_0.D.n88 Vbias 0.01557f
C7786 D_FlipFlop_0.D.t18 Vbias 0.07538f
C7787 D_FlipFlop_0.D.n89 Vbias 0.02171f
C7788 D_FlipFlop_0.D.n91 Vbias 0.01744f
C7789 D_FlipFlop_0.D.t25 Vbias 0.14499f
C7790 D_FlipFlop_6.3-input-nand_0.B Vbias -0.10555f
C7791 D_FlipFlop_0.D.n93 Vbias 0.14249f
C7792 D_FlipFlop_0.D.n94 Vbias 0.01557f
C7793 D_FlipFlop_0.D.t9 Vbias 0.07538f
C7794 D_FlipFlop_0.D.n95 Vbias 0.02171f
C7795 D_FlipFlop_0.D.n97 Vbias 0.01744f
C7796 D_FlipFlop_0.D.n98 Vbias 0.02184f
C7797 D_FlipFlop_0.D.n99 Vbias 0.07276f
C7798 D_FlipFlop_0.D.n100 Vbias 2.34064f
C7799 D_FlipFlop_0.D.n101 Vbias 1.45564f
C7800 D_FlipFlop_0.D.t5 Vbias 0.14499f
C7801 D_FlipFlop_5.Inverter_0.Vin Vbias -0.10555f
C7802 D_FlipFlop_0.D.n102 Vbias 0.14249f
C7803 D_FlipFlop_0.D.n103 Vbias 0.01557f
C7804 D_FlipFlop_0.D.t16 Vbias 0.07538f
C7805 D_FlipFlop_0.D.n104 Vbias 0.02171f
C7806 D_FlipFlop_0.D.n106 Vbias 0.01744f
C7807 D_FlipFlop_0.D.t10 Vbias 0.14499f
C7808 D_FlipFlop_5.3-input-nand_0.B Vbias -0.10555f
C7809 D_FlipFlop_0.D.n108 Vbias 0.14249f
C7810 D_FlipFlop_0.D.n109 Vbias 0.01557f
C7811 D_FlipFlop_0.D.t7 Vbias 0.07538f
C7812 D_FlipFlop_0.D.n110 Vbias 0.02171f
C7813 D_FlipFlop_0.D.n112 Vbias 0.01744f
C7814 D_FlipFlop_0.D.n113 Vbias 0.02184f
C7815 D_FlipFlop_0.D.n114 Vbias 0.06753f
C7816 D_FlipFlop_0.D.n115 Vbias 0.1788f
C7817 D_FlipFlop_0.D.n116 Vbias 0.99323f
C7818 D_FlipFlop_0.D.n117 Vbias 0.49764f
C7819 D_FlipFlop_1.3-input-nand_2.C.t6 Vbias 0.3425f
C7820 D_FlipFlop_1.3-input-nand_2.C.n0 Vbias 0.3551f
C7821 D_FlipFlop_1.3-input-nand_2.C.n1 Vbias 0.03842f
C7822 D_FlipFlop_1.3-input-nand_2.C.t2 Vbias 0.04477f
C7823 D_FlipFlop_1.3-input-nand_2.C.n2 Vbias 0.11971f
C7824 D_FlipFlop_1.3-input-nand_2.C.n3 Vbias 0.09193f
C7825 D_FlipFlop_1.3-input-nand_2.C.t4 Vbias 0.17806f
C7826 D_FlipFlop_1.3-input-nand_2.C.t5 Vbias 0.34248f
C7827 D_FlipFlop_1.3-input-nand_2.C.n4 Vbias 0.10005f
C7828 D_FlipFlop_1.3-input-nand_2.C.n5 Vbias 0.04279f
C7829 D_FlipFlop_1.3-input-nand_2.C.n6 Vbias 0.079f
C7830 D_FlipFlop_1.3-input-nand_2.C.n7 Vbias 0.13677f
C7831 D_FlipFlop_1.3-input-nand_2.C.n8 Vbias 0.10181f
C7832 D_FlipFlop_1.3-input-nand_2.C.n9 Vbias 0.04823f
C7833 D_FlipFlop_1.3-input-nand_2.C.n10 Vbias 0.124f
C7834 D_FlipFlop_1.3-input-nand_2.C.t0 Vbias 0.04742f
C7835 D_FlipFlop_1.3-input-nand_2.C.t1 Vbias 0.04645f
C7836 D_FlipFlop_1.3-input-nand_2.C.n11 Vbias 0.26418f
C7837 D_FlipFlop_1.3-input-nand_2.C.n12 Vbias 0.08722f
C7838 D_FlipFlop_1.3-input-nand_2.C.t3 Vbias 0.04645f
C7839 D_FlipFlop_1.3-input-nand_2.C.n13 Vbias 0.293f
C7840 D_FlipFlop_1.3-input-nand_2.C.t7 Vbias 0.17045f
C7841 D_FlipFlop_1.3-input-nand_2.C.n14 Vbias 0.05129f
C7842 D_FlipFlop_1.3-input-nand_2.Vout.t6 Vbias 0.35515f
C7843 D_FlipFlop_1.3-input-nand_2.Vout.n0 Vbias 0.10375f
C7844 D_FlipFlop_1.3-input-nand_2.Vout.n1 Vbias 0.04502f
C7845 D_FlipFlop_1.3-input-nand_2.Vout.n2 Vbias 0.19793f
C7846 D_FlipFlop_1.3-input-nand_2.Vout.t4 Vbias 0.17747f
C7847 D_FlipFlop_1.3-input-nand_2.Vout.t1 Vbias 0.04817f
C7848 D_FlipFlop_1.3-input-nand_2.Vout.n3 Vbias 0.30324f
C7849 D_FlipFlop_1.3-input-nand_2.Vout.t3 Vbias 0.04918f
C7850 D_FlipFlop_1.3-input-nand_2.Vout.t2 Vbias 0.04817f
C7851 D_FlipFlop_1.3-input-nand_2.Vout.n4 Vbias 0.27396f
C7852 D_FlipFlop_1.3-input-nand_2.Vout.n5 Vbias 0.09115f
C7853 D_FlipFlop_1.3-input-nand_2.Vout.n6 Vbias 0.01454f
C7854 D_FlipFlop_1.3-input-nand_2.Vout.n7 Vbias 0.01331f
C7855 D_FlipFlop_1.3-input-nand_2.Vout.t5 Vbias 0.35517f
C7856 D_FlipFlop_1.3-input-nand_2.Vout.n8 Vbias 0.36759f
C7857 D_FlipFlop_1.3-input-nand_2.Vout.t7 Vbias 0.18465f
C7858 D_FlipFlop_1.3-input-nand_2.Vout.n9 Vbias 0.18106f
C7859 D_FlipFlop_1.3-input-nand_2.Vout.n10 Vbias 0.10557f
C7860 D_FlipFlop_1.3-input-nand_2.Vout.n11 Vbias 0.05002f
C7861 D_FlipFlop_1.3-input-nand_2.Vout.t0 Vbias 0.04632f
C7862 D_FlipFlop_1.3-input-nand_2.Vout.n12 Vbias 0.22028f
C7863 CDAC8_0.switch_6.Z.t3 Vbias 0.03493f
C7864 CDAC8_0.switch_6.Z.t2 Vbias 0.0333f
C7865 CDAC8_0.switch_6.Z.t1 Vbias 0.0333f
C7866 CDAC8_0.switch_6.Z.n0 Vbias 0.1203f
C7867 CDAC8_0.switch_6.Z.n1 Vbias 0.27648f
C7868 CDAC8_0.switch_6.Z.n2 Vbias 0.03601f
C7869 CDAC8_0.switch_6.Z.n3 Vbias 1.50056f
C7870 CDAC8_0.switch_6.Z.n4 Vbias 1.08953f
C7871 CDAC8_0.switch_6.Z.t41 Vbias 5.88262f
C7872 CDAC8_0.switch_6.Z.n5 Vbias 1.36404f
C7873 CDAC8_0.switch_6.Z.t10 Vbias 5.88262f
C7874 CDAC8_0.switch_6.Z.n6 Vbias 1.36404f
C7875 CDAC8_0.switch_6.Z.t29 Vbias 5.88262f
C7876 CDAC8_0.switch_6.Z.n7 Vbias 1.36404f
C7877 CDAC8_0.switch_6.Z.t63 Vbias 5.96794f
C7878 CDAC8_0.switch_6.Z.t32 Vbias 5.96794f
C7879 CDAC8_0.switch_6.Z.n8 Vbias 2.23974f
C7880 CDAC8_0.switch_6.Z.n9 Vbias 2.23974f
C7881 CDAC8_0.switch_6.Z.t62 Vbias 5.88262f
C7882 CDAC8_0.switch_6.Z.n10 Vbias 1.36404f
C7883 CDAC8_0.switch_6.Z.n11 Vbias 1.12959f
C7884 CDAC8_0.switch_6.Z.n12 Vbias 1.12959f
C7885 CDAC8_0.switch_6.Z.t45 Vbias 5.88262f
C7886 CDAC8_0.switch_6.Z.n13 Vbias 1.36404f
C7887 CDAC8_0.switch_6.Z.n14 Vbias 1.12959f
C7888 CDAC8_0.switch_6.Z.n15 Vbias 1.12959f
C7889 CDAC8_0.switch_6.Z.t7 Vbias 5.88262f
C7890 CDAC8_0.switch_6.Z.n16 Vbias 1.36404f
C7891 CDAC8_0.switch_6.Z.t34 Vbias 5.88262f
C7892 CDAC8_0.switch_6.Z.n17 Vbias 1.36404f
C7893 CDAC8_0.switch_6.Z.n18 Vbias 1.12959f
C7894 CDAC8_0.switch_6.Z.n19 Vbias 1.12959f
C7895 CDAC8_0.switch_6.Z.t67 Vbias 5.88262f
C7896 CDAC8_0.switch_6.Z.n20 Vbias 1.36404f
C7897 CDAC8_0.switch_6.Z.t9 Vbias 5.88262f
C7898 CDAC8_0.switch_6.Z.n21 Vbias 1.36404f
C7899 CDAC8_0.switch_6.Z.t46 Vbias 5.88262f
C7900 CDAC8_0.switch_6.Z.n22 Vbias 1.36404f
C7901 CDAC8_0.switch_6.Z.t53 Vbias 5.88262f
C7902 CDAC8_0.switch_6.Z.n23 Vbias 1.36404f
C7903 CDAC8_0.switch_6.Z.t17 Vbias 5.88262f
C7904 CDAC8_0.switch_6.Z.n24 Vbias 1.36404f
C7905 CDAC8_0.switch_6.Z.t15 Vbias 5.88262f
C7906 CDAC8_0.switch_6.Z.n25 Vbias 1.36404f
C7907 CDAC8_0.switch_6.Z.t58 Vbias 5.88262f
C7908 CDAC8_0.switch_6.Z.n26 Vbias 1.36404f
C7909 CDAC8_0.switch_6.Z.t22 Vbias 5.88262f
C7910 CDAC8_0.switch_6.Z.n27 Vbias 1.36404f
C7911 CDAC8_0.switch_6.Z.t65 Vbias 5.88262f
C7912 CDAC8_0.switch_6.Z.n28 Vbias 1.36404f
C7913 CDAC8_0.switch_6.Z.t61 Vbias 5.88262f
C7914 CDAC8_0.switch_6.Z.n29 Vbias 1.36404f
C7915 CDAC8_0.switch_6.Z.t25 Vbias 5.88262f
C7916 CDAC8_0.switch_6.Z.n30 Vbias 1.36404f
C7917 CDAC8_0.switch_6.Z.t5 Vbias 6.12449f
C7918 CDAC8_0.switch_6.Z.t37 Vbias 6.12449f
C7919 CDAC8_0.switch_6.Z.n31 Vbias 2.41525f
C7920 CDAC8_0.switch_6.Z.n32 Vbias 2.41525f
C7921 CDAC8_0.switch_6.Z.t59 Vbias 5.88262f
C7922 CDAC8_0.switch_6.Z.n33 Vbias 1.36404f
C7923 CDAC8_0.switch_6.Z.n34 Vbias 1.12959f
C7924 CDAC8_0.switch_6.Z.n35 Vbias 1.12959f
C7925 CDAC8_0.switch_6.Z.t27 Vbias 5.88262f
C7926 CDAC8_0.switch_6.Z.n36 Vbias 1.36404f
C7927 CDAC8_0.switch_6.Z.n37 Vbias 1.12959f
C7928 CDAC8_0.switch_6.Z.n38 Vbias 1.12959f
C7929 CDAC8_0.switch_6.Z.t33 Vbias 5.88262f
C7930 CDAC8_0.switch_6.Z.n39 Vbias 1.36404f
C7931 CDAC8_0.switch_6.Z.n40 Vbias 1.12959f
C7932 CDAC8_0.switch_6.Z.n41 Vbias 1.12959f
C7933 CDAC8_0.switch_6.Z.t56 Vbias 5.88262f
C7934 CDAC8_0.switch_6.Z.n42 Vbias 1.24121f
C7935 CDAC8_0.switch_6.Z.n43 Vbias 0.7957f
C7936 CDAC8_0.switch_6.Z.t13 Vbias 5.88262f
C7937 CDAC8_0.switch_6.Z.n44 Vbias 1.36404f
C7938 CDAC8_0.switch_6.Z.t48 Vbias 5.88262f
C7939 CDAC8_0.switch_6.Z.n45 Vbias 1.36404f
C7940 CDAC8_0.switch_6.Z.t30 Vbias 5.88262f
C7941 CDAC8_0.switch_6.Z.n46 Vbias 1.36404f
C7942 CDAC8_0.switch_6.Z.t19 Vbias 5.88262f
C7943 CDAC8_0.switch_6.Z.n47 Vbias 1.36404f
C7944 CDAC8_0.switch_6.Z.t18 Vbias 5.88262f
C7945 CDAC8_0.switch_6.Z.n48 Vbias 1.36404f
C7946 CDAC8_0.switch_6.Z.t11 Vbias 5.88262f
C7947 CDAC8_0.switch_6.Z.n49 Vbias 1.36404f
C7948 CDAC8_0.switch_6.Z.t52 Vbias 5.88262f
C7949 CDAC8_0.switch_6.Z.n50 Vbias 1.36404f
C7950 CDAC8_0.switch_6.Z.t44 Vbias 5.88262f
C7951 CDAC8_0.switch_6.Z.n51 Vbias 1.36404f
C7952 CDAC8_0.switch_6.Z.t43 Vbias 5.88262f
C7953 CDAC8_0.switch_6.Z.n52 Vbias 1.36404f
C7954 CDAC8_0.switch_6.Z.t31 Vbias 5.96794f
C7955 CDAC8_0.switch_6.Z.t47 Vbias 5.96794f
C7956 CDAC8_0.switch_6.Z.n53 Vbias 2.23974f
C7957 CDAC8_0.switch_6.Z.n54 Vbias 2.23974f
C7958 CDAC8_0.switch_6.Z.t28 Vbias 5.88262f
C7959 CDAC8_0.switch_6.Z.n55 Vbias 1.36404f
C7960 CDAC8_0.switch_6.Z.n56 Vbias 1.12959f
C7961 CDAC8_0.switch_6.Z.n57 Vbias 1.12959f
C7962 CDAC8_0.switch_6.Z.t54 Vbias 5.88262f
C7963 CDAC8_0.switch_6.Z.n58 Vbias 1.36404f
C7964 CDAC8_0.switch_6.Z.n59 Vbias 1.24989f
C7965 CDAC8_0.switch_6.Z.n60 Vbias 1.24989f
C7966 CDAC8_0.switch_6.Z.t40 Vbias 5.88262f
C7967 CDAC8_0.switch_6.Z.n61 Vbias 1.36404f
C7968 CDAC8_0.switch_6.Z.n62 Vbias 1.08953f
C7969 CDAC8_0.switch_6.Z.t66 Vbias 5.88262f
C7970 CDAC8_0.switch_6.Z.n63 Vbias 1.36404f
C7971 CDAC8_0.switch_6.Z.n64 Vbias 1.12959f
C7972 CDAC8_0.switch_6.Z.n65 Vbias 1.12959f
C7973 CDAC8_0.switch_6.Z.t14 Vbias 5.88262f
C7974 CDAC8_0.switch_6.Z.n66 Vbias 1.36404f
C7975 CDAC8_0.switch_6.Z.n67 Vbias 0.6433f
C7976 CDAC8_0.switch_6.Z.t21 Vbias 5.88262f
C7977 CDAC8_0.switch_6.Z.n68 Vbias 1.36404f
C7978 CDAC8_0.switch_6.Z.n69 Vbias 1.12959f
C7979 CDAC8_0.switch_6.Z.n70 Vbias 1.12959f
C7980 CDAC8_0.switch_6.Z.t8 Vbias 5.88262f
C7981 CDAC8_0.switch_6.Z.n71 Vbias 1.36404f
C7982 CDAC8_0.switch_6.Z.n72 Vbias 1.12959f
C7983 CDAC8_0.switch_6.Z.n73 Vbias 1.12959f
C7984 CDAC8_0.switch_6.Z.t35 Vbias 5.88262f
C7985 CDAC8_0.switch_6.Z.n74 Vbias 1.36404f
C7986 CDAC8_0.switch_6.Z.n75 Vbias 1.12959f
C7987 CDAC8_0.switch_6.Z.n76 Vbias 1.12959f
C7988 CDAC8_0.switch_6.Z.t16 Vbias 5.88262f
C7989 CDAC8_0.switch_6.Z.n77 Vbias 1.36404f
C7990 CDAC8_0.switch_6.Z.n78 Vbias 1.12959f
C7991 CDAC8_0.switch_6.Z.n79 Vbias 1.12959f
C7992 CDAC8_0.switch_6.Z.t60 Vbias 5.88262f
C7993 CDAC8_0.switch_6.Z.n80 Vbias 1.36404f
C7994 CDAC8_0.switch_6.Z.t6 Vbias 5.88262f
C7995 CDAC8_0.switch_6.Z.n81 Vbias 1.36404f
C7996 CDAC8_0.switch_6.Z.n82 Vbias 1.12959f
C7997 CDAC8_0.switch_6.Z.n83 Vbias 1.12959f
C7998 CDAC8_0.switch_6.Z.t57 Vbias 5.88262f
C7999 CDAC8_0.switch_6.Z.n84 Vbias 1.36404f
C8000 CDAC8_0.switch_6.Z.n85 Vbias 1.12959f
C8001 CDAC8_0.switch_6.Z.t55 Vbias 5.88262f
C8002 CDAC8_0.switch_6.Z.n86 Vbias 1.36404f
C8003 CDAC8_0.switch_6.Z.t26 Vbias 5.88262f
C8004 CDAC8_0.switch_6.Z.n87 Vbias 1.36404f
C8005 CDAC8_0.switch_6.Z.t38 Vbias 5.88262f
C8006 CDAC8_0.switch_6.Z.n88 Vbias 1.36404f
C8007 CDAC8_0.switch_6.Z.t36 Vbias 6.12449f
C8008 CDAC8_0.switch_6.Z.t50 Vbias 6.12449f
C8009 CDAC8_0.switch_6.Z.n89 Vbias 2.41525f
C8010 CDAC8_0.switch_6.Z.n90 Vbias 2.41525f
C8011 CDAC8_0.switch_6.Z.t24 Vbias 5.88262f
C8012 CDAC8_0.switch_6.Z.n91 Vbias 1.36404f
C8013 CDAC8_0.switch_6.Z.n92 Vbias 1.12959f
C8014 CDAC8_0.switch_6.Z.n93 Vbias 1.12959f
C8015 CDAC8_0.switch_6.Z.t39 Vbias 5.88262f
C8016 CDAC8_0.switch_6.Z.n94 Vbias 1.36404f
C8017 CDAC8_0.switch_6.Z.n95 Vbias 1.12959f
C8018 CDAC8_0.switch_6.Z.n96 Vbias 1.12959f
C8019 CDAC8_0.switch_6.Z.t64 Vbias 5.88262f
C8020 CDAC8_0.switch_6.Z.n97 Vbias 1.36404f
C8021 CDAC8_0.switch_6.Z.n98 Vbias 1.12959f
C8022 CDAC8_0.switch_6.Z.n99 Vbias 1.12959f
C8023 CDAC8_0.switch_6.Z.t4 Vbias 5.88262f
C8024 CDAC8_0.switch_6.Z.n100 Vbias 1.24121f
C8025 CDAC8_0.switch_6.Z.n101 Vbias 2.49363f
C8026 CDAC8_0.switch_6.Z.n102 Vbias 2.49363f
C8027 CDAC8_0.switch_6.Z.n103 Vbias 0.7957f
C8028 CDAC8_0.switch_6.Z.n104 Vbias 1.12959f
C8029 CDAC8_0.switch_6.Z.t23 Vbias 5.88262f
C8030 CDAC8_0.switch_6.Z.n105 Vbias 1.36404f
C8031 CDAC8_0.switch_6.Z.n106 Vbias 1.12959f
C8032 CDAC8_0.switch_6.Z.n107 Vbias 1.12959f
C8033 CDAC8_0.switch_6.Z.t49 Vbias 5.88262f
C8034 CDAC8_0.switch_6.Z.n108 Vbias 1.36404f
C8035 CDAC8_0.switch_6.Z.n109 Vbias 1.12959f
C8036 CDAC8_0.switch_6.Z.n110 Vbias 1.12959f
C8037 CDAC8_0.switch_6.Z.t51 Vbias 5.88262f
C8038 CDAC8_0.switch_6.Z.n111 Vbias 1.36404f
C8039 CDAC8_0.switch_6.Z.n112 Vbias 1.12959f
C8040 CDAC8_0.switch_6.Z.n113 Vbias 1.12959f
C8041 CDAC8_0.switch_6.Z.t20 Vbias 5.88262f
C8042 CDAC8_0.switch_6.Z.n114 Vbias 1.36404f
C8043 CDAC8_0.switch_6.Z.n115 Vbias 1.12959f
C8044 CDAC8_0.switch_6.Z.n116 Vbias 1.12959f
C8045 CDAC8_0.switch_6.Z.t42 Vbias 5.88262f
C8046 CDAC8_0.switch_6.Z.n117 Vbias 1.36404f
C8047 CDAC8_0.switch_6.Z.n118 Vbias 1.12959f
C8048 CDAC8_0.switch_6.Z.n119 Vbias 1.12959f
C8049 CDAC8_0.switch_6.Z.t12 Vbias 5.88262f
C8050 CDAC8_0.switch_6.Z.n120 Vbias 1.36404f
C8051 CDAC8_0.switch_6.Z.n121 Vbias 0.6433f
C8052 CDAC8_0.switch_6.Z.n122 Vbias 1.45909f
C8053 CDAC8_0.switch_6.Z.n123 Vbias 1.93832f
C8054 CDAC8_0.switch_6.Z.n124 Vbias 0.01787f
C8055 CDAC8_0.switch_6.Z.t0 Vbias 0.03493f
C8056 CDAC8_0.switch_6.Z.n125 Vbias 0.14424f
C8057 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t1 Vbias 0.0608f
C8058 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n0 Vbias 0.13827f
C8059 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n1 Vbias 0.06674f
C8060 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t4 Vbias 0.24183f
C8061 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n2 Vbias 0.23689f
C8062 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n3 Vbias 0.04996f
C8063 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t3 Vbias 0.46511f
C8064 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n4 Vbias 0.13587f
C8065 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n5 Vbias 0.03381f
C8066 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n6 Vbias 0.04918f
C8067 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n7 Vbias 0.12602f
C8068 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n8 Vbias 0.12602f
C8069 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n9 Vbias 0.0655f
C8070 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t2 Vbias 0.06323f
C8071 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.t0 Vbias 0.07525f
C8072 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n10 Vbias 0.38033f
C8073 RingCounter_0.D_FlipFlop_15.Nand_Gate_1.Vout.n11 Vbias 0.1927f
C8074 CDAC8_0.switch_8.Z.t3 Vbias 0.03182f
C8075 CDAC8_0.switch_8.Z.t2 Vbias 0.03182f
C8076 CDAC8_0.switch_8.Z.n0 Vbias 0.11498f
C8077 CDAC8_0.switch_8.Z.n1 Vbias 0.24282f
C8078 CDAC8_0.switch_8.Z.n2 Vbias 0.03442f
C8079 CDAC8_0.switch_8.Z.t14 Vbias 5.70386f
C8080 CDAC8_0.switch_8.Z.n3 Vbias 1.9642f
C8081 CDAC8_0.switch_8.Z.t6 Vbias 5.70386f
C8082 CDAC8_0.switch_8.Z.t4 Vbias 5.9531f
C8083 CDAC8_0.switch_8.Z.t17 Vbias 5.62231f
C8084 CDAC8_0.switch_8.Z.n4 Vbias 3.16681f
C8085 CDAC8_0.switch_8.Z.t19 Vbias 5.62231f
C8086 CDAC8_0.switch_8.Z.n5 Vbias 1.91851f
C8087 CDAC8_0.switch_8.Z.t15 Vbias 5.62231f
C8088 CDAC8_0.switch_8.Z.n6 Vbias 1.91851f
C8089 CDAC8_0.switch_8.Z.t9 Vbias 5.62231f
C8090 CDAC8_0.switch_8.Z.n7 Vbias 1.6228f
C8091 CDAC8_0.switch_8.Z.t13 Vbias 5.62231f
C8092 CDAC8_0.switch_8.Z.n8 Vbias 1.74019f
C8093 CDAC8_0.switch_8.Z.t18 Vbias 5.62231f
C8094 CDAC8_0.switch_8.Z.n9 Vbias 1.59939f
C8095 CDAC8_0.switch_8.Z.t12 Vbias 5.9531f
C8096 CDAC8_0.switch_8.Z.t8 Vbias 5.62231f
C8097 CDAC8_0.switch_8.Z.n10 Vbias 3.16681f
C8098 CDAC8_0.switch_8.Z.t10 Vbias 5.62231f
C8099 CDAC8_0.switch_8.Z.n11 Vbias 1.91851f
C8100 CDAC8_0.switch_8.Z.t7 Vbias 5.62231f
C8101 CDAC8_0.switch_8.Z.n12 Vbias 1.91851f
C8102 CDAC8_0.switch_8.Z.t16 Vbias 5.62231f
C8103 CDAC8_0.switch_8.Z.n13 Vbias 1.6228f
C8104 CDAC8_0.switch_8.Z.n14 Vbias 1.12092f
C8105 CDAC8_0.switch_8.Z.n15 Vbias 1.12092f
C8106 CDAC8_0.switch_8.Z.t11 Vbias 5.62231f
C8107 CDAC8_0.switch_8.Z.n16 Vbias 1.59939f
C8108 CDAC8_0.switch_8.Z.t5 Vbias 5.62231f
C8109 CDAC8_0.switch_8.Z.n17 Vbias 1.74019f
C8110 CDAC8_0.switch_8.Z.n18 Vbias 1.92246f
C8111 CDAC8_0.switch_8.Z.n19 Vbias 0.48531f
C8112 CDAC8_0.switch_8.Z.n20 Vbias 0.01245f
C8113 CDAC8_0.switch_8.Z.n21 Vbias 0.0507f
C8114 CDAC8_0.switch_8.Z.t0 Vbias 0.03342f
C8115 CDAC8_0.switch_8.Z.n22 Vbias 0.09316f
C8116 CDAC8_0.switch_8.Z.t1 Vbias 0.0334f
C8117 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t2 Vbias 0.07037f
C8118 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n0 Vbias 0.16004f
C8119 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n1 Vbias 0.07725f
C8120 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t4 Vbias 0.2799f
C8121 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n2 Vbias 0.27418f
C8122 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n3 Vbias 0.05783f
C8123 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t5 Vbias 0.53832f
C8124 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n4 Vbias 0.15726f
C8125 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n5 Vbias 0.03913f
C8126 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n6 Vbias 0.05692f
C8127 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n7 Vbias 0.14585f
C8128 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n8 Vbias 0.14585f
C8129 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n9 Vbias 0.07581f
C8130 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t3 Vbias 0.07318f
C8131 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t0 Vbias 0.07454f
C8132 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.t1 Vbias 0.07302f
C8133 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n10 Vbias 0.41525f
C8134 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n11 Vbias 0.23391f
C8135 RingCounter_0.D_FlipFlop_11.3-input-nand_1.Vout.n12 Vbias 0.22303f
C8136 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t6 Vbias 0.45666f
C8137 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n0 Vbias 0.47347f
C8138 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n1 Vbias 0.05122f
C8139 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n2 Vbias 0.06839f
C8140 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t4 Vbias 0.22727f
C8141 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t1 Vbias 0.06194f
C8142 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n3 Vbias 0.39067f
C8143 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t3 Vbias 0.06323f
C8144 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t2 Vbias 0.06194f
C8145 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n4 Vbias 0.35224f
C8146 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n5 Vbias 0.11629f
C8147 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n6 Vbias 0.16533f
C8148 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n7 Vbias 0.06431f
C8149 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t7 Vbias 0.23742f
C8150 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t5 Vbias 0.45664f
C8151 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n8 Vbias 0.1334f
C8152 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n9 Vbias 0.05705f
C8153 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n10 Vbias 0.10533f
C8154 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n11 Vbias 0.18236f
C8155 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n12 Vbias 0.13574f
C8156 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n13 Vbias 0.12257f
C8157 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.n14 Vbias 0.0577f
C8158 RingCounter_0.D_FlipFlop_3.3-input-nand_2.C.t0 Vbias 0.05958f
C8159 D_FlipFlop_6.3-input-nand_2.C.t6 Vbias 0.3425f
C8160 D_FlipFlop_6.3-input-nand_2.C.n0 Vbias 0.3551f
C8161 D_FlipFlop_6.3-input-nand_2.C.n1 Vbias 0.03842f
C8162 D_FlipFlop_6.3-input-nand_2.C.n2 Vbias 0.05129f
C8163 D_FlipFlop_6.3-input-nand_2.C.t5 Vbias 0.17045f
C8164 D_FlipFlop_6.3-input-nand_2.C.t3 Vbias 0.04645f
C8165 D_FlipFlop_6.3-input-nand_2.C.n3 Vbias 0.293f
C8166 D_FlipFlop_6.3-input-nand_2.C.t1 Vbias 0.04742f
C8167 D_FlipFlop_6.3-input-nand_2.C.t2 Vbias 0.04645f
C8168 D_FlipFlop_6.3-input-nand_2.C.n4 Vbias 0.26418f
C8169 D_FlipFlop_6.3-input-nand_2.C.n5 Vbias 0.08722f
C8170 D_FlipFlop_6.3-input-nand_2.C.n6 Vbias 0.124f
C8171 D_FlipFlop_6.3-input-nand_2.C.n7 Vbias 0.04823f
C8172 D_FlipFlop_6.3-input-nand_2.C.t7 Vbias 0.17806f
C8173 D_FlipFlop_6.3-input-nand_2.C.t4 Vbias 0.34248f
C8174 D_FlipFlop_6.3-input-nand_2.C.n8 Vbias 0.10005f
C8175 D_FlipFlop_6.3-input-nand_2.C.n9 Vbias 0.04279f
C8176 D_FlipFlop_6.3-input-nand_2.C.n10 Vbias 0.079f
C8177 D_FlipFlop_6.3-input-nand_2.C.n11 Vbias 0.13677f
C8178 D_FlipFlop_6.3-input-nand_2.C.n12 Vbias 0.10181f
C8179 D_FlipFlop_6.3-input-nand_2.C.n13 Vbias 0.09193f
C8180 D_FlipFlop_6.3-input-nand_2.C.t0 Vbias 0.04477f
C8181 D_FlipFlop_6.3-input-nand_2.C.n14 Vbias 0.11971f
C8182 VDD.t944 Vbias 0.017f
C8183 VDD.t835 Vbias 0.017f
C8184 VDD.n0 Vbias 0.05322f
C8185 VDD.n1 Vbias 0.01999f
C8186 VDD.n2 Vbias 0.03694f
C8187 VDD.n3 Vbias 0.0216f
C8188 VDD.n4 Vbias 0.03694f
C8189 VDD.n5 Vbias 0.26017f
C8190 VDD.t834 Vbias 0.24595f
C8191 VDD.t1092 Vbias 0.22551f
C8192 VDD.n7 Vbias 0.03694f
C8193 VDD.n8 Vbias 0.03694f
C8194 VDD.n9 Vbias 0.06648f
C8195 VDD.t539 Vbias 0.24595f
C8196 VDD.n10 Vbias 0.03694f
C8197 VDD.n11 Vbias 0.03694f
C8198 VDD.t1093 Vbias 0.0169f
C8199 VDD.t540 Vbias 0.0169f
C8200 VDD.n12 Vbias 0.07902f
C8201 VDD.n13 Vbias 0.01699f
C8202 VDD.n14 Vbias 0.0228f
C8203 VDD.t911 Vbias 0.0169f
C8204 VDD.t202 Vbias 0.0169f
C8205 VDD.n15 Vbias 0.07902f
C8206 VDD.n16 Vbias 0.0228f
C8207 VDD.n17 Vbias 0.01999f
C8208 VDD.n18 Vbias 0.03694f
C8209 VDD.n19 Vbias 0.0216f
C8210 VDD.n20 Vbias 0.03694f
C8211 VDD.n21 Vbias 0.26017f
C8212 VDD.t910 Vbias 0.24595f
C8213 VDD.t201 Vbias 0.24595f
C8214 VDD.n23 Vbias 0.03694f
C8215 VDD.n24 Vbias 0.03694f
C8216 VDD.t638 Vbias 0.017f
C8217 VDD.n25 Vbias 0.05322f
C8218 VDD.n26 Vbias 0.01999f
C8219 VDD.n27 Vbias 0.03694f
C8220 VDD.n28 Vbias 0.0216f
C8221 VDD.n29 Vbias 0.03694f
C8222 VDD.n30 Vbias 0.26017f
C8223 VDD.t637 Vbias 0.24595f
C8224 VDD.t1065 Vbias 0.22551f
C8225 VDD.n32 Vbias 0.03694f
C8226 VDD.n33 Vbias 0.03694f
C8227 VDD.n34 Vbias 0.06648f
C8228 VDD.t821 Vbias 0.24595f
C8229 VDD.n35 Vbias 0.03694f
C8230 VDD.n36 Vbias 0.03694f
C8231 VDD.t1066 Vbias 0.0169f
C8232 VDD.t822 Vbias 0.0169f
C8233 VDD.n37 Vbias 0.07902f
C8234 VDD.n38 Vbias 0.01699f
C8235 VDD.n39 Vbias 0.0228f
C8236 VDD.t569 Vbias 0.0169f
C8237 VDD.t154 Vbias 0.0169f
C8238 VDD.n40 Vbias 0.07902f
C8239 VDD.n41 Vbias 0.0228f
C8240 VDD.n42 Vbias 0.01999f
C8241 VDD.n43 Vbias 0.03694f
C8242 VDD.n44 Vbias 0.0216f
C8243 VDD.n45 Vbias 0.03694f
C8244 VDD.n46 Vbias 0.26017f
C8245 VDD.t568 Vbias 0.24595f
C8246 VDD.t153 Vbias 0.24595f
C8247 VDD.n48 Vbias 0.03694f
C8248 VDD.n49 Vbias 0.03694f
C8249 VDD.t327 Vbias 0.017f
C8250 VDD.n50 Vbias 0.05322f
C8251 VDD.n51 Vbias 0.01999f
C8252 VDD.n52 Vbias 0.03694f
C8253 VDD.n53 Vbias 0.0216f
C8254 VDD.n54 Vbias 0.03694f
C8255 VDD.n55 Vbias 0.26017f
C8256 VDD.t326 Vbias 0.24595f
C8257 VDD.t1026 Vbias 0.22551f
C8258 VDD.n57 Vbias 0.03694f
C8259 VDD.n58 Vbias 0.03694f
C8260 VDD.n59 Vbias 0.06648f
C8261 VDD.t7 Vbias 0.24595f
C8262 VDD.n60 Vbias 0.03694f
C8263 VDD.n61 Vbias 0.03694f
C8264 VDD.t1027 Vbias 0.0169f
C8265 VDD.t8 Vbias 0.0169f
C8266 VDD.n62 Vbias 0.07902f
C8267 VDD.n63 Vbias 0.01699f
C8268 VDD.n64 Vbias 0.0228f
C8269 VDD.t994 Vbias 0.0169f
C8270 VDD.t828 Vbias 0.0169f
C8271 VDD.n65 Vbias 0.07902f
C8272 VDD.n66 Vbias 0.0228f
C8273 VDD.n67 Vbias 0.01999f
C8274 VDD.n68 Vbias 0.03694f
C8275 VDD.n69 Vbias 0.0216f
C8276 VDD.n70 Vbias 0.03694f
C8277 VDD.n71 Vbias 0.26017f
C8278 VDD.t993 Vbias 0.24595f
C8279 VDD.t827 Vbias 0.24595f
C8280 VDD.n73 Vbias 0.03694f
C8281 VDD.n74 Vbias 0.03694f
C8282 VDD.t860 Vbias 0.017f
C8283 VDD.n75 Vbias 0.05322f
C8284 VDD.n76 Vbias 0.01999f
C8285 VDD.n77 Vbias 0.03694f
C8286 VDD.n78 Vbias 0.0216f
C8287 VDD.n79 Vbias 0.03694f
C8288 VDD.n80 Vbias 0.26017f
C8289 VDD.t859 Vbias 0.24595f
C8290 VDD.t1071 Vbias 0.22551f
C8291 VDD.n82 Vbias 0.03694f
C8292 VDD.n83 Vbias 0.03694f
C8293 VDD.n84 Vbias 0.06648f
C8294 VDD.t250 Vbias 0.24595f
C8295 VDD.n85 Vbias 0.03694f
C8296 VDD.n86 Vbias 0.03694f
C8297 VDD.t1072 Vbias 0.0169f
C8298 VDD.t251 Vbias 0.0169f
C8299 VDD.n87 Vbias 0.07902f
C8300 VDD.n88 Vbias 0.01699f
C8301 VDD.n89 Vbias 0.0228f
C8302 VDD.t380 Vbias 0.0169f
C8303 VDD.t198 Vbias 0.0169f
C8304 VDD.n90 Vbias 0.07902f
C8305 VDD.n91 Vbias 0.0228f
C8306 VDD.n92 Vbias 0.01999f
C8307 VDD.n93 Vbias 0.03694f
C8308 VDD.n94 Vbias 0.0216f
C8309 VDD.n95 Vbias 0.03694f
C8310 VDD.n96 Vbias 0.26017f
C8311 VDD.t379 Vbias 0.24595f
C8312 VDD.t197 Vbias 0.24595f
C8313 VDD.n98 Vbias 0.03694f
C8314 VDD.n99 Vbias 0.03694f
C8315 VDD.n100 Vbias 0.01699f
C8316 VDD.n101 Vbias 0.06648f
C8317 VDD.n103 Vbias 0.26017f
C8318 VDD.n104 Vbias 0.01999f
C8319 VDD.n105 Vbias 0.0216f
C8320 VDD.n106 Vbias 0.01999f
C8321 VDD.n107 Vbias 0.03639f
C8322 VDD.n108 Vbias 0.18185f
C8323 VDD.n109 Vbias 0.18185f
C8324 VDD.n110 Vbias 0.03639f
C8325 VDD.n111 Vbias 0.01999f
C8326 VDD.n112 Vbias 0.06648f
C8327 VDD.n113 Vbias 0.24997f
C8328 VDD.n114 Vbias 0.01699f
C8329 VDD.n115 Vbias 0.06648f
C8330 VDD.n117 Vbias 0.26017f
C8331 VDD.n118 Vbias 0.01999f
C8332 VDD.n119 Vbias 0.0216f
C8333 VDD.n120 Vbias 0.01999f
C8334 VDD.n121 Vbias 0.03639f
C8335 VDD.n122 Vbias 0.18185f
C8336 VDD.n123 Vbias 0.18185f
C8337 VDD.n124 Vbias 0.03639f
C8338 VDD.n125 Vbias 0.01999f
C8339 VDD.n126 Vbias 0.0216f
C8340 VDD.n127 Vbias 0.01999f
C8341 VDD.n128 Vbias 0.03639f
C8342 VDD.n129 Vbias 0.24422f
C8343 VDD.n130 Vbias 0.24422f
C8344 VDD.n131 Vbias 0.03639f
C8345 VDD.n132 Vbias 0.01999f
C8346 VDD.n133 Vbias 0.06648f
C8347 VDD.n134 Vbias 0.24606f
C8348 VDD.n135 Vbias 0.01699f
C8349 VDD.n136 Vbias 0.06648f
C8350 VDD.n138 Vbias 0.26017f
C8351 VDD.n139 Vbias 0.01999f
C8352 VDD.n140 Vbias 0.0216f
C8353 VDD.n141 Vbias 0.01999f
C8354 VDD.n142 Vbias 0.03639f
C8355 VDD.n143 Vbias 0.18185f
C8356 VDD.n144 Vbias 0.18185f
C8357 VDD.n145 Vbias 0.03639f
C8358 VDD.n146 Vbias 0.01999f
C8359 VDD.n147 Vbias 0.06648f
C8360 VDD.n148 Vbias 0.24997f
C8361 VDD.n149 Vbias 0.01699f
C8362 VDD.n150 Vbias 0.06648f
C8363 VDD.n152 Vbias 0.26017f
C8364 VDD.n153 Vbias 0.01999f
C8365 VDD.n154 Vbias 0.0216f
C8366 VDD.n155 Vbias 0.01999f
C8367 VDD.n156 Vbias 0.03639f
C8368 VDD.n157 Vbias 0.18185f
C8369 VDD.n158 Vbias 0.18185f
C8370 VDD.n159 Vbias 0.03639f
C8371 VDD.n160 Vbias 0.01999f
C8372 VDD.n161 Vbias 0.0216f
C8373 VDD.n162 Vbias 0.01999f
C8374 VDD.n163 Vbias 0.03639f
C8375 VDD.n164 Vbias 0.24422f
C8376 VDD.n165 Vbias 0.24422f
C8377 VDD.n166 Vbias 0.03639f
C8378 VDD.n167 Vbias 0.01999f
C8379 VDD.n168 Vbias 0.06648f
C8380 VDD.n169 Vbias 0.24606f
C8381 VDD.n170 Vbias 0.01699f
C8382 VDD.n171 Vbias 0.06648f
C8383 VDD.n173 Vbias 0.26017f
C8384 VDD.n174 Vbias 0.01999f
C8385 VDD.n175 Vbias 0.0216f
C8386 VDD.n176 Vbias 0.01999f
C8387 VDD.n177 Vbias 0.03639f
C8388 VDD.n178 Vbias 0.18185f
C8389 VDD.n179 Vbias 0.18185f
C8390 VDD.n180 Vbias 0.03639f
C8391 VDD.n181 Vbias 0.01999f
C8392 VDD.n182 Vbias 0.06648f
C8393 VDD.n183 Vbias 0.24997f
C8394 VDD.n184 Vbias 0.01699f
C8395 VDD.n185 Vbias 0.06648f
C8396 VDD.n187 Vbias 0.26017f
C8397 VDD.n188 Vbias 0.01999f
C8398 VDD.n189 Vbias 0.0216f
C8399 VDD.n190 Vbias 0.01999f
C8400 VDD.n191 Vbias 0.03639f
C8401 VDD.n192 Vbias 0.18185f
C8402 VDD.n193 Vbias 0.18185f
C8403 VDD.n194 Vbias 0.03639f
C8404 VDD.n195 Vbias 0.01999f
C8405 VDD.n196 Vbias 0.0216f
C8406 VDD.n197 Vbias 0.01999f
C8407 VDD.n198 Vbias 0.03639f
C8408 VDD.n199 Vbias 0.24422f
C8409 VDD.n200 Vbias 0.24422f
C8410 VDD.n201 Vbias 0.03639f
C8411 VDD.n202 Vbias 0.01999f
C8412 VDD.n203 Vbias 0.06648f
C8413 VDD.n204 Vbias 0.24606f
C8414 VDD.n205 Vbias 0.01699f
C8415 VDD.n206 Vbias 0.06648f
C8416 VDD.n208 Vbias 0.26017f
C8417 VDD.n209 Vbias 0.01999f
C8418 VDD.n210 Vbias 0.0216f
C8419 VDD.n211 Vbias 0.01999f
C8420 VDD.n212 Vbias 0.03639f
C8421 VDD.n213 Vbias 0.18185f
C8422 VDD.n214 Vbias 0.18185f
C8423 VDD.n215 Vbias 0.03639f
C8424 VDD.n216 Vbias 0.01999f
C8425 VDD.n217 Vbias 0.06648f
C8426 VDD.n218 Vbias 0.24997f
C8427 VDD.n219 Vbias 0.01699f
C8428 VDD.n220 Vbias 0.06648f
C8429 VDD.n222 Vbias 0.26017f
C8430 VDD.n223 Vbias 0.01999f
C8431 VDD.n224 Vbias 0.0216f
C8432 VDD.n225 Vbias 0.01999f
C8433 VDD.n226 Vbias 0.03639f
C8434 VDD.n227 Vbias 0.18185f
C8435 VDD.n228 Vbias 0.18185f
C8436 VDD.n229 Vbias 0.03639f
C8437 VDD.n230 Vbias 0.01999f
C8438 VDD.n231 Vbias 0.0216f
C8439 VDD.n232 Vbias 0.01999f
C8440 VDD.n233 Vbias 0.03639f
C8441 VDD.n234 Vbias 0.24422f
C8442 VDD.n235 Vbias 0.24422f
C8443 VDD.n236 Vbias 0.03639f
C8444 VDD.n237 Vbias 0.01999f
C8445 VDD.n238 Vbias 0.06648f
C8446 VDD.n239 Vbias 0.01156f
C8447 VDD.n240 Vbias 0.27159f
C8448 VDD.t463 Vbias 1.48288f
C8449 VDD.t700 Vbias 1.17927f
C8450 VDD.t702 Vbias 1.17927f
C8451 VDD.n241 Vbias 0.66348f
C8452 VDD.t703 Vbias 0.18415f
C8453 VDD.n242 Vbias 2.42007f
C8454 VDD.n243 Vbias 1.39105f
C8455 VDD.n244 Vbias 0.82392f
C8456 VDD.n245 Vbias 0.1918f
C8457 VDD.n246 Vbias 0.16533f
C8458 VDD.n247 Vbias 0.19801f
C8459 VDD.n248 Vbias 0.17982f
C8460 VDD.n249 Vbias 2.825f
C8461 VDD.n250 Vbias 3.03142f
C8462 VDD.n251 Vbias 0.32644f
C8463 VDD.n252 Vbias 0.17982f
C8464 VDD.n253 Vbias 0.19801f
C8465 VDD.n254 Vbias 2.825f
C8466 VDD.n255 Vbias 0.18156f
C8467 VDD.t699 Vbias 3.16035f
C8468 VDD.n257 Vbias 0.18156f
C8469 VDD.n258 Vbias 0.10623f
C8470 VDD.n259 Vbias 0.10563f
C8471 VDD.n260 Vbias 0.10623f
C8472 VDD.n261 Vbias 0.18156f
C8473 VDD.t701 Vbias 3.16035f
C8474 VDD.n263 Vbias 0.18156f
C8475 VDD.n264 Vbias 0.16533f
C8476 VDD.n265 Vbias 0.14111f
C8477 VDD.n266 Vbias 0.08068f
C8478 VDD.n267 Vbias 0.37138f
C8479 VDD.n268 Vbias 0.23495f
C8480 VDD.n269 Vbias 0.40965f
C8481 VDD.n270 Vbias 0.23973f
C8482 VDD.t462 Vbias 3.90944f
C8483 VDD.n272 Vbias 3.357f
C8484 VDD.n273 Vbias 0.40965f
C8485 VDD.n275 Vbias 3.357f
C8486 VDD.n276 Vbias 0.23495f
C8487 VDD.n277 Vbias 0.32253f
C8488 VDD.n278 Vbias 0.01191f
C8489 VDD.n279 Vbias 0.01007f
C8490 VDD.n280 Vbias 0.03825f
C8491 VDD.n281 Vbias 0.44107f
C8492 VDD.t979 Vbias 0.017f
C8493 VDD.n282 Vbias 0.01999f
C8494 VDD.n283 Vbias 0.03694f
C8495 VDD.n284 Vbias 0.0216f
C8496 VDD.n285 Vbias 0.03694f
C8497 VDD.n286 Vbias 0.45845f
C8498 VDD.t978 Vbias 0.54191f
C8499 VDD.n288 Vbias 0.03639f
C8500 VDD.t933 Vbias 0.46278f
C8501 VDD.n289 Vbias 0.03694f
C8502 VDD.n290 Vbias 0.03694f
C8503 VDD.n291 Vbias 0.0216f
C8504 VDD.n292 Vbias 0.01836f
C8505 VDD.t984 Vbias 0.017f
C8506 VDD.t934 Vbias 0.017f
C8507 VDD.n293 Vbias 0.09713f
C8508 VDD.n294 Vbias 0.01914f
C8509 VDD.n295 Vbias 0.03902f
C8510 VDD.n296 Vbias 0.03694f
C8511 VDD.n297 Vbias 0.0216f
C8512 VDD.n298 Vbias 0.01836f
C8513 VDD.n299 Vbias 0.03639f
C8514 VDD.t335 Vbias 0.46278f
C8515 VDD.n300 Vbias 0.03694f
C8516 VDD.n301 Vbias 0.03694f
C8517 VDD.n302 Vbias 0.0216f
C8518 VDD.n303 Vbias 0.01836f
C8519 VDD.n304 Vbias 0.02305f
C8520 VDD.n305 Vbias 0.03902f
C8521 VDD.n306 Vbias 0.03694f
C8522 VDD.n307 Vbias 0.0216f
C8523 VDD.n308 Vbias 0.01836f
C8524 VDD.n309 Vbias 0.03639f
C8525 VDD.t411 Vbias 0.46278f
C8526 VDD.n310 Vbias 0.03694f
C8527 VDD.n311 Vbias 0.03694f
C8528 VDD.n312 Vbias 0.0216f
C8529 VDD.n313 Vbias 0.01836f
C8530 VDD.t546 Vbias 0.0169f
C8531 VDD.t413 Vbias 0.0169f
C8532 VDD.n314 Vbias 0.07902f
C8533 VDD.t336 Vbias 0.0169f
C8534 VDD.t412 Vbias 0.0169f
C8535 VDD.n315 Vbias 0.07902f
C8536 VDD.n316 Vbias 0.03023f
C8537 VDD.n317 Vbias 0.01699f
C8538 VDD.n318 Vbias 0.03902f
C8539 VDD.n319 Vbias 0.03694f
C8540 VDD.n320 Vbias 0.0216f
C8541 VDD.n321 Vbias 0.01836f
C8542 VDD.n322 Vbias 0.03639f
C8543 VDD.t394 Vbias 0.46278f
C8544 VDD.n323 Vbias 0.03694f
C8545 VDD.n324 Vbias 0.03694f
C8546 VDD.n325 Vbias 0.0216f
C8547 VDD.n326 Vbias 0.01836f
C8548 VDD.t932 Vbias 0.017f
C8549 VDD.t395 Vbias 0.017f
C8550 VDD.n327 Vbias 0.09713f
C8551 VDD.n328 Vbias 0.01914f
C8552 VDD.n329 Vbias 0.03902f
C8553 VDD.n330 Vbias 0.03694f
C8554 VDD.n331 Vbias 0.0216f
C8555 VDD.n332 Vbias 0.01836f
C8556 VDD.n333 Vbias 0.03639f
C8557 VDD.t596 Vbias 0.46278f
C8558 VDD.n334 Vbias 0.03694f
C8559 VDD.n335 Vbias 0.03694f
C8560 VDD.n336 Vbias 0.0216f
C8561 VDD.n337 Vbias 0.01836f
C8562 VDD.n338 Vbias 0.02305f
C8563 VDD.n339 Vbias 0.03902f
C8564 VDD.n340 Vbias 0.03694f
C8565 VDD.n341 Vbias 0.0216f
C8566 VDD.n342 Vbias 0.01836f
C8567 VDD.n343 Vbias 0.03639f
C8568 VDD.t174 Vbias 0.46278f
C8569 VDD.n344 Vbias 0.03694f
C8570 VDD.n345 Vbias 0.03694f
C8571 VDD.n346 Vbias 0.0216f
C8572 VDD.n347 Vbias 0.01836f
C8573 VDD.t606 Vbias 0.0169f
C8574 VDD.t175 Vbias 0.0169f
C8575 VDD.n348 Vbias 0.07902f
C8576 VDD.t597 Vbias 0.0169f
C8577 VDD.t383 Vbias 0.0169f
C8578 VDD.n349 Vbias 0.07902f
C8579 VDD.n350 Vbias 0.03023f
C8580 VDD.n351 Vbias 0.01699f
C8581 VDD.n352 Vbias 0.03902f
C8582 VDD.n353 Vbias 0.03694f
C8583 VDD.n354 Vbias 0.0216f
C8584 VDD.n355 Vbias 0.01836f
C8585 VDD.t414 Vbias 0.46278f
C8586 VDD.n356 Vbias 0.03694f
C8587 VDD.n357 Vbias 0.03694f
C8588 VDD.n358 Vbias 0.06648f
C8589 VDD.n359 Vbias 0.03639f
C8590 VDD.t478 Vbias 0.46278f
C8591 VDD.n360 Vbias 0.03694f
C8592 VDD.n361 Vbias 0.03694f
C8593 VDD.n362 Vbias 0.0216f
C8594 VDD.n363 Vbias 0.01836f
C8595 VDD.t415 Vbias 0.017f
C8596 VDD.n364 Vbias 0.05322f
C8597 VDD.n365 Vbias 0.01309f
C8598 VDD.n366 Vbias 0.01699f
C8599 VDD.n367 Vbias 0.03902f
C8600 VDD.n368 Vbias 0.03694f
C8601 VDD.n369 Vbias 0.0216f
C8602 VDD.n370 Vbias 0.01836f
C8603 VDD.n371 Vbias 0.03639f
C8604 VDD.t628 Vbias 0.46278f
C8605 VDD.n372 Vbias 0.03694f
C8606 VDD.n373 Vbias 0.03694f
C8607 VDD.n374 Vbias 0.0216f
C8608 VDD.n375 Vbias 0.01836f
C8609 VDD.t674 Vbias 0.0169f
C8610 VDD.t630 Vbias 0.0169f
C8611 VDD.n376 Vbias 0.07902f
C8612 VDD.t479 Vbias 0.0169f
C8613 VDD.t629 Vbias 0.0169f
C8614 VDD.n377 Vbias 0.07902f
C8615 VDD.n378 Vbias 0.03023f
C8616 VDD.n379 Vbias 0.01699f
C8617 VDD.n380 Vbias 0.03902f
C8618 VDD.n381 Vbias 0.03694f
C8619 VDD.n382 Vbias 0.0216f
C8620 VDD.n383 Vbias 0.01836f
C8621 VDD.n384 Vbias 0.03639f
C8622 VDD.t466 Vbias 0.46278f
C8623 VDD.n385 Vbias 0.03694f
C8624 VDD.n386 Vbias 0.03694f
C8625 VDD.n387 Vbias 0.0216f
C8626 VDD.n388 Vbias 0.01836f
C8627 VDD.t936 Vbias 0.017f
C8628 VDD.t467 Vbias 0.017f
C8629 VDD.n389 Vbias 0.09713f
C8630 VDD.n390 Vbias 0.01914f
C8631 VDD.n391 Vbias 0.03902f
C8632 VDD.n392 Vbias 0.03694f
C8633 VDD.n393 Vbias 0.0216f
C8634 VDD.n394 Vbias 0.01836f
C8635 VDD.n395 Vbias 0.03639f
C8636 VDD.t192 Vbias 0.46278f
C8637 VDD.n396 Vbias 0.03694f
C8638 VDD.n397 Vbias 0.03694f
C8639 VDD.n398 Vbias 0.0216f
C8640 VDD.n399 Vbias 0.01836f
C8641 VDD.n400 Vbias 0.02305f
C8642 VDD.n401 Vbias 0.03902f
C8643 VDD.n402 Vbias 0.03694f
C8644 VDD.n403 Vbias 0.0216f
C8645 VDD.n404 Vbias 0.01836f
C8646 VDD.n405 Vbias 0.03639f
C8647 VDD.t214 Vbias 0.46278f
C8648 VDD.n406 Vbias 0.03694f
C8649 VDD.n407 Vbias 0.03694f
C8650 VDD.n408 Vbias 0.0216f
C8651 VDD.n409 Vbias 0.01836f
C8652 VDD.t193 Vbias 0.0169f
C8653 VDD.t218 Vbias 0.0169f
C8654 VDD.n410 Vbias 0.07902f
C8655 VDD.t964 Vbias 0.0169f
C8656 VDD.t215 Vbias 0.0169f
C8657 VDD.n411 Vbias 0.07902f
C8658 VDD.n412 Vbias 0.03023f
C8659 VDD.n413 Vbias 0.01699f
C8660 VDD.n414 Vbias 0.03902f
C8661 VDD.n415 Vbias 0.03694f
C8662 VDD.n416 Vbias 0.0216f
C8663 VDD.n417 Vbias 0.01836f
C8664 VDD.n418 Vbias 0.01836f
C8665 VDD.n419 Vbias 0.03639f
C8666 VDD.n420 Vbias 0.50118f
C8667 VDD.n421 Vbias 0.03639f
C8668 VDD.n422 Vbias 0.03694f
C8669 VDD.n423 Vbias 0.04583f
C8670 VDD.n424 Vbias 0.03902f
C8671 VDD.n425 Vbias 0.01836f
C8672 VDD.n426 Vbias 0.03639f
C8673 VDD.n427 Vbias 0.37318f
C8674 VDD.n428 Vbias 0.01836f
C8675 VDD.n429 Vbias 0.03639f
C8676 VDD.n430 Vbias 0.37318f
C8677 VDD.n431 Vbias 0.03639f
C8678 VDD.n432 Vbias 0.03694f
C8679 VDD.n433 Vbias 0.04583f
C8680 VDD.n434 Vbias 0.03902f
C8681 VDD.n435 Vbias 0.01836f
C8682 VDD.n436 Vbias 0.03639f
C8683 VDD.n437 Vbias 0.37318f
C8684 VDD.n438 Vbias 0.01836f
C8685 VDD.n439 Vbias 0.03639f
C8686 VDD.n440 Vbias 0.37318f
C8687 VDD.n441 Vbias 0.03639f
C8688 VDD.n442 Vbias 0.03694f
C8689 VDD.n443 Vbias 0.04583f
C8690 VDD.n444 Vbias 0.03902f
C8691 VDD.n445 Vbias 0.01836f
C8692 VDD.n446 Vbias 0.03639f
C8693 VDD.n447 Vbias 0.50118f
C8694 VDD.n448 Vbias 0.01836f
C8695 VDD.n449 Vbias 0.03639f
C8696 VDD.n450 Vbias 0.50118f
C8697 VDD.n451 Vbias 0.03639f
C8698 VDD.n452 Vbias 0.03694f
C8699 VDD.n453 Vbias 0.04583f
C8700 VDD.n454 Vbias 0.03902f
C8701 VDD.n455 Vbias 0.01836f
C8702 VDD.n456 Vbias 0.03639f
C8703 VDD.n457 Vbias 0.37318f
C8704 VDD.n458 Vbias 0.01836f
C8705 VDD.n459 Vbias 0.03639f
C8706 VDD.n460 Vbias 0.37318f
C8707 VDD.n461 Vbias 0.03639f
C8708 VDD.n462 Vbias 0.03694f
C8709 VDD.n463 Vbias 0.04583f
C8710 VDD.n464 Vbias 0.03902f
C8711 VDD.n465 Vbias 0.01836f
C8712 VDD.n466 Vbias 0.03639f
C8713 VDD.n467 Vbias 0.50118f
C8714 VDD.n468 Vbias 0.50118f
C8715 VDD.n469 Vbias 0.03639f
C8716 VDD.n470 Vbias 0.01999f
C8717 VDD.n471 Vbias 0.0216f
C8718 VDD.n472 Vbias 0.01999f
C8719 VDD.n473 Vbias 0.03639f
C8720 VDD.n474 Vbias 0.50118f
C8721 VDD.n475 Vbias 0.01836f
C8722 VDD.n476 Vbias 0.03639f
C8723 VDD.n477 Vbias 0.50118f
C8724 VDD.n478 Vbias 0.03639f
C8725 VDD.n479 Vbias 0.03694f
C8726 VDD.n480 Vbias 0.04583f
C8727 VDD.n481 Vbias 0.03902f
C8728 VDD.n482 Vbias 0.01836f
C8729 VDD.n483 Vbias 0.03639f
C8730 VDD.n484 Vbias 0.37318f
C8731 VDD.n485 Vbias 0.01836f
C8732 VDD.n486 Vbias 0.03639f
C8733 VDD.n487 Vbias 0.37318f
C8734 VDD.n488 Vbias 0.03639f
C8735 VDD.n489 Vbias 0.03694f
C8736 VDD.n490 Vbias 0.04583f
C8737 VDD.n491 Vbias 0.03902f
C8738 VDD.n492 Vbias 0.01836f
C8739 VDD.n493 Vbias 0.03639f
C8740 VDD.n494 Vbias 0.37318f
C8741 VDD.n495 Vbias 0.01836f
C8742 VDD.n496 Vbias 0.03639f
C8743 VDD.n497 Vbias 0.37318f
C8744 VDD.n498 Vbias 0.03639f
C8745 VDD.n499 Vbias 0.03694f
C8746 VDD.n500 Vbias 0.04583f
C8747 VDD.n501 Vbias 0.03902f
C8748 VDD.n502 Vbias 0.01836f
C8749 VDD.n503 Vbias 0.03639f
C8750 VDD.n504 Vbias 0.50118f
C8751 VDD.n505 Vbias 0.01836f
C8752 VDD.n506 Vbias 0.03639f
C8753 VDD.n507 Vbias 0.50118f
C8754 VDD.n508 Vbias 0.03639f
C8755 VDD.n509 Vbias 0.03694f
C8756 VDD.n510 Vbias 0.04583f
C8757 VDD.n511 Vbias 0.03902f
C8758 VDD.n512 Vbias 0.01836f
C8759 VDD.n513 Vbias 0.03639f
C8760 VDD.n514 Vbias 0.37318f
C8761 VDD.n515 Vbias 0.01836f
C8762 VDD.n516 Vbias 0.03639f
C8763 VDD.n517 Vbias 0.37318f
C8764 VDD.n518 Vbias 0.03639f
C8765 VDD.n519 Vbias 0.03694f
C8766 VDD.n520 Vbias 0.04583f
C8767 VDD.n521 Vbias 0.03902f
C8768 VDD.n522 Vbias 0.01836f
C8769 VDD.n523 Vbias 0.03639f
C8770 VDD.n524 Vbias 0.37318f
C8771 VDD.n525 Vbias 0.01836f
C8772 VDD.n526 Vbias 0.03639f
C8773 VDD.n527 Vbias 0.37318f
C8774 VDD.n528 Vbias 0.03639f
C8775 VDD.n529 Vbias 0.03694f
C8776 VDD.n530 Vbias 0.04583f
C8777 VDD.n531 Vbias 0.03902f
C8778 VDD.n532 Vbias 0.01836f
C8779 VDD.n533 Vbias 0.03639f
C8780 VDD.n534 Vbias 0.50118f
C8781 VDD.n535 Vbias 0.50118f
C8782 VDD.n536 Vbias 0.03639f
C8783 VDD.n537 Vbias 0.01999f
C8784 VDD.n538 Vbias 0.06648f
C8785 VDD.n539 Vbias 0.01309f
C8786 VDD.n540 Vbias 0.07184f
C8787 VDD.n541 Vbias 0.19384f
C8788 VDD.t849 Vbias 0.017f
C8789 VDD.n542 Vbias 0.01999f
C8790 VDD.n543 Vbias 0.03694f
C8791 VDD.n544 Vbias 0.0216f
C8792 VDD.n545 Vbias 0.03694f
C8793 VDD.n546 Vbias 0.45845f
C8794 VDD.t848 Vbias 0.54191f
C8795 VDD.n548 Vbias 0.03639f
C8796 VDD.t648 Vbias 0.46278f
C8797 VDD.n549 Vbias 0.03694f
C8798 VDD.n550 Vbias 0.03694f
C8799 VDD.n551 Vbias 0.0216f
C8800 VDD.n552 Vbias 0.01836f
C8801 VDD.t649 Vbias 0.017f
C8802 VDD.t709 Vbias 0.017f
C8803 VDD.n553 Vbias 0.09713f
C8804 VDD.n554 Vbias 0.01914f
C8805 VDD.n555 Vbias 0.03902f
C8806 VDD.n556 Vbias 0.03694f
C8807 VDD.n557 Vbias 0.0216f
C8808 VDD.n558 Vbias 0.01836f
C8809 VDD.n559 Vbias 0.03639f
C8810 VDD.t316 Vbias 0.46278f
C8811 VDD.n560 Vbias 0.03694f
C8812 VDD.n561 Vbias 0.03694f
C8813 VDD.n562 Vbias 0.0216f
C8814 VDD.n563 Vbias 0.01836f
C8815 VDD.n564 Vbias 0.02305f
C8816 VDD.n565 Vbias 0.03902f
C8817 VDD.n566 Vbias 0.03694f
C8818 VDD.n567 Vbias 0.0216f
C8819 VDD.n568 Vbias 0.01836f
C8820 VDD.n569 Vbias 0.03639f
C8821 VDD.t514 Vbias 0.46278f
C8822 VDD.n570 Vbias 0.03694f
C8823 VDD.n571 Vbias 0.03694f
C8824 VDD.n572 Vbias 0.0216f
C8825 VDD.n573 Vbias 0.01836f
C8826 VDD.t980 Vbias 0.0169f
C8827 VDD.t515 Vbias 0.0169f
C8828 VDD.n574 Vbias 0.07902f
C8829 VDD.t317 Vbias 0.0169f
C8830 VDD.t518 Vbias 0.0169f
C8831 VDD.n575 Vbias 0.07902f
C8832 VDD.n576 Vbias 0.03023f
C8833 VDD.n577 Vbias 0.01699f
C8834 VDD.n578 Vbias 0.03902f
C8835 VDD.n579 Vbias 0.03694f
C8836 VDD.n580 Vbias 0.0216f
C8837 VDD.n581 Vbias 0.01836f
C8838 VDD.n582 Vbias 0.03639f
C8839 VDD.t484 Vbias 0.46278f
C8840 VDD.n583 Vbias 0.03694f
C8841 VDD.n584 Vbias 0.03694f
C8842 VDD.n585 Vbias 0.0216f
C8843 VDD.n586 Vbias 0.01836f
C8844 VDD.t708 Vbias 0.017f
C8845 VDD.t485 Vbias 0.017f
C8846 VDD.n587 Vbias 0.09713f
C8847 VDD.n588 Vbias 0.01914f
C8848 VDD.n589 Vbias 0.03902f
C8849 VDD.n590 Vbias 0.03694f
C8850 VDD.n591 Vbias 0.0216f
C8851 VDD.n592 Vbias 0.01836f
C8852 VDD.n593 Vbias 0.03639f
C8853 VDD.t635 Vbias 0.46278f
C8854 VDD.n594 Vbias 0.03694f
C8855 VDD.n595 Vbias 0.03694f
C8856 VDD.n596 Vbias 0.0216f
C8857 VDD.n597 Vbias 0.01836f
C8858 VDD.n598 Vbias 0.02305f
C8859 VDD.n599 Vbias 0.03902f
C8860 VDD.n600 Vbias 0.03694f
C8861 VDD.n601 Vbias 0.0216f
C8862 VDD.n602 Vbias 0.01836f
C8863 VDD.n603 Vbias 0.03639f
C8864 VDD.t176 Vbias 0.46278f
C8865 VDD.n604 Vbias 0.03694f
C8866 VDD.n605 Vbias 0.03694f
C8867 VDD.n606 Vbias 0.0216f
C8868 VDD.n607 Vbias 0.01836f
C8869 VDD.t982 Vbias 0.0169f
C8870 VDD.t177 Vbias 0.0169f
C8871 VDD.n608 Vbias 0.07902f
C8872 VDD.t636 Vbias 0.0169f
C8873 VDD.t288 Vbias 0.0169f
C8874 VDD.n609 Vbias 0.07902f
C8875 VDD.n610 Vbias 0.03023f
C8876 VDD.n611 Vbias 0.01699f
C8877 VDD.n612 Vbias 0.03902f
C8878 VDD.n613 Vbias 0.03694f
C8879 VDD.n614 Vbias 0.0216f
C8880 VDD.n615 Vbias 0.01836f
C8881 VDD.t516 Vbias 0.46278f
C8882 VDD.n616 Vbias 0.03694f
C8883 VDD.n617 Vbias 0.03694f
C8884 VDD.n618 Vbias 0.06648f
C8885 VDD.n619 Vbias 0.03639f
C8886 VDD.t216 Vbias 0.46278f
C8887 VDD.n620 Vbias 0.03694f
C8888 VDD.n621 Vbias 0.03694f
C8889 VDD.n622 Vbias 0.0216f
C8890 VDD.n623 Vbias 0.01836f
C8891 VDD.t517 Vbias 0.017f
C8892 VDD.n624 Vbias 0.05322f
C8893 VDD.n625 Vbias 0.01309f
C8894 VDD.n626 Vbias 0.01699f
C8895 VDD.n627 Vbias 0.03902f
C8896 VDD.n628 Vbias 0.03694f
C8897 VDD.n629 Vbias 0.0216f
C8898 VDD.n630 Vbias 0.01836f
C8899 VDD.n631 Vbias 0.03639f
C8900 VDD.t266 Vbias 0.46278f
C8901 VDD.n632 Vbias 0.03694f
C8902 VDD.n633 Vbias 0.03694f
C8903 VDD.n634 Vbias 0.0216f
C8904 VDD.n635 Vbias 0.01836f
C8905 VDD.t287 Vbias 0.0169f
C8906 VDD.t268 Vbias 0.0169f
C8907 VDD.n636 Vbias 0.07902f
C8908 VDD.t217 Vbias 0.0169f
C8909 VDD.t267 Vbias 0.0169f
C8910 VDD.n637 Vbias 0.07902f
C8911 VDD.n638 Vbias 0.03023f
C8912 VDD.n639 Vbias 0.01699f
C8913 VDD.n640 Vbias 0.03902f
C8914 VDD.n641 Vbias 0.03694f
C8915 VDD.n642 Vbias 0.0216f
C8916 VDD.n643 Vbias 0.01836f
C8917 VDD.n644 Vbias 0.03639f
C8918 VDD.t652 Vbias 0.46278f
C8919 VDD.n645 Vbias 0.03694f
C8920 VDD.n646 Vbias 0.03694f
C8921 VDD.n647 Vbias 0.0216f
C8922 VDD.n648 Vbias 0.01836f
C8923 VDD.t710 Vbias 0.017f
C8924 VDD.t653 Vbias 0.017f
C8925 VDD.n649 Vbias 0.09713f
C8926 VDD.n650 Vbias 0.01914f
C8927 VDD.n651 Vbias 0.03902f
C8928 VDD.n652 Vbias 0.03694f
C8929 VDD.n653 Vbias 0.0216f
C8930 VDD.n654 Vbias 0.01836f
C8931 VDD.n655 Vbias 0.03639f
C8932 VDD.t252 Vbias 0.46278f
C8933 VDD.n656 Vbias 0.03694f
C8934 VDD.n657 Vbias 0.03694f
C8935 VDD.n658 Vbias 0.0216f
C8936 VDD.n659 Vbias 0.01836f
C8937 VDD.n660 Vbias 0.02305f
C8938 VDD.n661 Vbias 0.03902f
C8939 VDD.n662 Vbias 0.03694f
C8940 VDD.n663 Vbias 0.0216f
C8941 VDD.n664 Vbias 0.01836f
C8942 VDD.n665 Vbias 0.03639f
C8943 VDD.t240 Vbias 0.46278f
C8944 VDD.n666 Vbias 0.03694f
C8945 VDD.n667 Vbias 0.03694f
C8946 VDD.n668 Vbias 0.0216f
C8947 VDD.n669 Vbias 0.01836f
C8948 VDD.t253 Vbias 0.0169f
C8949 VDD.t241 Vbias 0.0169f
C8950 VDD.n670 Vbias 0.07902f
C8951 VDD.t350 Vbias 0.0169f
C8952 VDD.t896 Vbias 0.0169f
C8953 VDD.n671 Vbias 0.07902f
C8954 VDD.n672 Vbias 0.03023f
C8955 VDD.n673 Vbias 0.01699f
C8956 VDD.n674 Vbias 0.03902f
C8957 VDD.n675 Vbias 0.03694f
C8958 VDD.n676 Vbias 0.0216f
C8959 VDD.n677 Vbias 0.01836f
C8960 VDD.n678 Vbias 0.01836f
C8961 VDD.n679 Vbias 0.03639f
C8962 VDD.n680 Vbias 0.50118f
C8963 VDD.n681 Vbias 0.03639f
C8964 VDD.n682 Vbias 0.03694f
C8965 VDD.n683 Vbias 0.04583f
C8966 VDD.n684 Vbias 0.03902f
C8967 VDD.n685 Vbias 0.01836f
C8968 VDD.n686 Vbias 0.03639f
C8969 VDD.n687 Vbias 0.37318f
C8970 VDD.n688 Vbias 0.01836f
C8971 VDD.n689 Vbias 0.03639f
C8972 VDD.n690 Vbias 0.37318f
C8973 VDD.n691 Vbias 0.03639f
C8974 VDD.n692 Vbias 0.03694f
C8975 VDD.n693 Vbias 0.04583f
C8976 VDD.n694 Vbias 0.03902f
C8977 VDD.n695 Vbias 0.01836f
C8978 VDD.n696 Vbias 0.03639f
C8979 VDD.n697 Vbias 0.37318f
C8980 VDD.n698 Vbias 0.01836f
C8981 VDD.n699 Vbias 0.03639f
C8982 VDD.n700 Vbias 0.37318f
C8983 VDD.n701 Vbias 0.03639f
C8984 VDD.n702 Vbias 0.03694f
C8985 VDD.n703 Vbias 0.04583f
C8986 VDD.n704 Vbias 0.03902f
C8987 VDD.n705 Vbias 0.01836f
C8988 VDD.n706 Vbias 0.03639f
C8989 VDD.n707 Vbias 0.50118f
C8990 VDD.n708 Vbias 0.01836f
C8991 VDD.n709 Vbias 0.03639f
C8992 VDD.n710 Vbias 0.50118f
C8993 VDD.n711 Vbias 0.03639f
C8994 VDD.n712 Vbias 0.03694f
C8995 VDD.n713 Vbias 0.04583f
C8996 VDD.n714 Vbias 0.03902f
C8997 VDD.n715 Vbias 0.01836f
C8998 VDD.n716 Vbias 0.03639f
C8999 VDD.n717 Vbias 0.37318f
C9000 VDD.n718 Vbias 0.01836f
C9001 VDD.n719 Vbias 0.03639f
C9002 VDD.n720 Vbias 0.37318f
C9003 VDD.n721 Vbias 0.03639f
C9004 VDD.n722 Vbias 0.03694f
C9005 VDD.n723 Vbias 0.04583f
C9006 VDD.n724 Vbias 0.03902f
C9007 VDD.n725 Vbias 0.01836f
C9008 VDD.n726 Vbias 0.03639f
C9009 VDD.n727 Vbias 0.50118f
C9010 VDD.n728 Vbias 0.50118f
C9011 VDD.n729 Vbias 0.03639f
C9012 VDD.n730 Vbias 0.01999f
C9013 VDD.n731 Vbias 0.0216f
C9014 VDD.n732 Vbias 0.01999f
C9015 VDD.n733 Vbias 0.03639f
C9016 VDD.n734 Vbias 0.50118f
C9017 VDD.n735 Vbias 0.01836f
C9018 VDD.n736 Vbias 0.03639f
C9019 VDD.n737 Vbias 0.50118f
C9020 VDD.n738 Vbias 0.03639f
C9021 VDD.n739 Vbias 0.03694f
C9022 VDD.n740 Vbias 0.04583f
C9023 VDD.n741 Vbias 0.03902f
C9024 VDD.n742 Vbias 0.01836f
C9025 VDD.n743 Vbias 0.03639f
C9026 VDD.n744 Vbias 0.37318f
C9027 VDD.n745 Vbias 0.01836f
C9028 VDD.n746 Vbias 0.03639f
C9029 VDD.n747 Vbias 0.37318f
C9030 VDD.n748 Vbias 0.03639f
C9031 VDD.n749 Vbias 0.03694f
C9032 VDD.n750 Vbias 0.04583f
C9033 VDD.n751 Vbias 0.03902f
C9034 VDD.n752 Vbias 0.01836f
C9035 VDD.n753 Vbias 0.03639f
C9036 VDD.n754 Vbias 0.37318f
C9037 VDD.n755 Vbias 0.01836f
C9038 VDD.n756 Vbias 0.03639f
C9039 VDD.n757 Vbias 0.37318f
C9040 VDD.n758 Vbias 0.03639f
C9041 VDD.n759 Vbias 0.03694f
C9042 VDD.n760 Vbias 0.04583f
C9043 VDD.n761 Vbias 0.03902f
C9044 VDD.n762 Vbias 0.01836f
C9045 VDD.n763 Vbias 0.03639f
C9046 VDD.n764 Vbias 0.50118f
C9047 VDD.n765 Vbias 0.01836f
C9048 VDD.n766 Vbias 0.03639f
C9049 VDD.n767 Vbias 0.50118f
C9050 VDD.n768 Vbias 0.03639f
C9051 VDD.n769 Vbias 0.03694f
C9052 VDD.n770 Vbias 0.04583f
C9053 VDD.n771 Vbias 0.03902f
C9054 VDD.n772 Vbias 0.01836f
C9055 VDD.n773 Vbias 0.03639f
C9056 VDD.n774 Vbias 0.37318f
C9057 VDD.n775 Vbias 0.01836f
C9058 VDD.n776 Vbias 0.03639f
C9059 VDD.n777 Vbias 0.37318f
C9060 VDD.n778 Vbias 0.03639f
C9061 VDD.n779 Vbias 0.03694f
C9062 VDD.n780 Vbias 0.04583f
C9063 VDD.n781 Vbias 0.03902f
C9064 VDD.n782 Vbias 0.01836f
C9065 VDD.n783 Vbias 0.03639f
C9066 VDD.n784 Vbias 0.37318f
C9067 VDD.n785 Vbias 0.01836f
C9068 VDD.n786 Vbias 0.03639f
C9069 VDD.n787 Vbias 0.37318f
C9070 VDD.n788 Vbias 0.03639f
C9071 VDD.n789 Vbias 0.03694f
C9072 VDD.n790 Vbias 0.04583f
C9073 VDD.n791 Vbias 0.03902f
C9074 VDD.n792 Vbias 0.01836f
C9075 VDD.n793 Vbias 0.03639f
C9076 VDD.n794 Vbias 0.50118f
C9077 VDD.n795 Vbias 0.50118f
C9078 VDD.n796 Vbias 0.03639f
C9079 VDD.n797 Vbias 0.01999f
C9080 VDD.n798 Vbias 0.06648f
C9081 VDD.n799 Vbias 0.01309f
C9082 VDD.n800 Vbias 0.07184f
C9083 VDD.n801 Vbias 0.23842f
C9084 VDD.t942 Vbias 0.017f
C9085 VDD.n802 Vbias 0.01999f
C9086 VDD.n803 Vbias 0.03694f
C9087 VDD.n804 Vbias 0.0216f
C9088 VDD.n805 Vbias 0.03694f
C9089 VDD.n806 Vbias 0.45845f
C9090 VDD.t941 Vbias 0.54191f
C9091 VDD.n808 Vbias 0.03639f
C9092 VDD.t392 Vbias 0.46278f
C9093 VDD.n809 Vbias 0.03694f
C9094 VDD.n810 Vbias 0.03694f
C9095 VDD.n811 Vbias 0.0216f
C9096 VDD.n812 Vbias 0.01836f
C9097 VDD.t393 Vbias 0.017f
C9098 VDD.t573 Vbias 0.017f
C9099 VDD.n813 Vbias 0.09713f
C9100 VDD.n814 Vbias 0.01914f
C9101 VDD.n815 Vbias 0.03902f
C9102 VDD.n816 Vbias 0.03694f
C9103 VDD.n817 Vbias 0.0216f
C9104 VDD.n818 Vbias 0.01836f
C9105 VDD.n819 Vbias 0.03639f
C9106 VDD.t585 Vbias 0.46278f
C9107 VDD.n820 Vbias 0.03694f
C9108 VDD.n821 Vbias 0.03694f
C9109 VDD.n822 Vbias 0.0216f
C9110 VDD.n823 Vbias 0.01836f
C9111 VDD.n824 Vbias 0.02305f
C9112 VDD.n825 Vbias 0.03902f
C9113 VDD.n826 Vbias 0.03694f
C9114 VDD.n827 Vbias 0.0216f
C9115 VDD.n828 Vbias 0.01836f
C9116 VDD.n829 Vbias 0.03639f
C9117 VDD.t612 Vbias 0.46278f
C9118 VDD.n830 Vbias 0.03694f
C9119 VDD.n831 Vbias 0.03694f
C9120 VDD.n832 Vbias 0.0216f
C9121 VDD.n833 Vbias 0.01836f
C9122 VDD.t845 Vbias 0.0169f
C9123 VDD.t614 Vbias 0.0169f
C9124 VDD.n834 Vbias 0.07902f
C9125 VDD.t586 Vbias 0.0169f
C9126 VDD.t613 Vbias 0.0169f
C9127 VDD.n835 Vbias 0.07902f
C9128 VDD.n836 Vbias 0.03023f
C9129 VDD.n837 Vbias 0.01699f
C9130 VDD.n838 Vbias 0.03902f
C9131 VDD.n839 Vbias 0.03694f
C9132 VDD.n840 Vbias 0.0216f
C9133 VDD.n841 Vbias 0.01836f
C9134 VDD.n842 Vbias 0.03639f
C9135 VDD.t434 Vbias 0.46278f
C9136 VDD.n843 Vbias 0.03694f
C9137 VDD.n844 Vbias 0.03694f
C9138 VDD.n845 Vbias 0.0216f
C9139 VDD.n846 Vbias 0.01836f
C9140 VDD.t826 Vbias 0.017f
C9141 VDD.t435 Vbias 0.017f
C9142 VDD.n847 Vbias 0.09713f
C9143 VDD.n848 Vbias 0.01914f
C9144 VDD.n849 Vbias 0.03902f
C9145 VDD.n850 Vbias 0.03694f
C9146 VDD.n851 Vbias 0.0216f
C9147 VDD.n852 Vbias 0.01836f
C9148 VDD.n853 Vbias 0.03639f
C9149 VDD.t168 Vbias 0.46278f
C9150 VDD.n854 Vbias 0.03694f
C9151 VDD.n855 Vbias 0.03694f
C9152 VDD.n856 Vbias 0.0216f
C9153 VDD.n857 Vbias 0.01836f
C9154 VDD.n858 Vbias 0.02305f
C9155 VDD.n859 Vbias 0.03902f
C9156 VDD.n860 Vbias 0.03694f
C9157 VDD.n861 Vbias 0.0216f
C9158 VDD.n862 Vbias 0.01836f
C9159 VDD.n863 Vbias 0.03639f
C9160 VDD.t138 Vbias 0.46278f
C9161 VDD.n864 Vbias 0.03694f
C9162 VDD.n865 Vbias 0.03694f
C9163 VDD.n866 Vbias 0.0216f
C9164 VDD.n867 Vbias 0.01836f
C9165 VDD.t169 Vbias 0.0169f
C9166 VDD.t139 Vbias 0.0169f
C9167 VDD.n868 Vbias 0.07902f
C9168 VDD.t558 Vbias 0.0169f
C9169 VDD.t962 Vbias 0.0169f
C9170 VDD.n869 Vbias 0.07902f
C9171 VDD.n870 Vbias 0.03023f
C9172 VDD.n871 Vbias 0.01699f
C9173 VDD.n872 Vbias 0.03902f
C9174 VDD.n873 Vbias 0.03694f
C9175 VDD.n874 Vbias 0.0216f
C9176 VDD.n875 Vbias 0.01836f
C9177 VDD.t178 Vbias 0.46278f
C9178 VDD.n876 Vbias 0.03694f
C9179 VDD.n877 Vbias 0.03694f
C9180 VDD.n878 Vbias 0.06648f
C9181 VDD.n879 Vbias 0.03639f
C9182 VDD.t136 Vbias 0.46278f
C9183 VDD.n880 Vbias 0.03694f
C9184 VDD.n881 Vbias 0.03694f
C9185 VDD.n882 Vbias 0.0216f
C9186 VDD.n883 Vbias 0.01836f
C9187 VDD.t179 Vbias 0.017f
C9188 VDD.n884 Vbias 0.05322f
C9189 VDD.n885 Vbias 0.01309f
C9190 VDD.n886 Vbias 0.01699f
C9191 VDD.n887 Vbias 0.03902f
C9192 VDD.n888 Vbias 0.03694f
C9193 VDD.n889 Vbias 0.0216f
C9194 VDD.n890 Vbias 0.01836f
C9195 VDD.n891 Vbias 0.03639f
C9196 VDD.t675 Vbias 0.46278f
C9197 VDD.n892 Vbias 0.03694f
C9198 VDD.n893 Vbias 0.03694f
C9199 VDD.n894 Vbias 0.0216f
C9200 VDD.n895 Vbias 0.01836f
C9201 VDD.t961 Vbias 0.0169f
C9202 VDD.t676 Vbias 0.0169f
C9203 VDD.n896 Vbias 0.07902f
C9204 VDD.t137 Vbias 0.0169f
C9205 VDD.t677 Vbias 0.0169f
C9206 VDD.n897 Vbias 0.07902f
C9207 VDD.n898 Vbias 0.03023f
C9208 VDD.n899 Vbias 0.01699f
C9209 VDD.n900 Vbias 0.03902f
C9210 VDD.n901 Vbias 0.03694f
C9211 VDD.n902 Vbias 0.0216f
C9212 VDD.n903 Vbias 0.01836f
C9213 VDD.n904 Vbias 0.03639f
C9214 VDD.t574 Vbias 0.46278f
C9215 VDD.n905 Vbias 0.03694f
C9216 VDD.n906 Vbias 0.03694f
C9217 VDD.n907 Vbias 0.0216f
C9218 VDD.n908 Vbias 0.01836f
C9219 VDD.t575 Vbias 0.017f
C9220 VDD.t983 Vbias 0.017f
C9221 VDD.n909 Vbias 0.09713f
C9222 VDD.n910 Vbias 0.01914f
C9223 VDD.n911 Vbias 0.03902f
C9224 VDD.n912 Vbias 0.03694f
C9225 VDD.n913 Vbias 0.0216f
C9226 VDD.n914 Vbias 0.01836f
C9227 VDD.n915 Vbias 0.03639f
C9228 VDD.t313 Vbias 0.46278f
C9229 VDD.n916 Vbias 0.03694f
C9230 VDD.n917 Vbias 0.03694f
C9231 VDD.n918 Vbias 0.0216f
C9232 VDD.n919 Vbias 0.01836f
C9233 VDD.n920 Vbias 0.02305f
C9234 VDD.n921 Vbias 0.03902f
C9235 VDD.n922 Vbias 0.03694f
C9236 VDD.n923 Vbias 0.0216f
C9237 VDD.n924 Vbias 0.01836f
C9238 VDD.n925 Vbias 0.03639f
C9239 VDD.t885 Vbias 0.46278f
C9240 VDD.n926 Vbias 0.03694f
C9241 VDD.n927 Vbias 0.03694f
C9242 VDD.n928 Vbias 0.0216f
C9243 VDD.n929 Vbias 0.01836f
C9244 VDD.t314 Vbias 0.0169f
C9245 VDD.t886 Vbias 0.0169f
C9246 VDD.n930 Vbias 0.07902f
C9247 VDD.t328 Vbias 0.0169f
C9248 VDD.t989 Vbias 0.0169f
C9249 VDD.n931 Vbias 0.07902f
C9250 VDD.n932 Vbias 0.03023f
C9251 VDD.n933 Vbias 0.01699f
C9252 VDD.n934 Vbias 0.03902f
C9253 VDD.n935 Vbias 0.03694f
C9254 VDD.n936 Vbias 0.0216f
C9255 VDD.n937 Vbias 0.01836f
C9256 VDD.n938 Vbias 0.01836f
C9257 VDD.n939 Vbias 0.03639f
C9258 VDD.n940 Vbias 0.50118f
C9259 VDD.n941 Vbias 0.03639f
C9260 VDD.n942 Vbias 0.03694f
C9261 VDD.n943 Vbias 0.04583f
C9262 VDD.n944 Vbias 0.03902f
C9263 VDD.n945 Vbias 0.01836f
C9264 VDD.n946 Vbias 0.03639f
C9265 VDD.n947 Vbias 0.37318f
C9266 VDD.n948 Vbias 0.01836f
C9267 VDD.n949 Vbias 0.03639f
C9268 VDD.n950 Vbias 0.37318f
C9269 VDD.n951 Vbias 0.03639f
C9270 VDD.n952 Vbias 0.03694f
C9271 VDD.n953 Vbias 0.04583f
C9272 VDD.n954 Vbias 0.03902f
C9273 VDD.n955 Vbias 0.01836f
C9274 VDD.n956 Vbias 0.03639f
C9275 VDD.n957 Vbias 0.37318f
C9276 VDD.n958 Vbias 0.01836f
C9277 VDD.n959 Vbias 0.03639f
C9278 VDD.n960 Vbias 0.37318f
C9279 VDD.n961 Vbias 0.03639f
C9280 VDD.n962 Vbias 0.03694f
C9281 VDD.n963 Vbias 0.04583f
C9282 VDD.n964 Vbias 0.03902f
C9283 VDD.n965 Vbias 0.01836f
C9284 VDD.n966 Vbias 0.03639f
C9285 VDD.n967 Vbias 0.50118f
C9286 VDD.n968 Vbias 0.01836f
C9287 VDD.n969 Vbias 0.03639f
C9288 VDD.n970 Vbias 0.50118f
C9289 VDD.n971 Vbias 0.03639f
C9290 VDD.n972 Vbias 0.03694f
C9291 VDD.n973 Vbias 0.04583f
C9292 VDD.n974 Vbias 0.03902f
C9293 VDD.n975 Vbias 0.01836f
C9294 VDD.n976 Vbias 0.03639f
C9295 VDD.n977 Vbias 0.37318f
C9296 VDD.n978 Vbias 0.01836f
C9297 VDD.n979 Vbias 0.03639f
C9298 VDD.n980 Vbias 0.37318f
C9299 VDD.n981 Vbias 0.03639f
C9300 VDD.n982 Vbias 0.03694f
C9301 VDD.n983 Vbias 0.04583f
C9302 VDD.n984 Vbias 0.03902f
C9303 VDD.n985 Vbias 0.01836f
C9304 VDD.n986 Vbias 0.03639f
C9305 VDD.n987 Vbias 0.50118f
C9306 VDD.n988 Vbias 0.50118f
C9307 VDD.n989 Vbias 0.03639f
C9308 VDD.n990 Vbias 0.01999f
C9309 VDD.n991 Vbias 0.0216f
C9310 VDD.n992 Vbias 0.01999f
C9311 VDD.n993 Vbias 0.03639f
C9312 VDD.n994 Vbias 0.50118f
C9313 VDD.n995 Vbias 0.01836f
C9314 VDD.n996 Vbias 0.03639f
C9315 VDD.n997 Vbias 0.50118f
C9316 VDD.n998 Vbias 0.03639f
C9317 VDD.n999 Vbias 0.03694f
C9318 VDD.n1000 Vbias 0.04583f
C9319 VDD.n1001 Vbias 0.03902f
C9320 VDD.n1002 Vbias 0.01836f
C9321 VDD.n1003 Vbias 0.03639f
C9322 VDD.n1004 Vbias 0.37318f
C9323 VDD.n1005 Vbias 0.01836f
C9324 VDD.n1006 Vbias 0.03639f
C9325 VDD.n1007 Vbias 0.37318f
C9326 VDD.n1008 Vbias 0.03639f
C9327 VDD.n1009 Vbias 0.03694f
C9328 VDD.n1010 Vbias 0.04583f
C9329 VDD.n1011 Vbias 0.03902f
C9330 VDD.n1012 Vbias 0.01836f
C9331 VDD.n1013 Vbias 0.03639f
C9332 VDD.n1014 Vbias 0.37318f
C9333 VDD.n1015 Vbias 0.01836f
C9334 VDD.n1016 Vbias 0.03639f
C9335 VDD.n1017 Vbias 0.37318f
C9336 VDD.n1018 Vbias 0.03639f
C9337 VDD.n1019 Vbias 0.03694f
C9338 VDD.n1020 Vbias 0.04583f
C9339 VDD.n1021 Vbias 0.03902f
C9340 VDD.n1022 Vbias 0.01836f
C9341 VDD.n1023 Vbias 0.03639f
C9342 VDD.n1024 Vbias 0.50118f
C9343 VDD.n1025 Vbias 0.01836f
C9344 VDD.n1026 Vbias 0.03639f
C9345 VDD.n1027 Vbias 0.50118f
C9346 VDD.n1028 Vbias 0.03639f
C9347 VDD.n1029 Vbias 0.03694f
C9348 VDD.n1030 Vbias 0.04583f
C9349 VDD.n1031 Vbias 0.03902f
C9350 VDD.n1032 Vbias 0.01836f
C9351 VDD.n1033 Vbias 0.03639f
C9352 VDD.n1034 Vbias 0.37318f
C9353 VDD.n1035 Vbias 0.01836f
C9354 VDD.n1036 Vbias 0.03639f
C9355 VDD.n1037 Vbias 0.37318f
C9356 VDD.n1038 Vbias 0.03639f
C9357 VDD.n1039 Vbias 0.03694f
C9358 VDD.n1040 Vbias 0.04583f
C9359 VDD.n1041 Vbias 0.03902f
C9360 VDD.n1042 Vbias 0.01836f
C9361 VDD.n1043 Vbias 0.03639f
C9362 VDD.n1044 Vbias 0.37318f
C9363 VDD.n1045 Vbias 0.01836f
C9364 VDD.n1046 Vbias 0.03639f
C9365 VDD.n1047 Vbias 0.37318f
C9366 VDD.n1048 Vbias 0.03639f
C9367 VDD.n1049 Vbias 0.03694f
C9368 VDD.n1050 Vbias 0.04583f
C9369 VDD.n1051 Vbias 0.03902f
C9370 VDD.n1052 Vbias 0.01836f
C9371 VDD.n1053 Vbias 0.03639f
C9372 VDD.n1054 Vbias 0.50118f
C9373 VDD.n1055 Vbias 0.50118f
C9374 VDD.n1056 Vbias 0.03639f
C9375 VDD.n1057 Vbias 0.01999f
C9376 VDD.n1058 Vbias 0.06648f
C9377 VDD.n1059 Vbias 0.01309f
C9378 VDD.n1060 Vbias 0.07184f
C9379 VDD.n1061 Vbias 0.23842f
C9380 VDD.t977 Vbias 0.017f
C9381 VDD.n1062 Vbias 0.01999f
C9382 VDD.n1063 Vbias 0.03694f
C9383 VDD.n1064 Vbias 0.0216f
C9384 VDD.n1065 Vbias 0.03694f
C9385 VDD.n1066 Vbias 0.45845f
C9386 VDD.t976 Vbias 0.54191f
C9387 VDD.n1068 Vbias 0.03639f
C9388 VDD.t71 Vbias 0.46278f
C9389 VDD.n1069 Vbias 0.03694f
C9390 VDD.n1070 Vbias 0.03694f
C9391 VDD.n1071 Vbias 0.0216f
C9392 VDD.n1072 Vbias 0.01836f
C9393 VDD.t72 Vbias 0.017f
C9394 VDD.t948 Vbias 0.017f
C9395 VDD.n1073 Vbias 0.09713f
C9396 VDD.n1074 Vbias 0.01914f
C9397 VDD.n1075 Vbias 0.03902f
C9398 VDD.n1076 Vbias 0.03694f
C9399 VDD.n1077 Vbias 0.0216f
C9400 VDD.n1078 Vbias 0.01836f
C9401 VDD.n1079 Vbias 0.03639f
C9402 VDD.t226 Vbias 0.46278f
C9403 VDD.n1080 Vbias 0.03694f
C9404 VDD.n1081 Vbias 0.03694f
C9405 VDD.n1082 Vbias 0.0216f
C9406 VDD.n1083 Vbias 0.01836f
C9407 VDD.n1084 Vbias 0.02305f
C9408 VDD.n1085 Vbias 0.03902f
C9409 VDD.n1086 Vbias 0.03694f
C9410 VDD.n1087 Vbias 0.0216f
C9411 VDD.n1088 Vbias 0.01836f
C9412 VDD.n1089 Vbias 0.03639f
C9413 VDD.t140 Vbias 0.46278f
C9414 VDD.n1090 Vbias 0.03694f
C9415 VDD.n1091 Vbias 0.03694f
C9416 VDD.n1092 Vbias 0.0216f
C9417 VDD.n1093 Vbias 0.01836f
C9418 VDD.t545 Vbias 0.0169f
C9419 VDD.t141 Vbias 0.0169f
C9420 VDD.n1094 Vbias 0.07902f
C9421 VDD.t227 Vbias 0.0169f
C9422 VDD.t458 Vbias 0.0169f
C9423 VDD.n1095 Vbias 0.07902f
C9424 VDD.n1096 Vbias 0.03023f
C9425 VDD.n1097 Vbias 0.01699f
C9426 VDD.n1098 Vbias 0.03902f
C9427 VDD.n1099 Vbias 0.03694f
C9428 VDD.n1100 Vbias 0.0216f
C9429 VDD.n1101 Vbias 0.01836f
C9430 VDD.n1102 Vbias 0.03639f
C9431 VDD.t129 Vbias 0.46278f
C9432 VDD.n1103 Vbias 0.03694f
C9433 VDD.n1104 Vbias 0.03694f
C9434 VDD.n1105 Vbias 0.0216f
C9435 VDD.n1106 Vbias 0.01836f
C9436 VDD.t945 Vbias 0.017f
C9437 VDD.t130 Vbias 0.017f
C9438 VDD.n1107 Vbias 0.09713f
C9439 VDD.n1108 Vbias 0.01914f
C9440 VDD.n1109 Vbias 0.03902f
C9441 VDD.n1110 Vbias 0.03694f
C9442 VDD.n1111 Vbias 0.0216f
C9443 VDD.n1112 Vbias 0.01836f
C9444 VDD.n1113 Vbias 0.03639f
C9445 VDD.t190 Vbias 0.46278f
C9446 VDD.n1114 Vbias 0.03694f
C9447 VDD.n1115 Vbias 0.03694f
C9448 VDD.n1116 Vbias 0.0216f
C9449 VDD.n1117 Vbias 0.01836f
C9450 VDD.n1118 Vbias 0.02305f
C9451 VDD.n1119 Vbias 0.03902f
C9452 VDD.n1120 Vbias 0.03694f
C9453 VDD.n1121 Vbias 0.0216f
C9454 VDD.n1122 Vbias 0.01836f
C9455 VDD.n1123 Vbias 0.03639f
C9456 VDD.t238 Vbias 0.46278f
C9457 VDD.n1124 Vbias 0.03694f
C9458 VDD.n1125 Vbias 0.03694f
C9459 VDD.n1126 Vbias 0.0216f
C9460 VDD.n1127 Vbias 0.01836f
C9461 VDD.t682 Vbias 0.0169f
C9462 VDD.t284 Vbias 0.0169f
C9463 VDD.n1128 Vbias 0.07902f
C9464 VDD.t191 Vbias 0.0169f
C9465 VDD.t239 Vbias 0.0169f
C9466 VDD.n1129 Vbias 0.07902f
C9467 VDD.n1130 Vbias 0.03023f
C9468 VDD.n1131 Vbias 0.01699f
C9469 VDD.n1132 Vbias 0.03902f
C9470 VDD.n1133 Vbias 0.03694f
C9471 VDD.n1134 Vbias 0.0216f
C9472 VDD.n1135 Vbias 0.01836f
C9473 VDD.t142 Vbias 0.46278f
C9474 VDD.n1136 Vbias 0.03694f
C9475 VDD.n1137 Vbias 0.03694f
C9476 VDD.n1138 Vbias 0.06648f
C9477 VDD.n1139 Vbias 0.03639f
C9478 VDD.t230 Vbias 0.46278f
C9479 VDD.n1140 Vbias 0.03694f
C9480 VDD.n1141 Vbias 0.03694f
C9481 VDD.n1142 Vbias 0.0216f
C9482 VDD.n1143 Vbias 0.01836f
C9483 VDD.t143 Vbias 0.017f
C9484 VDD.n1144 Vbias 0.05322f
C9485 VDD.n1145 Vbias 0.01309f
C9486 VDD.n1146 Vbias 0.01699f
C9487 VDD.n1147 Vbias 0.03902f
C9488 VDD.n1148 Vbias 0.03694f
C9489 VDD.n1149 Vbias 0.0216f
C9490 VDD.n1150 Vbias 0.01836f
C9491 VDD.n1151 Vbias 0.03639f
C9492 VDD.t442 Vbias 0.46278f
C9493 VDD.n1152 Vbias 0.03694f
C9494 VDD.n1153 Vbias 0.03694f
C9495 VDD.n1154 Vbias 0.0216f
C9496 VDD.n1155 Vbias 0.01836f
C9497 VDD.t503 Vbias 0.0169f
C9498 VDD.t444 Vbias 0.0169f
C9499 VDD.n1156 Vbias 0.07902f
C9500 VDD.t231 Vbias 0.0169f
C9501 VDD.t443 Vbias 0.0169f
C9502 VDD.n1157 Vbias 0.07902f
C9503 VDD.n1158 Vbias 0.03023f
C9504 VDD.n1159 Vbias 0.01699f
C9505 VDD.n1160 Vbias 0.03902f
C9506 VDD.n1161 Vbias 0.03694f
C9507 VDD.n1162 Vbias 0.0216f
C9508 VDD.n1163 Vbias 0.01836f
C9509 VDD.n1164 Vbias 0.03639f
C9510 VDD.t67 Vbias 0.46278f
C9511 VDD.n1165 Vbias 0.03694f
C9512 VDD.n1166 Vbias 0.03694f
C9513 VDD.n1167 Vbias 0.0216f
C9514 VDD.n1168 Vbias 0.01836f
C9515 VDD.t196 Vbias 0.017f
C9516 VDD.t68 Vbias 0.017f
C9517 VDD.n1169 Vbias 0.09713f
C9518 VDD.n1170 Vbias 0.01914f
C9519 VDD.n1171 Vbias 0.03902f
C9520 VDD.n1172 Vbias 0.03694f
C9521 VDD.n1173 Vbias 0.0216f
C9522 VDD.n1174 Vbias 0.01836f
C9523 VDD.n1175 Vbias 0.03639f
C9524 VDD.t13 Vbias 0.46278f
C9525 VDD.n1176 Vbias 0.03694f
C9526 VDD.n1177 Vbias 0.03694f
C9527 VDD.n1178 Vbias 0.0216f
C9528 VDD.n1179 Vbias 0.01836f
C9529 VDD.n1180 Vbias 0.02305f
C9530 VDD.n1181 Vbias 0.03902f
C9531 VDD.n1182 Vbias 0.03694f
C9532 VDD.n1183 Vbias 0.0216f
C9533 VDD.n1184 Vbias 0.01836f
C9534 VDD.n1185 Vbias 0.03639f
C9535 VDD.t188 Vbias 0.46278f
C9536 VDD.n1186 Vbias 0.03694f
C9537 VDD.n1187 Vbias 0.03694f
C9538 VDD.n1188 Vbias 0.0216f
C9539 VDD.n1189 Vbias 0.01836f
C9540 VDD.t362 Vbias 0.0169f
C9541 VDD.t189 Vbias 0.0169f
C9542 VDD.n1190 Vbias 0.07902f
C9543 VDD.t14 Vbias 0.0169f
C9544 VDD.t973 Vbias 0.0169f
C9545 VDD.n1191 Vbias 0.07902f
C9546 VDD.n1192 Vbias 0.03023f
C9547 VDD.n1193 Vbias 0.01699f
C9548 VDD.n1194 Vbias 0.03902f
C9549 VDD.n1195 Vbias 0.03694f
C9550 VDD.n1196 Vbias 0.0216f
C9551 VDD.n1197 Vbias 0.01836f
C9552 VDD.n1198 Vbias 0.01836f
C9553 VDD.n1199 Vbias 0.03639f
C9554 VDD.n1200 Vbias 0.50118f
C9555 VDD.n1201 Vbias 0.03639f
C9556 VDD.n1202 Vbias 0.03694f
C9557 VDD.n1203 Vbias 0.04583f
C9558 VDD.n1204 Vbias 0.03902f
C9559 VDD.n1205 Vbias 0.01836f
C9560 VDD.n1206 Vbias 0.03639f
C9561 VDD.n1207 Vbias 0.37318f
C9562 VDD.n1208 Vbias 0.01836f
C9563 VDD.n1209 Vbias 0.03639f
C9564 VDD.n1210 Vbias 0.37318f
C9565 VDD.n1211 Vbias 0.03639f
C9566 VDD.n1212 Vbias 0.03694f
C9567 VDD.n1213 Vbias 0.04583f
C9568 VDD.n1214 Vbias 0.03902f
C9569 VDD.n1215 Vbias 0.01836f
C9570 VDD.n1216 Vbias 0.03639f
C9571 VDD.n1217 Vbias 0.37318f
C9572 VDD.n1218 Vbias 0.01836f
C9573 VDD.n1219 Vbias 0.03639f
C9574 VDD.n1220 Vbias 0.37318f
C9575 VDD.n1221 Vbias 0.03639f
C9576 VDD.n1222 Vbias 0.03694f
C9577 VDD.n1223 Vbias 0.04583f
C9578 VDD.n1224 Vbias 0.03902f
C9579 VDD.n1225 Vbias 0.01836f
C9580 VDD.n1226 Vbias 0.03639f
C9581 VDD.n1227 Vbias 0.50118f
C9582 VDD.n1228 Vbias 0.01836f
C9583 VDD.n1229 Vbias 0.03639f
C9584 VDD.n1230 Vbias 0.50118f
C9585 VDD.n1231 Vbias 0.03639f
C9586 VDD.n1232 Vbias 0.03694f
C9587 VDD.n1233 Vbias 0.04583f
C9588 VDD.n1234 Vbias 0.03902f
C9589 VDD.n1235 Vbias 0.01836f
C9590 VDD.n1236 Vbias 0.03639f
C9591 VDD.n1237 Vbias 0.37318f
C9592 VDD.n1238 Vbias 0.01836f
C9593 VDD.n1239 Vbias 0.03639f
C9594 VDD.n1240 Vbias 0.37318f
C9595 VDD.n1241 Vbias 0.03639f
C9596 VDD.n1242 Vbias 0.03694f
C9597 VDD.n1243 Vbias 0.04583f
C9598 VDD.n1244 Vbias 0.03902f
C9599 VDD.n1245 Vbias 0.01836f
C9600 VDD.n1246 Vbias 0.03639f
C9601 VDD.n1247 Vbias 0.50118f
C9602 VDD.n1248 Vbias 0.50118f
C9603 VDD.n1249 Vbias 0.03639f
C9604 VDD.n1250 Vbias 0.01999f
C9605 VDD.n1251 Vbias 0.0216f
C9606 VDD.n1252 Vbias 0.01999f
C9607 VDD.n1253 Vbias 0.03639f
C9608 VDD.n1254 Vbias 0.50118f
C9609 VDD.n1255 Vbias 0.01836f
C9610 VDD.n1256 Vbias 0.03639f
C9611 VDD.n1257 Vbias 0.50118f
C9612 VDD.n1258 Vbias 0.03639f
C9613 VDD.n1259 Vbias 0.03694f
C9614 VDD.n1260 Vbias 0.04583f
C9615 VDD.n1261 Vbias 0.03902f
C9616 VDD.n1262 Vbias 0.01836f
C9617 VDD.n1263 Vbias 0.03639f
C9618 VDD.n1264 Vbias 0.37318f
C9619 VDD.n1265 Vbias 0.01836f
C9620 VDD.n1266 Vbias 0.03639f
C9621 VDD.n1267 Vbias 0.37318f
C9622 VDD.n1268 Vbias 0.03639f
C9623 VDD.n1269 Vbias 0.03694f
C9624 VDD.n1270 Vbias 0.04583f
C9625 VDD.n1271 Vbias 0.03902f
C9626 VDD.n1272 Vbias 0.01836f
C9627 VDD.n1273 Vbias 0.03639f
C9628 VDD.n1274 Vbias 0.37318f
C9629 VDD.n1275 Vbias 0.01836f
C9630 VDD.n1276 Vbias 0.03639f
C9631 VDD.n1277 Vbias 0.37318f
C9632 VDD.n1278 Vbias 0.03639f
C9633 VDD.n1279 Vbias 0.03694f
C9634 VDD.n1280 Vbias 0.04583f
C9635 VDD.n1281 Vbias 0.03902f
C9636 VDD.n1282 Vbias 0.01836f
C9637 VDD.n1283 Vbias 0.03639f
C9638 VDD.n1284 Vbias 0.50118f
C9639 VDD.n1285 Vbias 0.01836f
C9640 VDD.n1286 Vbias 0.03639f
C9641 VDD.n1287 Vbias 0.50118f
C9642 VDD.n1288 Vbias 0.03639f
C9643 VDD.n1289 Vbias 0.03694f
C9644 VDD.n1290 Vbias 0.04583f
C9645 VDD.n1291 Vbias 0.03902f
C9646 VDD.n1292 Vbias 0.01836f
C9647 VDD.n1293 Vbias 0.03639f
C9648 VDD.n1294 Vbias 0.37318f
C9649 VDD.n1295 Vbias 0.01836f
C9650 VDD.n1296 Vbias 0.03639f
C9651 VDD.n1297 Vbias 0.37318f
C9652 VDD.n1298 Vbias 0.03639f
C9653 VDD.n1299 Vbias 0.03694f
C9654 VDD.n1300 Vbias 0.04583f
C9655 VDD.n1301 Vbias 0.03902f
C9656 VDD.n1302 Vbias 0.01836f
C9657 VDD.n1303 Vbias 0.03639f
C9658 VDD.n1304 Vbias 0.37318f
C9659 VDD.n1305 Vbias 0.01836f
C9660 VDD.n1306 Vbias 0.03639f
C9661 VDD.n1307 Vbias 0.37318f
C9662 VDD.n1308 Vbias 0.03639f
C9663 VDD.n1309 Vbias 0.03694f
C9664 VDD.n1310 Vbias 0.04583f
C9665 VDD.n1311 Vbias 0.03902f
C9666 VDD.n1312 Vbias 0.01836f
C9667 VDD.n1313 Vbias 0.03639f
C9668 VDD.n1314 Vbias 0.50118f
C9669 VDD.n1315 Vbias 0.50118f
C9670 VDD.n1316 Vbias 0.03639f
C9671 VDD.n1317 Vbias 0.01999f
C9672 VDD.n1318 Vbias 0.06648f
C9673 VDD.n1319 Vbias 0.01309f
C9674 VDD.n1320 Vbias 0.07184f
C9675 VDD.n1321 Vbias 0.30746f
C9676 VDD.t853 Vbias 0.017f
C9677 VDD.n1322 Vbias 0.01999f
C9678 VDD.n1323 Vbias 0.03694f
C9679 VDD.n1324 Vbias 0.0216f
C9680 VDD.n1325 Vbias 0.03694f
C9681 VDD.n1326 Vbias 0.45845f
C9682 VDD.t852 Vbias 0.54191f
C9683 VDD.n1328 Vbias 0.03639f
C9684 VDD.t432 Vbias 0.46278f
C9685 VDD.n1329 Vbias 0.03694f
C9686 VDD.n1330 Vbias 0.03694f
C9687 VDD.n1331 Vbias 0.0216f
C9688 VDD.n1332 Vbias 0.01836f
C9689 VDD.t433 Vbias 0.017f
C9690 VDD.t883 Vbias 0.017f
C9691 VDD.n1333 Vbias 0.09713f
C9692 VDD.n1334 Vbias 0.01914f
C9693 VDD.n1335 Vbias 0.03902f
C9694 VDD.n1336 Vbias 0.03694f
C9695 VDD.n1337 Vbias 0.0216f
C9696 VDD.n1338 Vbias 0.01836f
C9697 VDD.n1339 Vbias 0.03639f
C9698 VDD.t264 Vbias 0.46278f
C9699 VDD.n1340 Vbias 0.03694f
C9700 VDD.n1341 Vbias 0.03694f
C9701 VDD.n1342 Vbias 0.0216f
C9702 VDD.n1343 Vbias 0.01836f
C9703 VDD.n1344 Vbias 0.02305f
C9704 VDD.n1345 Vbias 0.03902f
C9705 VDD.n1346 Vbias 0.03694f
C9706 VDD.n1347 Vbias 0.0216f
C9707 VDD.n1348 Vbias 0.01836f
C9708 VDD.n1349 Vbias 0.03639f
C9709 VDD.t416 Vbias 0.46278f
C9710 VDD.n1350 Vbias 0.03694f
C9711 VDD.n1351 Vbias 0.03694f
C9712 VDD.n1352 Vbias 0.0216f
C9713 VDD.n1353 Vbias 0.01836f
C9714 VDD.t631 Vbias 0.0169f
C9715 VDD.t417 Vbias 0.0169f
C9716 VDD.n1354 Vbias 0.07902f
C9717 VDD.t265 Vbias 0.0169f
C9718 VDD.t420 Vbias 0.0169f
C9719 VDD.n1355 Vbias 0.07902f
C9720 VDD.n1356 Vbias 0.03023f
C9721 VDD.n1357 Vbias 0.01699f
C9722 VDD.n1358 Vbias 0.03902f
C9723 VDD.n1359 Vbias 0.03694f
C9724 VDD.n1360 Vbias 0.0216f
C9725 VDD.n1361 Vbias 0.01836f
C9726 VDD.n1362 Vbias 0.03639f
C9727 VDD.t881 Vbias 0.46278f
C9728 VDD.n1363 Vbias 0.03694f
C9729 VDD.n1364 Vbias 0.03694f
C9730 VDD.n1365 Vbias 0.0216f
C9731 VDD.n1366 Vbias 0.01836f
C9732 VDD.t882 Vbias 0.017f
C9733 VDD.t987 Vbias 0.017f
C9734 VDD.n1367 Vbias 0.09713f
C9735 VDD.n1368 Vbias 0.01914f
C9736 VDD.n1369 Vbias 0.03902f
C9737 VDD.n1370 Vbias 0.03694f
C9738 VDD.n1371 Vbias 0.0216f
C9739 VDD.n1372 Vbias 0.01836f
C9740 VDD.n1373 Vbias 0.03639f
C9741 VDD.t523 Vbias 0.46278f
C9742 VDD.n1374 Vbias 0.03694f
C9743 VDD.n1375 Vbias 0.03694f
C9744 VDD.n1376 Vbias 0.0216f
C9745 VDD.n1377 Vbias 0.01836f
C9746 VDD.n1378 Vbias 0.02305f
C9747 VDD.n1379 Vbias 0.03902f
C9748 VDD.n1380 Vbias 0.03694f
C9749 VDD.n1381 Vbias 0.0216f
C9750 VDD.n1382 Vbias 0.01836f
C9751 VDD.n1383 Vbias 0.03639f
C9752 VDD.t687 Vbias 0.46278f
C9753 VDD.n1384 Vbias 0.03694f
C9754 VDD.n1385 Vbias 0.03694f
C9755 VDD.n1386 Vbias 0.0216f
C9756 VDD.n1387 Vbias 0.01836f
C9757 VDD.t524 Vbias 0.0169f
C9758 VDD.t864 Vbias 0.0169f
C9759 VDD.n1388 Vbias 0.07902f
C9760 VDD.t691 Vbias 0.0169f
C9761 VDD.t688 Vbias 0.0169f
C9762 VDD.n1389 Vbias 0.07902f
C9763 VDD.n1390 Vbias 0.03023f
C9764 VDD.n1391 Vbias 0.01699f
C9765 VDD.n1392 Vbias 0.03902f
C9766 VDD.n1393 Vbias 0.03694f
C9767 VDD.n1394 Vbias 0.0216f
C9768 VDD.n1395 Vbias 0.01836f
C9769 VDD.t418 Vbias 0.46278f
C9770 VDD.n1396 Vbias 0.03694f
C9771 VDD.n1397 Vbias 0.03694f
C9772 VDD.n1398 Vbias 0.06648f
C9773 VDD.n1399 Vbias 0.03639f
C9774 VDD.t360 Vbias 0.46278f
C9775 VDD.n1400 Vbias 0.03694f
C9776 VDD.n1401 Vbias 0.03694f
C9777 VDD.n1402 Vbias 0.0216f
C9778 VDD.n1403 Vbias 0.01836f
C9779 VDD.t419 Vbias 0.017f
C9780 VDD.n1404 Vbias 0.05322f
C9781 VDD.n1405 Vbias 0.01309f
C9782 VDD.n1406 Vbias 0.01699f
C9783 VDD.n1407 Vbias 0.03902f
C9784 VDD.n1408 Vbias 0.03694f
C9785 VDD.n1409 Vbias 0.0216f
C9786 VDD.n1410 Vbias 0.01836f
C9787 VDD.n1411 Vbias 0.03639f
C9788 VDD.t504 Vbias 0.46278f
C9789 VDD.n1412 Vbias 0.03694f
C9790 VDD.n1413 Vbias 0.03694f
C9791 VDD.n1414 Vbias 0.0216f
C9792 VDD.n1415 Vbias 0.01836f
C9793 VDD.t680 Vbias 0.0169f
C9794 VDD.t506 Vbias 0.0169f
C9795 VDD.n1416 Vbias 0.07902f
C9796 VDD.t361 Vbias 0.0169f
C9797 VDD.t505 Vbias 0.0169f
C9798 VDD.n1417 Vbias 0.07902f
C9799 VDD.n1418 Vbias 0.03023f
C9800 VDD.n1419 Vbias 0.01699f
C9801 VDD.n1420 Vbias 0.03902f
C9802 VDD.n1421 Vbias 0.03694f
C9803 VDD.n1422 Vbias 0.0216f
C9804 VDD.n1423 Vbias 0.01836f
C9805 VDD.n1424 Vbias 0.03639f
C9806 VDD.t436 Vbias 0.46278f
C9807 VDD.n1425 Vbias 0.03694f
C9808 VDD.n1426 Vbias 0.03694f
C9809 VDD.n1427 Vbias 0.0216f
C9810 VDD.n1428 Vbias 0.01836f
C9811 VDD.t535 Vbias 0.017f
C9812 VDD.t437 Vbias 0.017f
C9813 VDD.n1429 Vbias 0.09713f
C9814 VDD.n1430 Vbias 0.01914f
C9815 VDD.n1431 Vbias 0.03902f
C9816 VDD.n1432 Vbias 0.03694f
C9817 VDD.n1433 Vbias 0.0216f
C9818 VDD.n1434 Vbias 0.01836f
C9819 VDD.n1435 Vbias 0.03639f
C9820 VDD.t887 Vbias 0.46278f
C9821 VDD.n1436 Vbias 0.03694f
C9822 VDD.n1437 Vbias 0.03694f
C9823 VDD.n1438 Vbias 0.0216f
C9824 VDD.n1439 Vbias 0.01836f
C9825 VDD.n1440 Vbias 0.02305f
C9826 VDD.n1441 Vbias 0.03902f
C9827 VDD.n1442 Vbias 0.03694f
C9828 VDD.n1443 Vbias 0.0216f
C9829 VDD.n1444 Vbias 0.01836f
C9830 VDD.n1445 Vbias 0.03639f
C9831 VDD.t403 Vbias 0.46278f
C9832 VDD.n1446 Vbias 0.03694f
C9833 VDD.n1447 Vbias 0.03694f
C9834 VDD.n1448 Vbias 0.0216f
C9835 VDD.n1449 Vbias 0.01836f
C9836 VDD.t996 Vbias 0.0169f
C9837 VDD.t901 Vbias 0.0169f
C9838 VDD.n1450 Vbias 0.07902f
C9839 VDD.t888 Vbias 0.0169f
C9840 VDD.t404 Vbias 0.0169f
C9841 VDD.n1451 Vbias 0.07902f
C9842 VDD.n1452 Vbias 0.03023f
C9843 VDD.n1453 Vbias 0.01699f
C9844 VDD.n1454 Vbias 0.03902f
C9845 VDD.n1455 Vbias 0.03694f
C9846 VDD.n1456 Vbias 0.0216f
C9847 VDD.n1457 Vbias 0.01836f
C9848 VDD.n1458 Vbias 0.01836f
C9849 VDD.n1459 Vbias 0.03639f
C9850 VDD.n1460 Vbias 0.50118f
C9851 VDD.n1461 Vbias 0.03639f
C9852 VDD.n1462 Vbias 0.03694f
C9853 VDD.n1463 Vbias 0.04583f
C9854 VDD.n1464 Vbias 0.03902f
C9855 VDD.n1465 Vbias 0.01836f
C9856 VDD.n1466 Vbias 0.03639f
C9857 VDD.n1467 Vbias 0.37318f
C9858 VDD.n1468 Vbias 0.01836f
C9859 VDD.n1469 Vbias 0.03639f
C9860 VDD.n1470 Vbias 0.37318f
C9861 VDD.n1471 Vbias 0.03639f
C9862 VDD.n1472 Vbias 0.03694f
C9863 VDD.n1473 Vbias 0.04583f
C9864 VDD.n1474 Vbias 0.03902f
C9865 VDD.n1475 Vbias 0.01836f
C9866 VDD.n1476 Vbias 0.03639f
C9867 VDD.n1477 Vbias 0.37318f
C9868 VDD.n1478 Vbias 0.01836f
C9869 VDD.n1479 Vbias 0.03639f
C9870 VDD.n1480 Vbias 0.37318f
C9871 VDD.n1481 Vbias 0.03639f
C9872 VDD.n1482 Vbias 0.03694f
C9873 VDD.n1483 Vbias 0.04583f
C9874 VDD.n1484 Vbias 0.03902f
C9875 VDD.n1485 Vbias 0.01836f
C9876 VDD.n1486 Vbias 0.03639f
C9877 VDD.n1487 Vbias 0.50118f
C9878 VDD.n1488 Vbias 0.01836f
C9879 VDD.n1489 Vbias 0.03639f
C9880 VDD.n1490 Vbias 0.50118f
C9881 VDD.n1491 Vbias 0.03639f
C9882 VDD.n1492 Vbias 0.03694f
C9883 VDD.n1493 Vbias 0.04583f
C9884 VDD.n1494 Vbias 0.03902f
C9885 VDD.n1495 Vbias 0.01836f
C9886 VDD.n1496 Vbias 0.03639f
C9887 VDD.n1497 Vbias 0.37318f
C9888 VDD.n1498 Vbias 0.01836f
C9889 VDD.n1499 Vbias 0.03639f
C9890 VDD.n1500 Vbias 0.37318f
C9891 VDD.n1501 Vbias 0.03639f
C9892 VDD.n1502 Vbias 0.03694f
C9893 VDD.n1503 Vbias 0.04583f
C9894 VDD.n1504 Vbias 0.03902f
C9895 VDD.n1505 Vbias 0.01836f
C9896 VDD.n1506 Vbias 0.03639f
C9897 VDD.n1507 Vbias 0.50118f
C9898 VDD.n1508 Vbias 0.50118f
C9899 VDD.n1509 Vbias 0.03639f
C9900 VDD.n1510 Vbias 0.01999f
C9901 VDD.n1511 Vbias 0.0216f
C9902 VDD.n1512 Vbias 0.01999f
C9903 VDD.n1513 Vbias 0.03639f
C9904 VDD.n1514 Vbias 0.50118f
C9905 VDD.n1515 Vbias 0.01836f
C9906 VDD.n1516 Vbias 0.03639f
C9907 VDD.n1517 Vbias 0.50118f
C9908 VDD.n1518 Vbias 0.03639f
C9909 VDD.n1519 Vbias 0.03694f
C9910 VDD.n1520 Vbias 0.04583f
C9911 VDD.n1521 Vbias 0.03902f
C9912 VDD.n1522 Vbias 0.01836f
C9913 VDD.n1523 Vbias 0.03639f
C9914 VDD.n1524 Vbias 0.37318f
C9915 VDD.n1525 Vbias 0.01836f
C9916 VDD.n1526 Vbias 0.03639f
C9917 VDD.n1527 Vbias 0.37318f
C9918 VDD.n1528 Vbias 0.03639f
C9919 VDD.n1529 Vbias 0.03694f
C9920 VDD.n1530 Vbias 0.04583f
C9921 VDD.n1531 Vbias 0.03902f
C9922 VDD.n1532 Vbias 0.01836f
C9923 VDD.n1533 Vbias 0.03639f
C9924 VDD.n1534 Vbias 0.37318f
C9925 VDD.n1535 Vbias 0.01836f
C9926 VDD.n1536 Vbias 0.03639f
C9927 VDD.n1537 Vbias 0.37318f
C9928 VDD.n1538 Vbias 0.03639f
C9929 VDD.n1539 Vbias 0.03694f
C9930 VDD.n1540 Vbias 0.04583f
C9931 VDD.n1541 Vbias 0.03902f
C9932 VDD.n1542 Vbias 0.01836f
C9933 VDD.n1543 Vbias 0.03639f
C9934 VDD.n1544 Vbias 0.50118f
C9935 VDD.n1545 Vbias 0.01836f
C9936 VDD.n1546 Vbias 0.03639f
C9937 VDD.n1547 Vbias 0.50118f
C9938 VDD.n1548 Vbias 0.03639f
C9939 VDD.n1549 Vbias 0.03694f
C9940 VDD.n1550 Vbias 0.04583f
C9941 VDD.n1551 Vbias 0.03902f
C9942 VDD.n1552 Vbias 0.01836f
C9943 VDD.n1553 Vbias 0.03639f
C9944 VDD.n1554 Vbias 0.37318f
C9945 VDD.n1555 Vbias 0.01836f
C9946 VDD.n1556 Vbias 0.03639f
C9947 VDD.n1557 Vbias 0.37318f
C9948 VDD.n1558 Vbias 0.03639f
C9949 VDD.n1559 Vbias 0.03694f
C9950 VDD.n1560 Vbias 0.04583f
C9951 VDD.n1561 Vbias 0.03902f
C9952 VDD.n1562 Vbias 0.01836f
C9953 VDD.n1563 Vbias 0.03639f
C9954 VDD.n1564 Vbias 0.37318f
C9955 VDD.n1565 Vbias 0.01836f
C9956 VDD.n1566 Vbias 0.03639f
C9957 VDD.n1567 Vbias 0.37318f
C9958 VDD.n1568 Vbias 0.03639f
C9959 VDD.n1569 Vbias 0.03694f
C9960 VDD.n1570 Vbias 0.04583f
C9961 VDD.n1571 Vbias 0.03902f
C9962 VDD.n1572 Vbias 0.01836f
C9963 VDD.n1573 Vbias 0.03639f
C9964 VDD.n1574 Vbias 0.50118f
C9965 VDD.n1575 Vbias 0.50118f
C9966 VDD.n1576 Vbias 0.03639f
C9967 VDD.n1577 Vbias 0.01999f
C9968 VDD.n1578 Vbias 0.06648f
C9969 VDD.n1579 Vbias 0.01309f
C9970 VDD.n1580 Vbias 0.07184f
C9971 VDD.n1581 Vbias 0.30746f
C9972 VDD.t940 Vbias 0.017f
C9973 VDD.n1582 Vbias 0.01999f
C9974 VDD.n1583 Vbias 0.03694f
C9975 VDD.n1584 Vbias 0.0216f
C9976 VDD.n1585 Vbias 0.03694f
C9977 VDD.n1586 Vbias 0.45845f
C9978 VDD.t939 Vbias 0.54191f
C9979 VDD.n1588 Vbias 0.03639f
C9980 VDD.t289 Vbias 0.46278f
C9981 VDD.n1589 Vbias 0.03694f
C9982 VDD.n1590 Vbias 0.03694f
C9983 VDD.n1591 Vbias 0.0216f
C9984 VDD.n1592 Vbias 0.01836f
C9985 VDD.t389 Vbias 0.017f
C9986 VDD.t290 Vbias 0.017f
C9987 VDD.n1593 Vbias 0.09713f
C9988 VDD.n1594 Vbias 0.01914f
C9989 VDD.n1595 Vbias 0.03902f
C9990 VDD.n1596 Vbias 0.03694f
C9991 VDD.n1597 Vbias 0.0216f
C9992 VDD.n1598 Vbias 0.01836f
C9993 VDD.n1599 Vbias 0.03639f
C9994 VDD.t843 Vbias 0.46278f
C9995 VDD.n1600 Vbias 0.03694f
C9996 VDD.n1601 Vbias 0.03694f
C9997 VDD.n1602 Vbias 0.0216f
C9998 VDD.n1603 Vbias 0.01836f
C9999 VDD.n1604 Vbias 0.02305f
C10000 VDD.n1605 Vbias 0.03902f
C10001 VDD.n1606 Vbias 0.03694f
C10002 VDD.n1607 Vbias 0.0216f
C10003 VDD.n1608 Vbias 0.01836f
C10004 VDD.n1609 Vbias 0.03639f
C10005 VDD.t131 Vbias 0.46278f
C10006 VDD.n1610 Vbias 0.03694f
C10007 VDD.n1611 Vbias 0.03694f
C10008 VDD.n1612 Vbias 0.0216f
C10009 VDD.n1613 Vbias 0.01836f
C10010 VDD.t844 Vbias 0.0169f
C10011 VDD.t132 Vbias 0.0169f
C10012 VDD.n1614 Vbias 0.07902f
C10013 VDD.t917 Vbias 0.0169f
C10014 VDD.t135 Vbias 0.0169f
C10015 VDD.n1615 Vbias 0.07902f
C10016 VDD.n1616 Vbias 0.03023f
C10017 VDD.n1617 Vbias 0.01699f
C10018 VDD.n1618 Vbias 0.03902f
C10019 VDD.n1619 Vbias 0.03694f
C10020 VDD.n1620 Vbias 0.0216f
C10021 VDD.n1621 Vbias 0.01836f
C10022 VDD.n1622 Vbias 0.03639f
C10023 VDD.t580 Vbias 0.46278f
C10024 VDD.n1623 Vbias 0.03694f
C10025 VDD.n1624 Vbias 0.03694f
C10026 VDD.n1625 Vbias 0.0216f
C10027 VDD.n1626 Vbias 0.01836f
C10028 VDD.t581 Vbias 0.017f
C10029 VDD.t654 Vbias 0.017f
C10030 VDD.n1627 Vbias 0.09713f
C10031 VDD.n1628 Vbias 0.01914f
C10032 VDD.n1629 Vbias 0.03902f
C10033 VDD.n1630 Vbias 0.03694f
C10034 VDD.n1631 Vbias 0.0216f
C10035 VDD.n1632 Vbias 0.01836f
C10036 VDD.n1633 Vbias 0.03639f
C10037 VDD.t593 Vbias 0.46278f
C10038 VDD.n1634 Vbias 0.03694f
C10039 VDD.n1635 Vbias 0.03694f
C10040 VDD.n1636 Vbias 0.0216f
C10041 VDD.n1637 Vbias 0.01836f
C10042 VDD.n1638 Vbias 0.02305f
C10043 VDD.n1639 Vbias 0.03902f
C10044 VDD.n1640 Vbias 0.03694f
C10045 VDD.n1641 Vbias 0.0216f
C10046 VDD.n1642 Vbias 0.01836f
C10047 VDD.n1643 Vbias 0.03639f
C10048 VDD.t371 Vbias 0.46278f
C10049 VDD.n1644 Vbias 0.03694f
C10050 VDD.n1645 Vbias 0.03694f
C10051 VDD.n1646 Vbias 0.0216f
C10052 VDD.n1647 Vbias 0.01836f
C10053 VDD.t681 Vbias 0.0169f
C10054 VDD.t400 Vbias 0.0169f
C10055 VDD.n1648 Vbias 0.07902f
C10056 VDD.t594 Vbias 0.0169f
C10057 VDD.t372 Vbias 0.0169f
C10058 VDD.n1649 Vbias 0.07902f
C10059 VDD.n1650 Vbias 0.03023f
C10060 VDD.n1651 Vbias 0.01699f
C10061 VDD.n1652 Vbias 0.03902f
C10062 VDD.n1653 Vbias 0.03694f
C10063 VDD.n1654 Vbias 0.0216f
C10064 VDD.n1655 Vbias 0.01836f
C10065 VDD.t133 Vbias 0.46278f
C10066 VDD.n1656 Vbias 0.03694f
C10067 VDD.n1657 Vbias 0.03694f
C10068 VDD.n1658 Vbias 0.06648f
C10069 VDD.n1659 Vbias 0.03639f
C10070 VDD.t369 Vbias 0.46278f
C10071 VDD.n1660 Vbias 0.03694f
C10072 VDD.n1661 Vbias 0.03694f
C10073 VDD.n1662 Vbias 0.0216f
C10074 VDD.n1663 Vbias 0.01836f
C10075 VDD.t134 Vbias 0.017f
C10076 VDD.n1664 Vbias 0.05322f
C10077 VDD.n1665 Vbias 0.01309f
C10078 VDD.n1666 Vbias 0.01699f
C10079 VDD.n1667 Vbias 0.03902f
C10080 VDD.n1668 Vbias 0.03694f
C10081 VDD.n1669 Vbias 0.0216f
C10082 VDD.n1670 Vbias 0.01836f
C10083 VDD.n1671 Vbias 0.03639f
C10084 VDD.t670 Vbias 0.46278f
C10085 VDD.n1672 Vbias 0.03694f
C10086 VDD.n1673 Vbias 0.03694f
C10087 VDD.n1674 Vbias 0.0216f
C10088 VDD.n1675 Vbias 0.01836f
C10089 VDD.t370 Vbias 0.0169f
C10090 VDD.t671 Vbias 0.0169f
C10091 VDD.n1676 Vbias 0.07902f
C10092 VDD.t401 Vbias 0.0169f
C10093 VDD.t672 Vbias 0.0169f
C10094 VDD.n1677 Vbias 0.07902f
C10095 VDD.n1678 Vbias 0.03023f
C10096 VDD.n1679 Vbias 0.01699f
C10097 VDD.n1680 Vbias 0.03902f
C10098 VDD.n1681 Vbias 0.03694f
C10099 VDD.n1682 Vbias 0.0216f
C10100 VDD.n1683 Vbias 0.01836f
C10101 VDD.n1684 Vbias 0.03639f
C10102 VDD.t293 Vbias 0.46278f
C10103 VDD.n1685 Vbias 0.03694f
C10104 VDD.n1686 Vbias 0.03694f
C10105 VDD.n1687 Vbias 0.0216f
C10106 VDD.n1688 Vbias 0.01836f
C10107 VDD.t294 Vbias 0.017f
C10108 VDD.t483 Vbias 0.017f
C10109 VDD.n1689 Vbias 0.09713f
C10110 VDD.n1690 Vbias 0.01914f
C10111 VDD.n1691 Vbias 0.03902f
C10112 VDD.n1692 Vbias 0.03694f
C10113 VDD.n1693 Vbias 0.0216f
C10114 VDD.n1694 Vbias 0.01836f
C10115 VDD.n1695 Vbias 0.03639f
C10116 VDD.t587 Vbias 0.46278f
C10117 VDD.n1696 Vbias 0.03694f
C10118 VDD.n1697 Vbias 0.03694f
C10119 VDD.n1698 Vbias 0.0216f
C10120 VDD.n1699 Vbias 0.01836f
C10121 VDD.n1700 Vbias 0.02305f
C10122 VDD.n1701 Vbias 0.03902f
C10123 VDD.n1702 Vbias 0.03694f
C10124 VDD.n1703 Vbias 0.0216f
C10125 VDD.n1704 Vbias 0.01836f
C10126 VDD.n1705 Vbias 0.03639f
C10127 VDD.t5 Vbias 0.46278f
C10128 VDD.n1706 Vbias 0.03694f
C10129 VDD.n1707 Vbias 0.03694f
C10130 VDD.n1708 Vbias 0.0216f
C10131 VDD.n1709 Vbias 0.01836f
C10132 VDD.t588 Vbias 0.0169f
C10133 VDD.t425 Vbias 0.0169f
C10134 VDD.n1710 Vbias 0.07902f
C10135 VDD.t963 Vbias 0.0169f
C10136 VDD.t6 Vbias 0.0169f
C10137 VDD.n1711 Vbias 0.07902f
C10138 VDD.n1712 Vbias 0.03023f
C10139 VDD.n1713 Vbias 0.01699f
C10140 VDD.n1714 Vbias 0.03902f
C10141 VDD.n1715 Vbias 0.03694f
C10142 VDD.n1716 Vbias 0.0216f
C10143 VDD.n1717 Vbias 0.01836f
C10144 VDD.n1718 Vbias 0.01836f
C10145 VDD.n1719 Vbias 0.03639f
C10146 VDD.n1720 Vbias 0.50118f
C10147 VDD.n1721 Vbias 0.03639f
C10148 VDD.n1722 Vbias 0.03694f
C10149 VDD.n1723 Vbias 0.04583f
C10150 VDD.n1724 Vbias 0.03902f
C10151 VDD.n1725 Vbias 0.01836f
C10152 VDD.n1726 Vbias 0.03639f
C10153 VDD.n1727 Vbias 0.37318f
C10154 VDD.n1728 Vbias 0.01836f
C10155 VDD.n1729 Vbias 0.03639f
C10156 VDD.n1730 Vbias 0.37318f
C10157 VDD.n1731 Vbias 0.03639f
C10158 VDD.n1732 Vbias 0.03694f
C10159 VDD.n1733 Vbias 0.04583f
C10160 VDD.n1734 Vbias 0.03902f
C10161 VDD.n1735 Vbias 0.01836f
C10162 VDD.n1736 Vbias 0.03639f
C10163 VDD.n1737 Vbias 0.37318f
C10164 VDD.n1738 Vbias 0.01836f
C10165 VDD.n1739 Vbias 0.03639f
C10166 VDD.n1740 Vbias 0.37318f
C10167 VDD.n1741 Vbias 0.03639f
C10168 VDD.n1742 Vbias 0.03694f
C10169 VDD.n1743 Vbias 0.04583f
C10170 VDD.n1744 Vbias 0.03902f
C10171 VDD.n1745 Vbias 0.01836f
C10172 VDD.n1746 Vbias 0.03639f
C10173 VDD.n1747 Vbias 0.50118f
C10174 VDD.n1748 Vbias 0.01836f
C10175 VDD.n1749 Vbias 0.03639f
C10176 VDD.n1750 Vbias 0.50118f
C10177 VDD.n1751 Vbias 0.03639f
C10178 VDD.n1752 Vbias 0.03694f
C10179 VDD.n1753 Vbias 0.04583f
C10180 VDD.n1754 Vbias 0.03902f
C10181 VDD.n1755 Vbias 0.01836f
C10182 VDD.n1756 Vbias 0.03639f
C10183 VDD.n1757 Vbias 0.37318f
C10184 VDD.n1758 Vbias 0.01836f
C10185 VDD.n1759 Vbias 0.03639f
C10186 VDD.n1760 Vbias 0.37318f
C10187 VDD.n1761 Vbias 0.03639f
C10188 VDD.n1762 Vbias 0.03694f
C10189 VDD.n1763 Vbias 0.04583f
C10190 VDD.n1764 Vbias 0.03902f
C10191 VDD.n1765 Vbias 0.01836f
C10192 VDD.n1766 Vbias 0.03639f
C10193 VDD.n1767 Vbias 0.50118f
C10194 VDD.n1768 Vbias 0.50118f
C10195 VDD.n1769 Vbias 0.03639f
C10196 VDD.n1770 Vbias 0.01999f
C10197 VDD.n1771 Vbias 0.0216f
C10198 VDD.n1772 Vbias 0.01999f
C10199 VDD.n1773 Vbias 0.03639f
C10200 VDD.n1774 Vbias 0.50118f
C10201 VDD.n1775 Vbias 0.01836f
C10202 VDD.n1776 Vbias 0.03639f
C10203 VDD.n1777 Vbias 0.50118f
C10204 VDD.n1778 Vbias 0.03639f
C10205 VDD.n1779 Vbias 0.03694f
C10206 VDD.n1780 Vbias 0.04583f
C10207 VDD.n1781 Vbias 0.03902f
C10208 VDD.n1782 Vbias 0.01836f
C10209 VDD.n1783 Vbias 0.03639f
C10210 VDD.n1784 Vbias 0.37318f
C10211 VDD.n1785 Vbias 0.01836f
C10212 VDD.n1786 Vbias 0.03639f
C10213 VDD.n1787 Vbias 0.37318f
C10214 VDD.n1788 Vbias 0.03639f
C10215 VDD.n1789 Vbias 0.03694f
C10216 VDD.n1790 Vbias 0.04583f
C10217 VDD.n1791 Vbias 0.03902f
C10218 VDD.n1792 Vbias 0.01836f
C10219 VDD.n1793 Vbias 0.03639f
C10220 VDD.n1794 Vbias 0.37318f
C10221 VDD.n1795 Vbias 0.01836f
C10222 VDD.n1796 Vbias 0.03639f
C10223 VDD.n1797 Vbias 0.37318f
C10224 VDD.n1798 Vbias 0.03639f
C10225 VDD.n1799 Vbias 0.03694f
C10226 VDD.n1800 Vbias 0.04583f
C10227 VDD.n1801 Vbias 0.03902f
C10228 VDD.n1802 Vbias 0.01836f
C10229 VDD.n1803 Vbias 0.03639f
C10230 VDD.n1804 Vbias 0.50118f
C10231 VDD.n1805 Vbias 0.01836f
C10232 VDD.n1806 Vbias 0.03639f
C10233 VDD.n1807 Vbias 0.50118f
C10234 VDD.n1808 Vbias 0.03639f
C10235 VDD.n1809 Vbias 0.03694f
C10236 VDD.n1810 Vbias 0.04583f
C10237 VDD.n1811 Vbias 0.03902f
C10238 VDD.n1812 Vbias 0.01836f
C10239 VDD.n1813 Vbias 0.03639f
C10240 VDD.n1814 Vbias 0.37318f
C10241 VDD.n1815 Vbias 0.01836f
C10242 VDD.n1816 Vbias 0.03639f
C10243 VDD.n1817 Vbias 0.37318f
C10244 VDD.n1818 Vbias 0.03639f
C10245 VDD.n1819 Vbias 0.03694f
C10246 VDD.n1820 Vbias 0.04583f
C10247 VDD.n1821 Vbias 0.03902f
C10248 VDD.n1822 Vbias 0.01836f
C10249 VDD.n1823 Vbias 0.03639f
C10250 VDD.n1824 Vbias 0.37318f
C10251 VDD.n1825 Vbias 0.01836f
C10252 VDD.n1826 Vbias 0.03639f
C10253 VDD.n1827 Vbias 0.37318f
C10254 VDD.n1828 Vbias 0.03639f
C10255 VDD.n1829 Vbias 0.03694f
C10256 VDD.n1830 Vbias 0.04583f
C10257 VDD.n1831 Vbias 0.03902f
C10258 VDD.n1832 Vbias 0.01836f
C10259 VDD.n1833 Vbias 0.03639f
C10260 VDD.n1834 Vbias 0.50118f
C10261 VDD.n1835 Vbias 0.50118f
C10262 VDD.n1836 Vbias 0.03639f
C10263 VDD.n1837 Vbias 0.01999f
C10264 VDD.n1838 Vbias 0.06648f
C10265 VDD.n1839 Vbias 0.01309f
C10266 VDD.n1840 Vbias 0.07184f
C10267 VDD.n1841 Vbias 0.23842f
C10268 VDD.t914 Vbias 0.017f
C10269 VDD.n1842 Vbias 0.01999f
C10270 VDD.n1843 Vbias 0.03694f
C10271 VDD.n1844 Vbias 0.0216f
C10272 VDD.n1845 Vbias 0.03694f
C10273 VDD.n1846 Vbias 0.45845f
C10274 VDD.t913 Vbias 0.54191f
C10275 VDD.n1848 Vbias 0.03639f
C10276 VDD.t29 Vbias 0.46278f
C10277 VDD.n1849 Vbias 0.03694f
C10278 VDD.n1850 Vbias 0.03694f
C10279 VDD.n1851 Vbias 0.0216f
C10280 VDD.n1852 Vbias 0.01836f
C10281 VDD.t785 Vbias 0.017f
C10282 VDD.t30 Vbias 0.017f
C10283 VDD.n1853 Vbias 0.09713f
C10284 VDD.n1854 Vbias 0.01914f
C10285 VDD.n1855 Vbias 0.03902f
C10286 VDD.n1856 Vbias 0.03694f
C10287 VDD.n1857 Vbias 0.0216f
C10288 VDD.n1858 Vbias 0.01836f
C10289 VDD.n1859 Vbias 0.03639f
C10290 VDD.t455 Vbias 0.46278f
C10291 VDD.n1860 Vbias 0.03694f
C10292 VDD.n1861 Vbias 0.03694f
C10293 VDD.n1862 Vbias 0.0216f
C10294 VDD.n1863 Vbias 0.01836f
C10295 VDD.n1864 Vbias 0.02305f
C10296 VDD.n1865 Vbias 0.03902f
C10297 VDD.n1866 Vbias 0.03694f
C10298 VDD.n1867 Vbias 0.0216f
C10299 VDD.n1868 Vbias 0.01836f
C10300 VDD.n1869 Vbias 0.03639f
C10301 VDD.t1020 Vbias 0.46278f
C10302 VDD.n1870 Vbias 0.03694f
C10303 VDD.n1871 Vbias 0.03694f
C10304 VDD.n1872 Vbias 0.0216f
C10305 VDD.n1873 Vbias 0.01836f
C10306 VDD.t902 Vbias 0.0169f
C10307 VDD.t1021 Vbias 0.0169f
C10308 VDD.n1874 Vbias 0.07902f
C10309 VDD.t456 Vbias 0.0169f
C10310 VDD.t1067 Vbias 0.0169f
C10311 VDD.n1875 Vbias 0.07902f
C10312 VDD.n1876 Vbias 0.03023f
C10313 VDD.n1877 Vbias 0.01699f
C10314 VDD.n1878 Vbias 0.03902f
C10315 VDD.n1879 Vbias 0.03694f
C10316 VDD.n1880 Vbias 0.0216f
C10317 VDD.n1881 Vbias 0.01836f
C10318 VDD.n1882 Vbias 0.03639f
C10319 VDD.t91 Vbias 0.46278f
C10320 VDD.n1883 Vbias 0.03694f
C10321 VDD.n1884 Vbias 0.03694f
C10322 VDD.n1885 Vbias 0.0216f
C10323 VDD.n1886 Vbias 0.01836f
C10324 VDD.t92 Vbias 0.017f
C10325 VDD.t723 Vbias 0.017f
C10326 VDD.n1887 Vbias 0.09633f
C10327 VDD.n1888 Vbias 0.04493f
C10328 VDD.n1890 Vbias 0.03902f
C10329 VDD.n1891 Vbias 0.03694f
C10330 VDD.n1892 Vbias 0.0216f
C10331 VDD.n1893 Vbias 0.01836f
C10332 VDD.n1894 Vbias 0.03639f
C10333 VDD.t228 Vbias 0.46278f
C10334 VDD.n1895 Vbias 0.03694f
C10335 VDD.n1896 Vbias 0.03694f
C10336 VDD.n1897 Vbias 0.0216f
C10337 VDD.n1898 Vbias 0.01836f
C10338 VDD.n1899 Vbias 0.03902f
C10339 VDD.n1900 Vbias 0.03694f
C10340 VDD.n1901 Vbias 0.07027f
C10341 VDD.t229 Vbias 0.0169f
C10342 VDD.t929 Vbias 0.0169f
C10343 VDD.n1902 Vbias 0.07902f
C10344 VDD.t261 Vbias 0.0169f
C10345 VDD.t424 Vbias 0.0169f
C10346 VDD.n1903 Vbias 0.07902f
C10347 VDD.n1904 Vbias 0.03902f
C10348 VDD.n1905 Vbias 0.03694f
C10349 VDD.n1906 Vbias 0.03902f
C10350 VDD.n1907 Vbias 0.03639f
C10351 VDD.n1908 Vbias 0.03639f
C10352 VDD.n1909 Vbias 0.03694f
C10353 VDD.n1910 Vbias 0.0216f
C10354 VDD.n1911 Vbias 0.01836f
C10355 VDD.n1912 Vbias 0.03639f
C10356 VDD.n1913 Vbias 0.01836f
C10357 VDD.n1914 Vbias 0.03639f
C10358 VDD.n1915 Vbias 0.37318f
C10359 VDD.n1916 Vbias 0.37318f
C10360 VDD.n1917 Vbias 0.01836f
C10361 VDD.n1918 Vbias 0.01836f
C10362 VDD.n1919 Vbias 0.0216f
C10363 VDD.n1920 Vbias 0.03694f
C10364 VDD.t1074 Vbias 0.46278f
C10365 VDD.n1921 Vbias 0.03694f
C10366 VDD.n1922 Vbias 0.03694f
C10367 VDD.n1923 Vbias 0.06648f
C10368 VDD.n1924 Vbias 0.03639f
C10369 VDD.t305 Vbias 0.46278f
C10370 VDD.n1925 Vbias 0.03694f
C10371 VDD.n1926 Vbias 0.03694f
C10372 VDD.n1927 Vbias 0.0216f
C10373 VDD.n1928 Vbias 0.01836f
C10374 VDD.t1075 Vbias 0.017f
C10375 VDD.n1929 Vbias 0.05322f
C10376 VDD.n1930 Vbias 0.01309f
C10377 VDD.n1931 Vbias 0.01699f
C10378 VDD.n1932 Vbias 0.03902f
C10379 VDD.n1933 Vbias 0.03694f
C10380 VDD.n1934 Vbias 0.0216f
C10381 VDD.n1935 Vbias 0.01836f
C10382 VDD.n1936 Vbias 0.03639f
C10383 VDD.t969 Vbias 0.46278f
C10384 VDD.n1937 Vbias 0.03694f
C10385 VDD.n1938 Vbias 0.03694f
C10386 VDD.n1939 Vbias 0.0216f
C10387 VDD.n1940 Vbias 0.01836f
C10388 VDD.t306 Vbias 0.0169f
C10389 VDD.t970 Vbias 0.0169f
C10390 VDD.n1941 Vbias 0.07902f
C10391 VDD.t495 Vbias 0.0169f
C10392 VDD.t971 Vbias 0.0169f
C10393 VDD.n1942 Vbias 0.07902f
C10394 VDD.n1943 Vbias 0.03023f
C10395 VDD.n1944 Vbias 0.01699f
C10396 VDD.n1945 Vbias 0.03902f
C10397 VDD.n1946 Vbias 0.03694f
C10398 VDD.n1947 Vbias 0.0216f
C10399 VDD.n1948 Vbias 0.01836f
C10400 VDD.n1949 Vbias 0.03639f
C10401 VDD.t113 Vbias 0.46278f
C10402 VDD.n1950 Vbias 0.03694f
C10403 VDD.n1951 Vbias 0.03694f
C10404 VDD.n1952 Vbias 0.0216f
C10405 VDD.n1953 Vbias 0.01836f
C10406 VDD.t114 Vbias 0.017f
C10407 VDD.t747 Vbias 0.017f
C10408 VDD.n1954 Vbias 0.09713f
C10409 VDD.n1955 Vbias 0.01914f
C10410 VDD.n1956 Vbias 0.03902f
C10411 VDD.n1957 Vbias 0.03694f
C10412 VDD.n1958 Vbias 0.0216f
C10413 VDD.n1959 Vbias 0.01836f
C10414 VDD.n1960 Vbias 0.03639f
C10415 VDD.t897 Vbias 0.46278f
C10416 VDD.n1961 Vbias 0.03694f
C10417 VDD.n1962 Vbias 0.03694f
C10418 VDD.n1963 Vbias 0.0216f
C10419 VDD.n1964 Vbias 0.01836f
C10420 VDD.n1965 Vbias 0.02305f
C10421 VDD.n1966 Vbias 0.03902f
C10422 VDD.n1967 Vbias 0.03694f
C10423 VDD.n1968 Vbias 0.0216f
C10424 VDD.n1969 Vbias 0.01836f
C10425 VDD.n1970 Vbias 0.03639f
C10426 VDD.t480 Vbias 0.46278f
C10427 VDD.n1971 Vbias 0.03694f
C10428 VDD.n1972 Vbias 0.03694f
C10429 VDD.n1973 Vbias 0.0216f
C10430 VDD.n1974 Vbias 0.01836f
C10431 VDD.t927 Vbias 0.0169f
C10432 VDD.t481 Vbias 0.0169f
C10433 VDD.n1975 Vbias 0.07902f
C10434 VDD.t898 Vbias 0.0169f
C10435 VDD.t536 Vbias 0.0169f
C10436 VDD.n1976 Vbias 0.07902f
C10437 VDD.n1977 Vbias 0.03023f
C10438 VDD.t3 Vbias 0.017f
C10439 VDD.n1978 Vbias 0.01999f
C10440 VDD.n1979 Vbias 0.03694f
C10441 VDD.n1980 Vbias 0.0216f
C10442 VDD.n1981 Vbias 0.03694f
C10443 VDD.n1982 Vbias 0.45845f
C10444 VDD.t2 Vbias 0.54191f
C10445 VDD.n1984 Vbias 0.03639f
C10446 VDD.t51 Vbias 0.46278f
C10447 VDD.n1985 Vbias 0.03694f
C10448 VDD.n1986 Vbias 0.03694f
C10449 VDD.n1987 Vbias 0.0216f
C10450 VDD.n1988 Vbias 0.01836f
C10451 VDD.t801 Vbias 0.017f
C10452 VDD.t52 Vbias 0.017f
C10453 VDD.n1989 Vbias 0.09713f
C10454 VDD.n1990 Vbias 0.01914f
C10455 VDD.n1991 Vbias 0.03902f
C10456 VDD.n1992 Vbias 0.03694f
C10457 VDD.n1993 Vbias 0.0216f
C10458 VDD.n1994 Vbias 0.01836f
C10459 VDD.n1995 Vbias 0.03639f
C10460 VDD.t646 Vbias 0.46278f
C10461 VDD.n1996 Vbias 0.03694f
C10462 VDD.n1997 Vbias 0.03694f
C10463 VDD.n1998 Vbias 0.0216f
C10464 VDD.n1999 Vbias 0.01836f
C10465 VDD.n2000 Vbias 0.02305f
C10466 VDD.n2001 Vbias 0.03902f
C10467 VDD.n2002 Vbias 0.03694f
C10468 VDD.n2003 Vbias 0.0216f
C10469 VDD.n2004 Vbias 0.01836f
C10470 VDD.n2005 Vbias 0.03639f
C10471 VDD.t1016 Vbias 0.46278f
C10472 VDD.n2006 Vbias 0.03694f
C10473 VDD.n2007 Vbias 0.03694f
C10474 VDD.n2008 Vbias 0.0216f
C10475 VDD.n2009 Vbias 0.01836f
C10476 VDD.t880 Vbias 0.0169f
C10477 VDD.t1086 Vbias 0.0169f
C10478 VDD.n2010 Vbias 0.07902f
C10479 VDD.t647 Vbias 0.0169f
C10480 VDD.t1017 Vbias 0.0169f
C10481 VDD.n2011 Vbias 0.07902f
C10482 VDD.n2012 Vbias 0.03023f
C10483 VDD.n2013 Vbias 0.01699f
C10484 VDD.n2014 Vbias 0.03902f
C10485 VDD.n2015 Vbias 0.03694f
C10486 VDD.n2016 Vbias 0.0216f
C10487 VDD.n2017 Vbias 0.01836f
C10488 VDD.n2018 Vbias 0.03639f
C10489 VDD.t117 Vbias 0.46278f
C10490 VDD.n2019 Vbias 0.03694f
C10491 VDD.n2020 Vbias 0.03694f
C10492 VDD.n2021 Vbias 0.0216f
C10493 VDD.n2022 Vbias 0.01836f
C10494 VDD.t118 Vbias 0.017f
C10495 VDD.t753 Vbias 0.017f
C10496 VDD.n2023 Vbias 0.09633f
C10497 VDD.n2024 Vbias 0.04493f
C10498 VDD.n2026 Vbias 0.03902f
C10499 VDD.n2027 Vbias 0.03694f
C10500 VDD.n2028 Vbias 0.0216f
C10501 VDD.n2029 Vbias 0.01836f
C10502 VDD.n2030 Vbias 0.03639f
C10503 VDD.t256 Vbias 0.46278f
C10504 VDD.n2031 Vbias 0.03694f
C10505 VDD.n2032 Vbias 0.03694f
C10506 VDD.n2033 Vbias 0.0216f
C10507 VDD.n2034 Vbias 0.01836f
C10508 VDD.n2035 Vbias 0.03902f
C10509 VDD.n2036 Vbias 0.03694f
C10510 VDD.n2037 Vbias 0.07027f
C10511 VDD.t257 Vbias 0.0169f
C10512 VDD.t18 Vbias 0.0169f
C10513 VDD.n2038 Vbias 0.07902f
C10514 VDD.t919 Vbias 0.0169f
C10515 VDD.t388 Vbias 0.0169f
C10516 VDD.n2039 Vbias 0.07902f
C10517 VDD.n2040 Vbias 0.03902f
C10518 VDD.n2041 Vbias 0.03694f
C10519 VDD.n2042 Vbias 0.03902f
C10520 VDD.n2043 Vbias 0.03639f
C10521 VDD.n2044 Vbias 0.03639f
C10522 VDD.n2045 Vbias 0.03694f
C10523 VDD.n2046 Vbias 0.0216f
C10524 VDD.n2047 Vbias 0.01836f
C10525 VDD.n2048 Vbias 0.03639f
C10526 VDD.n2049 Vbias 0.01836f
C10527 VDD.n2050 Vbias 0.03639f
C10528 VDD.n2051 Vbias 0.37318f
C10529 VDD.n2052 Vbias 0.37318f
C10530 VDD.n2053 Vbias 0.01836f
C10531 VDD.n2054 Vbias 0.01836f
C10532 VDD.n2055 Vbias 0.0216f
C10533 VDD.n2056 Vbias 0.03694f
C10534 VDD.t1068 Vbias 0.46278f
C10535 VDD.n2057 Vbias 0.03694f
C10536 VDD.n2058 Vbias 0.03694f
C10537 VDD.n2059 Vbias 0.06648f
C10538 VDD.n2060 Vbias 0.03639f
C10539 VDD.t19 Vbias 0.46278f
C10540 VDD.n2061 Vbias 0.03694f
C10541 VDD.n2062 Vbias 0.03694f
C10542 VDD.n2063 Vbias 0.0216f
C10543 VDD.n2064 Vbias 0.01836f
C10544 VDD.t1069 Vbias 0.017f
C10545 VDD.n2065 Vbias 0.05322f
C10546 VDD.n2066 Vbias 0.01309f
C10547 VDD.n2067 Vbias 0.01699f
C10548 VDD.n2068 Vbias 0.03902f
C10549 VDD.n2069 Vbias 0.03694f
C10550 VDD.n2070 Vbias 0.0216f
C10551 VDD.n2071 Vbias 0.01836f
C10552 VDD.n2072 Vbias 0.03639f
C10553 VDD.t607 Vbias 0.46278f
C10554 VDD.n2073 Vbias 0.03694f
C10555 VDD.n2074 Vbias 0.03694f
C10556 VDD.n2075 Vbias 0.0216f
C10557 VDD.n2076 Vbias 0.01836f
C10558 VDD.t639 Vbias 0.0169f
C10559 VDD.t609 Vbias 0.0169f
C10560 VDD.n2077 Vbias 0.07902f
C10561 VDD.t20 Vbias 0.0169f
C10562 VDD.t608 Vbias 0.0169f
C10563 VDD.n2078 Vbias 0.07902f
C10564 VDD.n2079 Vbias 0.03023f
C10565 VDD.n2080 Vbias 0.01699f
C10566 VDD.n2081 Vbias 0.03902f
C10567 VDD.n2082 Vbias 0.03694f
C10568 VDD.n2083 Vbias 0.0216f
C10569 VDD.n2084 Vbias 0.01836f
C10570 VDD.n2085 Vbias 0.03639f
C10571 VDD.t57 Vbias 0.46278f
C10572 VDD.n2086 Vbias 0.03694f
C10573 VDD.n2087 Vbias 0.03694f
C10574 VDD.n2088 Vbias 0.0216f
C10575 VDD.n2089 Vbias 0.01836f
C10576 VDD.t58 Vbias 0.017f
C10577 VDD.t795 Vbias 0.017f
C10578 VDD.n2090 Vbias 0.09713f
C10579 VDD.n2091 Vbias 0.01914f
C10580 VDD.n2092 Vbias 0.03902f
C10581 VDD.n2093 Vbias 0.03694f
C10582 VDD.n2094 Vbias 0.0216f
C10583 VDD.n2095 Vbias 0.01836f
C10584 VDD.n2096 Vbias 0.03639f
C10585 VDD.t232 Vbias 0.46278f
C10586 VDD.n2097 Vbias 0.03694f
C10587 VDD.n2098 Vbias 0.03694f
C10588 VDD.n2099 Vbias 0.0216f
C10589 VDD.n2100 Vbias 0.01836f
C10590 VDD.n2101 Vbias 0.02305f
C10591 VDD.n2102 Vbias 0.03902f
C10592 VDD.n2103 Vbias 0.03694f
C10593 VDD.n2104 Vbias 0.0216f
C10594 VDD.n2105 Vbias 0.01836f
C10595 VDD.n2106 Vbias 0.03639f
C10596 VDD.t602 Vbias 0.46278f
C10597 VDD.n2107 Vbias 0.03694f
C10598 VDD.n2108 Vbias 0.03694f
C10599 VDD.n2109 Vbias 0.0216f
C10600 VDD.n2110 Vbias 0.01836f
C10601 VDD.t233 Vbias 0.0169f
C10602 VDD.t603 Vbias 0.0169f
C10603 VDD.n2111 Vbias 0.07902f
C10604 VDD.t999 Vbias 0.0169f
C10605 VDD.t872 Vbias 0.0169f
C10606 VDD.n2112 Vbias 0.07902f
C10607 VDD.n2113 Vbias 0.03023f
C10608 VDD.t921 Vbias 0.017f
C10609 VDD.n2114 Vbias 0.01999f
C10610 VDD.n2115 Vbias 0.03694f
C10611 VDD.n2116 Vbias 0.0216f
C10612 VDD.n2117 Vbias 0.03694f
C10613 VDD.n2118 Vbias 0.45845f
C10614 VDD.t920 Vbias 0.54191f
C10615 VDD.n2120 Vbias 0.03639f
C10616 VDD.t89 Vbias 0.46278f
C10617 VDD.n2121 Vbias 0.03694f
C10618 VDD.n2122 Vbias 0.03694f
C10619 VDD.n2123 Vbias 0.0216f
C10620 VDD.n2124 Vbias 0.01836f
C10621 VDD.t737 Vbias 0.017f
C10622 VDD.t90 Vbias 0.017f
C10623 VDD.n2125 Vbias 0.09713f
C10624 VDD.n2126 Vbias 0.01914f
C10625 VDD.n2127 Vbias 0.03902f
C10626 VDD.n2128 Vbias 0.03694f
C10627 VDD.n2129 Vbias 0.0216f
C10628 VDD.n2130 Vbias 0.01836f
C10629 VDD.n2131 Vbias 0.03639f
C10630 VDD.t186 Vbias 0.46278f
C10631 VDD.n2132 Vbias 0.03694f
C10632 VDD.n2133 Vbias 0.03694f
C10633 VDD.n2134 Vbias 0.0216f
C10634 VDD.n2135 Vbias 0.01836f
C10635 VDD.n2136 Vbias 0.02305f
C10636 VDD.n2137 Vbias 0.03902f
C10637 VDD.n2138 Vbias 0.03694f
C10638 VDD.n2139 Vbias 0.0216f
C10639 VDD.n2140 Vbias 0.01836f
C10640 VDD.n2141 Vbias 0.03639f
C10641 VDD.t1042 Vbias 0.46278f
C10642 VDD.n2142 Vbias 0.03694f
C10643 VDD.n2143 Vbias 0.03694f
C10644 VDD.n2144 Vbias 0.0216f
C10645 VDD.n2145 Vbias 0.01836f
C10646 VDD.t884 Vbias 0.0169f
C10647 VDD.t1098 Vbias 0.0169f
C10648 VDD.n2146 Vbias 0.07902f
C10649 VDD.t187 Vbias 0.0169f
C10650 VDD.t1043 Vbias 0.0169f
C10651 VDD.n2147 Vbias 0.07902f
C10652 VDD.n2148 Vbias 0.03023f
C10653 VDD.n2149 Vbias 0.01699f
C10654 VDD.n2150 Vbias 0.03902f
C10655 VDD.n2151 Vbias 0.03694f
C10656 VDD.n2152 Vbias 0.0216f
C10657 VDD.n2153 Vbias 0.01836f
C10658 VDD.n2154 Vbias 0.03639f
C10659 VDD.t39 Vbias 0.46278f
C10660 VDD.n2155 Vbias 0.03694f
C10661 VDD.n2156 Vbias 0.03694f
C10662 VDD.n2157 Vbias 0.0216f
C10663 VDD.n2158 Vbias 0.01836f
C10664 VDD.t40 Vbias 0.017f
C10665 VDD.t777 Vbias 0.017f
C10666 VDD.n2159 Vbias 0.09633f
C10667 VDD.n2160 Vbias 0.04493f
C10668 VDD.n2162 Vbias 0.03902f
C10669 VDD.n2163 Vbias 0.03694f
C10670 VDD.n2164 Vbias 0.0216f
C10671 VDD.n2165 Vbias 0.01836f
C10672 VDD.n2166 Vbias 0.03639f
C10673 VDD.t512 Vbias 0.46278f
C10674 VDD.n2167 Vbias 0.03694f
C10675 VDD.n2168 Vbias 0.03694f
C10676 VDD.n2169 Vbias 0.0216f
C10677 VDD.n2170 Vbias 0.01836f
C10678 VDD.n2171 Vbias 0.03902f
C10679 VDD.n2172 Vbias 0.03694f
C10680 VDD.n2173 Vbias 0.07027f
C10681 VDD.t957 Vbias 0.0169f
C10682 VDD.t1105 Vbias 0.0169f
C10683 VDD.n2174 Vbias 0.07902f
C10684 VDD.t513 Vbias 0.0169f
C10685 VDD.t222 Vbias 0.0169f
C10686 VDD.n2175 Vbias 0.07902f
C10687 VDD.n2176 Vbias 0.03902f
C10688 VDD.n2177 Vbias 0.03694f
C10689 VDD.n2178 Vbias 0.03902f
C10690 VDD.n2179 Vbias 0.03639f
C10691 VDD.n2180 Vbias 0.03639f
C10692 VDD.n2181 Vbias 0.03694f
C10693 VDD.n2182 Vbias 0.0216f
C10694 VDD.n2183 Vbias 0.01836f
C10695 VDD.n2184 Vbias 0.03639f
C10696 VDD.n2185 Vbias 0.01836f
C10697 VDD.n2186 Vbias 0.03639f
C10698 VDD.n2187 Vbias 0.37318f
C10699 VDD.n2188 Vbias 0.37318f
C10700 VDD.n2189 Vbias 0.01836f
C10701 VDD.n2190 Vbias 0.01836f
C10702 VDD.n2191 Vbias 0.0216f
C10703 VDD.n2192 Vbias 0.03694f
C10704 VDD.t1082 Vbias 0.46278f
C10705 VDD.n2193 Vbias 0.03694f
C10706 VDD.n2194 Vbias 0.03694f
C10707 VDD.n2195 Vbias 0.06648f
C10708 VDD.n2196 Vbias 0.03639f
C10709 VDD.t223 Vbias 0.46278f
C10710 VDD.n2197 Vbias 0.03694f
C10711 VDD.n2198 Vbias 0.03694f
C10712 VDD.n2199 Vbias 0.0216f
C10713 VDD.n2200 Vbias 0.01836f
C10714 VDD.t1083 Vbias 0.017f
C10715 VDD.n2201 Vbias 0.05322f
C10716 VDD.n2202 Vbias 0.01309f
C10717 VDD.n2203 Vbias 0.01699f
C10718 VDD.n2204 Vbias 0.03902f
C10719 VDD.n2205 Vbias 0.03694f
C10720 VDD.n2206 Vbias 0.0216f
C10721 VDD.n2207 Vbias 0.01836f
C10722 VDD.n2208 Vbias 0.03639f
C10723 VDD.t685 Vbias 0.46278f
C10724 VDD.n2209 Vbias 0.03694f
C10725 VDD.n2210 Vbias 0.03694f
C10726 VDD.n2211 Vbias 0.0216f
C10727 VDD.n2212 Vbias 0.01836f
C10728 VDD.t224 Vbias 0.0169f
C10729 VDD.t686 Vbias 0.0169f
C10730 VDD.n2213 Vbias 0.07902f
C10731 VDD.t430 Vbias 0.0169f
C10732 VDD.t836 Vbias 0.0169f
C10733 VDD.n2214 Vbias 0.07902f
C10734 VDD.n2215 Vbias 0.03023f
C10735 VDD.n2216 Vbias 0.01699f
C10736 VDD.n2217 Vbias 0.03902f
C10737 VDD.n2218 Vbias 0.03694f
C10738 VDD.n2219 Vbias 0.0216f
C10739 VDD.n2220 Vbias 0.01836f
C10740 VDD.n2221 Vbias 0.03639f
C10741 VDD.t63 Vbias 0.46278f
C10742 VDD.n2222 Vbias 0.03694f
C10743 VDD.n2223 Vbias 0.03694f
C10744 VDD.n2224 Vbias 0.0216f
C10745 VDD.n2225 Vbias 0.01836f
C10746 VDD.t64 Vbias 0.017f
C10747 VDD.t803 Vbias 0.017f
C10748 VDD.n2226 Vbias 0.09713f
C10749 VDD.n2227 Vbias 0.01914f
C10750 VDD.n2228 Vbias 0.03902f
C10751 VDD.n2229 Vbias 0.03694f
C10752 VDD.n2230 Vbias 0.0216f
C10753 VDD.n2231 Vbias 0.01836f
C10754 VDD.n2232 Vbias 0.03639f
C10755 VDD.t460 Vbias 0.46278f
C10756 VDD.n2233 Vbias 0.03694f
C10757 VDD.n2234 Vbias 0.03694f
C10758 VDD.n2235 Vbias 0.0216f
C10759 VDD.n2236 Vbias 0.01836f
C10760 VDD.n2237 Vbias 0.02305f
C10761 VDD.n2238 Vbias 0.03902f
C10762 VDD.n2239 Vbias 0.03694f
C10763 VDD.n2240 Vbias 0.0216f
C10764 VDD.n2241 Vbias 0.01836f
C10765 VDD.n2242 Vbias 0.03639f
C10766 VDD.t578 Vbias 0.46278f
C10767 VDD.n2243 Vbias 0.03694f
C10768 VDD.n2244 Vbias 0.03694f
C10769 VDD.n2245 Vbias 0.0216f
C10770 VDD.n2246 Vbias 0.01836f
C10771 VDD.t538 Vbias 0.0169f
C10772 VDD.t617 Vbias 0.0169f
C10773 VDD.n2247 Vbias 0.07902f
C10774 VDD.t461 Vbias 0.0169f
C10775 VDD.t579 Vbias 0.0169f
C10776 VDD.n2248 Vbias 0.07902f
C10777 VDD.n2249 Vbias 0.03023f
C10778 VDD.t292 Vbias 0.017f
C10779 VDD.n2250 Vbias 0.01999f
C10780 VDD.n2251 Vbias 0.03694f
C10781 VDD.n2252 Vbias 0.0216f
C10782 VDD.n2253 Vbias 0.03694f
C10783 VDD.n2254 Vbias 0.45845f
C10784 VDD.t291 Vbias 0.54191f
C10785 VDD.n2256 Vbias 0.03639f
C10786 VDD.t97 Vbias 0.46278f
C10787 VDD.n2257 Vbias 0.03694f
C10788 VDD.n2258 Vbias 0.03694f
C10789 VDD.n2259 Vbias 0.0216f
C10790 VDD.n2260 Vbias 0.01836f
C10791 VDD.t749 Vbias 0.017f
C10792 VDD.t98 Vbias 0.017f
C10793 VDD.n2261 Vbias 0.09713f
C10794 VDD.n2262 Vbias 0.01914f
C10795 VDD.n2263 Vbias 0.03902f
C10796 VDD.n2264 Vbias 0.03694f
C10797 VDD.n2265 Vbias 0.0216f
C10798 VDD.n2266 Vbias 0.01836f
C10799 VDD.n2267 Vbias 0.03639f
C10800 VDD.t564 Vbias 0.46278f
C10801 VDD.n2268 Vbias 0.03694f
C10802 VDD.n2269 Vbias 0.03694f
C10803 VDD.n2270 Vbias 0.0216f
C10804 VDD.n2271 Vbias 0.01836f
C10805 VDD.n2272 Vbias 0.02305f
C10806 VDD.n2273 Vbias 0.03902f
C10807 VDD.n2274 Vbias 0.03694f
C10808 VDD.n2275 Vbias 0.0216f
C10809 VDD.n2276 Vbias 0.01836f
C10810 VDD.n2277 Vbias 0.03639f
C10811 VDD.t1050 Vbias 0.46278f
C10812 VDD.n2278 Vbias 0.03694f
C10813 VDD.n2279 Vbias 0.03694f
C10814 VDD.n2280 Vbias 0.0216f
C10815 VDD.n2281 Vbias 0.01836f
C10816 VDD.t931 Vbias 0.0169f
C10817 VDD.t1051 Vbias 0.0169f
C10818 VDD.n2282 Vbias 0.07902f
C10819 VDD.t565 Vbias 0.0169f
C10820 VDD.t1091 Vbias 0.0169f
C10821 VDD.n2283 Vbias 0.07902f
C10822 VDD.n2284 Vbias 0.03023f
C10823 VDD.n2285 Vbias 0.01699f
C10824 VDD.n2286 Vbias 0.03902f
C10825 VDD.n2287 Vbias 0.03694f
C10826 VDD.n2288 Vbias 0.0216f
C10827 VDD.n2289 Vbias 0.01836f
C10828 VDD.n2290 Vbias 0.03639f
C10829 VDD.t109 Vbias 0.46278f
C10830 VDD.n2291 Vbias 0.03694f
C10831 VDD.n2292 Vbias 0.03694f
C10832 VDD.n2293 Vbias 0.0216f
C10833 VDD.n2294 Vbias 0.01836f
C10834 VDD.t110 Vbias 0.017f
C10835 VDD.t741 Vbias 0.017f
C10836 VDD.n2295 Vbias 0.09633f
C10837 VDD.n2296 Vbias 0.04493f
C10838 VDD.n2298 Vbias 0.03902f
C10839 VDD.n2299 Vbias 0.03694f
C10840 VDD.n2300 Vbias 0.0216f
C10841 VDD.n2301 Vbias 0.01836f
C10842 VDD.n2302 Vbias 0.03639f
C10843 VDD.t451 Vbias 0.46278f
C10844 VDD.n2303 Vbias 0.03694f
C10845 VDD.n2304 Vbias 0.03694f
C10846 VDD.n2305 Vbias 0.0216f
C10847 VDD.n2306 Vbias 0.01836f
C10848 VDD.n2307 Vbias 0.03902f
C10849 VDD.n2308 Vbias 0.03694f
C10850 VDD.n2309 Vbias 0.07027f
C10851 VDD.t875 Vbias 0.0169f
C10852 VDD.t968 Vbias 0.0169f
C10853 VDD.n2310 Vbias 0.07902f
C10854 VDD.t452 Vbias 0.0169f
C10855 VDD.t955 Vbias 0.0169f
C10856 VDD.n2311 Vbias 0.07902f
C10857 VDD.n2312 Vbias 0.03902f
C10858 VDD.n2313 Vbias 0.03694f
C10859 VDD.n2314 Vbias 0.03902f
C10860 VDD.n2315 Vbias 0.03639f
C10861 VDD.n2316 Vbias 0.03639f
C10862 VDD.n2317 Vbias 0.03694f
C10863 VDD.n2318 Vbias 0.0216f
C10864 VDD.n2319 Vbias 0.01836f
C10865 VDD.n2320 Vbias 0.03639f
C10866 VDD.n2321 Vbias 0.01836f
C10867 VDD.n2322 Vbias 0.03639f
C10868 VDD.n2323 Vbias 0.37318f
C10869 VDD.n2324 Vbias 0.37318f
C10870 VDD.n2325 Vbias 0.01836f
C10871 VDD.n2326 Vbias 0.01836f
C10872 VDD.n2327 Vbias 0.0216f
C10873 VDD.n2328 Vbias 0.03694f
C10874 VDD.t1010 Vbias 0.46278f
C10875 VDD.n2329 Vbias 0.03694f
C10876 VDD.n2330 Vbias 0.03694f
C10877 VDD.n2331 Vbias 0.06648f
C10878 VDD.n2332 Vbias 0.03639f
C10879 VDD.t660 Vbias 0.46278f
C10880 VDD.n2333 Vbias 0.03694f
C10881 VDD.n2334 Vbias 0.03694f
C10882 VDD.n2335 Vbias 0.0216f
C10883 VDD.n2336 Vbias 0.01836f
C10884 VDD.t1011 Vbias 0.017f
C10885 VDD.n2337 Vbias 0.05322f
C10886 VDD.n2338 Vbias 0.01309f
C10887 VDD.n2339 Vbias 0.01699f
C10888 VDD.n2340 Vbias 0.03902f
C10889 VDD.n2341 Vbias 0.03694f
C10890 VDD.n2342 Vbias 0.0216f
C10891 VDD.n2343 Vbias 0.01836f
C10892 VDD.n2344 Vbias 0.03639f
C10893 VDD.t337 Vbias 0.46278f
C10894 VDD.n2345 Vbias 0.03694f
C10895 VDD.n2346 Vbias 0.03694f
C10896 VDD.n2347 Vbias 0.0216f
C10897 VDD.n2348 Vbias 0.01836f
C10898 VDD.t661 Vbias 0.0169f
C10899 VDD.t338 Vbias 0.0169f
C10900 VDD.n2349 Vbias 0.07902f
C10901 VDD.t998 Vbias 0.0169f
C10902 VDD.t956 Vbias 0.0169f
C10903 VDD.n2350 Vbias 0.07902f
C10904 VDD.n2351 Vbias 0.03023f
C10905 VDD.n2352 Vbias 0.01699f
C10906 VDD.n2353 Vbias 0.03902f
C10907 VDD.n2354 Vbias 0.03694f
C10908 VDD.n2355 Vbias 0.0216f
C10909 VDD.n2356 Vbias 0.01836f
C10910 VDD.n2357 Vbias 0.03639f
C10911 VDD.t123 Vbias 0.46278f
C10912 VDD.n2358 Vbias 0.03694f
C10913 VDD.n2359 Vbias 0.03694f
C10914 VDD.n2360 Vbias 0.0216f
C10915 VDD.n2361 Vbias 0.01836f
C10916 VDD.t124 Vbias 0.017f
C10917 VDD.t755 Vbias 0.017f
C10918 VDD.n2362 Vbias 0.09713f
C10919 VDD.n2363 Vbias 0.01914f
C10920 VDD.n2364 Vbias 0.03902f
C10921 VDD.n2365 Vbias 0.03694f
C10922 VDD.n2366 Vbias 0.0216f
C10923 VDD.n2367 Vbias 0.01836f
C10924 VDD.n2368 Vbias 0.03639f
C10925 VDD.t625 Vbias 0.46278f
C10926 VDD.n2369 Vbias 0.03694f
C10927 VDD.n2370 Vbias 0.03694f
C10928 VDD.n2371 Vbias 0.0216f
C10929 VDD.n2372 Vbias 0.01836f
C10930 VDD.n2373 Vbias 0.02305f
C10931 VDD.n2374 Vbias 0.03902f
C10932 VDD.n2375 Vbias 0.03694f
C10933 VDD.n2376 Vbias 0.0216f
C10934 VDD.n2377 Vbias 0.01836f
C10935 VDD.n2378 Vbias 0.03639f
C10936 VDD.t453 Vbias 0.46278f
C10937 VDD.n2379 Vbias 0.03694f
C10938 VDD.n2380 Vbias 0.03694f
C10939 VDD.n2381 Vbias 0.0216f
C10940 VDD.n2382 Vbias 0.01836f
C10941 VDD.t626 Vbias 0.0169f
C10942 VDD.t454 Vbias 0.0169f
C10943 VDD.n2383 Vbias 0.07902f
C10944 VDD.t823 Vbias 0.0169f
C10945 VDD.t908 Vbias 0.0169f
C10946 VDD.n2384 Vbias 0.07902f
C10947 VDD.n2385 Vbias 0.03023f
C10948 VDD.t904 Vbias 0.017f
C10949 VDD.n2386 Vbias 0.01999f
C10950 VDD.n2387 Vbias 0.03694f
C10951 VDD.n2388 Vbias 0.0216f
C10952 VDD.n2389 Vbias 0.03694f
C10953 VDD.n2390 Vbias 0.45845f
C10954 VDD.t903 Vbias 0.54191f
C10955 VDD.n2392 Vbias 0.03639f
C10956 VDD.t95 Vbias 0.46278f
C10957 VDD.n2393 Vbias 0.03694f
C10958 VDD.n2394 Vbias 0.03694f
C10959 VDD.n2395 Vbias 0.0216f
C10960 VDD.n2396 Vbias 0.01836f
C10961 VDD.t743 Vbias 0.017f
C10962 VDD.t96 Vbias 0.017f
C10963 VDD.n2397 Vbias 0.09713f
C10964 VDD.n2398 Vbias 0.01914f
C10965 VDD.n2399 Vbias 0.03902f
C10966 VDD.n2400 Vbias 0.03694f
C10967 VDD.n2401 Vbias 0.0216f
C10968 VDD.n2402 Vbias 0.01836f
C10969 VDD.n2403 Vbias 0.03639f
C10970 VDD.t591 Vbias 0.46278f
C10971 VDD.n2404 Vbias 0.03694f
C10972 VDD.n2405 Vbias 0.03694f
C10973 VDD.n2406 Vbias 0.0216f
C10974 VDD.n2407 Vbias 0.01836f
C10975 VDD.n2408 Vbias 0.02305f
C10976 VDD.n2409 Vbias 0.03902f
C10977 VDD.n2410 Vbias 0.03694f
C10978 VDD.n2411 Vbias 0.0216f
C10979 VDD.n2412 Vbias 0.01836f
C10980 VDD.n2413 Vbias 0.03639f
C10981 VDD.t1048 Vbias 0.46278f
C10982 VDD.n2414 Vbias 0.03694f
C10983 VDD.n2415 Vbias 0.03694f
C10984 VDD.n2416 Vbias 0.0216f
C10985 VDD.n2417 Vbias 0.01836f
C10986 VDD.t907 Vbias 0.0169f
C10987 VDD.t1100 Vbias 0.0169f
C10988 VDD.n2418 Vbias 0.07902f
C10989 VDD.t592 Vbias 0.0169f
C10990 VDD.t1049 Vbias 0.0169f
C10991 VDD.n2419 Vbias 0.07902f
C10992 VDD.n2420 Vbias 0.03023f
C10993 VDD.n2421 Vbias 0.01699f
C10994 VDD.n2422 Vbias 0.03902f
C10995 VDD.n2423 Vbias 0.03694f
C10996 VDD.n2424 Vbias 0.0216f
C10997 VDD.n2425 Vbias 0.01836f
C10998 VDD.n2426 Vbias 0.03639f
C10999 VDD.t31 Vbias 0.46278f
C11000 VDD.n2427 Vbias 0.03694f
C11001 VDD.n2428 Vbias 0.03694f
C11002 VDD.n2429 Vbias 0.0216f
C11003 VDD.n2430 Vbias 0.01836f
C11004 VDD.t32 Vbias 0.017f
C11005 VDD.t767 Vbias 0.017f
C11006 VDD.n2431 Vbias 0.09633f
C11007 VDD.n2432 Vbias 0.04493f
C11008 VDD.n2434 Vbias 0.03902f
C11009 VDD.n2435 Vbias 0.03694f
C11010 VDD.n2436 Vbias 0.0216f
C11011 VDD.n2437 Vbias 0.01836f
C11012 VDD.n2438 Vbias 0.03639f
C11013 VDD.t426 Vbias 0.46278f
C11014 VDD.n2439 Vbias 0.03694f
C11015 VDD.n2440 Vbias 0.03694f
C11016 VDD.n2441 Vbias 0.0216f
C11017 VDD.n2442 Vbias 0.01836f
C11018 VDD.n2443 Vbias 0.03902f
C11019 VDD.n2444 Vbias 0.03694f
C11020 VDD.n2445 Vbias 0.07027f
C11021 VDD.t894 Vbias 0.0169f
C11022 VDD.t497 Vbias 0.0169f
C11023 VDD.n2446 Vbias 0.07902f
C11024 VDD.t427 Vbias 0.0169f
C11025 VDD.t237 Vbias 0.0169f
C11026 VDD.n2447 Vbias 0.07902f
C11027 VDD.n2448 Vbias 0.03902f
C11028 VDD.n2449 Vbias 0.03694f
C11029 VDD.n2450 Vbias 0.03902f
C11030 VDD.n2451 Vbias 0.03639f
C11031 VDD.n2452 Vbias 0.03639f
C11032 VDD.n2453 Vbias 0.03694f
C11033 VDD.n2454 Vbias 0.0216f
C11034 VDD.n2455 Vbias 0.01836f
C11035 VDD.n2456 Vbias 0.03639f
C11036 VDD.n2457 Vbias 0.01836f
C11037 VDD.n2458 Vbias 0.03639f
C11038 VDD.n2459 Vbias 0.37318f
C11039 VDD.n2460 Vbias 0.37318f
C11040 VDD.n2461 Vbias 0.01836f
C11041 VDD.n2462 Vbias 0.01836f
C11042 VDD.n2463 Vbias 0.0216f
C11043 VDD.n2464 Vbias 0.03694f
C11044 VDD.t1038 Vbias 0.46278f
C11045 VDD.n2465 Vbias 0.03694f
C11046 VDD.n2466 Vbias 0.03694f
C11047 VDD.n2467 Vbias 0.06648f
C11048 VDD.n2468 Vbias 0.03639f
C11049 VDD.t234 Vbias 0.46278f
C11050 VDD.n2469 Vbias 0.03694f
C11051 VDD.n2470 Vbias 0.03694f
C11052 VDD.n2471 Vbias 0.0216f
C11053 VDD.n2472 Vbias 0.01836f
C11054 VDD.t1039 Vbias 0.017f
C11055 VDD.n2473 Vbias 0.05322f
C11056 VDD.n2474 Vbias 0.01309f
C11057 VDD.n2475 Vbias 0.01699f
C11058 VDD.n2476 Vbias 0.03902f
C11059 VDD.n2477 Vbias 0.03694f
C11060 VDD.n2478 Vbias 0.0216f
C11061 VDD.n2479 Vbias 0.01836f
C11062 VDD.n2480 Vbias 0.03639f
C11063 VDD.t262 Vbias 0.46278f
C11064 VDD.n2481 Vbias 0.03694f
C11065 VDD.n2482 Vbias 0.03694f
C11066 VDD.n2483 Vbias 0.0216f
C11067 VDD.n2484 Vbias 0.01836f
C11068 VDD.t235 Vbias 0.0169f
C11069 VDD.t263 Vbias 0.0169f
C11070 VDD.n2485 Vbias 0.07902f
C11071 VDD.t645 Vbias 0.0169f
C11072 VDD.t496 Vbias 0.0169f
C11073 VDD.n2486 Vbias 0.07902f
C11074 VDD.n2487 Vbias 0.03023f
C11075 VDD.n2488 Vbias 0.01699f
C11076 VDD.n2489 Vbias 0.03902f
C11077 VDD.n2490 Vbias 0.03694f
C11078 VDD.n2491 Vbias 0.0216f
C11079 VDD.n2492 Vbias 0.01836f
C11080 VDD.n2493 Vbias 0.03639f
C11081 VDD.t41 Vbias 0.46278f
C11082 VDD.n2494 Vbias 0.03694f
C11083 VDD.n2495 Vbias 0.03694f
C11084 VDD.n2496 Vbias 0.0216f
C11085 VDD.n2497 Vbias 0.01836f
C11086 VDD.t42 Vbias 0.017f
C11087 VDD.t783 Vbias 0.017f
C11088 VDD.n2498 Vbias 0.09713f
C11089 VDD.n2499 Vbias 0.01914f
C11090 VDD.n2500 Vbias 0.03902f
C11091 VDD.n2501 Vbias 0.03694f
C11092 VDD.n2502 Vbias 0.0216f
C11093 VDD.n2503 Vbias 0.01836f
C11094 VDD.n2504 Vbias 0.03639f
C11095 VDD.t322 Vbias 0.46278f
C11096 VDD.n2505 Vbias 0.03694f
C11097 VDD.n2506 Vbias 0.03694f
C11098 VDD.n2507 Vbias 0.0216f
C11099 VDD.n2508 Vbias 0.01836f
C11100 VDD.n2509 Vbias 0.02305f
C11101 VDD.n2510 Vbias 0.03902f
C11102 VDD.n2511 Vbias 0.03694f
C11103 VDD.n2512 Vbias 0.0216f
C11104 VDD.n2513 Vbias 0.01836f
C11105 VDD.n2514 Vbias 0.03639f
C11106 VDD.t355 Vbias 0.46278f
C11107 VDD.n2515 Vbias 0.03694f
C11108 VDD.n2516 Vbias 0.03694f
C11109 VDD.n2517 Vbias 0.0216f
C11110 VDD.n2518 Vbias 0.01836f
C11111 VDD.t494 Vbias 0.0169f
C11112 VDD.t519 Vbias 0.0169f
C11113 VDD.n2519 Vbias 0.07902f
C11114 VDD.t323 Vbias 0.0169f
C11115 VDD.t356 Vbias 0.0169f
C11116 VDD.n2520 Vbias 0.07902f
C11117 VDD.n2521 Vbias 0.03023f
C11118 VDD.t572 Vbias 0.017f
C11119 VDD.n2522 Vbias 0.01999f
C11120 VDD.n2523 Vbias 0.03694f
C11121 VDD.n2524 Vbias 0.0216f
C11122 VDD.n2525 Vbias 0.03694f
C11123 VDD.n2526 Vbias 0.45845f
C11124 VDD.t571 Vbias 0.54191f
C11125 VDD.n2528 Vbias 0.03639f
C11126 VDD.t127 Vbias 0.46278f
C11127 VDD.n2529 Vbias 0.03694f
C11128 VDD.n2530 Vbias 0.03694f
C11129 VDD.n2531 Vbias 0.0216f
C11130 VDD.n2532 Vbias 0.01836f
C11131 VDD.t769 Vbias 0.017f
C11132 VDD.t128 Vbias 0.017f
C11133 VDD.n2533 Vbias 0.09713f
C11134 VDD.n2534 Vbias 0.01914f
C11135 VDD.n2535 Vbias 0.03902f
C11136 VDD.n2536 Vbias 0.03694f
C11137 VDD.n2537 Vbias 0.0216f
C11138 VDD.n2538 Vbias 0.01836f
C11139 VDD.n2539 Vbias 0.03639f
C11140 VDD.t353 Vbias 0.46278f
C11141 VDD.n2540 Vbias 0.03694f
C11142 VDD.n2541 Vbias 0.03694f
C11143 VDD.n2542 Vbias 0.0216f
C11144 VDD.n2543 Vbias 0.01836f
C11145 VDD.n2544 Vbias 0.02305f
C11146 VDD.n2545 Vbias 0.03902f
C11147 VDD.n2546 Vbias 0.03694f
C11148 VDD.n2547 Vbias 0.0216f
C11149 VDD.n2548 Vbias 0.01836f
C11150 VDD.n2549 Vbias 0.03639f
C11151 VDD.t1022 Vbias 0.46278f
C11152 VDD.n2550 Vbias 0.03694f
C11153 VDD.n2551 Vbias 0.03694f
C11154 VDD.n2552 Vbias 0.0216f
C11155 VDD.n2553 Vbias 0.01836f
C11156 VDD.t354 Vbias 0.0169f
C11157 VDD.t1023 Vbias 0.0169f
C11158 VDD.n2554 Vbias 0.07902f
C11159 VDD.t595 Vbias 0.0169f
C11160 VDD.t1073 Vbias 0.0169f
C11161 VDD.n2555 Vbias 0.07902f
C11162 VDD.n2556 Vbias 0.03023f
C11163 VDD.n2557 Vbias 0.01699f
C11164 VDD.n2558 Vbias 0.03902f
C11165 VDD.n2559 Vbias 0.03694f
C11166 VDD.n2560 Vbias 0.0216f
C11167 VDD.n2561 Vbias 0.01836f
C11168 VDD.n2562 Vbias 0.03639f
C11169 VDD.t79 Vbias 0.46278f
C11170 VDD.n2563 Vbias 0.03694f
C11171 VDD.n2564 Vbias 0.03694f
C11172 VDD.n2565 Vbias 0.0216f
C11173 VDD.n2566 Vbias 0.01836f
C11174 VDD.t80 Vbias 0.017f
C11175 VDD.t721 Vbias 0.017f
C11176 VDD.n2567 Vbias 0.09633f
C11177 VDD.n2568 Vbias 0.04493f
C11178 VDD.n2570 Vbias 0.03902f
C11179 VDD.n2571 Vbias 0.03694f
C11180 VDD.n2572 Vbias 0.0216f
C11181 VDD.n2573 Vbias 0.01836f
C11182 VDD.n2574 Vbias 0.03639f
C11183 VDD.t476 Vbias 0.46278f
C11184 VDD.n2575 Vbias 0.03694f
C11185 VDD.n2576 Vbias 0.03694f
C11186 VDD.n2577 Vbias 0.0216f
C11187 VDD.n2578 Vbias 0.01836f
C11188 VDD.n2579 Vbias 0.03902f
C11189 VDD.n2580 Vbias 0.03694f
C11190 VDD.n2581 Vbias 0.07027f
C11191 VDD.t854 Vbias 0.0169f
C11192 VDD.t622 Vbias 0.0169f
C11193 VDD.n2582 Vbias 0.07902f
C11194 VDD.t477 Vbias 0.0169f
C11195 VDD.t439 Vbias 0.0169f
C11196 VDD.n2583 Vbias 0.07902f
C11197 VDD.n2584 Vbias 0.03902f
C11198 VDD.n2585 Vbias 0.03694f
C11199 VDD.n2586 Vbias 0.03902f
C11200 VDD.n2587 Vbias 0.03639f
C11201 VDD.n2588 Vbias 0.03639f
C11202 VDD.n2589 Vbias 0.03694f
C11203 VDD.n2590 Vbias 0.0216f
C11204 VDD.n2591 Vbias 0.01836f
C11205 VDD.n2592 Vbias 0.03639f
C11206 VDD.n2593 Vbias 0.01836f
C11207 VDD.n2594 Vbias 0.03639f
C11208 VDD.n2595 Vbias 0.37318f
C11209 VDD.n2596 Vbias 0.37318f
C11210 VDD.n2597 Vbias 0.01836f
C11211 VDD.n2598 Vbias 0.01836f
C11212 VDD.n2599 Vbias 0.0216f
C11213 VDD.n2600 Vbias 0.03694f
C11214 VDD.t1062 Vbias 0.46278f
C11215 VDD.n2601 Vbias 0.03694f
C11216 VDD.n2602 Vbias 0.03694f
C11217 VDD.n2603 Vbias 0.06648f
C11218 VDD.n2604 Vbias 0.03639f
C11219 VDD.t440 Vbias 0.46278f
C11220 VDD.n2605 Vbias 0.03694f
C11221 VDD.n2606 Vbias 0.03694f
C11222 VDD.n2607 Vbias 0.0216f
C11223 VDD.n2608 Vbias 0.01836f
C11224 VDD.t1063 Vbias 0.017f
C11225 VDD.n2609 Vbias 0.05322f
C11226 VDD.n2610 Vbias 0.01309f
C11227 VDD.n2611 Vbias 0.01699f
C11228 VDD.n2612 Vbias 0.03902f
C11229 VDD.n2613 Vbias 0.03694f
C11230 VDD.n2614 Vbias 0.0216f
C11231 VDD.n2615 Vbias 0.01836f
C11232 VDD.n2616 Vbias 0.03639f
C11233 VDD.t817 Vbias 0.46278f
C11234 VDD.n2617 Vbias 0.03694f
C11235 VDD.n2618 Vbias 0.03694f
C11236 VDD.n2619 Vbias 0.0216f
C11237 VDD.n2620 Vbias 0.01836f
C11238 VDD.t441 Vbias 0.0169f
C11239 VDD.t819 Vbias 0.0169f
C11240 VDD.n2621 Vbias 0.07902f
C11241 VDD.t623 Vbias 0.0169f
C11242 VDD.t818 Vbias 0.0169f
C11243 VDD.n2622 Vbias 0.07902f
C11244 VDD.n2623 Vbias 0.03023f
C11245 VDD.n2624 Vbias 0.01699f
C11246 VDD.n2625 Vbias 0.03902f
C11247 VDD.n2626 Vbias 0.03694f
C11248 VDD.n2627 Vbias 0.0216f
C11249 VDD.n2628 Vbias 0.01836f
C11250 VDD.n2629 Vbias 0.03639f
C11251 VDD.t59 Vbias 0.46278f
C11252 VDD.n2630 Vbias 0.03694f
C11253 VDD.n2631 Vbias 0.03694f
C11254 VDD.n2632 Vbias 0.0216f
C11255 VDD.n2633 Vbias 0.01836f
C11256 VDD.t60 Vbias 0.017f
C11257 VDD.t799 Vbias 0.017f
C11258 VDD.n2634 Vbias 0.09713f
C11259 VDD.n2635 Vbias 0.01914f
C11260 VDD.n2636 Vbias 0.03902f
C11261 VDD.n2637 Vbias 0.03694f
C11262 VDD.n2638 Vbias 0.0216f
C11263 VDD.n2639 Vbias 0.01836f
C11264 VDD.n2640 Vbias 0.03639f
C11265 VDD.t474 Vbias 0.46278f
C11266 VDD.n2641 Vbias 0.03694f
C11267 VDD.n2642 Vbias 0.03694f
C11268 VDD.n2643 Vbias 0.0216f
C11269 VDD.n2644 Vbias 0.01836f
C11270 VDD.n2645 Vbias 0.02305f
C11271 VDD.n2646 Vbias 0.03902f
C11272 VDD.n2647 Vbias 0.03694f
C11273 VDD.n2648 Vbias 0.0216f
C11274 VDD.n2649 Vbias 0.01836f
C11275 VDD.n2650 Vbias 0.03639f
C11276 VDD.t320 Vbias 0.46278f
C11277 VDD.n2651 Vbias 0.03694f
C11278 VDD.n2652 Vbias 0.03694f
C11279 VDD.n2653 Vbias 0.0216f
C11280 VDD.n2654 Vbias 0.01836f
C11281 VDD.t482 Vbias 0.0169f
C11282 VDD.t457 Vbias 0.0169f
C11283 VDD.n2655 Vbias 0.07902f
C11284 VDD.t475 Vbias 0.0169f
C11285 VDD.t321 Vbias 0.0169f
C11286 VDD.n2656 Vbias 0.07902f
C11287 VDD.n2657 Vbias 0.03023f
C11288 VDD.t877 Vbias 0.017f
C11289 VDD.n2658 Vbias 0.01999f
C11290 VDD.n2659 Vbias 0.03694f
C11291 VDD.n2660 Vbias 0.0216f
C11292 VDD.n2661 Vbias 0.03694f
C11293 VDD.n2662 Vbias 0.45845f
C11294 VDD.t876 Vbias 0.54191f
C11295 VDD.n2664 Vbias 0.03639f
C11296 VDD.t45 Vbias 0.46278f
C11297 VDD.n2665 Vbias 0.03694f
C11298 VDD.n2666 Vbias 0.03694f
C11299 VDD.n2667 Vbias 0.0216f
C11300 VDD.n2668 Vbias 0.01836f
C11301 VDD.t791 Vbias 0.017f
C11302 VDD.t46 Vbias 0.017f
C11303 VDD.n2669 Vbias 0.09713f
C11304 VDD.n2670 Vbias 0.01914f
C11305 VDD.n2671 Vbias 0.03902f
C11306 VDD.n2672 Vbias 0.03694f
C11307 VDD.n2673 Vbias 0.0216f
C11308 VDD.n2674 Vbias 0.01836f
C11309 VDD.n2675 Vbias 0.03639f
C11310 VDD.t318 Vbias 0.46278f
C11311 VDD.n2676 Vbias 0.03694f
C11312 VDD.n2677 Vbias 0.03694f
C11313 VDD.n2678 Vbias 0.0216f
C11314 VDD.n2679 Vbias 0.01836f
C11315 VDD.n2680 Vbias 0.02305f
C11316 VDD.n2681 Vbias 0.03902f
C11317 VDD.n2682 Vbias 0.03694f
C11318 VDD.n2683 Vbias 0.0216f
C11319 VDD.n2684 Vbias 0.01836f
C11320 VDD.n2685 Vbias 0.03639f
C11321 VDD.t1018 Vbias 0.46278f
C11322 VDD.n2686 Vbias 0.03694f
C11323 VDD.n2687 Vbias 0.03694f
C11324 VDD.n2688 Vbias 0.0216f
C11325 VDD.n2689 Vbias 0.01836f
C11326 VDD.t319 Vbias 0.0169f
C11327 VDD.t1087 Vbias 0.0169f
C11328 VDD.n2690 Vbias 0.07902f
C11329 VDD.t632 Vbias 0.0169f
C11330 VDD.t1019 Vbias 0.0169f
C11331 VDD.n2691 Vbias 0.07902f
C11332 VDD.n2692 Vbias 0.03023f
C11333 VDD.n2693 Vbias 0.01699f
C11334 VDD.n2694 Vbias 0.03902f
C11335 VDD.n2695 Vbias 0.03694f
C11336 VDD.n2696 Vbias 0.0216f
C11337 VDD.n2697 Vbias 0.01836f
C11338 VDD.n2698 Vbias 0.03639f
C11339 VDD.t105 Vbias 0.46278f
C11340 VDD.n2699 Vbias 0.03694f
C11341 VDD.n2700 Vbias 0.03694f
C11342 VDD.n2701 Vbias 0.0216f
C11343 VDD.n2702 Vbias 0.01836f
C11344 VDD.t106 Vbias 0.017f
C11345 VDD.t735 Vbias 0.017f
C11346 VDD.n2703 Vbias 0.09633f
C11347 VDD.n2704 Vbias 0.04493f
C11348 VDD.n2706 Vbias 0.03902f
C11349 VDD.n2707 Vbias 0.03694f
C11350 VDD.n2708 Vbias 0.0216f
C11351 VDD.n2709 Vbias 0.01836f
C11352 VDD.n2710 Vbias 0.03639f
C11353 VDD.t925 Vbias 0.46278f
C11354 VDD.n2711 Vbias 0.03694f
C11355 VDD.n2712 Vbias 0.03694f
C11356 VDD.n2713 Vbias 0.0216f
C11357 VDD.n2714 Vbias 0.01836f
C11358 VDD.n2715 Vbias 0.03902f
C11359 VDD.n2716 Vbias 0.03694f
C11360 VDD.n2717 Vbias 0.07027f
C11361 VDD.t953 Vbias 0.0169f
C11362 VDD.t559 Vbias 0.0169f
C11363 VDD.n2718 Vbias 0.07902f
C11364 VDD.t926 Vbias 0.0169f
C11365 VDD.t526 Vbias 0.0169f
C11366 VDD.n2719 Vbias 0.07902f
C11367 VDD.n2720 Vbias 0.03902f
C11368 VDD.n2721 Vbias 0.03694f
C11369 VDD.n2722 Vbias 0.03902f
C11370 VDD.n2723 Vbias 0.03639f
C11371 VDD.n2724 Vbias 0.03639f
C11372 VDD.n2725 Vbias 0.03694f
C11373 VDD.n2726 Vbias 0.0216f
C11374 VDD.n2727 Vbias 0.01836f
C11375 VDD.n2728 Vbias 0.03639f
C11376 VDD.n2729 Vbias 0.01836f
C11377 VDD.n2730 Vbias 0.03639f
C11378 VDD.n2731 Vbias 0.37318f
C11379 VDD.n2732 Vbias 0.37318f
C11380 VDD.n2733 Vbias 0.01836f
C11381 VDD.n2734 Vbias 0.01836f
C11382 VDD.n2735 Vbias 0.0216f
C11383 VDD.n2736 Vbias 0.03694f
C11384 VDD.t1006 Vbias 0.46278f
C11385 VDD.n2737 Vbias 0.03694f
C11386 VDD.n2738 Vbias 0.03694f
C11387 VDD.n2739 Vbias 0.06648f
C11388 VDD.n2740 Vbias 0.03639f
C11389 VDD.t527 Vbias 0.46278f
C11390 VDD.n2741 Vbias 0.03694f
C11391 VDD.n2742 Vbias 0.03694f
C11392 VDD.n2743 Vbias 0.0216f
C11393 VDD.n2744 Vbias 0.01836f
C11394 VDD.t1007 Vbias 0.017f
C11395 VDD.n2745 Vbias 0.05322f
C11396 VDD.n2746 Vbias 0.01309f
C11397 VDD.n2747 Vbias 0.01699f
C11398 VDD.n2748 Vbias 0.03902f
C11399 VDD.n2749 Vbias 0.03694f
C11400 VDD.n2750 Vbias 0.0216f
C11401 VDD.n2751 Vbias 0.01836f
C11402 VDD.n2752 Vbias 0.03639f
C11403 VDD.t295 Vbias 0.46278f
C11404 VDD.n2753 Vbias 0.03694f
C11405 VDD.n2754 Vbias 0.03694f
C11406 VDD.n2755 Vbias 0.0216f
C11407 VDD.n2756 Vbias 0.01836f
C11408 VDD.t528 Vbias 0.0169f
C11409 VDD.t296 Vbias 0.0169f
C11410 VDD.n2757 Vbias 0.07902f
C11411 VDD.t560 Vbias 0.0169f
C11412 VDD.t839 Vbias 0.0169f
C11413 VDD.n2758 Vbias 0.07902f
C11414 VDD.n2759 Vbias 0.03023f
C11415 VDD.n2760 Vbias 0.01699f
C11416 VDD.n2761 Vbias 0.03902f
C11417 VDD.n2762 Vbias 0.03694f
C11418 VDD.n2763 Vbias 0.0216f
C11419 VDD.n2764 Vbias 0.01836f
C11420 VDD.n2765 Vbias 0.03639f
C11421 VDD.t115 Vbias 0.46278f
C11422 VDD.n2766 Vbias 0.03694f
C11423 VDD.n2767 Vbias 0.03694f
C11424 VDD.n2768 Vbias 0.0216f
C11425 VDD.n2769 Vbias 0.01836f
C11426 VDD.t116 Vbias 0.017f
C11427 VDD.t751 Vbias 0.017f
C11428 VDD.n2770 Vbias 0.09713f
C11429 VDD.n2771 Vbias 0.01914f
C11430 VDD.n2772 Vbias 0.03902f
C11431 VDD.n2773 Vbias 0.03694f
C11432 VDD.n2774 Vbias 0.0216f
C11433 VDD.n2775 Vbias 0.01836f
C11434 VDD.n2776 Vbias 0.03639f
C11435 VDD.t0 Vbias 0.46278f
C11436 VDD.n2777 Vbias 0.03694f
C11437 VDD.n2778 Vbias 0.03694f
C11438 VDD.n2779 Vbias 0.0216f
C11439 VDD.n2780 Vbias 0.01836f
C11440 VDD.n2781 Vbias 0.02305f
C11441 VDD.n2782 Vbias 0.03902f
C11442 VDD.n2783 Vbias 0.03694f
C11443 VDD.n2784 Vbias 0.0216f
C11444 VDD.n2785 Vbias 0.01836f
C11445 VDD.n2786 Vbias 0.03639f
C11446 VDD.t182 Vbias 0.46278f
C11447 VDD.n2787 Vbias 0.03694f
C11448 VDD.n2788 Vbias 0.03694f
C11449 VDD.n2789 Vbias 0.0216f
C11450 VDD.n2790 Vbias 0.01836f
C11451 VDD.t1 Vbias 0.0169f
C11452 VDD.t627 Vbias 0.0169f
C11453 VDD.n2791 Vbias 0.07902f
C11454 VDD.t842 Vbias 0.0169f
C11455 VDD.t183 Vbias 0.0169f
C11456 VDD.n2792 Vbias 0.07902f
C11457 VDD.n2793 Vbias 0.03023f
C11458 VDD.t1103 Vbias 0.017f
C11459 VDD.n2794 Vbias 0.01999f
C11460 VDD.n2795 Vbias 0.03694f
C11461 VDD.n2796 Vbias 0.0216f
C11462 VDD.n2797 Vbias 0.03694f
C11463 VDD.n2798 Vbias 0.45845f
C11464 VDD.t1102 Vbias 0.54191f
C11465 VDD.n2800 Vbias 0.03639f
C11466 VDD.t93 Vbias 0.46278f
C11467 VDD.n2801 Vbias 0.03694f
C11468 VDD.n2802 Vbias 0.03694f
C11469 VDD.n2803 Vbias 0.0216f
C11470 VDD.n2804 Vbias 0.01836f
C11471 VDD.t739 Vbias 0.017f
C11472 VDD.t94 Vbias 0.017f
C11473 VDD.n2805 Vbias 0.09713f
C11474 VDD.n2806 Vbias 0.01914f
C11475 VDD.n2807 Vbias 0.03902f
C11476 VDD.n2808 Vbias 0.03694f
C11477 VDD.n2809 Vbias 0.0216f
C11478 VDD.n2810 Vbias 0.01836f
C11479 VDD.n2811 Vbias 0.03639f
C11480 VDD.t180 Vbias 0.46278f
C11481 VDD.n2812 Vbias 0.03694f
C11482 VDD.n2813 Vbias 0.03694f
C11483 VDD.n2814 Vbias 0.0216f
C11484 VDD.n2815 Vbias 0.01836f
C11485 VDD.n2816 Vbias 0.02305f
C11486 VDD.n2817 Vbias 0.03902f
C11487 VDD.n2818 Vbias 0.03694f
C11488 VDD.n2819 Vbias 0.0216f
C11489 VDD.n2820 Vbias 0.01836f
C11490 VDD.n2821 Vbias 0.03639f
C11491 VDD.t1045 Vbias 0.46278f
C11492 VDD.n2822 Vbias 0.03694f
C11493 VDD.n2823 Vbias 0.03694f
C11494 VDD.n2824 Vbias 0.0216f
C11495 VDD.n2825 Vbias 0.01836f
C11496 VDD.t181 Vbias 0.0169f
C11497 VDD.t1099 Vbias 0.0169f
C11498 VDD.n2826 Vbias 0.07902f
C11499 VDD.t547 Vbias 0.0169f
C11500 VDD.t1046 Vbias 0.0169f
C11501 VDD.n2827 Vbias 0.07902f
C11502 VDD.n2828 Vbias 0.03023f
C11503 VDD.n2829 Vbias 0.01699f
C11504 VDD.n2830 Vbias 0.03902f
C11505 VDD.n2831 Vbias 0.03694f
C11506 VDD.n2832 Vbias 0.0216f
C11507 VDD.n2833 Vbias 0.01836f
C11508 VDD.n2834 Vbias 0.03639f
C11509 VDD.t27 Vbias 0.46278f
C11510 VDD.n2835 Vbias 0.03694f
C11511 VDD.n2836 Vbias 0.03694f
C11512 VDD.n2837 Vbias 0.0216f
C11513 VDD.n2838 Vbias 0.01836f
C11514 VDD.t28 Vbias 0.017f
C11515 VDD.t763 Vbias 0.017f
C11516 VDD.n2839 Vbias 0.09633f
C11517 VDD.n2840 Vbias 0.04493f
C11518 VDD.n2842 Vbias 0.03902f
C11519 VDD.n2843 Vbias 0.03694f
C11520 VDD.n2844 Vbias 0.0216f
C11521 VDD.n2845 Vbias 0.01836f
C11522 VDD.n2846 Vbias 0.03639f
C11523 VDD.t373 Vbias 0.46278f
C11524 VDD.n2847 Vbias 0.03694f
C11525 VDD.n2848 Vbias 0.03694f
C11526 VDD.n2849 Vbias 0.0216f
C11527 VDD.n2850 Vbias 0.01836f
C11528 VDD.n2851 Vbias 0.03902f
C11529 VDD.n2852 Vbias 0.03694f
C11530 VDD.n2853 Vbias 0.07027f
C11531 VDD.t374 Vbias 0.0169f
C11532 VDD.t511 Vbias 0.0169f
C11533 VDD.n2854 Vbias 0.07902f
C11534 VDD.t1106 Vbias 0.0169f
C11535 VDD.t542 Vbias 0.0169f
C11536 VDD.n2855 Vbias 0.07902f
C11537 VDD.n2856 Vbias 0.03902f
C11538 VDD.n2857 Vbias 0.03694f
C11539 VDD.n2858 Vbias 0.03902f
C11540 VDD.n2859 Vbias 0.03639f
C11541 VDD.n2860 Vbias 0.03639f
C11542 VDD.n2861 Vbias 0.03694f
C11543 VDD.n2862 Vbias 0.0216f
C11544 VDD.n2863 Vbias 0.01836f
C11545 VDD.n2864 Vbias 0.03639f
C11546 VDD.n2865 Vbias 0.01836f
C11547 VDD.n2866 Vbias 0.03639f
C11548 VDD.n2867 Vbias 0.37318f
C11549 VDD.n2868 Vbias 0.37318f
C11550 VDD.n2869 Vbias 0.01836f
C11551 VDD.n2870 Vbias 0.01836f
C11552 VDD.n2871 Vbias 0.0216f
C11553 VDD.n2872 Vbias 0.03694f
C11554 VDD.t1034 Vbias 0.46278f
C11555 VDD.n2873 Vbias 0.03694f
C11556 VDD.n2874 Vbias 0.03694f
C11557 VDD.n2875 Vbias 0.06648f
C11558 VDD.n2876 Vbias 0.03639f
C11559 VDD.t543 Vbias 0.46278f
C11560 VDD.n2877 Vbias 0.03694f
C11561 VDD.n2878 Vbias 0.03694f
C11562 VDD.n2879 Vbias 0.0216f
C11563 VDD.n2880 Vbias 0.01836f
C11564 VDD.t1035 Vbias 0.017f
C11565 VDD.n2881 Vbias 0.05322f
C11566 VDD.n2882 Vbias 0.01309f
C11567 VDD.n2883 Vbias 0.01699f
C11568 VDD.n2884 Vbias 0.03902f
C11569 VDD.n2885 Vbias 0.03694f
C11570 VDD.n2886 Vbias 0.0216f
C11571 VDD.n2887 Vbias 0.01836f
C11572 VDD.n2888 Vbias 0.03639f
C11573 VDD.t166 Vbias 0.46278f
C11574 VDD.n2889 Vbias 0.03694f
C11575 VDD.n2890 Vbias 0.03694f
C11576 VDD.n2891 Vbias 0.0216f
C11577 VDD.n2892 Vbias 0.01836f
C11578 VDD.t544 Vbias 0.0169f
C11579 VDD.t334 Vbias 0.0169f
C11580 VDD.n2893 Vbias 0.07902f
C11581 VDD.t930 Vbias 0.0169f
C11582 VDD.t167 Vbias 0.0169f
C11583 VDD.n2894 Vbias 0.07902f
C11584 VDD.n2895 Vbias 0.03023f
C11585 VDD.n2896 Vbias 0.01699f
C11586 VDD.n2897 Vbias 0.03902f
C11587 VDD.n2898 Vbias 0.03694f
C11588 VDD.n2899 Vbias 0.0216f
C11589 VDD.n2900 Vbias 0.01836f
C11590 VDD.n2901 Vbias 0.03639f
C11591 VDD.t37 Vbias 0.46278f
C11592 VDD.n2902 Vbias 0.03694f
C11593 VDD.n2903 Vbias 0.03694f
C11594 VDD.n2904 Vbias 0.0216f
C11595 VDD.n2905 Vbias 0.01836f
C11596 VDD.t38 Vbias 0.017f
C11597 VDD.t775 Vbias 0.017f
C11598 VDD.n2906 Vbias 0.09713f
C11599 VDD.n2907 Vbias 0.01914f
C11600 VDD.n2908 Vbias 0.03902f
C11601 VDD.n2909 Vbias 0.03694f
C11602 VDD.n2910 Vbias 0.0216f
C11603 VDD.n2911 Vbias 0.01836f
C11604 VDD.n2912 Vbias 0.03639f
C11605 VDD.t704 Vbias 0.46278f
C11606 VDD.n2913 Vbias 0.03694f
C11607 VDD.n2914 Vbias 0.03694f
C11608 VDD.n2915 Vbias 0.0216f
C11609 VDD.n2916 Vbias 0.01836f
C11610 VDD.n2917 Vbias 0.02305f
C11611 VDD.n2918 Vbias 0.03902f
C11612 VDD.n2919 Vbias 0.03694f
C11613 VDD.n2920 Vbias 0.0216f
C11614 VDD.n2921 Vbias 0.01836f
C11615 VDD.n2922 Vbias 0.03639f
C11616 VDD.t689 Vbias 0.46278f
C11617 VDD.n2923 Vbias 0.03694f
C11618 VDD.n2924 Vbias 0.03694f
C11619 VDD.n2925 Vbias 0.0216f
C11620 VDD.n2926 Vbias 0.01836f
C11621 VDD.t705 Vbias 0.0169f
C11622 VDD.t690 Vbias 0.0169f
C11623 VDD.n2927 Vbias 0.07902f
C11624 VDD.t840 Vbias 0.0169f
C11625 VDD.t698 Vbias 0.0169f
C11626 VDD.n2928 Vbias 0.07902f
C11627 VDD.n2929 Vbias 0.03023f
C11628 VDD.t697 Vbias 0.017f
C11629 VDD.n2930 Vbias 0.01999f
C11630 VDD.n2931 Vbias 0.03694f
C11631 VDD.n2932 Vbias 0.0216f
C11632 VDD.n2933 Vbias 0.03694f
C11633 VDD.n2934 Vbias 0.45845f
C11634 VDD.t696 Vbias 0.54191f
C11635 VDD.n2936 Vbias 0.03639f
C11636 VDD.t119 Vbias 0.46278f
C11637 VDD.n2937 Vbias 0.03694f
C11638 VDD.n2938 Vbias 0.03694f
C11639 VDD.n2939 Vbias 0.0216f
C11640 VDD.n2940 Vbias 0.01836f
C11641 VDD.t765 Vbias 0.017f
C11642 VDD.t120 Vbias 0.017f
C11643 VDD.n2941 Vbias 0.09713f
C11644 VDD.n2942 Vbias 0.01914f
C11645 VDD.n2943 Vbias 0.03902f
C11646 VDD.n2944 Vbias 0.03694f
C11647 VDD.n2945 Vbias 0.0216f
C11648 VDD.n2946 Vbias 0.01836f
C11649 VDD.n2947 Vbias 0.03639f
C11650 VDD.t692 Vbias 0.46278f
C11651 VDD.n2948 Vbias 0.03694f
C11652 VDD.n2949 Vbias 0.03694f
C11653 VDD.n2950 Vbias 0.0216f
C11654 VDD.n2951 Vbias 0.01836f
C11655 VDD.n2952 Vbias 0.02305f
C11656 VDD.n2953 Vbias 0.03902f
C11657 VDD.n2954 Vbias 0.03694f
C11658 VDD.n2955 Vbias 0.0216f
C11659 VDD.n2956 Vbias 0.01836f
C11660 VDD.n2957 Vbias 0.03639f
C11661 VDD.t1014 Vbias 0.46278f
C11662 VDD.n2958 Vbias 0.03694f
C11663 VDD.n2959 Vbias 0.03694f
C11664 VDD.n2960 Vbias 0.0216f
C11665 VDD.n2961 Vbias 0.01836f
C11666 VDD.t693 Vbias 0.0169f
C11667 VDD.t1015 Vbias 0.0169f
C11668 VDD.n2962 Vbias 0.07902f
C11669 VDD.t975 Vbias 0.0169f
C11670 VDD.t1064 Vbias 0.0169f
C11671 VDD.n2963 Vbias 0.07902f
C11672 VDD.n2964 Vbias 0.03023f
C11673 VDD.n2965 Vbias 0.01699f
C11674 VDD.n2966 Vbias 0.03902f
C11675 VDD.n2967 Vbias 0.03694f
C11676 VDD.n2968 Vbias 0.0216f
C11677 VDD.n2969 Vbias 0.01836f
C11678 VDD.n2970 Vbias 0.03639f
C11679 VDD.t75 Vbias 0.46278f
C11680 VDD.n2971 Vbias 0.03694f
C11681 VDD.n2972 Vbias 0.03694f
C11682 VDD.n2973 Vbias 0.0216f
C11683 VDD.n2974 Vbias 0.01836f
C11684 VDD.t76 Vbias 0.017f
C11685 VDD.t717 Vbias 0.017f
C11686 VDD.n2975 Vbias 0.09633f
C11687 VDD.n2976 Vbias 0.04493f
C11688 VDD.n2977 Vbias 0.55479f
C11689 VDD.t1140 Vbias 0.12359f
C11690 VDD.n2978 Vbias 0.12446f
C11691 VDD.n2979 Vbias 0.01328f
C11692 VDD.t778 Vbias 0.06426f
C11693 VDD.n2980 Vbias 0.01851f
C11694 VDD.n2983 Vbias 0.02099f
C11695 VDD.t1134 Vbias 0.12359f
C11696 VDD.n2984 Vbias 0.0361f
C11697 VDD.n2985 Vbias 0.01567f
C11698 VDD.n2986 Vbias 0.06888f
C11699 VDD.t718 Vbias 0.05748f
C11700 VDD.n2987 Vbias 0.03298f
C11701 VDD.n2988 Vbias 0.10227f
C11702 VDD.t1120 Vbias 0.12359f
C11703 VDD.n2989 Vbias 0.12446f
C11704 VDD.n2990 Vbias 0.01328f
C11705 VDD.t780 Vbias 0.06426f
C11706 VDD.n2991 Vbias 0.01851f
C11707 VDD.n2995 Vbias 0.13128f
C11708 VDD.n2996 Vbias 0.16f
C11709 VDD.n2997 Vbias 0.55479f
C11710 VDD.t730 Vbias 0.06426f
C11711 VDD.n2998 Vbias 0.05994f
C11712 VDD.n2999 Vbias 0.01328f
C11713 VDD.t1126 Vbias 0.12359f
C11714 VDD.n3000 Vbias 0.0361f
C11715 VDD.n3001 Vbias 0.01199f
C11716 VDD.n3002 Vbias 0.02025f
C11717 VDD.n3003 Vbias 0.02099f
C11718 VDD.t1157 Vbias 0.12359f
C11719 VDD.n3004 Vbias 0.12814f
C11720 VDD.n3005 Vbias 0.01386f
C11721 VDD.n3006 Vbias 0.01851f
C11722 VDD.t806 Vbias 0.05773f
C11723 VDD.n3007 Vbias 0.11603f
C11724 VDD.n3008 Vbias 0.03298f
C11725 VDD.t772 Vbias 0.06426f
C11726 VDD.n3009 Vbias 0.05994f
C11727 VDD.n3010 Vbias 0.01328f
C11728 VDD.t1125 Vbias 0.12359f
C11729 VDD.n3011 Vbias 0.0361f
C11730 VDD.n3012 Vbias 0.01199f
C11731 VDD.n3013 Vbias 0.02025f
C11732 VDD.n3015 Vbias 0.12697f
C11733 VDD.n3016 Vbias 0.13295f
C11734 VDD.t1158 Vbias 0.12359f
C11735 VDD.n3017 Vbias 0.0361f
C11736 VDD.n3018 Vbias 0.01199f
C11737 VDD.n3019 Vbias 0.02025f
C11738 VDD.t1119 Vbias 0.12359f
C11739 VDD.n3020 Vbias 0.12814f
C11740 VDD.n3021 Vbias 0.01386f
C11741 VDD.n3022 Vbias 0.01851f
C11742 VDD.t768 Vbias 0.05773f
C11743 VDD.n3023 Vbias 0.11603f
C11744 VDD.n3024 Vbias 0.03298f
C11745 VDD.t798 Vbias 0.06426f
C11746 VDD.n3025 Vbias 0.05994f
C11747 VDD.n3026 Vbias 0.01328f
C11748 VDD.t1139 Vbias 0.12359f
C11749 VDD.n3027 Vbias 0.0361f
C11750 VDD.n3028 Vbias 0.01199f
C11751 VDD.n3029 Vbias 0.02025f
C11752 VDD.n3030 Vbias 0.07665f
C11753 VDD.n3031 Vbias 0.19471f
C11754 VDD.n3033 Vbias 0.01328f
C11755 VDD.n3034 Vbias 0.05994f
C11756 VDD.t720 Vbias 0.05693f
C11757 VDD.n3035 Vbias 0.10524f
C11758 VDD.n3036 Vbias 0.55479f
C11759 VDD.t714 Vbias 0.06426f
C11760 VDD.n3037 Vbias 0.05994f
C11761 VDD.n3038 Vbias 0.01328f
C11762 VDD.t1135 Vbias 0.12359f
C11763 VDD.n3039 Vbias 0.0361f
C11764 VDD.n3040 Vbias 0.01199f
C11765 VDD.n3041 Vbias 0.02025f
C11766 VDD.n3042 Vbias 0.02099f
C11767 VDD.t1143 Vbias 0.12359f
C11768 VDD.n3043 Vbias 0.12814f
C11769 VDD.n3044 Vbias 0.01386f
C11770 VDD.n3045 Vbias 0.01851f
C11771 VDD.t724 Vbias 0.05773f
C11772 VDD.n3046 Vbias 0.11603f
C11773 VDD.n3047 Vbias 0.03298f
C11774 VDD.t796 Vbias 0.06426f
C11775 VDD.n3048 Vbias 0.05994f
C11776 VDD.n3049 Vbias 0.01328f
C11777 VDD.t1111 Vbias 0.12359f
C11778 VDD.n3050 Vbias 0.0361f
C11779 VDD.n3051 Vbias 0.01199f
C11780 VDD.n3052 Vbias 0.02025f
C11781 VDD.n3054 Vbias 0.12697f
C11782 VDD.n3055 Vbias 0.13295f
C11783 VDD.t728 Vbias 0.06426f
C11784 VDD.n3056 Vbias 0.05994f
C11785 VDD.n3057 Vbias 0.01328f
C11786 VDD.t1127 Vbias 0.12359f
C11787 VDD.n3058 Vbias 0.0361f
C11788 VDD.n3059 Vbias 0.01199f
C11789 VDD.n3060 Vbias 0.02025f
C11790 VDD.n3061 Vbias 0.02099f
C11791 VDD.t1136 Vbias 0.12359f
C11792 VDD.n3062 Vbias 0.12814f
C11793 VDD.n3063 Vbias 0.01386f
C11794 VDD.n3064 Vbias 0.01851f
C11795 VDD.t744 Vbias 0.05773f
C11796 VDD.n3065 Vbias 0.11603f
C11797 VDD.n3066 Vbias 0.03298f
C11798 VDD.t812 Vbias 0.06426f
C11799 VDD.n3067 Vbias 0.05994f
C11800 VDD.n3068 Vbias 0.01328f
C11801 VDD.t1153 Vbias 0.12359f
C11802 VDD.n3069 Vbias 0.0361f
C11803 VDD.n3070 Vbias 0.01199f
C11804 VDD.n3071 Vbias 0.02025f
C11805 VDD.n3073 Vbias 0.12697f
C11806 VDD.n3074 Vbias 0.13295f
C11807 VDD.n3075 Vbias 1.39487f
C11808 VDD.t756 Vbias 0.06426f
C11809 VDD.n3076 Vbias 0.05994f
C11810 VDD.n3077 Vbias 0.01328f
C11811 VDD.t1113 Vbias 0.12359f
C11812 VDD.n3078 Vbias 0.0361f
C11813 VDD.n3079 Vbias 0.01199f
C11814 VDD.n3080 Vbias 0.02025f
C11815 VDD.n3081 Vbias 0.02099f
C11816 VDD.t1124 Vbias 0.12359f
C11817 VDD.n3082 Vbias 0.12814f
C11818 VDD.n3083 Vbias 0.01386f
C11819 VDD.n3084 Vbias 0.01851f
C11820 VDD.t804 Vbias 0.05773f
C11821 VDD.n3085 Vbias 0.11603f
C11822 VDD.n3086 Vbias 0.03298f
C11823 VDD.t726 Vbias 0.06426f
C11824 VDD.n3087 Vbias 0.05994f
C11825 VDD.n3088 Vbias 0.01328f
C11826 VDD.t1128 Vbias 0.12359f
C11827 VDD.n3089 Vbias 0.0361f
C11828 VDD.n3090 Vbias 0.01199f
C11829 VDD.n3091 Vbias 0.02025f
C11830 VDD.n3093 Vbias 0.12697f
C11831 VDD.n3094 Vbias 0.13295f
C11832 VDD.t1132 Vbias 0.12359f
C11833 VDD.n3095 Vbias 0.0361f
C11834 VDD.n3096 Vbias 0.01199f
C11835 VDD.n3097 Vbias 0.02025f
C11836 VDD.t1110 Vbias 0.12359f
C11837 VDD.n3098 Vbias 0.12814f
C11838 VDD.n3099 Vbias 0.01386f
C11839 VDD.n3100 Vbias 0.01851f
C11840 VDD.t800 Vbias 0.05773f
C11841 VDD.n3101 Vbias 0.11603f
C11842 VDD.n3102 Vbias 0.03298f
C11843 VDD.t794 Vbias 0.06426f
C11844 VDD.n3103 Vbias 0.05994f
C11845 VDD.n3104 Vbias 0.01328f
C11846 VDD.t1141 Vbias 0.12359f
C11847 VDD.n3105 Vbias 0.0361f
C11848 VDD.n3106 Vbias 0.01199f
C11849 VDD.n3107 Vbias 0.02025f
C11850 VDD.n3108 Vbias 0.07665f
C11851 VDD.n3109 Vbias 0.19471f
C11852 VDD.n3111 Vbias 0.01328f
C11853 VDD.n3112 Vbias 0.05994f
C11854 VDD.t752 Vbias 0.05693f
C11855 VDD.n3113 Vbias 0.10524f
C11856 VDD.t1149 Vbias 0.12359f
C11857 VDD.n3114 Vbias 0.0361f
C11858 VDD.n3115 Vbias 0.01199f
C11859 VDD.n3116 Vbias 0.02025f
C11860 VDD.t1121 Vbias 0.12359f
C11861 VDD.n3117 Vbias 0.12814f
C11862 VDD.n3118 Vbias 0.01386f
C11863 VDD.n3119 Vbias 0.01851f
C11864 VDD.t784 Vbias 0.05773f
C11865 VDD.n3120 Vbias 0.11603f
C11866 VDD.n3121 Vbias 0.03298f
C11867 VDD.t746 Vbias 0.06426f
C11868 VDD.n3122 Vbias 0.05994f
C11869 VDD.n3123 Vbias 0.01328f
C11870 VDD.t1116 Vbias 0.12359f
C11871 VDD.n3124 Vbias 0.0361f
C11872 VDD.n3125 Vbias 0.01199f
C11873 VDD.n3126 Vbias 0.02025f
C11874 VDD.n3127 Vbias 0.07665f
C11875 VDD.n3128 Vbias 0.19471f
C11876 VDD.n3130 Vbias 0.01328f
C11877 VDD.n3131 Vbias 0.05994f
C11878 VDD.t722 Vbias 0.05693f
C11879 VDD.n3132 Vbias 0.10524f
C11880 VDD.n3133 Vbias 1.13968f
C11881 VDD.n3134 Vbias 0.7221f
C11882 VDD.n3135 Vbias 0.275f
C11883 VDD.n3136 Vbias 0.27852f
C11884 VDD.n3137 Vbias 1.1396f
C11885 VDD.n3138 Vbias 1.14318f
C11886 VDD.n3139 Vbias 0.58347f
C11887 VDD.t808 Vbias 0.06426f
C11888 VDD.n3140 Vbias 0.05994f
C11889 VDD.n3141 Vbias 0.01328f
C11890 VDD.t1156 Vbias 0.12359f
C11891 VDD.n3142 Vbias 0.0361f
C11892 VDD.n3143 Vbias 0.01199f
C11893 VDD.n3144 Vbias 0.02025f
C11894 VDD.n3145 Vbias 0.02099f
C11895 VDD.t1154 Vbias 0.12359f
C11896 VDD.n3146 Vbias 0.12814f
C11897 VDD.n3147 Vbias 0.01386f
C11898 VDD.n3148 Vbias 0.01851f
C11899 VDD.t810 Vbias 0.05773f
C11900 VDD.n3149 Vbias 0.11603f
C11901 VDD.n3150 Vbias 0.03298f
C11902 VDD.t732 Vbias 0.06426f
C11903 VDD.n3151 Vbias 0.05994f
C11904 VDD.n3152 Vbias 0.01328f
C11905 VDD.t1122 Vbias 0.12359f
C11906 VDD.n3153 Vbias 0.0361f
C11907 VDD.n3154 Vbias 0.01199f
C11908 VDD.n3155 Vbias 0.02025f
C11909 VDD.n3157 Vbias 0.12697f
C11910 VDD.n3158 Vbias 0.13295f
C11911 VDD.t1155 Vbias 0.12359f
C11912 VDD.n3159 Vbias 0.0361f
C11913 VDD.n3160 Vbias 0.01199f
C11914 VDD.n3161 Vbias 0.02025f
C11915 VDD.t1151 Vbias 0.12359f
C11916 VDD.n3162 Vbias 0.12814f
C11917 VDD.n3163 Vbias 0.01386f
C11918 VDD.n3164 Vbias 0.01851f
C11919 VDD.t736 Vbias 0.05773f
C11920 VDD.n3165 Vbias 0.11603f
C11921 VDD.n3166 Vbias 0.03298f
C11922 VDD.t802 Vbias 0.06426f
C11923 VDD.n3167 Vbias 0.05994f
C11924 VDD.n3168 Vbias 0.01328f
C11925 VDD.t1138 Vbias 0.12359f
C11926 VDD.n3169 Vbias 0.0361f
C11927 VDD.n3170 Vbias 0.01199f
C11928 VDD.n3171 Vbias 0.02025f
C11929 VDD.n3172 Vbias 0.07665f
C11930 VDD.n3173 Vbias 0.19471f
C11931 VDD.n3175 Vbias 0.01328f
C11932 VDD.n3176 Vbias 0.05994f
C11933 VDD.t776 Vbias 0.05693f
C11934 VDD.n3177 Vbias 0.10524f
C11935 VDD.n3178 Vbias 1.1396f
C11936 VDD.n3179 Vbias 1.14318f
C11937 VDD.n3180 Vbias 0.55479f
C11938 VDD.n3181 Vbias 0.55479f
C11939 VDD.n3182 Vbias 1.14318f
C11940 VDD.t1130 Vbias 0.12359f
C11941 VDD.n3183 Vbias 0.0361f
C11942 VDD.n3184 Vbias 0.01199f
C11943 VDD.n3185 Vbias 0.02025f
C11944 VDD.t1133 Vbias 0.12359f
C11945 VDD.n3186 Vbias 0.12814f
C11946 VDD.n3187 Vbias 0.01386f
C11947 VDD.n3188 Vbias 0.01851f
C11948 VDD.t748 Vbias 0.05773f
C11949 VDD.n3189 Vbias 0.11603f
C11950 VDD.n3190 Vbias 0.03298f
C11951 VDD.t754 Vbias 0.06426f
C11952 VDD.n3191 Vbias 0.05994f
C11953 VDD.n3192 Vbias 0.01328f
C11954 VDD.t1129 Vbias 0.12359f
C11955 VDD.n3193 Vbias 0.0361f
C11956 VDD.n3194 Vbias 0.01199f
C11957 VDD.n3195 Vbias 0.02025f
C11958 VDD.n3196 Vbias 0.07665f
C11959 VDD.n3197 Vbias 0.19471f
C11960 VDD.n3199 Vbias 0.01328f
C11961 VDD.n3200 Vbias 0.05994f
C11962 VDD.t740 Vbias 0.05693f
C11963 VDD.n3201 Vbias 0.10524f
C11964 VDD.n3202 Vbias 1.1396f
C11965 VDD.n3203 Vbias 0.55479f
C11966 VDD.n3204 Vbias 0.24851f
C11967 VDD.t161 Vbias 0.01699f
C11968 VDD.t673 Vbias 0.01699f
C11969 VDD.n3205 Vbias 0.10299f
C11970 VDD.n3206 Vbias 0.03902f
C11971 VDD.n3207 Vbias 0.03694f
C11972 VDD.n3208 Vbias 0.03902f
C11973 VDD.n3209 Vbias 0.03639f
C11974 VDD.n3210 Vbias 0.03639f
C11975 VDD.n3211 Vbias 0.50118f
C11976 VDD.n3212 Vbias 0.01836f
C11977 VDD.n3213 Vbias 0.01836f
C11978 VDD.n3214 Vbias 0.0216f
C11979 VDD.n3215 Vbias 0.03694f
C11980 VDD.n3216 Vbias 0.03639f
C11981 VDD.t315 Vbias 0.46278f
C11982 VDD.n3217 Vbias 0.03694f
C11983 VDD.n3218 Vbias 0.03694f
C11984 VDD.n3219 Vbias 0.0216f
C11985 VDD.n3220 Vbias 0.01836f
C11986 VDD.n3221 Vbias 0.02215f
C11987 VDD.n3222 Vbias 0.03902f
C11988 VDD.n3223 Vbias 0.03694f
C11989 VDD.n3224 Vbias 0.0216f
C11990 VDD.n3225 Vbias 0.01836f
C11991 VDD.n3226 Vbias 0.03639f
C11992 VDD.t282 Vbias 0.46278f
C11993 VDD.n3227 Vbias 0.03694f
C11994 VDD.n3228 Vbias 0.03694f
C11995 VDD.n3229 Vbias 0.0216f
C11996 VDD.n3230 Vbias 0.01836f
C11997 VDD.n3231 Vbias 0.03902f
C11998 VDD.n3232 Vbias 0.03694f
C11999 VDD.n3233 Vbias 0.0216f
C12000 VDD.n3234 Vbias 0.01836f
C12001 VDD.n3235 Vbias 0.01836f
C12002 VDD.n3236 Vbias 0.03639f
C12003 VDD.n3237 Vbias 0.50118f
C12004 VDD.n3238 Vbias 0.03639f
C12005 VDD.n3239 Vbias 0.03694f
C12006 VDD.n3240 Vbias 0.14151f
C12007 VDD.n3241 Vbias 0.02579f
C12008 VDD.t967 Vbias 0.01858f
C12009 VDD.n3242 Vbias 0.06635f
C12010 VDD.n3243 Vbias 0.02581f
C12011 VDD.n3245 Vbias 0.40967f
C12012 VDD.n3246 Vbias 0.01999f
C12013 VDD.n3247 Vbias 0.03694f
C12014 VDD.n3248 Vbias 0.0216f
C12015 VDD.n3249 Vbias 0.03694f
C12016 VDD.t407 Vbias 0.22551f
C12017 VDD.n3250 Vbias 0.03694f
C12018 VDD.n3251 Vbias 0.03694f
C12019 VDD.n3252 Vbias 0.0216f
C12020 VDD.n3253 Vbias 0.01999f
C12021 VDD.t406 Vbias 0.01699f
C12022 VDD.n3254 Vbias 0.24838f
C12023 VDD.t465 Vbias 0.01699f
C12024 VDD.n3255 Vbias 0.05918f
C12025 VDD.n3256 Vbias 0.01999f
C12026 VDD.n3257 Vbias 0.03694f
C12027 VDD.n3258 Vbias 0.0216f
C12028 VDD.n3259 Vbias 0.03694f
C12029 VDD.n3260 Vbias 0.26017f
C12030 VDD.t464 Vbias 0.24595f
C12031 VDD.t225 Vbias 0.22551f
C12032 VDD.n3262 Vbias 0.03694f
C12033 VDD.n3263 Vbias 0.03694f
C12034 VDD.n3264 Vbias 0.0216f
C12035 VDD.n3265 Vbias 0.01999f
C12036 VDD.n3266 Vbias 0.01999f
C12037 VDD.n3267 Vbias 0.03694f
C12038 VDD.n3268 Vbias 0.0216f
C12039 VDD.n3269 Vbias 0.03694f
C12040 VDD.n3270 Vbias 0.03639f
C12041 VDD.n3271 Vbias 0.18185f
C12042 VDD.n3272 Vbias 0.03639f
C12043 VDD.n3273 Vbias 0.18185f
C12044 VDD.t381 Vbias 0.24595f
C12045 VDD.n3275 Vbias 0.26017f
C12046 VDD.n3276 Vbias 0.01999f
C12047 VDD.n3277 Vbias 0.06648f
C12048 VDD.n3278 Vbias 0.03346f
C12049 VDD.t619 Vbias 0.01858f
C12050 VDD.n3279 Vbias 0.06636f
C12051 VDD.n3280 Vbias 0.02579f
C12052 VDD.n3282 Vbias 0.66679f
C12053 VDD.n3283 Vbias 0.01999f
C12054 VDD.n3284 Vbias 0.03694f
C12055 VDD.n3285 Vbias 0.0216f
C12056 VDD.n3286 Vbias 0.03694f
C12057 VDD.t386 Vbias 0.22551f
C12058 VDD.n3287 Vbias 0.03694f
C12059 VDD.n3288 Vbias 0.03694f
C12060 VDD.n3289 Vbias 0.0216f
C12061 VDD.n3290 Vbias 0.01999f
C12062 VDD.t385 Vbias 0.01699f
C12063 VDD.t786 Vbias 0.06426f
C12064 VDD.n3291 Vbias 0.05994f
C12065 VDD.n3292 Vbias 0.01328f
C12066 VDD.t1152 Vbias 0.12359f
C12067 VDD.n3293 Vbias 0.0361f
C12068 VDD.n3294 Vbias 0.01199f
C12069 VDD.n3295 Vbias 0.02025f
C12070 VDD.n3296 Vbias 0.02099f
C12071 VDD.t1114 Vbias 0.12359f
C12072 VDD.n3297 Vbias 0.12814f
C12073 VDD.n3298 Vbias 0.01386f
C12074 VDD.n3299 Vbias 0.01851f
C12075 VDD.t788 Vbias 0.05773f
C12076 VDD.n3300 Vbias 0.11603f
C12077 VDD.n3301 Vbias 0.03298f
C12078 VDD.t814 Vbias 0.06426f
C12079 VDD.n3302 Vbias 0.05994f
C12080 VDD.n3303 Vbias 0.01328f
C12081 VDD.t1137 Vbias 0.12359f
C12082 VDD.n3304 Vbias 0.0361f
C12083 VDD.n3305 Vbias 0.01199f
C12084 VDD.n3306 Vbias 0.02025f
C12085 VDD.n3308 Vbias 0.12697f
C12086 VDD.n3309 Vbias 0.13295f
C12087 VDD.n3310 Vbias 0.21255f
C12088 VDD.t212 Vbias 0.01699f
C12089 VDD.n3311 Vbias 0.05918f
C12090 VDD.n3312 Vbias 0.01999f
C12091 VDD.n3313 Vbias 0.03694f
C12092 VDD.n3314 Vbias 0.0216f
C12093 VDD.n3315 Vbias 0.03694f
C12094 VDD.n3316 Vbias 0.26017f
C12095 VDD.t211 Vbias 0.24595f
C12096 VDD.t213 Vbias 0.22551f
C12097 VDD.n3318 Vbias 0.03694f
C12098 VDD.n3319 Vbias 0.03694f
C12099 VDD.n3320 Vbias 0.0216f
C12100 VDD.n3321 Vbias 0.01999f
C12101 VDD.n3322 Vbias 0.01999f
C12102 VDD.n3323 Vbias 0.03694f
C12103 VDD.n3324 Vbias 0.0216f
C12104 VDD.n3325 Vbias 0.03694f
C12105 VDD.n3326 Vbias 0.03639f
C12106 VDD.n3327 Vbias 0.18185f
C12107 VDD.n3328 Vbias 0.03639f
C12108 VDD.n3329 Vbias 0.18185f
C12109 VDD.t533 Vbias 0.24595f
C12110 VDD.n3331 Vbias 0.26017f
C12111 VDD.n3332 Vbias 0.01999f
C12112 VDD.n3333 Vbias 0.06648f
C12113 VDD.n3334 Vbias 0.79053f
C12114 VDD.t916 Vbias 0.02233f
C12115 VDD.n3335 Vbias 0.10253f
C12116 VDD.n3336 Vbias 0.02734f
C12117 VDD.t534 Vbias 0.01858f
C12118 VDD.n3337 Vbias 0.06636f
C12119 VDD.n3338 Vbias 0.02734f
C12120 VDD.n3339 Vbias 0.05805f
C12121 VDD.t988 Vbias 0.02232f
C12122 VDD.n3340 Vbias 0.13076f
C12123 VDD.n3341 Vbias 0.09126f
C12124 VDD.t308 Vbias 0.01858f
C12125 VDD.n3342 Vbias 0.06636f
C12126 VDD.n3343 Vbias 0.02734f
C12127 VDD.n3344 Vbias 0.05805f
C12128 VDD.t895 Vbias 0.02232f
C12129 VDD.n3345 Vbias 0.11637f
C12130 VDD.n3346 Vbias 0.07687f
C12131 VDD.n3348 Vbias 0.02579f
C12132 VDD.n3349 Vbias 0.02215f
C12133 VDD.n3350 Vbias 0.06648f
C12134 VDD.n3351 Vbias 0.01999f
C12135 VDD.n3352 Vbias 0.03639f
C12136 VDD.n3353 Vbias 0.18185f
C12137 VDD.n3354 Vbias 0.18185f
C12138 VDD.n3355 Vbias 0.03639f
C12139 VDD.n3356 Vbias 0.01999f
C12140 VDD.n3357 Vbias 0.06648f
C12141 VDD.n3358 Vbias 0.01151f
C12142 VDD.n3359 Vbias 0.08999f
C12143 VDD.n3360 Vbias 0.26476f
C12144 VDD.n3361 Vbias 0.23398f
C12145 VDD.n3362 Vbias 0.08999f
C12146 VDD.n3363 Vbias 0.01999f
C12147 VDD.n3364 Vbias 0.03694f
C12148 VDD.n3365 Vbias 0.0216f
C12149 VDD.n3366 Vbias 0.03694f
C12150 VDD.n3367 Vbias 0.26017f
C12151 VDD.t384 Vbias 0.24595f
C12152 VDD.n3369 Vbias 0.03639f
C12153 VDD.n3370 Vbias 0.18185f
C12154 VDD.n3371 Vbias 0.18185f
C12155 VDD.n3372 Vbias 0.03639f
C12156 VDD.n3373 Vbias 0.01999f
C12157 VDD.n3374 Vbias 0.06648f
C12158 VDD.n3375 Vbias 0.01151f
C12159 VDD.n3376 Vbias 0.05918f
C12160 VDD.n3377 Vbias 0.02579f
C12161 VDD.n3378 Vbias 0.02215f
C12162 VDD.n3379 Vbias 0.06648f
C12163 VDD.n3380 Vbias 0.01999f
C12164 VDD.n3381 Vbias 0.03639f
C12165 VDD.n3382 Vbias 0.18185f
C12166 VDD.n3383 Vbias 0.03639f
C12167 VDD.n3384 Vbias 0.18185f
C12168 VDD.t307 Vbias 0.24595f
C12169 VDD.n3386 Vbias 0.26017f
C12170 VDD.n3387 Vbias 0.01999f
C12171 VDD.n3388 Vbias 0.06648f
C12172 VDD.n3389 Vbias 0.03346f
C12173 VDD.n3390 Vbias 0.58844f
C12174 VDD.n3391 Vbias 0.49906f
C12175 VDD.n3392 Vbias 0.01999f
C12176 VDD.n3393 Vbias 0.03694f
C12177 VDD.n3394 Vbias 0.0216f
C12178 VDD.n3395 Vbias 0.03694f
C12179 VDD.t992 Vbias 0.22551f
C12180 VDD.n3396 Vbias 0.03694f
C12181 VDD.n3397 Vbias 0.03694f
C12182 VDD.n3398 Vbias 0.0216f
C12183 VDD.n3399 Vbias 0.01999f
C12184 VDD.t991 Vbias 0.01699f
C12185 VDD.n3400 Vbias 0.08999f
C12186 VDD.n3401 Vbias 0.01999f
C12187 VDD.n3402 Vbias 0.03694f
C12188 VDD.n3403 Vbias 0.0216f
C12189 VDD.n3404 Vbias 0.03694f
C12190 VDD.n3405 Vbias 0.26017f
C12191 VDD.t990 Vbias 0.24595f
C12192 VDD.n3407 Vbias 0.03639f
C12193 VDD.n3408 Vbias 0.18185f
C12194 VDD.n3409 Vbias 0.18185f
C12195 VDD.n3410 Vbias 0.03639f
C12196 VDD.n3411 Vbias 0.01999f
C12197 VDD.n3412 Vbias 0.06648f
C12198 VDD.n3413 Vbias 0.01151f
C12199 VDD.n3414 Vbias 0.05918f
C12200 VDD.n3415 Vbias 0.02215f
C12201 VDD.n3416 Vbias 0.06648f
C12202 VDD.n3417 Vbias 0.01999f
C12203 VDD.n3418 Vbias 0.03639f
C12204 VDD.n3419 Vbias 0.18185f
C12205 VDD.n3420 Vbias 0.03639f
C12206 VDD.n3421 Vbias 0.18185f
C12207 VDD.t618 Vbias 0.24595f
C12208 VDD.n3423 Vbias 0.26017f
C12209 VDD.n3424 Vbias 0.01999f
C12210 VDD.n3425 Vbias 0.06648f
C12211 VDD.n3426 Vbias 0.03346f
C12212 VDD.n3428 Vbias 0.09126f
C12213 VDD.t974 Vbias 0.02232f
C12214 VDD.n3429 Vbias 0.13076f
C12215 VDD.n3430 Vbias 0.05805f
C12216 VDD.n3431 Vbias 0.02734f
C12217 VDD.t382 Vbias 0.01858f
C12218 VDD.n3432 Vbias 0.06636f
C12219 VDD.n3433 Vbias 0.02734f
C12220 VDD.n3434 Vbias 0.05805f
C12221 VDD.t4 Vbias 0.02232f
C12222 VDD.n3435 Vbias 0.13076f
C12223 VDD.n3436 Vbias 0.09126f
C12224 VDD.t868 Vbias 0.01858f
C12225 VDD.n3437 Vbias 0.06636f
C12226 VDD.n3438 Vbias 0.02734f
C12227 VDD.n3439 Vbias 0.05805f
C12228 VDD.t402 Vbias 0.02232f
C12229 VDD.n3440 Vbias 0.24735f
C12230 VDD.n3441 Vbias 0.20785f
C12231 VDD.n3443 Vbias 0.02579f
C12232 VDD.n3444 Vbias 0.02215f
C12233 VDD.n3445 Vbias 0.06648f
C12234 VDD.n3446 Vbias 0.01999f
C12235 VDD.n3447 Vbias 0.03639f
C12236 VDD.n3448 Vbias 0.18185f
C12237 VDD.n3449 Vbias 0.18185f
C12238 VDD.n3450 Vbias 0.03639f
C12239 VDD.n3451 Vbias 0.01999f
C12240 VDD.n3452 Vbias 0.06648f
C12241 VDD.n3453 Vbias 0.01151f
C12242 VDD.n3454 Vbias 0.08999f
C12243 VDD.n3455 Vbias 0.36497f
C12244 VDD.n3456 Vbias 0.36497f
C12245 VDD.n3457 Vbias 0.08999f
C12246 VDD.n3458 Vbias 0.01999f
C12247 VDD.n3459 Vbias 0.03694f
C12248 VDD.n3460 Vbias 0.0216f
C12249 VDD.n3461 Vbias 0.03694f
C12250 VDD.n3462 Vbias 0.26017f
C12251 VDD.t405 Vbias 0.24595f
C12252 VDD.n3464 Vbias 0.03639f
C12253 VDD.n3465 Vbias 0.18185f
C12254 VDD.n3466 Vbias 0.18185f
C12255 VDD.n3467 Vbias 0.03639f
C12256 VDD.n3468 Vbias 0.01999f
C12257 VDD.n3469 Vbias 0.06648f
C12258 VDD.n3470 Vbias 0.01151f
C12259 VDD.n3471 Vbias 0.05918f
C12260 VDD.n3472 Vbias 0.02579f
C12261 VDD.n3473 Vbias 0.02215f
C12262 VDD.n3474 Vbias 0.06648f
C12263 VDD.n3475 Vbias 0.01999f
C12264 VDD.n3476 Vbias 0.03639f
C12265 VDD.n3477 Vbias 0.18185f
C12266 VDD.n3478 Vbias 0.03639f
C12267 VDD.n3479 Vbias 0.18185f
C12268 VDD.t867 Vbias 0.24595f
C12269 VDD.n3481 Vbias 0.26017f
C12270 VDD.n3482 Vbias 0.01999f
C12271 VDD.n3483 Vbias 0.06648f
C12272 VDD.n3484 Vbias 0.03346f
C12273 VDD.n3485 Vbias 0.2309f
C12274 VDD.n3486 Vbias 0.01999f
C12275 VDD.n3487 Vbias 0.03694f
C12276 VDD.n3488 Vbias 0.0216f
C12277 VDD.n3489 Vbias 0.03694f
C12278 VDD.t642 Vbias 0.22551f
C12279 VDD.n3490 Vbias 0.03694f
C12280 VDD.n3491 Vbias 0.03694f
C12281 VDD.n3492 Vbias 0.0216f
C12282 VDD.n3493 Vbias 0.01999f
C12283 VDD.t641 Vbias 0.01699f
C12284 VDD.n3494 Vbias 0.08999f
C12285 VDD.n3495 Vbias 0.01999f
C12286 VDD.n3496 Vbias 0.03694f
C12287 VDD.n3497 Vbias 0.0216f
C12288 VDD.n3498 Vbias 0.03694f
C12289 VDD.n3499 Vbias 0.26017f
C12290 VDD.t640 Vbias 0.24595f
C12291 VDD.n3501 Vbias 0.03639f
C12292 VDD.n3502 Vbias 0.18185f
C12293 VDD.n3503 Vbias 0.18185f
C12294 VDD.n3504 Vbias 0.03639f
C12295 VDD.n3505 Vbias 0.01999f
C12296 VDD.n3506 Vbias 0.06648f
C12297 VDD.n3507 Vbias 0.01151f
C12298 VDD.n3508 Vbias 0.05918f
C12299 VDD.n3509 Vbias 0.02215f
C12300 VDD.n3510 Vbias 0.06648f
C12301 VDD.n3511 Vbias 0.01999f
C12302 VDD.n3512 Vbias 0.03639f
C12303 VDD.n3513 Vbias 0.18185f
C12304 VDD.n3514 Vbias 0.03639f
C12305 VDD.n3515 Vbias 0.18185f
C12306 VDD.t966 Vbias 0.24595f
C12307 VDD.n3517 Vbias 0.26017f
C12308 VDD.n3518 Vbias 0.01999f
C12309 VDD.n3519 Vbias 0.06648f
C12310 VDD.n3520 Vbias 0.03375f
C12311 VDD.n3522 Vbias 0.0914f
C12312 VDD.t159 Vbias 0.02232f
C12313 VDD.n3523 Vbias 0.13089f
C12314 VDD.n3524 Vbias 0.05805f
C12315 VDD.n3525 Vbias 0.02734f
C12316 VDD.t557 Vbias 0.01858f
C12317 VDD.n3526 Vbias 0.06636f
C12318 VDD.t532 Vbias 0.02233f
C12319 VDD.n3527 Vbias 0.02734f
C12320 VDD.n3528 Vbias 0.05805f
C12321 VDD.t283 Vbias 0.01858f
C12322 VDD.n3529 Vbias 0.06654f
C12323 VDD.n3530 Vbias 0.04142f
C12324 VDD.n3532 Vbias 0.03346f
C12325 VDD.n3533 Vbias 0.04583f
C12326 VDD.n3534 Vbias 0.03902f
C12327 VDD.n3535 Vbias 0.01836f
C12328 VDD.n3536 Vbias 0.03639f
C12329 VDD.n3537 Vbias 0.37318f
C12330 VDD.n3538 Vbias 0.01836f
C12331 VDD.n3539 Vbias 0.03639f
C12332 VDD.n3540 Vbias 0.37318f
C12333 VDD.n3541 Vbias 0.03639f
C12334 VDD.n3542 Vbias 0.03694f
C12335 VDD.n3543 Vbias 0.04583f
C12336 VDD.n3544 Vbias 0.03902f
C12337 VDD.n3545 Vbias 0.01836f
C12338 VDD.n3546 Vbias 0.03639f
C12339 VDD.n3547 Vbias 0.37318f
C12340 VDD.n3548 Vbias 0.37318f
C12341 VDD.n3549 Vbias 0.03639f
C12342 VDD.n3550 Vbias 0.03639f
C12343 VDD.n3551 Vbias 0.01836f
C12344 VDD.n3552 Vbias 0.01836f
C12345 VDD.n3553 Vbias 0.0216f
C12346 VDD.n3554 Vbias 0.03694f
C12347 VDD.t160 Vbias 0.46278f
C12348 VDD.n3555 Vbias 0.03694f
C12349 VDD.n3556 Vbias 0.04583f
C12350 VDD.n3557 Vbias 0.01151f
C12351 VDD.n3558 Vbias 0.08999f
C12352 VDD.n3559 Vbias 0.26068f
C12353 VDD.t1115 Vbias 0.12359f
C12354 VDD.n3560 Vbias 0.0361f
C12355 VDD.n3561 Vbias 0.01199f
C12356 VDD.n3562 Vbias 0.02025f
C12357 VDD.t1147 Vbias 0.12359f
C12358 VDD.n3563 Vbias 0.12814f
C12359 VDD.n3564 Vbias 0.01386f
C12360 VDD.n3565 Vbias 0.01851f
C12361 VDD.t742 Vbias 0.05773f
C12362 VDD.n3566 Vbias 0.11603f
C12363 VDD.n3567 Vbias 0.03298f
C12364 VDD.t782 Vbias 0.06426f
C12365 VDD.n3568 Vbias 0.05994f
C12366 VDD.n3569 Vbias 0.01328f
C12367 VDD.t1146 Vbias 0.12359f
C12368 VDD.n3570 Vbias 0.0361f
C12369 VDD.n3571 Vbias 0.01199f
C12370 VDD.n3572 Vbias 0.02025f
C12371 VDD.n3573 Vbias 0.07665f
C12372 VDD.n3574 Vbias 0.19471f
C12373 VDD.n3576 Vbias 0.01328f
C12374 VDD.n3577 Vbias 0.05994f
C12375 VDD.t766 Vbias 0.05693f
C12376 VDD.n3578 Vbias 0.10524f
C12377 VDD.n3579 Vbias 0.19036f
C12378 VDD.n3580 Vbias 0.55479f
C12379 VDD.n3581 Vbias 0.55479f
C12380 VDD.n3582 Vbias 1.1396f
C12381 VDD.n3583 Vbias 1.14318f
C12382 VDD.n3584 Vbias 0.55479f
C12383 VDD.t758 Vbias 0.06426f
C12384 VDD.n3585 Vbias 0.05994f
C12385 VDD.n3586 Vbias 0.01328f
C12386 VDD.t1112 Vbias 0.12359f
C12387 VDD.n3587 Vbias 0.0361f
C12388 VDD.n3588 Vbias 0.01199f
C12389 VDD.n3589 Vbias 0.02025f
C12390 VDD.n3590 Vbias 0.02099f
C12391 VDD.t1144 Vbias 0.12359f
C12392 VDD.n3591 Vbias 0.12814f
C12393 VDD.n3592 Vbias 0.01386f
C12394 VDD.n3593 Vbias 0.01851f
C12395 VDD.t760 Vbias 0.05773f
C12396 VDD.n3594 Vbias 0.11603f
C12397 VDD.n3595 Vbias 0.03298f
C12398 VDD.t792 Vbias 0.06426f
C12399 VDD.n3596 Vbias 0.05994f
C12400 VDD.n3597 Vbias 0.01328f
C12401 VDD.t1145 Vbias 0.12359f
C12402 VDD.n3598 Vbias 0.0361f
C12403 VDD.n3599 Vbias 0.01199f
C12404 VDD.n3600 Vbias 0.02025f
C12405 VDD.n3602 Vbias 0.12697f
C12406 VDD.n3603 Vbias 0.13295f
C12407 VDD.t1131 Vbias 0.12359f
C12408 VDD.n3604 Vbias 0.0361f
C12409 VDD.n3605 Vbias 0.01199f
C12410 VDD.n3606 Vbias 0.02025f
C12411 VDD.t1109 Vbias 0.12359f
C12412 VDD.n3607 Vbias 0.12814f
C12413 VDD.n3608 Vbias 0.01386f
C12414 VDD.n3609 Vbias 0.01851f
C12415 VDD.t790 Vbias 0.05773f
C12416 VDD.n3610 Vbias 0.11603f
C12417 VDD.n3611 Vbias 0.03298f
C12418 VDD.t750 Vbias 0.06426f
C12419 VDD.n3612 Vbias 0.05994f
C12420 VDD.n3613 Vbias 0.01328f
C12421 VDD.t1108 Vbias 0.12359f
C12422 VDD.n3614 Vbias 0.0361f
C12423 VDD.n3615 Vbias 0.01199f
C12424 VDD.n3616 Vbias 0.02025f
C12425 VDD.n3617 Vbias 0.07665f
C12426 VDD.n3618 Vbias 0.19471f
C12427 VDD.n3620 Vbias 0.01328f
C12428 VDD.n3621 Vbias 0.05994f
C12429 VDD.t734 Vbias 0.05693f
C12430 VDD.n3622 Vbias 0.10524f
C12431 VDD.n3623 Vbias 1.1396f
C12432 VDD.n3624 Vbias 1.14318f
C12433 VDD.n3625 Vbias 0.58347f
C12434 VDD.n3626 Vbias 1.47357f
C12435 VDD.t1117 Vbias 0.12359f
C12436 VDD.n3627 Vbias 0.0361f
C12437 VDD.n3628 Vbias 0.01199f
C12438 VDD.n3629 Vbias 0.02025f
C12439 VDD.t1150 Vbias 0.12359f
C12440 VDD.n3630 Vbias 0.12814f
C12441 VDD.n3631 Vbias 0.01386f
C12442 VDD.n3632 Vbias 0.01851f
C12443 VDD.t738 Vbias 0.05773f
C12444 VDD.n3633 Vbias 0.11603f
C12445 VDD.n3634 Vbias 0.03298f
C12446 VDD.t774 Vbias 0.06426f
C12447 VDD.n3635 Vbias 0.05994f
C12448 VDD.n3636 Vbias 0.01328f
C12449 VDD.t1148 Vbias 0.12359f
C12450 VDD.n3637 Vbias 0.0361f
C12451 VDD.n3638 Vbias 0.01199f
C12452 VDD.n3639 Vbias 0.02025f
C12453 VDD.n3640 Vbias 0.07665f
C12454 VDD.n3641 Vbias 0.19471f
C12455 VDD.n3643 Vbias 0.01328f
C12456 VDD.n3644 Vbias 0.05994f
C12457 VDD.t762 Vbias 0.05693f
C12458 VDD.n3645 Vbias 0.10524f
C12459 VDD.n3646 Vbias 1.1396f
C12460 VDD.n3647 Vbias 0.59673f
C12461 VDD.t1142 Vbias 0.12359f
C12462 VDD.n3648 Vbias 0.0361f
C12463 VDD.n3649 Vbias 0.01199f
C12464 VDD.n3650 Vbias 0.02025f
C12465 VDD.t1123 Vbias 0.12359f
C12466 VDD.n3651 Vbias 0.12814f
C12467 VDD.n3652 Vbias 0.01386f
C12468 VDD.n3653 Vbias 0.01851f
C12469 VDD.t764 Vbias 0.05773f
C12470 VDD.n3654 Vbias 0.11603f
C12471 VDD.n3655 Vbias 0.03298f
C12472 VDD.t770 Vbias 0.06426f
C12473 VDD.n3656 Vbias 0.05994f
C12474 VDD.n3657 Vbias 0.01328f
C12475 VDD.t1118 Vbias 0.12359f
C12476 VDD.n3658 Vbias 0.0361f
C12477 VDD.n3659 Vbias 0.01199f
C12478 VDD.n3660 Vbias 0.02025f
C12479 VDD.n3661 Vbias 0.07665f
C12480 VDD.n3662 Vbias 0.19471f
C12481 VDD.n3664 Vbias 0.01328f
C12482 VDD.n3665 Vbias 0.05994f
C12483 VDD.t716 Vbias 0.05693f
C12484 VDD.n3666 Vbias 0.40742f
C12485 VDD.n3668 Vbias 0.03902f
C12486 VDD.n3669 Vbias 0.03694f
C12487 VDD.n3670 Vbias 0.0216f
C12488 VDD.n3671 Vbias 0.01836f
C12489 VDD.n3672 Vbias 0.03639f
C12490 VDD.t164 Vbias 0.46278f
C12491 VDD.n3673 Vbias 0.03694f
C12492 VDD.n3674 Vbias 0.03694f
C12493 VDD.n3675 Vbias 0.0216f
C12494 VDD.n3676 Vbias 0.01836f
C12495 VDD.n3677 Vbias 0.03902f
C12496 VDD.n3678 Vbias 0.03694f
C12497 VDD.n3679 Vbias 0.07027f
C12498 VDD.t584 Vbias 0.0169f
C12499 VDD.t683 Vbias 0.0169f
C12500 VDD.n3680 Vbias 0.07902f
C12501 VDD.t165 Vbias 0.0169f
C12502 VDD.t163 Vbias 0.0169f
C12503 VDD.n3681 Vbias 0.07902f
C12504 VDD.n3682 Vbias 0.03902f
C12505 VDD.n3683 Vbias 0.03694f
C12506 VDD.n3684 Vbias 0.03902f
C12507 VDD.n3685 Vbias 0.03639f
C12508 VDD.n3686 Vbias 0.03639f
C12509 VDD.n3687 Vbias 0.03694f
C12510 VDD.n3688 Vbias 0.0216f
C12511 VDD.n3689 Vbias 0.01836f
C12512 VDD.n3690 Vbias 0.03639f
C12513 VDD.n3691 Vbias 0.01836f
C12514 VDD.n3692 Vbias 0.03639f
C12515 VDD.n3693 Vbias 0.37318f
C12516 VDD.n3694 Vbias 0.37318f
C12517 VDD.n3695 Vbias 0.01836f
C12518 VDD.n3696 Vbias 0.01836f
C12519 VDD.n3697 Vbias 0.0216f
C12520 VDD.n3698 Vbias 0.03694f
C12521 VDD.t1094 Vbias 0.46278f
C12522 VDD.n3699 Vbias 0.03694f
C12523 VDD.n3700 Vbias 0.03694f
C12524 VDD.n3701 Vbias 0.06648f
C12525 VDD.n3702 Vbias 0.03639f
C12526 VDD.t246 Vbias 0.46278f
C12527 VDD.n3703 Vbias 0.03694f
C12528 VDD.n3704 Vbias 0.03694f
C12529 VDD.n3705 Vbias 0.0216f
C12530 VDD.n3706 Vbias 0.01836f
C12531 VDD.t1095 Vbias 0.017f
C12532 VDD.n3707 Vbias 0.05322f
C12533 VDD.n3708 Vbias 0.01309f
C12534 VDD.n3709 Vbias 0.01699f
C12535 VDD.n3710 Vbias 0.03902f
C12536 VDD.n3711 Vbias 0.03694f
C12537 VDD.n3712 Vbias 0.0216f
C12538 VDD.n3713 Vbias 0.01836f
C12539 VDD.n3714 Vbias 0.03639f
C12540 VDD.t550 Vbias 0.46278f
C12541 VDD.n3715 Vbias 0.03694f
C12542 VDD.n3716 Vbias 0.03694f
C12543 VDD.n3717 Vbias 0.0216f
C12544 VDD.n3718 Vbias 0.01836f
C12545 VDD.t247 Vbias 0.0169f
C12546 VDD.t552 Vbias 0.0169f
C12547 VDD.n3719 Vbias 0.07902f
C12548 VDD.t684 Vbias 0.0169f
C12549 VDD.t551 Vbias 0.0169f
C12550 VDD.n3720 Vbias 0.07902f
C12551 VDD.n3721 Vbias 0.03023f
C12552 VDD.n3722 Vbias 0.01699f
C12553 VDD.n3723 Vbias 0.03902f
C12554 VDD.n3724 Vbias 0.03694f
C12555 VDD.n3725 Vbias 0.0216f
C12556 VDD.n3726 Vbias 0.01836f
C12557 VDD.n3727 Vbias 0.03639f
C12558 VDD.t35 Vbias 0.46278f
C12559 VDD.n3728 Vbias 0.03694f
C12560 VDD.n3729 Vbias 0.03694f
C12561 VDD.n3730 Vbias 0.0216f
C12562 VDD.n3731 Vbias 0.01836f
C12563 VDD.t36 Vbias 0.017f
C12564 VDD.t771 Vbias 0.017f
C12565 VDD.n3732 Vbias 0.09713f
C12566 VDD.n3733 Vbias 0.01914f
C12567 VDD.n3734 Vbias 0.03902f
C12568 VDD.n3735 Vbias 0.03694f
C12569 VDD.n3736 Vbias 0.0216f
C12570 VDD.n3737 Vbias 0.01836f
C12571 VDD.n3738 Vbias 0.03639f
C12572 VDD.t633 Vbias 0.46278f
C12573 VDD.n3739 Vbias 0.03694f
C12574 VDD.n3740 Vbias 0.03694f
C12575 VDD.n3741 Vbias 0.0216f
C12576 VDD.n3742 Vbias 0.01836f
C12577 VDD.n3743 Vbias 0.02305f
C12578 VDD.n3744 Vbias 0.03902f
C12579 VDD.n3745 Vbias 0.03694f
C12580 VDD.n3746 Vbias 0.0216f
C12581 VDD.n3747 Vbias 0.01836f
C12582 VDD.n3748 Vbias 0.03639f
C12583 VDD.t347 Vbias 0.46278f
C12584 VDD.n3749 Vbias 0.03694f
C12585 VDD.n3750 Vbias 0.03694f
C12586 VDD.n3751 Vbias 0.0216f
C12587 VDD.n3752 Vbias 0.01836f
C12588 VDD.t909 Vbias 0.0169f
C12589 VDD.t537 Vbias 0.0169f
C12590 VDD.n3753 Vbias 0.07902f
C12591 VDD.t634 Vbias 0.0169f
C12592 VDD.t348 Vbias 0.0169f
C12593 VDD.n3754 Vbias 0.07902f
C12594 VDD.n3755 Vbias 0.03023f
C12595 VDD.n3756 Vbias 0.01699f
C12596 VDD.n3757 Vbias 0.03902f
C12597 VDD.n3758 Vbias 0.03694f
C12598 VDD.n3759 Vbias 0.0216f
C12599 VDD.n3760 Vbias 0.01836f
C12600 VDD.n3761 Vbias 0.01836f
C12601 VDD.n3762 Vbias 0.03639f
C12602 VDD.n3763 Vbias 0.50118f
C12603 VDD.n3764 Vbias 0.03639f
C12604 VDD.n3765 Vbias 0.03694f
C12605 VDD.n3766 Vbias 0.04583f
C12606 VDD.n3767 Vbias 0.03902f
C12607 VDD.n3768 Vbias 0.01836f
C12608 VDD.n3769 Vbias 0.03639f
C12609 VDD.n3770 Vbias 0.37318f
C12610 VDD.n3771 Vbias 0.01836f
C12611 VDD.n3772 Vbias 0.03639f
C12612 VDD.n3773 Vbias 0.37318f
C12613 VDD.n3774 Vbias 0.03639f
C12614 VDD.n3775 Vbias 0.03694f
C12615 VDD.n3776 Vbias 0.04583f
C12616 VDD.n3777 Vbias 0.03902f
C12617 VDD.n3778 Vbias 0.01836f
C12618 VDD.n3779 Vbias 0.03639f
C12619 VDD.n3780 Vbias 0.37318f
C12620 VDD.n3781 Vbias 0.01836f
C12621 VDD.n3782 Vbias 0.03639f
C12622 VDD.n3783 Vbias 0.37318f
C12623 VDD.n3784 Vbias 0.03639f
C12624 VDD.n3785 Vbias 0.03694f
C12625 VDD.n3786 Vbias 0.04583f
C12626 VDD.n3787 Vbias 0.03902f
C12627 VDD.n3788 Vbias 0.01836f
C12628 VDD.n3789 Vbias 0.03639f
C12629 VDD.n3790 Vbias 0.50118f
C12630 VDD.n3791 Vbias 0.01836f
C12631 VDD.n3792 Vbias 0.03639f
C12632 VDD.n3793 Vbias 0.50118f
C12633 VDD.n3794 Vbias 0.03639f
C12634 VDD.n3795 Vbias 0.03694f
C12635 VDD.n3796 Vbias 0.04583f
C12636 VDD.n3797 Vbias 0.03902f
C12637 VDD.n3798 Vbias 0.01836f
C12638 VDD.n3799 Vbias 0.03639f
C12639 VDD.n3800 Vbias 0.37318f
C12640 VDD.n3801 Vbias 0.01836f
C12641 VDD.n3802 Vbias 0.03639f
C12642 VDD.n3803 Vbias 0.37318f
C12643 VDD.n3804 Vbias 0.03639f
C12644 VDD.n3805 Vbias 0.03694f
C12645 VDD.n3806 Vbias 0.04583f
C12646 VDD.n3807 Vbias 0.03902f
C12647 VDD.n3808 Vbias 0.01836f
C12648 VDD.n3809 Vbias 0.03639f
C12649 VDD.n3810 Vbias 0.50118f
C12650 VDD.n3811 Vbias 0.50118f
C12651 VDD.n3812 Vbias 0.03639f
C12652 VDD.n3813 Vbias 0.01999f
C12653 VDD.n3814 Vbias 0.0216f
C12654 VDD.n3815 Vbias 0.01999f
C12655 VDD.n3816 Vbias 0.03639f
C12656 VDD.n3817 Vbias 0.50118f
C12657 VDD.n3818 Vbias 0.50118f
C12658 VDD.n3819 Vbias 0.03639f
C12659 VDD.n3820 Vbias 0.03639f
C12660 VDD.n3821 Vbias 0.01836f
C12661 VDD.n3822 Vbias 0.01836f
C12662 VDD.n3823 Vbias 0.0216f
C12663 VDD.n3824 Vbias 0.03694f
C12664 VDD.t162 Vbias 0.46278f
C12665 VDD.n3825 Vbias 0.03694f
C12666 VDD.n3826 Vbias 0.04583f
C12667 VDD.n3827 Vbias 0.01699f
C12668 VDD.n3828 Vbias 0.03023f
C12669 VDD.n3829 Vbias 0.02225f
C12670 VDD.n3830 Vbias 0.04583f
C12671 VDD.n3831 Vbias 0.03902f
C12672 VDD.n3832 Vbias 0.01836f
C12673 VDD.n3833 Vbias 0.03639f
C12674 VDD.n3834 Vbias 0.37318f
C12675 VDD.n3835 Vbias 0.01836f
C12676 VDD.n3836 Vbias 0.03639f
C12677 VDD.n3837 Vbias 0.37318f
C12678 VDD.n3838 Vbias 0.03639f
C12679 VDD.n3839 Vbias 0.03694f
C12680 VDD.n3840 Vbias 0.04583f
C12681 VDD.n3841 Vbias 0.03902f
C12682 VDD.n3842 Vbias 0.01836f
C12683 VDD.n3843 Vbias 0.03639f
C12684 VDD.n3844 Vbias 0.50118f
C12685 VDD.n3845 Vbias 0.01836f
C12686 VDD.n3846 Vbias 0.03639f
C12687 VDD.n3847 Vbias 0.50118f
C12688 VDD.n3848 Vbias 0.03639f
C12689 VDD.n3849 Vbias 0.03694f
C12690 VDD.n3850 Vbias 0.04583f
C12691 VDD.n3851 Vbias 0.03902f
C12692 VDD.n3852 Vbias 0.01836f
C12693 VDD.n3853 Vbias 0.03639f
C12694 VDD.n3854 Vbias 0.37318f
C12695 VDD.n3855 Vbias 0.01836f
C12696 VDD.n3856 Vbias 0.03639f
C12697 VDD.n3857 Vbias 0.37318f
C12698 VDD.n3858 Vbias 0.03639f
C12699 VDD.n3859 Vbias 0.03694f
C12700 VDD.n3860 Vbias 0.04583f
C12701 VDD.n3861 Vbias 0.03902f
C12702 VDD.n3862 Vbias 0.01836f
C12703 VDD.n3863 Vbias 0.03639f
C12704 VDD.n3864 Vbias 0.37318f
C12705 VDD.n3865 Vbias 0.01836f
C12706 VDD.n3866 Vbias 0.03639f
C12707 VDD.n3867 Vbias 0.37318f
C12708 VDD.n3868 Vbias 0.03639f
C12709 VDD.n3869 Vbias 0.03694f
C12710 VDD.n3870 Vbias 0.04583f
C12711 VDD.n3871 Vbias 0.03902f
C12712 VDD.n3872 Vbias 0.01836f
C12713 VDD.n3873 Vbias 0.03639f
C12714 VDD.n3874 Vbias 0.50118f
C12715 VDD.n3875 Vbias 0.50118f
C12716 VDD.n3876 Vbias 0.03639f
C12717 VDD.n3877 Vbias 0.01999f
C12718 VDD.n3878 Vbias 0.06648f
C12719 VDD.n3879 Vbias 0.01309f
C12720 VDD.n3880 Vbias 0.11022f
C12721 VDD.n3881 Vbias 0.01699f
C12722 VDD.n3882 Vbias 0.03902f
C12723 VDD.n3883 Vbias 0.03694f
C12724 VDD.n3884 Vbias 0.0216f
C12725 VDD.n3885 Vbias 0.01836f
C12726 VDD.n3886 Vbias 0.01836f
C12727 VDD.n3887 Vbias 0.03639f
C12728 VDD.n3888 Vbias 0.50118f
C12729 VDD.n3889 Vbias 0.03639f
C12730 VDD.n3890 Vbias 0.03694f
C12731 VDD.n3891 Vbias 0.04583f
C12732 VDD.n3892 Vbias 0.03902f
C12733 VDD.n3893 Vbias 0.01836f
C12734 VDD.n3894 Vbias 0.03639f
C12735 VDD.n3895 Vbias 0.37318f
C12736 VDD.n3896 Vbias 0.01836f
C12737 VDD.n3897 Vbias 0.03639f
C12738 VDD.n3898 Vbias 0.37318f
C12739 VDD.n3899 Vbias 0.03639f
C12740 VDD.n3900 Vbias 0.03694f
C12741 VDD.n3901 Vbias 0.04583f
C12742 VDD.n3902 Vbias 0.03902f
C12743 VDD.n3903 Vbias 0.01836f
C12744 VDD.n3904 Vbias 0.03639f
C12745 VDD.n3905 Vbias 0.37318f
C12746 VDD.n3906 Vbias 0.01836f
C12747 VDD.n3907 Vbias 0.03639f
C12748 VDD.n3908 Vbias 0.37318f
C12749 VDD.n3909 Vbias 0.03639f
C12750 VDD.n3910 Vbias 0.03694f
C12751 VDD.n3911 Vbias 0.04583f
C12752 VDD.n3912 Vbias 0.03902f
C12753 VDD.n3913 Vbias 0.01836f
C12754 VDD.n3914 Vbias 0.03639f
C12755 VDD.n3915 Vbias 0.50118f
C12756 VDD.n3916 Vbias 0.01836f
C12757 VDD.n3917 Vbias 0.03639f
C12758 VDD.n3918 Vbias 0.50118f
C12759 VDD.n3919 Vbias 0.03639f
C12760 VDD.n3920 Vbias 0.03694f
C12761 VDD.n3921 Vbias 0.04583f
C12762 VDD.n3922 Vbias 0.03902f
C12763 VDD.n3923 Vbias 0.01836f
C12764 VDD.n3924 Vbias 0.03639f
C12765 VDD.n3925 Vbias 0.37318f
C12766 VDD.n3926 Vbias 0.01836f
C12767 VDD.n3927 Vbias 0.03639f
C12768 VDD.n3928 Vbias 0.37318f
C12769 VDD.n3929 Vbias 0.03639f
C12770 VDD.n3930 Vbias 0.03694f
C12771 VDD.n3931 Vbias 0.04583f
C12772 VDD.n3932 Vbias 0.03902f
C12773 VDD.n3933 Vbias 0.01836f
C12774 VDD.n3934 Vbias 0.03639f
C12775 VDD.n3935 Vbias 0.50118f
C12776 VDD.n3936 Vbias 0.50118f
C12777 VDD.n3937 Vbias 0.03639f
C12778 VDD.n3938 Vbias 0.01999f
C12779 VDD.n3939 Vbias 0.0216f
C12780 VDD.n3940 Vbias 0.01999f
C12781 VDD.n3941 Vbias 0.03639f
C12782 VDD.n3942 Vbias 0.50118f
C12783 VDD.n3943 Vbias 0.50118f
C12784 VDD.n3944 Vbias 0.03639f
C12785 VDD.n3945 Vbias 0.03639f
C12786 VDD.n3946 Vbias 0.01836f
C12787 VDD.n3947 Vbias 0.01836f
C12788 VDD.n3948 Vbias 0.0216f
C12789 VDD.n3949 Vbias 0.03694f
C12790 VDD.t510 Vbias 0.46278f
C12791 VDD.n3950 Vbias 0.03694f
C12792 VDD.n3951 Vbias 0.04583f
C12793 VDD.n3952 Vbias 0.01699f
C12794 VDD.n3953 Vbias 0.03023f
C12795 VDD.n3954 Vbias 0.02225f
C12796 VDD.n3955 Vbias 0.04583f
C12797 VDD.n3956 Vbias 0.03902f
C12798 VDD.n3957 Vbias 0.01836f
C12799 VDD.n3958 Vbias 0.03639f
C12800 VDD.n3959 Vbias 0.37318f
C12801 VDD.n3960 Vbias 0.01836f
C12802 VDD.n3961 Vbias 0.03639f
C12803 VDD.n3962 Vbias 0.37318f
C12804 VDD.n3963 Vbias 0.03639f
C12805 VDD.n3964 Vbias 0.03694f
C12806 VDD.n3965 Vbias 0.04583f
C12807 VDD.n3966 Vbias 0.03902f
C12808 VDD.n3967 Vbias 0.01836f
C12809 VDD.n3968 Vbias 0.03639f
C12810 VDD.n3969 Vbias 0.50118f
C12811 VDD.n3970 Vbias 0.01836f
C12812 VDD.n3971 Vbias 0.03639f
C12813 VDD.n3972 Vbias 0.50118f
C12814 VDD.n3973 Vbias 0.03639f
C12815 VDD.n3974 Vbias 0.03694f
C12816 VDD.n3975 Vbias 0.04583f
C12817 VDD.n3976 Vbias 0.03902f
C12818 VDD.n3977 Vbias 0.01836f
C12819 VDD.n3978 Vbias 0.03639f
C12820 VDD.n3979 Vbias 0.37318f
C12821 VDD.n3980 Vbias 0.01836f
C12822 VDD.n3981 Vbias 0.03639f
C12823 VDD.n3982 Vbias 0.37318f
C12824 VDD.n3983 Vbias 0.03639f
C12825 VDD.n3984 Vbias 0.03694f
C12826 VDD.n3985 Vbias 0.04583f
C12827 VDD.n3986 Vbias 0.03902f
C12828 VDD.n3987 Vbias 0.01836f
C12829 VDD.n3988 Vbias 0.03639f
C12830 VDD.n3989 Vbias 0.37318f
C12831 VDD.n3990 Vbias 0.01836f
C12832 VDD.n3991 Vbias 0.03639f
C12833 VDD.n3992 Vbias 0.37318f
C12834 VDD.n3993 Vbias 0.03639f
C12835 VDD.n3994 Vbias 0.03694f
C12836 VDD.n3995 Vbias 0.04583f
C12837 VDD.n3996 Vbias 0.03902f
C12838 VDD.n3997 Vbias 0.01836f
C12839 VDD.n3998 Vbias 0.03639f
C12840 VDD.n3999 Vbias 0.50118f
C12841 VDD.n4000 Vbias 0.50118f
C12842 VDD.n4001 Vbias 0.03639f
C12843 VDD.n4002 Vbias 0.01999f
C12844 VDD.n4003 Vbias 0.06648f
C12845 VDD.n4004 Vbias 0.01309f
C12846 VDD.n4005 Vbias 0.11022f
C12847 VDD.n4006 Vbias 0.01699f
C12848 VDD.n4007 Vbias 0.03902f
C12849 VDD.n4008 Vbias 0.03694f
C12850 VDD.n4009 Vbias 0.0216f
C12851 VDD.n4010 Vbias 0.01836f
C12852 VDD.n4011 Vbias 0.01836f
C12853 VDD.n4012 Vbias 0.03639f
C12854 VDD.n4013 Vbias 0.50118f
C12855 VDD.n4014 Vbias 0.03639f
C12856 VDD.n4015 Vbias 0.03694f
C12857 VDD.n4016 Vbias 0.04583f
C12858 VDD.n4017 Vbias 0.03902f
C12859 VDD.n4018 Vbias 0.01836f
C12860 VDD.n4019 Vbias 0.03639f
C12861 VDD.n4020 Vbias 0.37318f
C12862 VDD.n4021 Vbias 0.01836f
C12863 VDD.n4022 Vbias 0.03639f
C12864 VDD.n4023 Vbias 0.37318f
C12865 VDD.n4024 Vbias 0.03639f
C12866 VDD.n4025 Vbias 0.03694f
C12867 VDD.n4026 Vbias 0.04583f
C12868 VDD.n4027 Vbias 0.03902f
C12869 VDD.n4028 Vbias 0.01836f
C12870 VDD.n4029 Vbias 0.03639f
C12871 VDD.n4030 Vbias 0.37318f
C12872 VDD.n4031 Vbias 0.01836f
C12873 VDD.n4032 Vbias 0.03639f
C12874 VDD.n4033 Vbias 0.37318f
C12875 VDD.n4034 Vbias 0.03639f
C12876 VDD.n4035 Vbias 0.03694f
C12877 VDD.n4036 Vbias 0.04583f
C12878 VDD.n4037 Vbias 0.03902f
C12879 VDD.n4038 Vbias 0.01836f
C12880 VDD.n4039 Vbias 0.03639f
C12881 VDD.n4040 Vbias 0.50118f
C12882 VDD.n4041 Vbias 0.01836f
C12883 VDD.n4042 Vbias 0.03639f
C12884 VDD.n4043 Vbias 0.50118f
C12885 VDD.n4044 Vbias 0.03639f
C12886 VDD.n4045 Vbias 0.03694f
C12887 VDD.n4046 Vbias 0.04583f
C12888 VDD.n4047 Vbias 0.03902f
C12889 VDD.n4048 Vbias 0.01836f
C12890 VDD.n4049 Vbias 0.03639f
C12891 VDD.n4050 Vbias 0.37318f
C12892 VDD.n4051 Vbias 0.01836f
C12893 VDD.n4052 Vbias 0.03639f
C12894 VDD.n4053 Vbias 0.37318f
C12895 VDD.n4054 Vbias 0.03639f
C12896 VDD.n4055 Vbias 0.03694f
C12897 VDD.n4056 Vbias 0.04583f
C12898 VDD.n4057 Vbias 0.03902f
C12899 VDD.n4058 Vbias 0.01836f
C12900 VDD.n4059 Vbias 0.03639f
C12901 VDD.n4060 Vbias 0.50118f
C12902 VDD.n4061 Vbias 0.50118f
C12903 VDD.n4062 Vbias 0.03639f
C12904 VDD.n4063 Vbias 0.01999f
C12905 VDD.n4064 Vbias 0.0216f
C12906 VDD.n4065 Vbias 0.01999f
C12907 VDD.n4066 Vbias 0.03639f
C12908 VDD.n4067 Vbias 0.50118f
C12909 VDD.n4068 Vbias 0.50118f
C12910 VDD.n4069 Vbias 0.03639f
C12911 VDD.n4070 Vbias 0.03639f
C12912 VDD.n4071 Vbias 0.01836f
C12913 VDD.n4072 Vbias 0.01836f
C12914 VDD.n4073 Vbias 0.0216f
C12915 VDD.n4074 Vbias 0.03694f
C12916 VDD.t525 Vbias 0.46278f
C12917 VDD.n4075 Vbias 0.03694f
C12918 VDD.n4076 Vbias 0.04583f
C12919 VDD.n4077 Vbias 0.01699f
C12920 VDD.n4078 Vbias 0.03023f
C12921 VDD.n4079 Vbias 0.02225f
C12922 VDD.n4080 Vbias 0.04583f
C12923 VDD.n4081 Vbias 0.03902f
C12924 VDD.n4082 Vbias 0.01836f
C12925 VDD.n4083 Vbias 0.03639f
C12926 VDD.n4084 Vbias 0.37318f
C12927 VDD.n4085 Vbias 0.01836f
C12928 VDD.n4086 Vbias 0.03639f
C12929 VDD.n4087 Vbias 0.37318f
C12930 VDD.n4088 Vbias 0.03639f
C12931 VDD.n4089 Vbias 0.03694f
C12932 VDD.n4090 Vbias 0.04583f
C12933 VDD.n4091 Vbias 0.03902f
C12934 VDD.n4092 Vbias 0.01836f
C12935 VDD.n4093 Vbias 0.03639f
C12936 VDD.n4094 Vbias 0.50118f
C12937 VDD.n4095 Vbias 0.01836f
C12938 VDD.n4096 Vbias 0.03639f
C12939 VDD.n4097 Vbias 0.50118f
C12940 VDD.n4098 Vbias 0.03639f
C12941 VDD.n4099 Vbias 0.03694f
C12942 VDD.n4100 Vbias 0.04583f
C12943 VDD.n4101 Vbias 0.03902f
C12944 VDD.n4102 Vbias 0.01836f
C12945 VDD.n4103 Vbias 0.03639f
C12946 VDD.n4104 Vbias 0.37318f
C12947 VDD.n4105 Vbias 0.01836f
C12948 VDD.n4106 Vbias 0.03639f
C12949 VDD.n4107 Vbias 0.37318f
C12950 VDD.n4108 Vbias 0.03639f
C12951 VDD.n4109 Vbias 0.03694f
C12952 VDD.n4110 Vbias 0.04583f
C12953 VDD.n4111 Vbias 0.03902f
C12954 VDD.n4112 Vbias 0.01836f
C12955 VDD.n4113 Vbias 0.03639f
C12956 VDD.n4114 Vbias 0.37318f
C12957 VDD.n4115 Vbias 0.01836f
C12958 VDD.n4116 Vbias 0.03639f
C12959 VDD.n4117 Vbias 0.37318f
C12960 VDD.n4118 Vbias 0.03639f
C12961 VDD.n4119 Vbias 0.03694f
C12962 VDD.n4120 Vbias 0.04583f
C12963 VDD.n4121 Vbias 0.03902f
C12964 VDD.n4122 Vbias 0.01836f
C12965 VDD.n4123 Vbias 0.03639f
C12966 VDD.n4124 Vbias 0.50118f
C12967 VDD.n4125 Vbias 0.50118f
C12968 VDD.n4126 Vbias 0.03639f
C12969 VDD.n4127 Vbias 0.01999f
C12970 VDD.n4128 Vbias 0.06648f
C12971 VDD.n4129 Vbias 0.01309f
C12972 VDD.n4130 Vbias 0.11022f
C12973 VDD.n4131 Vbias 0.01699f
C12974 VDD.n4132 Vbias 0.03902f
C12975 VDD.n4133 Vbias 0.03694f
C12976 VDD.n4134 Vbias 0.0216f
C12977 VDD.n4135 Vbias 0.01836f
C12978 VDD.n4136 Vbias 0.01836f
C12979 VDD.n4137 Vbias 0.03639f
C12980 VDD.n4138 Vbias 0.50118f
C12981 VDD.n4139 Vbias 0.03639f
C12982 VDD.n4140 Vbias 0.03694f
C12983 VDD.n4141 Vbias 0.04583f
C12984 VDD.n4142 Vbias 0.03902f
C12985 VDD.n4143 Vbias 0.01836f
C12986 VDD.n4144 Vbias 0.03639f
C12987 VDD.n4145 Vbias 0.37318f
C12988 VDD.n4146 Vbias 0.01836f
C12989 VDD.n4147 Vbias 0.03639f
C12990 VDD.n4148 Vbias 0.37318f
C12991 VDD.n4149 Vbias 0.03639f
C12992 VDD.n4150 Vbias 0.03694f
C12993 VDD.n4151 Vbias 0.04583f
C12994 VDD.n4152 Vbias 0.03902f
C12995 VDD.n4153 Vbias 0.01836f
C12996 VDD.n4154 Vbias 0.03639f
C12997 VDD.n4155 Vbias 0.37318f
C12998 VDD.n4156 Vbias 0.01836f
C12999 VDD.n4157 Vbias 0.03639f
C13000 VDD.n4158 Vbias 0.37318f
C13001 VDD.n4159 Vbias 0.03639f
C13002 VDD.n4160 Vbias 0.03694f
C13003 VDD.n4161 Vbias 0.04583f
C13004 VDD.n4162 Vbias 0.03902f
C13005 VDD.n4163 Vbias 0.01836f
C13006 VDD.n4164 Vbias 0.03639f
C13007 VDD.n4165 Vbias 0.50118f
C13008 VDD.n4166 Vbias 0.01836f
C13009 VDD.n4167 Vbias 0.03639f
C13010 VDD.n4168 Vbias 0.50118f
C13011 VDD.n4169 Vbias 0.03639f
C13012 VDD.n4170 Vbias 0.03694f
C13013 VDD.n4171 Vbias 0.04583f
C13014 VDD.n4172 Vbias 0.03902f
C13015 VDD.n4173 Vbias 0.01836f
C13016 VDD.n4174 Vbias 0.03639f
C13017 VDD.n4175 Vbias 0.37318f
C13018 VDD.n4176 Vbias 0.01836f
C13019 VDD.n4177 Vbias 0.03639f
C13020 VDD.n4178 Vbias 0.37318f
C13021 VDD.n4179 Vbias 0.03639f
C13022 VDD.n4180 Vbias 0.03694f
C13023 VDD.n4181 Vbias 0.04583f
C13024 VDD.n4182 Vbias 0.03902f
C13025 VDD.n4183 Vbias 0.01836f
C13026 VDD.n4184 Vbias 0.03639f
C13027 VDD.n4185 Vbias 0.50118f
C13028 VDD.n4186 Vbias 0.50118f
C13029 VDD.n4187 Vbias 0.03639f
C13030 VDD.n4188 Vbias 0.01999f
C13031 VDD.n4189 Vbias 0.0216f
C13032 VDD.n4190 Vbias 0.01999f
C13033 VDD.n4191 Vbias 0.03639f
C13034 VDD.n4192 Vbias 0.50118f
C13035 VDD.n4193 Vbias 0.50118f
C13036 VDD.n4194 Vbias 0.03639f
C13037 VDD.n4195 Vbias 0.03639f
C13038 VDD.n4196 Vbias 0.01836f
C13039 VDD.n4197 Vbias 0.01836f
C13040 VDD.n4198 Vbias 0.0216f
C13041 VDD.n4199 Vbias 0.03694f
C13042 VDD.t438 Vbias 0.46278f
C13043 VDD.n4200 Vbias 0.03694f
C13044 VDD.n4201 Vbias 0.04583f
C13045 VDD.n4202 Vbias 0.01699f
C13046 VDD.n4203 Vbias 0.03023f
C13047 VDD.n4204 Vbias 0.02225f
C13048 VDD.n4205 Vbias 0.04583f
C13049 VDD.n4206 Vbias 0.03902f
C13050 VDD.n4207 Vbias 0.01836f
C13051 VDD.n4208 Vbias 0.03639f
C13052 VDD.n4209 Vbias 0.37318f
C13053 VDD.n4210 Vbias 0.01836f
C13054 VDD.n4211 Vbias 0.03639f
C13055 VDD.n4212 Vbias 0.37318f
C13056 VDD.n4213 Vbias 0.03639f
C13057 VDD.n4214 Vbias 0.03694f
C13058 VDD.n4215 Vbias 0.04583f
C13059 VDD.n4216 Vbias 0.03902f
C13060 VDD.n4217 Vbias 0.01836f
C13061 VDD.n4218 Vbias 0.03639f
C13062 VDD.n4219 Vbias 0.50118f
C13063 VDD.n4220 Vbias 0.01836f
C13064 VDD.n4221 Vbias 0.03639f
C13065 VDD.n4222 Vbias 0.50118f
C13066 VDD.n4223 Vbias 0.03639f
C13067 VDD.n4224 Vbias 0.03694f
C13068 VDD.n4225 Vbias 0.04583f
C13069 VDD.n4226 Vbias 0.03902f
C13070 VDD.n4227 Vbias 0.01836f
C13071 VDD.n4228 Vbias 0.03639f
C13072 VDD.n4229 Vbias 0.37318f
C13073 VDD.n4230 Vbias 0.01836f
C13074 VDD.n4231 Vbias 0.03639f
C13075 VDD.n4232 Vbias 0.37318f
C13076 VDD.n4233 Vbias 0.03639f
C13077 VDD.n4234 Vbias 0.03694f
C13078 VDD.n4235 Vbias 0.04583f
C13079 VDD.n4236 Vbias 0.03902f
C13080 VDD.n4237 Vbias 0.01836f
C13081 VDD.n4238 Vbias 0.03639f
C13082 VDD.n4239 Vbias 0.37318f
C13083 VDD.n4240 Vbias 0.01836f
C13084 VDD.n4241 Vbias 0.03639f
C13085 VDD.n4242 Vbias 0.37318f
C13086 VDD.n4243 Vbias 0.03639f
C13087 VDD.n4244 Vbias 0.03694f
C13088 VDD.n4245 Vbias 0.04583f
C13089 VDD.n4246 Vbias 0.03902f
C13090 VDD.n4247 Vbias 0.01836f
C13091 VDD.n4248 Vbias 0.03639f
C13092 VDD.n4249 Vbias 0.50118f
C13093 VDD.n4250 Vbias 0.50118f
C13094 VDD.n4251 Vbias 0.03639f
C13095 VDD.n4252 Vbias 0.01999f
C13096 VDD.n4253 Vbias 0.06648f
C13097 VDD.n4254 Vbias 0.01309f
C13098 VDD.n4255 Vbias 0.11022f
C13099 VDD.n4256 Vbias 0.01699f
C13100 VDD.n4257 Vbias 0.03902f
C13101 VDD.n4258 Vbias 0.03694f
C13102 VDD.n4259 Vbias 0.0216f
C13103 VDD.n4260 Vbias 0.01836f
C13104 VDD.n4261 Vbias 0.01836f
C13105 VDD.n4262 Vbias 0.03639f
C13106 VDD.n4263 Vbias 0.50118f
C13107 VDD.n4264 Vbias 0.03639f
C13108 VDD.n4265 Vbias 0.03694f
C13109 VDD.n4266 Vbias 0.04583f
C13110 VDD.n4267 Vbias 0.03902f
C13111 VDD.n4268 Vbias 0.01836f
C13112 VDD.n4269 Vbias 0.03639f
C13113 VDD.n4270 Vbias 0.37318f
C13114 VDD.n4271 Vbias 0.01836f
C13115 VDD.n4272 Vbias 0.03639f
C13116 VDD.n4273 Vbias 0.37318f
C13117 VDD.n4274 Vbias 0.03639f
C13118 VDD.n4275 Vbias 0.03694f
C13119 VDD.n4276 Vbias 0.04583f
C13120 VDD.n4277 Vbias 0.03902f
C13121 VDD.n4278 Vbias 0.01836f
C13122 VDD.n4279 Vbias 0.03639f
C13123 VDD.n4280 Vbias 0.37318f
C13124 VDD.n4281 Vbias 0.01836f
C13125 VDD.n4282 Vbias 0.03639f
C13126 VDD.n4283 Vbias 0.37318f
C13127 VDD.n4284 Vbias 0.03639f
C13128 VDD.n4285 Vbias 0.03694f
C13129 VDD.n4286 Vbias 0.04583f
C13130 VDD.n4287 Vbias 0.03902f
C13131 VDD.n4288 Vbias 0.01836f
C13132 VDD.n4289 Vbias 0.03639f
C13133 VDD.n4290 Vbias 0.50118f
C13134 VDD.n4291 Vbias 0.01836f
C13135 VDD.n4292 Vbias 0.03639f
C13136 VDD.n4293 Vbias 0.50118f
C13137 VDD.n4294 Vbias 0.03639f
C13138 VDD.n4295 Vbias 0.03694f
C13139 VDD.n4296 Vbias 0.04583f
C13140 VDD.n4297 Vbias 0.03902f
C13141 VDD.n4298 Vbias 0.01836f
C13142 VDD.n4299 Vbias 0.03639f
C13143 VDD.n4300 Vbias 0.37318f
C13144 VDD.n4301 Vbias 0.01836f
C13145 VDD.n4302 Vbias 0.03639f
C13146 VDD.n4303 Vbias 0.37318f
C13147 VDD.n4304 Vbias 0.03639f
C13148 VDD.n4305 Vbias 0.03694f
C13149 VDD.n4306 Vbias 0.04583f
C13150 VDD.n4307 Vbias 0.03902f
C13151 VDD.n4308 Vbias 0.01836f
C13152 VDD.n4309 Vbias 0.03639f
C13153 VDD.n4310 Vbias 0.50118f
C13154 VDD.n4311 Vbias 0.50118f
C13155 VDD.n4312 Vbias 0.03639f
C13156 VDD.n4313 Vbias 0.01999f
C13157 VDD.n4314 Vbias 0.0216f
C13158 VDD.n4315 Vbias 0.01999f
C13159 VDD.n4316 Vbias 0.03639f
C13160 VDD.n4317 Vbias 0.50118f
C13161 VDD.n4318 Vbias 0.50118f
C13162 VDD.n4319 Vbias 0.03639f
C13163 VDD.n4320 Vbias 0.03639f
C13164 VDD.n4321 Vbias 0.01836f
C13165 VDD.n4322 Vbias 0.01836f
C13166 VDD.n4323 Vbias 0.0216f
C13167 VDD.n4324 Vbias 0.03694f
C13168 VDD.t236 Vbias 0.46278f
C13169 VDD.n4325 Vbias 0.03694f
C13170 VDD.n4326 Vbias 0.04583f
C13171 VDD.n4327 Vbias 0.01699f
C13172 VDD.n4328 Vbias 0.03023f
C13173 VDD.n4329 Vbias 0.02225f
C13174 VDD.n4330 Vbias 0.04583f
C13175 VDD.n4331 Vbias 0.03902f
C13176 VDD.n4332 Vbias 0.01836f
C13177 VDD.n4333 Vbias 0.03639f
C13178 VDD.n4334 Vbias 0.37318f
C13179 VDD.n4335 Vbias 0.01836f
C13180 VDD.n4336 Vbias 0.03639f
C13181 VDD.n4337 Vbias 0.37318f
C13182 VDD.n4338 Vbias 0.03639f
C13183 VDD.n4339 Vbias 0.03694f
C13184 VDD.n4340 Vbias 0.04583f
C13185 VDD.n4341 Vbias 0.03902f
C13186 VDD.n4342 Vbias 0.01836f
C13187 VDD.n4343 Vbias 0.03639f
C13188 VDD.n4344 Vbias 0.50118f
C13189 VDD.n4345 Vbias 0.01836f
C13190 VDD.n4346 Vbias 0.03639f
C13191 VDD.n4347 Vbias 0.50118f
C13192 VDD.n4348 Vbias 0.03639f
C13193 VDD.n4349 Vbias 0.03694f
C13194 VDD.n4350 Vbias 0.04583f
C13195 VDD.n4351 Vbias 0.03902f
C13196 VDD.n4352 Vbias 0.01836f
C13197 VDD.n4353 Vbias 0.03639f
C13198 VDD.n4354 Vbias 0.37318f
C13199 VDD.n4355 Vbias 0.01836f
C13200 VDD.n4356 Vbias 0.03639f
C13201 VDD.n4357 Vbias 0.37318f
C13202 VDD.n4358 Vbias 0.03639f
C13203 VDD.n4359 Vbias 0.03694f
C13204 VDD.n4360 Vbias 0.04583f
C13205 VDD.n4361 Vbias 0.03902f
C13206 VDD.n4362 Vbias 0.01836f
C13207 VDD.n4363 Vbias 0.03639f
C13208 VDD.n4364 Vbias 0.37318f
C13209 VDD.n4365 Vbias 0.01836f
C13210 VDD.n4366 Vbias 0.03639f
C13211 VDD.n4367 Vbias 0.37318f
C13212 VDD.n4368 Vbias 0.03639f
C13213 VDD.n4369 Vbias 0.03694f
C13214 VDD.n4370 Vbias 0.04583f
C13215 VDD.n4371 Vbias 0.03902f
C13216 VDD.n4372 Vbias 0.01836f
C13217 VDD.n4373 Vbias 0.03639f
C13218 VDD.n4374 Vbias 0.50118f
C13219 VDD.n4375 Vbias 0.50118f
C13220 VDD.n4376 Vbias 0.03639f
C13221 VDD.n4377 Vbias 0.01999f
C13222 VDD.n4378 Vbias 0.06648f
C13223 VDD.n4379 Vbias 0.01309f
C13224 VDD.n4380 Vbias 0.11022f
C13225 VDD.n4381 Vbias 0.01699f
C13226 VDD.n4382 Vbias 0.03902f
C13227 VDD.n4383 Vbias 0.03694f
C13228 VDD.n4384 Vbias 0.0216f
C13229 VDD.n4385 Vbias 0.01836f
C13230 VDD.n4386 Vbias 0.01836f
C13231 VDD.n4387 Vbias 0.03639f
C13232 VDD.n4388 Vbias 0.50118f
C13233 VDD.n4389 Vbias 0.03639f
C13234 VDD.n4390 Vbias 0.03694f
C13235 VDD.n4391 Vbias 0.04583f
C13236 VDD.n4392 Vbias 0.03902f
C13237 VDD.n4393 Vbias 0.01836f
C13238 VDD.n4394 Vbias 0.03639f
C13239 VDD.n4395 Vbias 0.37318f
C13240 VDD.n4396 Vbias 0.01836f
C13241 VDD.n4397 Vbias 0.03639f
C13242 VDD.n4398 Vbias 0.37318f
C13243 VDD.n4399 Vbias 0.03639f
C13244 VDD.n4400 Vbias 0.03694f
C13245 VDD.n4401 Vbias 0.04583f
C13246 VDD.n4402 Vbias 0.03902f
C13247 VDD.n4403 Vbias 0.01836f
C13248 VDD.n4404 Vbias 0.03639f
C13249 VDD.n4405 Vbias 0.37318f
C13250 VDD.n4406 Vbias 0.01836f
C13251 VDD.n4407 Vbias 0.03639f
C13252 VDD.n4408 Vbias 0.37318f
C13253 VDD.n4409 Vbias 0.03639f
C13254 VDD.n4410 Vbias 0.03694f
C13255 VDD.n4411 Vbias 0.04583f
C13256 VDD.n4412 Vbias 0.03902f
C13257 VDD.n4413 Vbias 0.01836f
C13258 VDD.n4414 Vbias 0.03639f
C13259 VDD.n4415 Vbias 0.50118f
C13260 VDD.n4416 Vbias 0.01836f
C13261 VDD.n4417 Vbias 0.03639f
C13262 VDD.n4418 Vbias 0.50118f
C13263 VDD.n4419 Vbias 0.03639f
C13264 VDD.n4420 Vbias 0.03694f
C13265 VDD.n4421 Vbias 0.04583f
C13266 VDD.n4422 Vbias 0.03902f
C13267 VDD.n4423 Vbias 0.01836f
C13268 VDD.n4424 Vbias 0.03639f
C13269 VDD.n4425 Vbias 0.37318f
C13270 VDD.n4426 Vbias 0.01836f
C13271 VDD.n4427 Vbias 0.03639f
C13272 VDD.n4428 Vbias 0.37318f
C13273 VDD.n4429 Vbias 0.03639f
C13274 VDD.n4430 Vbias 0.03694f
C13275 VDD.n4431 Vbias 0.04583f
C13276 VDD.n4432 Vbias 0.03902f
C13277 VDD.n4433 Vbias 0.01836f
C13278 VDD.n4434 Vbias 0.03639f
C13279 VDD.n4435 Vbias 0.50118f
C13280 VDD.n4436 Vbias 0.50118f
C13281 VDD.n4437 Vbias 0.03639f
C13282 VDD.n4438 Vbias 0.01999f
C13283 VDD.n4439 Vbias 0.0216f
C13284 VDD.n4440 Vbias 0.01999f
C13285 VDD.n4441 Vbias 0.03639f
C13286 VDD.n4442 Vbias 0.50118f
C13287 VDD.n4443 Vbias 0.50118f
C13288 VDD.n4444 Vbias 0.03639f
C13289 VDD.n4445 Vbias 0.03639f
C13290 VDD.n4446 Vbias 0.01836f
C13291 VDD.n4447 Vbias 0.01836f
C13292 VDD.n4448 Vbias 0.0216f
C13293 VDD.n4449 Vbias 0.03694f
C13294 VDD.t954 Vbias 0.46278f
C13295 VDD.n4450 Vbias 0.03694f
C13296 VDD.n4451 Vbias 0.04583f
C13297 VDD.n4452 Vbias 0.01699f
C13298 VDD.n4453 Vbias 0.03023f
C13299 VDD.n4454 Vbias 0.02225f
C13300 VDD.n4455 Vbias 0.04583f
C13301 VDD.n4456 Vbias 0.03902f
C13302 VDD.n4457 Vbias 0.01836f
C13303 VDD.n4458 Vbias 0.03639f
C13304 VDD.n4459 Vbias 0.37318f
C13305 VDD.n4460 Vbias 0.01836f
C13306 VDD.n4461 Vbias 0.03639f
C13307 VDD.n4462 Vbias 0.37318f
C13308 VDD.n4463 Vbias 0.03639f
C13309 VDD.n4464 Vbias 0.03694f
C13310 VDD.n4465 Vbias 0.04583f
C13311 VDD.n4466 Vbias 0.03902f
C13312 VDD.n4467 Vbias 0.01836f
C13313 VDD.n4468 Vbias 0.03639f
C13314 VDD.n4469 Vbias 0.50118f
C13315 VDD.n4470 Vbias 0.01836f
C13316 VDD.n4471 Vbias 0.03639f
C13317 VDD.n4472 Vbias 0.50118f
C13318 VDD.n4473 Vbias 0.03639f
C13319 VDD.n4474 Vbias 0.03694f
C13320 VDD.n4475 Vbias 0.04583f
C13321 VDD.n4476 Vbias 0.03902f
C13322 VDD.n4477 Vbias 0.01836f
C13323 VDD.n4478 Vbias 0.03639f
C13324 VDD.n4479 Vbias 0.37318f
C13325 VDD.n4480 Vbias 0.01836f
C13326 VDD.n4481 Vbias 0.03639f
C13327 VDD.n4482 Vbias 0.37318f
C13328 VDD.n4483 Vbias 0.03639f
C13329 VDD.n4484 Vbias 0.03694f
C13330 VDD.n4485 Vbias 0.04583f
C13331 VDD.n4486 Vbias 0.03902f
C13332 VDD.n4487 Vbias 0.01836f
C13333 VDD.n4488 Vbias 0.03639f
C13334 VDD.n4489 Vbias 0.37318f
C13335 VDD.n4490 Vbias 0.01836f
C13336 VDD.n4491 Vbias 0.03639f
C13337 VDD.n4492 Vbias 0.37318f
C13338 VDD.n4493 Vbias 0.03639f
C13339 VDD.n4494 Vbias 0.03694f
C13340 VDD.n4495 Vbias 0.04583f
C13341 VDD.n4496 Vbias 0.03902f
C13342 VDD.n4497 Vbias 0.01836f
C13343 VDD.n4498 Vbias 0.03639f
C13344 VDD.n4499 Vbias 0.50118f
C13345 VDD.n4500 Vbias 0.50118f
C13346 VDD.n4501 Vbias 0.03639f
C13347 VDD.n4502 Vbias 0.01999f
C13348 VDD.n4503 Vbias 0.06648f
C13349 VDD.n4504 Vbias 0.01309f
C13350 VDD.n4505 Vbias 0.11022f
C13351 VDD.n4506 Vbias 0.01699f
C13352 VDD.n4507 Vbias 0.03902f
C13353 VDD.n4508 Vbias 0.03694f
C13354 VDD.n4509 Vbias 0.0216f
C13355 VDD.n4510 Vbias 0.01836f
C13356 VDD.n4511 Vbias 0.01836f
C13357 VDD.n4512 Vbias 0.03639f
C13358 VDD.n4513 Vbias 0.50118f
C13359 VDD.n4514 Vbias 0.03639f
C13360 VDD.n4515 Vbias 0.03694f
C13361 VDD.n4516 Vbias 0.04583f
C13362 VDD.n4517 Vbias 0.03902f
C13363 VDD.n4518 Vbias 0.01836f
C13364 VDD.n4519 Vbias 0.03639f
C13365 VDD.n4520 Vbias 0.37318f
C13366 VDD.n4521 Vbias 0.01836f
C13367 VDD.n4522 Vbias 0.03639f
C13368 VDD.n4523 Vbias 0.37318f
C13369 VDD.n4524 Vbias 0.03639f
C13370 VDD.n4525 Vbias 0.03694f
C13371 VDD.n4526 Vbias 0.04583f
C13372 VDD.n4527 Vbias 0.03902f
C13373 VDD.n4528 Vbias 0.01836f
C13374 VDD.n4529 Vbias 0.03639f
C13375 VDD.n4530 Vbias 0.37318f
C13376 VDD.n4531 Vbias 0.01836f
C13377 VDD.n4532 Vbias 0.03639f
C13378 VDD.n4533 Vbias 0.37318f
C13379 VDD.n4534 Vbias 0.03639f
C13380 VDD.n4535 Vbias 0.03694f
C13381 VDD.n4536 Vbias 0.04583f
C13382 VDD.n4537 Vbias 0.03902f
C13383 VDD.n4538 Vbias 0.01836f
C13384 VDD.n4539 Vbias 0.03639f
C13385 VDD.n4540 Vbias 0.50118f
C13386 VDD.n4541 Vbias 0.01836f
C13387 VDD.n4542 Vbias 0.03639f
C13388 VDD.n4543 Vbias 0.50118f
C13389 VDD.n4544 Vbias 0.03639f
C13390 VDD.n4545 Vbias 0.03694f
C13391 VDD.n4546 Vbias 0.04583f
C13392 VDD.n4547 Vbias 0.03902f
C13393 VDD.n4548 Vbias 0.01836f
C13394 VDD.n4549 Vbias 0.03639f
C13395 VDD.n4550 Vbias 0.37318f
C13396 VDD.n4551 Vbias 0.01836f
C13397 VDD.n4552 Vbias 0.03639f
C13398 VDD.n4553 Vbias 0.37318f
C13399 VDD.n4554 Vbias 0.03639f
C13400 VDD.n4555 Vbias 0.03694f
C13401 VDD.n4556 Vbias 0.04583f
C13402 VDD.n4557 Vbias 0.03902f
C13403 VDD.n4558 Vbias 0.01836f
C13404 VDD.n4559 Vbias 0.03639f
C13405 VDD.n4560 Vbias 0.50118f
C13406 VDD.n4561 Vbias 0.50118f
C13407 VDD.n4562 Vbias 0.03639f
C13408 VDD.n4563 Vbias 0.01999f
C13409 VDD.n4564 Vbias 0.0216f
C13410 VDD.n4565 Vbias 0.01999f
C13411 VDD.n4566 Vbias 0.03639f
C13412 VDD.n4567 Vbias 0.50118f
C13413 VDD.n4568 Vbias 0.50118f
C13414 VDD.n4569 Vbias 0.03639f
C13415 VDD.n4570 Vbias 0.03639f
C13416 VDD.n4571 Vbias 0.01836f
C13417 VDD.n4572 Vbias 0.01836f
C13418 VDD.n4573 Vbias 0.0216f
C13419 VDD.n4574 Vbias 0.03694f
C13420 VDD.t221 Vbias 0.46278f
C13421 VDD.n4575 Vbias 0.03694f
C13422 VDD.n4576 Vbias 0.04583f
C13423 VDD.n4577 Vbias 0.01699f
C13424 VDD.n4578 Vbias 0.03023f
C13425 VDD.n4579 Vbias 0.02225f
C13426 VDD.n4580 Vbias 0.04583f
C13427 VDD.n4581 Vbias 0.03902f
C13428 VDD.n4582 Vbias 0.01836f
C13429 VDD.n4583 Vbias 0.03639f
C13430 VDD.n4584 Vbias 0.37318f
C13431 VDD.n4585 Vbias 0.01836f
C13432 VDD.n4586 Vbias 0.03639f
C13433 VDD.n4587 Vbias 0.37318f
C13434 VDD.n4588 Vbias 0.03639f
C13435 VDD.n4589 Vbias 0.03694f
C13436 VDD.n4590 Vbias 0.04583f
C13437 VDD.n4591 Vbias 0.03902f
C13438 VDD.n4592 Vbias 0.01836f
C13439 VDD.n4593 Vbias 0.03639f
C13440 VDD.n4594 Vbias 0.50118f
C13441 VDD.n4595 Vbias 0.01836f
C13442 VDD.n4596 Vbias 0.03639f
C13443 VDD.n4597 Vbias 0.50118f
C13444 VDD.n4598 Vbias 0.03639f
C13445 VDD.n4599 Vbias 0.03694f
C13446 VDD.n4600 Vbias 0.04583f
C13447 VDD.n4601 Vbias 0.03902f
C13448 VDD.n4602 Vbias 0.01836f
C13449 VDD.n4603 Vbias 0.03639f
C13450 VDD.n4604 Vbias 0.37318f
C13451 VDD.n4605 Vbias 0.01836f
C13452 VDD.n4606 Vbias 0.03639f
C13453 VDD.n4607 Vbias 0.37318f
C13454 VDD.n4608 Vbias 0.03639f
C13455 VDD.n4609 Vbias 0.03694f
C13456 VDD.n4610 Vbias 0.04583f
C13457 VDD.n4611 Vbias 0.03902f
C13458 VDD.n4612 Vbias 0.01836f
C13459 VDD.n4613 Vbias 0.03639f
C13460 VDD.n4614 Vbias 0.37318f
C13461 VDD.n4615 Vbias 0.01836f
C13462 VDD.n4616 Vbias 0.03639f
C13463 VDD.n4617 Vbias 0.37318f
C13464 VDD.n4618 Vbias 0.03639f
C13465 VDD.n4619 Vbias 0.03694f
C13466 VDD.n4620 Vbias 0.04583f
C13467 VDD.n4621 Vbias 0.03902f
C13468 VDD.n4622 Vbias 0.01836f
C13469 VDD.n4623 Vbias 0.03639f
C13470 VDD.n4624 Vbias 0.50118f
C13471 VDD.n4625 Vbias 0.50118f
C13472 VDD.n4626 Vbias 0.03639f
C13473 VDD.n4627 Vbias 0.01999f
C13474 VDD.n4628 Vbias 0.06648f
C13475 VDD.n4629 Vbias 0.01309f
C13476 VDD.n4630 Vbias 0.11022f
C13477 VDD.n4631 Vbias 0.01699f
C13478 VDD.n4632 Vbias 0.03902f
C13479 VDD.n4633 Vbias 0.03694f
C13480 VDD.n4634 Vbias 0.0216f
C13481 VDD.n4635 Vbias 0.01836f
C13482 VDD.n4636 Vbias 0.01836f
C13483 VDD.n4637 Vbias 0.03639f
C13484 VDD.n4638 Vbias 0.50118f
C13485 VDD.n4639 Vbias 0.03639f
C13486 VDD.n4640 Vbias 0.03694f
C13487 VDD.n4641 Vbias 0.04583f
C13488 VDD.n4642 Vbias 0.03902f
C13489 VDD.n4643 Vbias 0.01836f
C13490 VDD.n4644 Vbias 0.03639f
C13491 VDD.n4645 Vbias 0.37318f
C13492 VDD.n4646 Vbias 0.01836f
C13493 VDD.n4647 Vbias 0.03639f
C13494 VDD.n4648 Vbias 0.37318f
C13495 VDD.n4649 Vbias 0.03639f
C13496 VDD.n4650 Vbias 0.03694f
C13497 VDD.n4651 Vbias 0.04583f
C13498 VDD.n4652 Vbias 0.03902f
C13499 VDD.n4653 Vbias 0.01836f
C13500 VDD.n4654 Vbias 0.03639f
C13501 VDD.n4655 Vbias 0.37318f
C13502 VDD.n4656 Vbias 0.01836f
C13503 VDD.n4657 Vbias 0.03639f
C13504 VDD.n4658 Vbias 0.37318f
C13505 VDD.n4659 Vbias 0.03639f
C13506 VDD.n4660 Vbias 0.03694f
C13507 VDD.n4661 Vbias 0.04583f
C13508 VDD.n4662 Vbias 0.03902f
C13509 VDD.n4663 Vbias 0.01836f
C13510 VDD.n4664 Vbias 0.03639f
C13511 VDD.n4665 Vbias 0.50118f
C13512 VDD.n4666 Vbias 0.01836f
C13513 VDD.n4667 Vbias 0.03639f
C13514 VDD.n4668 Vbias 0.50118f
C13515 VDD.n4669 Vbias 0.03639f
C13516 VDD.n4670 Vbias 0.03694f
C13517 VDD.n4671 Vbias 0.04583f
C13518 VDD.n4672 Vbias 0.03902f
C13519 VDD.n4673 Vbias 0.01836f
C13520 VDD.n4674 Vbias 0.03639f
C13521 VDD.n4675 Vbias 0.37318f
C13522 VDD.n4676 Vbias 0.01836f
C13523 VDD.n4677 Vbias 0.03639f
C13524 VDD.n4678 Vbias 0.37318f
C13525 VDD.n4679 Vbias 0.03639f
C13526 VDD.n4680 Vbias 0.03694f
C13527 VDD.n4681 Vbias 0.04583f
C13528 VDD.n4682 Vbias 0.03902f
C13529 VDD.n4683 Vbias 0.01836f
C13530 VDD.n4684 Vbias 0.03639f
C13531 VDD.n4685 Vbias 0.50118f
C13532 VDD.n4686 Vbias 0.50118f
C13533 VDD.n4687 Vbias 0.03639f
C13534 VDD.n4688 Vbias 0.01999f
C13535 VDD.n4689 Vbias 0.0216f
C13536 VDD.n4690 Vbias 0.01999f
C13537 VDD.n4691 Vbias 0.03639f
C13538 VDD.n4692 Vbias 0.50118f
C13539 VDD.n4693 Vbias 0.50118f
C13540 VDD.n4694 Vbias 0.03639f
C13541 VDD.n4695 Vbias 0.03639f
C13542 VDD.n4696 Vbias 0.01836f
C13543 VDD.n4697 Vbias 0.01836f
C13544 VDD.n4698 Vbias 0.0216f
C13545 VDD.n4699 Vbias 0.03694f
C13546 VDD.t17 Vbias 0.46278f
C13547 VDD.n4700 Vbias 0.03694f
C13548 VDD.n4701 Vbias 0.04583f
C13549 VDD.n4702 Vbias 0.01699f
C13550 VDD.n4703 Vbias 0.03023f
C13551 VDD.n4704 Vbias 0.02225f
C13552 VDD.n4705 Vbias 0.04583f
C13553 VDD.n4706 Vbias 0.03902f
C13554 VDD.n4707 Vbias 0.01836f
C13555 VDD.n4708 Vbias 0.03639f
C13556 VDD.n4709 Vbias 0.37318f
C13557 VDD.n4710 Vbias 0.01836f
C13558 VDD.n4711 Vbias 0.03639f
C13559 VDD.n4712 Vbias 0.37318f
C13560 VDD.n4713 Vbias 0.03639f
C13561 VDD.n4714 Vbias 0.03694f
C13562 VDD.n4715 Vbias 0.04583f
C13563 VDD.n4716 Vbias 0.03902f
C13564 VDD.n4717 Vbias 0.01836f
C13565 VDD.n4718 Vbias 0.03639f
C13566 VDD.n4719 Vbias 0.50118f
C13567 VDD.n4720 Vbias 0.01836f
C13568 VDD.n4721 Vbias 0.03639f
C13569 VDD.n4722 Vbias 0.50118f
C13570 VDD.n4723 Vbias 0.03639f
C13571 VDD.n4724 Vbias 0.03694f
C13572 VDD.n4725 Vbias 0.04583f
C13573 VDD.n4726 Vbias 0.03902f
C13574 VDD.n4727 Vbias 0.01836f
C13575 VDD.n4728 Vbias 0.03639f
C13576 VDD.n4729 Vbias 0.37318f
C13577 VDD.n4730 Vbias 0.01836f
C13578 VDD.n4731 Vbias 0.03639f
C13579 VDD.n4732 Vbias 0.37318f
C13580 VDD.n4733 Vbias 0.03639f
C13581 VDD.n4734 Vbias 0.03694f
C13582 VDD.n4735 Vbias 0.04583f
C13583 VDD.n4736 Vbias 0.03902f
C13584 VDD.n4737 Vbias 0.01836f
C13585 VDD.n4738 Vbias 0.03639f
C13586 VDD.n4739 Vbias 0.37318f
C13587 VDD.n4740 Vbias 0.01836f
C13588 VDD.n4741 Vbias 0.03639f
C13589 VDD.n4742 Vbias 0.37318f
C13590 VDD.n4743 Vbias 0.03639f
C13591 VDD.n4744 Vbias 0.03694f
C13592 VDD.n4745 Vbias 0.04583f
C13593 VDD.n4746 Vbias 0.03902f
C13594 VDD.n4747 Vbias 0.01836f
C13595 VDD.n4748 Vbias 0.03639f
C13596 VDD.n4749 Vbias 0.50118f
C13597 VDD.n4750 Vbias 0.50118f
C13598 VDD.n4751 Vbias 0.03639f
C13599 VDD.n4752 Vbias 0.01999f
C13600 VDD.n4753 Vbias 0.06648f
C13601 VDD.n4754 Vbias 0.01309f
C13602 VDD.n4755 Vbias 0.08931f
C13603 VDD.t204 Vbias 0.017f
C13604 VDD.n4756 Vbias 0.01999f
C13605 VDD.n4757 Vbias 0.03694f
C13606 VDD.n4758 Vbias 0.0216f
C13607 VDD.n4759 Vbias 0.03694f
C13608 VDD.t87 Vbias 0.46278f
C13609 VDD.n4760 Vbias 0.03639f
C13610 VDD.n4761 Vbias 0.03694f
C13611 VDD.n4762 Vbias 0.03694f
C13612 VDD.n4763 Vbias 0.0216f
C13613 VDD.n4764 Vbias 0.01836f
C13614 VDD.n4765 Vbias 0.03902f
C13615 VDD.t745 Vbias 0.017f
C13616 VDD.t88 Vbias 0.017f
C13617 VDD.n4766 Vbias 0.09713f
C13618 VDD.n4767 Vbias 0.01914f
C13619 VDD.n4768 Vbias 0.03694f
C13620 VDD.n4769 Vbias 0.0216f
C13621 VDD.n4770 Vbias 0.01836f
C13622 VDD.t205 Vbias 0.46278f
C13623 VDD.n4771 Vbias 0.03639f
C13624 VDD.n4772 Vbias 0.03694f
C13625 VDD.n4773 Vbias 0.03694f
C13626 VDD.n4774 Vbias 0.0216f
C13627 VDD.n4775 Vbias 0.01836f
C13628 VDD.n4776 Vbias 0.03902f
C13629 VDD.n4777 Vbias 0.02305f
C13630 VDD.n4778 Vbias 0.03694f
C13631 VDD.n4779 Vbias 0.0216f
C13632 VDD.n4780 Vbias 0.01836f
C13633 VDD.t1004 Vbias 0.46278f
C13634 VDD.n4781 Vbias 0.03639f
C13635 VDD.n4782 Vbias 0.03694f
C13636 VDD.n4783 Vbias 0.03694f
C13637 VDD.n4784 Vbias 0.0216f
C13638 VDD.n4785 Vbias 0.01836f
C13639 VDD.n4786 Vbias 0.03902f
C13640 VDD.t1081 Vbias 0.0169f
C13641 VDD.t206 Vbias 0.0169f
C13642 VDD.n4787 Vbias 0.07902f
C13643 VDD.t1005 Vbias 0.0169f
C13644 VDD.t408 Vbias 0.0169f
C13645 VDD.n4788 Vbias 0.07902f
C13646 VDD.n4789 Vbias 0.03023f
C13647 VDD.n4790 Vbias 0.01699f
C13648 VDD.n4791 Vbias 0.03694f
C13649 VDD.n4792 Vbias 0.0216f
C13650 VDD.n4793 Vbias 0.01836f
C13651 VDD.t77 Vbias 0.46278f
C13652 VDD.n4794 Vbias 0.03639f
C13653 VDD.n4795 Vbias 0.03694f
C13654 VDD.n4796 Vbias 0.03694f
C13655 VDD.n4797 Vbias 0.0216f
C13656 VDD.n4798 Vbias 0.01836f
C13657 VDD.n4799 Vbias 0.03902f
C13658 VDD.t78 Vbias 0.017f
C13659 VDD.t813 Vbias 0.017f
C13660 VDD.n4800 Vbias 0.09713f
C13661 VDD.n4801 Vbias 0.01914f
C13662 VDD.n4802 Vbias 0.03694f
C13663 VDD.n4803 Vbias 0.0216f
C13664 VDD.n4804 Vbias 0.01836f
C13665 VDD.t445 Vbias 0.46278f
C13666 VDD.n4805 Vbias 0.03639f
C13667 VDD.n4806 Vbias 0.03694f
C13668 VDD.n4807 Vbias 0.03694f
C13669 VDD.n4808 Vbias 0.0216f
C13670 VDD.n4809 Vbias 0.01836f
C13671 VDD.n4810 Vbias 0.03902f
C13672 VDD.n4811 Vbias 0.02305f
C13673 VDD.n4812 Vbias 0.03694f
C13674 VDD.n4813 Vbias 0.0216f
C13675 VDD.n4814 Vbias 0.01836f
C13676 VDD.t244 Vbias 0.46278f
C13677 VDD.n4815 Vbias 0.03639f
C13678 VDD.n4816 Vbias 0.03694f
C13679 VDD.n4817 Vbias 0.03694f
C13680 VDD.n4818 Vbias 0.0216f
C13681 VDD.n4819 Vbias 0.01836f
C13682 VDD.n4820 Vbias 0.03902f
C13683 VDD.t422 Vbias 0.0169f
C13684 VDD.t446 Vbias 0.0169f
C13685 VDD.n4821 Vbias 0.07902f
C13686 VDD.t245 Vbias 0.0169f
C13687 VDD.t820 Vbias 0.0169f
C13688 VDD.n4822 Vbias 0.07902f
C13689 VDD.n4823 Vbias 0.03023f
C13690 VDD.n4824 Vbias 0.01699f
C13691 VDD.n4825 Vbias 0.03694f
C13692 VDD.n4826 Vbias 0.0216f
C13693 VDD.n4827 Vbias 0.01836f
C13694 VDD.t1052 Vbias 0.46278f
C13695 VDD.n4828 Vbias 0.03694f
C13696 VDD.n4829 Vbias 0.03694f
C13697 VDD.n4830 Vbias 0.06648f
C13698 VDD.t242 Vbias 0.46278f
C13699 VDD.n4831 Vbias 0.03639f
C13700 VDD.n4832 Vbias 0.03694f
C13701 VDD.n4833 Vbias 0.03694f
C13702 VDD.n4834 Vbias 0.0216f
C13703 VDD.n4835 Vbias 0.01836f
C13704 VDD.n4836 Vbias 0.03902f
C13705 VDD.t1053 Vbias 0.017f
C13706 VDD.n4837 Vbias 0.05322f
C13707 VDD.n4838 Vbias 0.01309f
C13708 VDD.n4839 Vbias 0.01699f
C13709 VDD.n4840 Vbias 0.03694f
C13710 VDD.n4841 Vbias 0.0216f
C13711 VDD.n4842 Vbias 0.01836f
C13712 VDD.t655 Vbias 0.46278f
C13713 VDD.n4843 Vbias 0.03639f
C13714 VDD.n4844 Vbias 0.03694f
C13715 VDD.n4845 Vbias 0.03694f
C13716 VDD.n4846 Vbias 0.0216f
C13717 VDD.n4847 Vbias 0.01836f
C13718 VDD.n4848 Vbias 0.03902f
C13719 VDD.t656 Vbias 0.0169f
C13720 VDD.t243 Vbias 0.0169f
C13721 VDD.n4849 Vbias 0.07902f
C13722 VDD.t657 Vbias 0.0169f
C13723 VDD.t421 Vbias 0.0169f
C13724 VDD.n4850 Vbias 0.07902f
C13725 VDD.n4851 Vbias 0.03023f
C13726 VDD.n4852 Vbias 0.01699f
C13727 VDD.n4853 Vbias 0.03694f
C13728 VDD.n4854 Vbias 0.0216f
C13729 VDD.n4855 Vbias 0.01836f
C13730 VDD.t101 Vbias 0.46278f
C13731 VDD.n4856 Vbias 0.03639f
C13732 VDD.n4857 Vbias 0.03694f
C13733 VDD.n4858 Vbias 0.03694f
C13734 VDD.n4859 Vbias 0.0216f
C13735 VDD.n4860 Vbias 0.01836f
C13736 VDD.n4861 Vbias 0.03902f
C13737 VDD.t102 Vbias 0.017f
C13738 VDD.t729 Vbias 0.017f
C13739 VDD.n4862 Vbias 0.09713f
C13740 VDD.n4863 Vbias 0.01914f
C13741 VDD.n4864 Vbias 0.03694f
C13742 VDD.n4865 Vbias 0.0216f
C13743 VDD.n4866 Vbias 0.01836f
C13744 VDD.t248 Vbias 0.46278f
C13745 VDD.n4867 Vbias 0.03639f
C13746 VDD.n4868 Vbias 0.03694f
C13747 VDD.n4869 Vbias 0.03694f
C13748 VDD.n4870 Vbias 0.0216f
C13749 VDD.n4871 Vbias 0.01836f
C13750 VDD.n4872 Vbias 0.03902f
C13751 VDD.n4873 Vbias 0.02305f
C13752 VDD.n4874 Vbias 0.03694f
C13753 VDD.n4875 Vbias 0.0216f
C13754 VDD.n4876 Vbias 0.01836f
C13755 VDD.t492 Vbias 0.46278f
C13756 VDD.n4877 Vbias 0.03639f
C13757 VDD.n4878 Vbias 0.03694f
C13758 VDD.n4879 Vbias 0.03694f
C13759 VDD.n4880 Vbias 0.0216f
C13760 VDD.n4881 Vbias 0.01836f
C13761 VDD.n4882 Vbias 0.03902f
C13762 VDD.n4883 Vbias 0.03694f
C13763 VDD.n4884 Vbias 0.0216f
C13764 VDD.n4885 Vbias 0.01836f
C13765 VDD.n4886 Vbias 0.01836f
C13766 VDD.n4887 Vbias 0.03639f
C13767 VDD.n4888 Vbias 0.50118f
C13768 VDD.n4889 Vbias 0.03639f
C13769 VDD.n4890 Vbias 0.03694f
C13770 VDD.t493 Vbias 0.0169f
C13771 VDD.t249 Vbias 0.0169f
C13772 VDD.n4891 Vbias 0.07902f
C13773 VDD.t912 Vbias 0.0169f
C13774 VDD.t349 Vbias 0.0169f
C13775 VDD.n4892 Vbias 0.07902f
C13776 VDD.n4893 Vbias 0.04958f
C13777 VDD.n4894 Vbias 0.05277f
C13778 VDD.n4895 Vbias 0.03902f
C13779 VDD.n4896 Vbias 0.01836f
C13780 VDD.n4897 Vbias 0.03639f
C13781 VDD.n4898 Vbias 0.37318f
C13782 VDD.n4899 Vbias 0.01836f
C13783 VDD.n4900 Vbias 0.03639f
C13784 VDD.n4901 Vbias 0.37318f
C13785 VDD.n4902 Vbias 0.03639f
C13786 VDD.n4903 Vbias 0.03694f
C13787 VDD.n4904 Vbias 0.04583f
C13788 VDD.n4905 Vbias 0.03902f
C13789 VDD.n4906 Vbias 0.01836f
C13790 VDD.n4907 Vbias 0.03639f
C13791 VDD.n4908 Vbias 0.37318f
C13792 VDD.n4909 Vbias 0.01836f
C13793 VDD.n4910 Vbias 0.03639f
C13794 VDD.n4911 Vbias 0.37318f
C13795 VDD.n4912 Vbias 0.03639f
C13796 VDD.n4913 Vbias 0.03694f
C13797 VDD.n4914 Vbias 0.04583f
C13798 VDD.n4915 Vbias 0.03902f
C13799 VDD.n4916 Vbias 0.01836f
C13800 VDD.n4917 Vbias 0.03639f
C13801 VDD.n4918 Vbias 0.50118f
C13802 VDD.n4919 Vbias 0.01836f
C13803 VDD.n4920 Vbias 0.03639f
C13804 VDD.n4921 Vbias 0.50118f
C13805 VDD.n4922 Vbias 0.03639f
C13806 VDD.n4923 Vbias 0.03694f
C13807 VDD.n4924 Vbias 0.04583f
C13808 VDD.n4925 Vbias 0.03902f
C13809 VDD.n4926 Vbias 0.01836f
C13810 VDD.n4927 Vbias 0.03639f
C13811 VDD.n4928 Vbias 0.37318f
C13812 VDD.n4929 Vbias 0.01836f
C13813 VDD.n4930 Vbias 0.03639f
C13814 VDD.n4931 Vbias 0.37318f
C13815 VDD.n4932 Vbias 0.03639f
C13816 VDD.n4933 Vbias 0.03694f
C13817 VDD.n4934 Vbias 0.04583f
C13818 VDD.n4935 Vbias 0.03902f
C13819 VDD.n4936 Vbias 0.01836f
C13820 VDD.n4937 Vbias 0.03639f
C13821 VDD.n4938 Vbias 0.50118f
C13822 VDD.n4939 Vbias 0.50118f
C13823 VDD.n4940 Vbias 0.03639f
C13824 VDD.n4941 Vbias 0.01999f
C13825 VDD.n4942 Vbias 0.0216f
C13826 VDD.n4943 Vbias 0.01999f
C13827 VDD.n4944 Vbias 0.03639f
C13828 VDD.n4945 Vbias 0.50118f
C13829 VDD.n4946 Vbias 0.01836f
C13830 VDD.n4947 Vbias 0.03639f
C13831 VDD.n4948 Vbias 0.50118f
C13832 VDD.n4949 Vbias 0.03639f
C13833 VDD.n4950 Vbias 0.03694f
C13834 VDD.n4951 Vbias 0.04583f
C13835 VDD.n4952 Vbias 0.03902f
C13836 VDD.n4953 Vbias 0.01836f
C13837 VDD.n4954 Vbias 0.03639f
C13838 VDD.n4955 Vbias 0.37318f
C13839 VDD.n4956 Vbias 0.01836f
C13840 VDD.n4957 Vbias 0.03639f
C13841 VDD.n4958 Vbias 0.37318f
C13842 VDD.n4959 Vbias 0.03639f
C13843 VDD.n4960 Vbias 0.03694f
C13844 VDD.n4961 Vbias 0.04583f
C13845 VDD.n4962 Vbias 0.03902f
C13846 VDD.n4963 Vbias 0.01836f
C13847 VDD.n4964 Vbias 0.03639f
C13848 VDD.n4965 Vbias 0.37318f
C13849 VDD.n4966 Vbias 0.01836f
C13850 VDD.n4967 Vbias 0.03639f
C13851 VDD.n4968 Vbias 0.37318f
C13852 VDD.n4969 Vbias 0.03639f
C13853 VDD.n4970 Vbias 0.03694f
C13854 VDD.n4971 Vbias 0.04583f
C13855 VDD.n4972 Vbias 0.03902f
C13856 VDD.n4973 Vbias 0.01836f
C13857 VDD.n4974 Vbias 0.03639f
C13858 VDD.n4975 Vbias 0.50118f
C13859 VDD.n4976 Vbias 0.01836f
C13860 VDD.n4977 Vbias 0.03639f
C13861 VDD.n4978 Vbias 0.50118f
C13862 VDD.n4979 Vbias 0.03639f
C13863 VDD.n4980 Vbias 0.03694f
C13864 VDD.n4981 Vbias 0.04583f
C13865 VDD.n4982 Vbias 0.03902f
C13866 VDD.n4983 Vbias 0.01836f
C13867 VDD.n4984 Vbias 0.03639f
C13868 VDD.n4985 Vbias 0.37318f
C13869 VDD.n4986 Vbias 0.01836f
C13870 VDD.n4987 Vbias 0.03639f
C13871 VDD.n4988 Vbias 0.37318f
C13872 VDD.n4989 Vbias 0.03639f
C13873 VDD.n4990 Vbias 0.03694f
C13874 VDD.n4991 Vbias 0.04583f
C13875 VDD.n4992 Vbias 0.03902f
C13876 VDD.n4993 Vbias 0.01836f
C13877 VDD.n4994 Vbias 0.03639f
C13878 VDD.n4995 Vbias 0.37318f
C13879 VDD.n4996 Vbias 0.01836f
C13880 VDD.n4997 Vbias 0.03639f
C13881 VDD.n4998 Vbias 0.37318f
C13882 VDD.n4999 Vbias 0.03639f
C13883 VDD.n5000 Vbias 0.03694f
C13884 VDD.n5001 Vbias 0.04583f
C13885 VDD.n5002 Vbias 0.03902f
C13886 VDD.n5003 Vbias 0.01836f
C13887 VDD.n5004 Vbias 0.03639f
C13888 VDD.n5005 Vbias 0.50118f
C13889 VDD.n5006 Vbias 0.03639f
C13890 VDD.n5007 Vbias 0.50118f
C13891 VDD.t203 Vbias 0.54191f
C13892 VDD.n5009 Vbias 0.45845f
C13893 VDD.n5010 Vbias 0.01999f
C13894 VDD.n5011 Vbias 0.06648f
C13895 VDD.n5012 Vbias 0.01309f
C13896 VDD.n5013 Vbias 0.05322f
C13897 VDD.t960 Vbias 0.0169f
C13898 VDD.t865 Vbias 0.0169f
C13899 VDD.n5014 Vbias 0.07902f
C13900 VDD.t938 Vbias 0.0169f
C13901 VDD.t145 Vbias 0.0169f
C13902 VDD.n5015 Vbias 0.07902f
C13903 VDD.n5016 Vbias 0.03023f
C13904 VDD.n5017 Vbias 0.03902f
C13905 VDD.n5018 Vbias 0.03694f
C13906 VDD.n5019 Vbias 0.03902f
C13907 VDD.n5020 Vbias 0.03639f
C13908 VDD.n5021 Vbias 0.03639f
C13909 VDD.n5022 Vbias 0.50118f
C13910 VDD.n5023 Vbias 0.01836f
C13911 VDD.n5024 Vbias 0.01836f
C13912 VDD.n5025 Vbias 0.0216f
C13913 VDD.n5026 Vbias 0.03694f
C13914 VDD.n5027 Vbias 0.03639f
C13915 VDD.t144 Vbias 0.46278f
C13916 VDD.n5028 Vbias 0.03694f
C13917 VDD.n5029 Vbias 0.03694f
C13918 VDD.n5030 Vbias 0.0216f
C13919 VDD.n5031 Vbias 0.01836f
C13920 VDD.n5032 Vbias 0.02305f
C13921 VDD.n5033 Vbias 0.03902f
C13922 VDD.n5034 Vbias 0.03694f
C13923 VDD.n5035 Vbias 0.0216f
C13924 VDD.n5036 Vbias 0.01836f
C13925 VDD.n5037 Vbias 0.03639f
C13926 VDD.t23 Vbias 0.46278f
C13927 VDD.n5038 Vbias 0.03694f
C13928 VDD.n5039 Vbias 0.03694f
C13929 VDD.n5040 Vbias 0.0216f
C13930 VDD.n5041 Vbias 0.01836f
C13931 VDD.n5042 Vbias 0.01914f
C13932 VDD.n5043 Vbias 0.03902f
C13933 VDD.n5044 Vbias 0.03694f
C13934 VDD.n5045 Vbias 0.0216f
C13935 VDD.n5046 Vbias 0.01836f
C13936 VDD.n5047 Vbias 0.03639f
C13937 VDD.t507 Vbias 0.46278f
C13938 VDD.n5048 Vbias 0.03694f
C13939 VDD.n5049 Vbias 0.03694f
C13940 VDD.n5050 Vbias 0.0216f
C13941 VDD.n5051 Vbias 0.01836f
C13942 VDD.t24 Vbias 0.017f
C13943 VDD.t757 Vbias 0.017f
C13944 VDD.n5052 Vbias 0.09713f
C13945 VDD.n5053 Vbias 0.01699f
C13946 VDD.n5054 Vbias 0.03902f
C13947 VDD.n5055 Vbias 0.03694f
C13948 VDD.n5056 Vbias 0.0216f
C13949 VDD.n5057 Vbias 0.01836f
C13950 VDD.n5058 Vbias 0.03639f
C13951 VDD.t9 Vbias 0.46278f
C13952 VDD.n5059 Vbias 0.03694f
C13953 VDD.n5060 Vbias 0.03694f
C13954 VDD.n5061 Vbias 0.0216f
C13955 VDD.n5062 Vbias 0.01836f
C13956 VDD.t509 Vbias 0.0169f
C13957 VDD.t668 Vbias 0.0169f
C13958 VDD.n5063 Vbias 0.07902f
C13959 VDD.t508 Vbias 0.0169f
C13960 VDD.t10 Vbias 0.0169f
C13961 VDD.n5064 Vbias 0.07902f
C13962 VDD.n5065 Vbias 0.03023f
C13963 VDD.n5066 Vbias 0.01699f
C13964 VDD.n5067 Vbias 0.03902f
C13965 VDD.n5068 Vbias 0.03694f
C13966 VDD.n5069 Vbias 0.0216f
C13967 VDD.n5070 Vbias 0.01836f
C13968 VDD.t1076 Vbias 0.46278f
C13969 VDD.n5071 Vbias 0.03694f
C13970 VDD.n5072 Vbias 0.03694f
C13971 VDD.n5073 Vbias 0.06648f
C13972 VDD.n5074 Vbias 0.03639f
C13973 VDD.t11 Vbias 0.46278f
C13974 VDD.n5075 Vbias 0.03694f
C13975 VDD.n5076 Vbias 0.03694f
C13976 VDD.n5077 Vbias 0.0216f
C13977 VDD.n5078 Vbias 0.01836f
C13978 VDD.t1077 Vbias 0.017f
C13979 VDD.n5079 Vbias 0.01309f
C13980 VDD.n5080 Vbias 0.05322f
C13981 VDD.n5081 Vbias 0.01699f
C13982 VDD.n5082 Vbias 0.03902f
C13983 VDD.n5083 Vbias 0.03694f
C13984 VDD.n5084 Vbias 0.0216f
C13985 VDD.n5085 Vbias 0.01836f
C13986 VDD.n5086 Vbias 0.03639f
C13987 VDD.t561 Vbias 0.46278f
C13988 VDD.n5087 Vbias 0.03694f
C13989 VDD.n5088 Vbias 0.03694f
C13990 VDD.n5089 Vbias 0.0216f
C13991 VDD.n5090 Vbias 0.01836f
C13992 VDD.t12 Vbias 0.0169f
C13993 VDD.t562 Vbias 0.0169f
C13994 VDD.n5091 Vbias 0.07902f
C13995 VDD.t667 Vbias 0.0169f
C13996 VDD.t824 Vbias 0.0169f
C13997 VDD.n5092 Vbias 0.07902f
C13998 VDD.n5093 Vbias 0.03023f
C13999 VDD.n5094 Vbias 0.02305f
C14000 VDD.n5095 Vbias 0.03902f
C14001 VDD.n5096 Vbias 0.03694f
C14002 VDD.n5097 Vbias 0.0216f
C14003 VDD.n5098 Vbias 0.01836f
C14004 VDD.n5099 Vbias 0.03639f
C14005 VDD.t99 Vbias 0.46278f
C14006 VDD.n5100 Vbias 0.03694f
C14007 VDD.n5101 Vbias 0.03694f
C14008 VDD.n5102 Vbias 0.0216f
C14009 VDD.n5103 Vbias 0.01836f
C14010 VDD.n5104 Vbias 0.01914f
C14011 VDD.n5105 Vbias 0.03902f
C14012 VDD.n5106 Vbias 0.03694f
C14013 VDD.n5107 Vbias 0.0216f
C14014 VDD.n5108 Vbias 0.01836f
C14015 VDD.n5109 Vbias 0.03639f
C14016 VDD.t1030 Vbias 0.46278f
C14017 VDD.n5110 Vbias 0.03694f
C14018 VDD.n5111 Vbias 0.03694f
C14019 VDD.n5112 Vbias 0.0216f
C14020 VDD.n5113 Vbias 0.01836f
C14021 VDD.t100 Vbias 0.017f
C14022 VDD.t727 Vbias 0.017f
C14023 VDD.n5114 Vbias 0.09713f
C14024 VDD.n5115 Vbias 0.01699f
C14025 VDD.n5116 Vbias 0.03902f
C14026 VDD.n5117 Vbias 0.03694f
C14027 VDD.n5118 Vbias 0.0216f
C14028 VDD.n5119 Vbias 0.01836f
C14029 VDD.n5120 Vbias 0.03639f
C14030 VDD.t598 Vbias 0.46278f
C14031 VDD.n5121 Vbias 0.03694f
C14032 VDD.n5122 Vbias 0.03694f
C14033 VDD.n5123 Vbias 0.0216f
C14034 VDD.n5124 Vbias 0.01836f
C14035 VDD.t1097 Vbias 0.0169f
C14036 VDD.t861 Vbias 0.0169f
C14037 VDD.n5125 Vbias 0.07902f
C14038 VDD.t1031 Vbias 0.0169f
C14039 VDD.t599 Vbias 0.0169f
C14040 VDD.n5126 Vbias 0.07902f
C14041 VDD.n5127 Vbias 0.03023f
C14042 VDD.n5128 Vbias 0.02305f
C14043 VDD.n5129 Vbias 0.03902f
C14044 VDD.n5130 Vbias 0.03694f
C14045 VDD.n5131 Vbias 0.0216f
C14046 VDD.n5132 Vbias 0.01836f
C14047 VDD.n5133 Vbias 0.03639f
C14048 VDD.t47 Vbias 0.46278f
C14049 VDD.n5134 Vbias 0.03694f
C14050 VDD.n5135 Vbias 0.03694f
C14051 VDD.n5136 Vbias 0.0216f
C14052 VDD.n5137 Vbias 0.01836f
C14053 VDD.n5138 Vbias 0.01914f
C14054 VDD.n5139 Vbias 0.03902f
C14055 VDD.n5140 Vbias 0.03694f
C14056 VDD.n5141 Vbias 0.0216f
C14057 VDD.n5142 Vbias 0.01836f
C14058 VDD.t566 Vbias 0.54191f
C14059 VDD.n5143 Vbias 0.03694f
C14060 VDD.n5144 Vbias 0.03694f
C14061 VDD.n5145 Vbias 0.0216f
C14062 VDD.n5147 Vbias 0.45845f
C14063 VDD.n5148 Vbias 0.01999f
C14064 VDD.t805 Vbias 0.017f
C14065 VDD.t48 Vbias 0.017f
C14066 VDD.n5149 Vbias 0.09713f
C14067 VDD.t567 Vbias 0.017f
C14068 VDD.t869 Vbias 0.0169f
C14069 VDD.t286 Vbias 0.0169f
C14070 VDD.n5150 Vbias 0.07902f
C14071 VDD.t863 Vbias 0.0169f
C14072 VDD.t459 Vbias 0.0169f
C14073 VDD.n5151 Vbias 0.07902f
C14074 VDD.n5152 Vbias 0.03023f
C14075 VDD.n5153 Vbias 0.03902f
C14076 VDD.n5154 Vbias 0.03694f
C14077 VDD.n5155 Vbias 0.03902f
C14078 VDD.n5156 Vbias 0.03639f
C14079 VDD.n5157 Vbias 0.03639f
C14080 VDD.n5158 Vbias 0.50118f
C14081 VDD.n5159 Vbias 0.01836f
C14082 VDD.n5160 Vbias 0.01836f
C14083 VDD.n5161 Vbias 0.0216f
C14084 VDD.n5162 Vbias 0.03694f
C14085 VDD.n5163 Vbias 0.03639f
C14086 VDD.t285 Vbias 0.46278f
C14087 VDD.n5164 Vbias 0.03694f
C14088 VDD.n5165 Vbias 0.03694f
C14089 VDD.n5166 Vbias 0.0216f
C14090 VDD.n5167 Vbias 0.01836f
C14091 VDD.n5168 Vbias 0.02305f
C14092 VDD.n5169 Vbias 0.03902f
C14093 VDD.n5170 Vbias 0.03694f
C14094 VDD.n5171 Vbias 0.0216f
C14095 VDD.n5172 Vbias 0.01836f
C14096 VDD.n5173 Vbias 0.03639f
C14097 VDD.t73 Vbias 0.46278f
C14098 VDD.n5174 Vbias 0.03694f
C14099 VDD.n5175 Vbias 0.03694f
C14100 VDD.n5176 Vbias 0.0216f
C14101 VDD.n5177 Vbias 0.01836f
C14102 VDD.n5178 Vbias 0.01914f
C14103 VDD.n5179 Vbias 0.03902f
C14104 VDD.n5180 Vbias 0.03694f
C14105 VDD.n5181 Vbias 0.0216f
C14106 VDD.n5182 Vbias 0.01836f
C14107 VDD.n5183 Vbias 0.03639f
C14108 VDD.t341 Vbias 0.46278f
C14109 VDD.n5184 Vbias 0.03694f
C14110 VDD.n5185 Vbias 0.03694f
C14111 VDD.n5186 Vbias 0.0216f
C14112 VDD.n5187 Vbias 0.01836f
C14113 VDD.t74 Vbias 0.017f
C14114 VDD.t809 Vbias 0.017f
C14115 VDD.n5188 Vbias 0.09713f
C14116 VDD.n5189 Vbias 0.01699f
C14117 VDD.n5190 Vbias 0.03902f
C14118 VDD.n5191 Vbias 0.03694f
C14119 VDD.n5192 Vbias 0.0216f
C14120 VDD.n5193 Vbias 0.01836f
C14121 VDD.n5194 Vbias 0.03639f
C14122 VDD.t665 Vbias 0.46278f
C14123 VDD.n5195 Vbias 0.03694f
C14124 VDD.n5196 Vbias 0.03694f
C14125 VDD.n5197 Vbias 0.0216f
C14126 VDD.n5198 Vbias 0.01836f
C14127 VDD.t711 Vbias 0.0169f
C14128 VDD.t832 Vbias 0.0169f
C14129 VDD.n5199 Vbias 0.07902f
C14130 VDD.t342 Vbias 0.0169f
C14131 VDD.t666 Vbias 0.0169f
C14132 VDD.n5200 Vbias 0.07902f
C14133 VDD.n5201 Vbias 0.03023f
C14134 VDD.n5202 Vbias 0.01699f
C14135 VDD.n5203 Vbias 0.03902f
C14136 VDD.n5204 Vbias 0.03694f
C14137 VDD.n5205 Vbias 0.0216f
C14138 VDD.n5206 Vbias 0.01836f
C14139 VDD.t1058 Vbias 0.46278f
C14140 VDD.n5207 Vbias 0.03694f
C14141 VDD.n5208 Vbias 0.03694f
C14142 VDD.n5209 Vbias 0.06648f
C14143 VDD.n5210 Vbias 0.03639f
C14144 VDD.t643 Vbias 0.46278f
C14145 VDD.n5211 Vbias 0.03694f
C14146 VDD.n5212 Vbias 0.03694f
C14147 VDD.n5213 Vbias 0.0216f
C14148 VDD.n5214 Vbias 0.01836f
C14149 VDD.t1059 Vbias 0.017f
C14150 VDD.n5215 Vbias 0.01309f
C14151 VDD.n5216 Vbias 0.05322f
C14152 VDD.n5217 Vbias 0.01699f
C14153 VDD.n5218 Vbias 0.03902f
C14154 VDD.n5219 Vbias 0.03694f
C14155 VDD.n5220 Vbias 0.0216f
C14156 VDD.n5221 Vbias 0.01836f
C14157 VDD.n5222 Vbias 0.03639f
C14158 VDD.t486 Vbias 0.46278f
C14159 VDD.n5223 Vbias 0.03694f
C14160 VDD.n5224 Vbias 0.03694f
C14161 VDD.n5225 Vbias 0.0216f
C14162 VDD.n5226 Vbias 0.01836f
C14163 VDD.t664 Vbias 0.0169f
C14164 VDD.t487 Vbias 0.0169f
C14165 VDD.n5227 Vbias 0.07902f
C14166 VDD.t644 Vbias 0.0169f
C14167 VDD.t522 Vbias 0.0169f
C14168 VDD.n5228 Vbias 0.07902f
C14169 VDD.n5229 Vbias 0.03023f
C14170 VDD.n5230 Vbias 0.02305f
C14171 VDD.n5231 Vbias 0.03902f
C14172 VDD.n5232 Vbias 0.03694f
C14173 VDD.n5233 Vbias 0.0216f
C14174 VDD.n5234 Vbias 0.01836f
C14175 VDD.n5235 Vbias 0.03639f
C14176 VDD.t111 Vbias 0.46278f
C14177 VDD.n5236 Vbias 0.03694f
C14178 VDD.n5237 Vbias 0.03694f
C14179 VDD.n5238 Vbias 0.0216f
C14180 VDD.n5239 Vbias 0.01836f
C14181 VDD.n5240 Vbias 0.01914f
C14182 VDD.n5241 Vbias 0.03902f
C14183 VDD.n5242 Vbias 0.03694f
C14184 VDD.n5243 Vbias 0.0216f
C14185 VDD.n5244 Vbias 0.01836f
C14186 VDD.n5245 Vbias 0.03639f
C14187 VDD.t1032 Vbias 0.46278f
C14188 VDD.n5246 Vbias 0.03694f
C14189 VDD.n5247 Vbias 0.03694f
C14190 VDD.n5248 Vbias 0.0216f
C14191 VDD.n5249 Vbias 0.01836f
C14192 VDD.t112 Vbias 0.017f
C14193 VDD.t733 Vbias 0.017f
C14194 VDD.n5250 Vbias 0.09713f
C14195 VDD.n5251 Vbias 0.01699f
C14196 VDD.n5252 Vbias 0.03902f
C14197 VDD.n5253 Vbias 0.03694f
C14198 VDD.n5254 Vbias 0.0216f
C14199 VDD.n5255 Vbias 0.01836f
C14200 VDD.n5256 Vbias 0.03639f
C14201 VDD.t398 Vbias 0.46278f
C14202 VDD.n5257 Vbias 0.03694f
C14203 VDD.n5258 Vbias 0.03694f
C14204 VDD.n5259 Vbias 0.0216f
C14205 VDD.n5260 Vbias 0.01836f
C14206 VDD.t1033 Vbias 0.0169f
C14207 VDD.t399 Vbias 0.0169f
C14208 VDD.n5261 Vbias 0.07902f
C14209 VDD.t1078 Vbias 0.0169f
C14210 VDD.t1107 Vbias 0.0169f
C14211 VDD.n5262 Vbias 0.07902f
C14212 VDD.n5263 Vbias 0.03023f
C14213 VDD.n5264 Vbias 0.02305f
C14214 VDD.n5265 Vbias 0.03902f
C14215 VDD.n5266 Vbias 0.03694f
C14216 VDD.n5267 Vbias 0.0216f
C14217 VDD.n5268 Vbias 0.01836f
C14218 VDD.n5269 Vbias 0.03639f
C14219 VDD.t55 Vbias 0.46278f
C14220 VDD.n5270 Vbias 0.03694f
C14221 VDD.n5271 Vbias 0.03694f
C14222 VDD.n5272 Vbias 0.0216f
C14223 VDD.n5273 Vbias 0.01836f
C14224 VDD.n5274 Vbias 0.01914f
C14225 VDD.n5275 Vbias 0.03902f
C14226 VDD.n5276 Vbias 0.03694f
C14227 VDD.n5277 Vbias 0.0216f
C14228 VDD.n5278 Vbias 0.01836f
C14229 VDD.t155 Vbias 0.54191f
C14230 VDD.n5279 Vbias 0.03694f
C14231 VDD.n5280 Vbias 0.03694f
C14232 VDD.n5281 Vbias 0.0216f
C14233 VDD.n5283 Vbias 0.45845f
C14234 VDD.n5284 Vbias 0.01999f
C14235 VDD.t811 Vbias 0.017f
C14236 VDD.t56 Vbias 0.017f
C14237 VDD.n5285 Vbias 0.09713f
C14238 VDD.t156 Vbias 0.017f
C14239 VDD.t488 Vbias 0.0169f
C14240 VDD.t610 Vbias 0.0169f
C14241 VDD.n5286 Vbias 0.07902f
C14242 VDD.t152 Vbias 0.0169f
C14243 VDD.t448 Vbias 0.0169f
C14244 VDD.n5287 Vbias 0.07902f
C14245 VDD.n5288 Vbias 0.03023f
C14246 VDD.n5289 Vbias 0.03902f
C14247 VDD.n5290 Vbias 0.03694f
C14248 VDD.n5291 Vbias 0.03902f
C14249 VDD.n5292 Vbias 0.03639f
C14250 VDD.n5293 Vbias 0.03639f
C14251 VDD.n5294 Vbias 0.50118f
C14252 VDD.n5295 Vbias 0.01836f
C14253 VDD.n5296 Vbias 0.01836f
C14254 VDD.n5297 Vbias 0.0216f
C14255 VDD.n5298 Vbias 0.03694f
C14256 VDD.n5299 Vbias 0.03639f
C14257 VDD.t447 Vbias 0.46278f
C14258 VDD.n5300 Vbias 0.03694f
C14259 VDD.n5301 Vbias 0.03694f
C14260 VDD.n5302 Vbias 0.0216f
C14261 VDD.n5303 Vbias 0.01836f
C14262 VDD.n5304 Vbias 0.02305f
C14263 VDD.n5305 Vbias 0.03902f
C14264 VDD.n5306 Vbias 0.03694f
C14265 VDD.n5307 Vbias 0.0216f
C14266 VDD.n5308 Vbias 0.01836f
C14267 VDD.n5309 Vbias 0.03639f
C14268 VDD.t83 Vbias 0.46278f
C14269 VDD.n5310 Vbias 0.03694f
C14270 VDD.n5311 Vbias 0.03694f
C14271 VDD.n5312 Vbias 0.0216f
C14272 VDD.n5313 Vbias 0.01836f
C14273 VDD.n5314 Vbias 0.01914f
C14274 VDD.n5315 Vbias 0.03902f
C14275 VDD.n5316 Vbias 0.03694f
C14276 VDD.n5317 Vbias 0.0216f
C14277 VDD.n5318 Vbias 0.01836f
C14278 VDD.n5319 Vbias 0.03639f
C14279 VDD.t363 Vbias 0.46278f
C14280 VDD.n5320 Vbias 0.03694f
C14281 VDD.n5321 Vbias 0.03694f
C14282 VDD.n5322 Vbias 0.0216f
C14283 VDD.n5323 Vbias 0.01836f
C14284 VDD.t84 Vbias 0.017f
C14285 VDD.t715 Vbias 0.017f
C14286 VDD.n5324 Vbias 0.09713f
C14287 VDD.n5325 Vbias 0.01699f
C14288 VDD.n5326 Vbias 0.03902f
C14289 VDD.n5327 Vbias 0.03694f
C14290 VDD.n5328 Vbias 0.0216f
C14291 VDD.n5329 Vbias 0.01836f
C14292 VDD.n5330 Vbias 0.03639f
C14293 VDD.t15 Vbias 0.46278f
C14294 VDD.n5331 Vbias 0.03694f
C14295 VDD.n5332 Vbias 0.03694f
C14296 VDD.n5333 Vbias 0.0216f
C14297 VDD.n5334 Vbias 0.01836f
C14298 VDD.t833 Vbias 0.0169f
C14299 VDD.t679 Vbias 0.0169f
C14300 VDD.n5335 Vbias 0.07902f
C14301 VDD.t364 Vbias 0.0169f
C14302 VDD.t16 Vbias 0.0169f
C14303 VDD.n5336 Vbias 0.07902f
C14304 VDD.n5337 Vbias 0.03023f
C14305 VDD.n5338 Vbias 0.01699f
C14306 VDD.n5339 Vbias 0.03902f
C14307 VDD.n5340 Vbias 0.03694f
C14308 VDD.n5341 Vbias 0.0216f
C14309 VDD.n5342 Vbias 0.01836f
C14310 VDD.t1084 Vbias 0.46278f
C14311 VDD.n5343 Vbias 0.03694f
C14312 VDD.n5344 Vbias 0.03694f
C14313 VDD.n5345 Vbias 0.06648f
C14314 VDD.n5346 Vbias 0.03639f
C14315 VDD.t21 Vbias 0.46278f
C14316 VDD.n5347 Vbias 0.03694f
C14317 VDD.n5348 Vbias 0.03694f
C14318 VDD.n5349 Vbias 0.0216f
C14319 VDD.n5350 Vbias 0.01836f
C14320 VDD.t1085 Vbias 0.017f
C14321 VDD.n5351 Vbias 0.01309f
C14322 VDD.n5352 Vbias 0.05322f
C14323 VDD.n5353 Vbias 0.01699f
C14324 VDD.n5354 Vbias 0.03902f
C14325 VDD.n5355 Vbias 0.03694f
C14326 VDD.n5356 Vbias 0.0216f
C14327 VDD.n5357 Vbias 0.01836f
C14328 VDD.n5358 Vbias 0.03639f
C14329 VDD.t615 Vbias 0.46278f
C14330 VDD.n5359 Vbias 0.03694f
C14331 VDD.n5360 Vbias 0.03694f
C14332 VDD.n5361 Vbias 0.0216f
C14333 VDD.n5362 Vbias 0.01836f
C14334 VDD.t22 Vbias 0.0169f
C14335 VDD.t616 Vbias 0.0169f
C14336 VDD.n5363 Vbias 0.07902f
C14337 VDD.t678 Vbias 0.0169f
C14338 VDD.t935 Vbias 0.0169f
C14339 VDD.n5364 Vbias 0.07902f
C14340 VDD.n5365 Vbias 0.03023f
C14341 VDD.n5366 Vbias 0.02305f
C14342 VDD.n5367 Vbias 0.03902f
C14343 VDD.n5368 Vbias 0.03694f
C14344 VDD.n5369 Vbias 0.0216f
C14345 VDD.n5370 Vbias 0.01836f
C14346 VDD.n5371 Vbias 0.03639f
C14347 VDD.t65 Vbias 0.46278f
C14348 VDD.n5372 Vbias 0.03694f
C14349 VDD.n5373 Vbias 0.03694f
C14350 VDD.n5374 Vbias 0.0216f
C14351 VDD.n5375 Vbias 0.01836f
C14352 VDD.n5376 Vbias 0.01914f
C14353 VDD.n5377 Vbias 0.03902f
C14354 VDD.n5378 Vbias 0.03694f
C14355 VDD.n5379 Vbias 0.0216f
C14356 VDD.n5380 Vbias 0.01836f
C14357 VDD.n5381 Vbias 0.03639f
C14358 VDD.t1060 Vbias 0.46278f
C14359 VDD.n5382 Vbias 0.03694f
C14360 VDD.n5383 Vbias 0.03694f
C14361 VDD.n5384 Vbias 0.0216f
C14362 VDD.n5385 Vbias 0.01836f
C14363 VDD.t66 Vbias 0.017f
C14364 VDD.t797 Vbias 0.017f
C14365 VDD.n5386 Vbias 0.09713f
C14366 VDD.n5387 Vbias 0.01699f
C14367 VDD.n5388 Vbias 0.03902f
C14368 VDD.n5389 Vbias 0.03694f
C14369 VDD.n5390 Vbias 0.0216f
C14370 VDD.n5391 Vbias 0.01836f
C14371 VDD.n5392 Vbias 0.03639f
C14372 VDD.t172 Vbias 0.46278f
C14373 VDD.n5393 Vbias 0.03694f
C14374 VDD.n5394 Vbias 0.03694f
C14375 VDD.n5395 Vbias 0.0216f
C14376 VDD.n5396 Vbias 0.01836f
C14377 VDD.t1061 Vbias 0.0169f
C14378 VDD.t173 Vbias 0.0169f
C14379 VDD.n5397 Vbias 0.07902f
C14380 VDD.t1096 Vbias 0.0169f
C14381 VDD.t858 Vbias 0.0169f
C14382 VDD.n5398 Vbias 0.07902f
C14383 VDD.n5399 Vbias 0.03023f
C14384 VDD.n5400 Vbias 0.02305f
C14385 VDD.n5401 Vbias 0.03902f
C14386 VDD.n5402 Vbias 0.03694f
C14387 VDD.n5403 Vbias 0.0216f
C14388 VDD.n5404 Vbias 0.01836f
C14389 VDD.n5405 Vbias 0.03639f
C14390 VDD.t69 Vbias 0.46278f
C14391 VDD.n5406 Vbias 0.03694f
C14392 VDD.n5407 Vbias 0.03694f
C14393 VDD.n5408 Vbias 0.0216f
C14394 VDD.n5409 Vbias 0.01836f
C14395 VDD.n5410 Vbias 0.01914f
C14396 VDD.n5411 Vbias 0.03902f
C14397 VDD.n5412 Vbias 0.03694f
C14398 VDD.n5413 Vbias 0.0216f
C14399 VDD.n5414 Vbias 0.01836f
C14400 VDD.t837 Vbias 0.54191f
C14401 VDD.n5415 Vbias 0.03694f
C14402 VDD.n5416 Vbias 0.03694f
C14403 VDD.n5417 Vbias 0.0216f
C14404 VDD.n5419 Vbias 0.45845f
C14405 VDD.n5420 Vbias 0.01999f
C14406 VDD.t725 Vbias 0.017f
C14407 VDD.t70 Vbias 0.017f
C14408 VDD.n5421 Vbias 0.09713f
C14409 VDD.t838 Vbias 0.017f
C14410 VDD.t659 Vbias 0.0169f
C14411 VDD.t541 Vbias 0.0169f
C14412 VDD.n5422 Vbias 0.07902f
C14413 VDD.t995 Vbias 0.0169f
C14414 VDD.t200 Vbias 0.0169f
C14415 VDD.n5423 Vbias 0.07902f
C14416 VDD.n5424 Vbias 0.03023f
C14417 VDD.n5425 Vbias 0.03902f
C14418 VDD.n5426 Vbias 0.03694f
C14419 VDD.n5427 Vbias 0.03902f
C14420 VDD.n5428 Vbias 0.03639f
C14421 VDD.n5429 Vbias 0.03639f
C14422 VDD.n5430 Vbias 0.50118f
C14423 VDD.n5431 Vbias 0.01836f
C14424 VDD.n5432 Vbias 0.01836f
C14425 VDD.n5433 Vbias 0.0216f
C14426 VDD.n5434 Vbias 0.03694f
C14427 VDD.n5435 Vbias 0.03639f
C14428 VDD.t199 Vbias 0.46278f
C14429 VDD.n5436 Vbias 0.03694f
C14430 VDD.n5437 Vbias 0.03694f
C14431 VDD.n5438 Vbias 0.0216f
C14432 VDD.n5439 Vbias 0.01836f
C14433 VDD.n5440 Vbias 0.02305f
C14434 VDD.n5441 Vbias 0.03902f
C14435 VDD.n5442 Vbias 0.03694f
C14436 VDD.n5443 Vbias 0.0216f
C14437 VDD.n5444 Vbias 0.01836f
C14438 VDD.n5445 Vbias 0.03639f
C14439 VDD.t49 Vbias 0.46278f
C14440 VDD.n5446 Vbias 0.03694f
C14441 VDD.n5447 Vbias 0.03694f
C14442 VDD.n5448 Vbias 0.0216f
C14443 VDD.n5449 Vbias 0.01836f
C14444 VDD.n5450 Vbias 0.01914f
C14445 VDD.n5451 Vbias 0.03902f
C14446 VDD.n5452 Vbias 0.03694f
C14447 VDD.n5453 Vbias 0.0216f
C14448 VDD.n5454 Vbias 0.01836f
C14449 VDD.n5455 Vbias 0.03639f
C14450 VDD.t428 Vbias 0.46278f
C14451 VDD.n5456 Vbias 0.03694f
C14452 VDD.n5457 Vbias 0.03694f
C14453 VDD.n5458 Vbias 0.0216f
C14454 VDD.n5459 Vbias 0.01836f
C14455 VDD.t50 Vbias 0.017f
C14456 VDD.t787 Vbias 0.017f
C14457 VDD.n5460 Vbias 0.09713f
C14458 VDD.n5461 Vbias 0.01699f
C14459 VDD.n5462 Vbias 0.03902f
C14460 VDD.n5463 Vbias 0.03694f
C14461 VDD.n5464 Vbias 0.0216f
C14462 VDD.n5465 Vbias 0.01836f
C14463 VDD.n5466 Vbias 0.03639f
C14464 VDD.t170 Vbias 0.46278f
C14465 VDD.n5467 Vbias 0.03694f
C14466 VDD.n5468 Vbias 0.03694f
C14467 VDD.n5469 Vbias 0.0216f
C14468 VDD.n5470 Vbias 0.01836f
C14469 VDD.t429 Vbias 0.0169f
C14470 VDD.t279 Vbias 0.0169f
C14471 VDD.n5471 Vbias 0.07902f
C14472 VDD.t972 Vbias 0.0169f
C14473 VDD.t171 Vbias 0.0169f
C14474 VDD.n5472 Vbias 0.07902f
C14475 VDD.n5473 Vbias 0.03023f
C14476 VDD.n5474 Vbias 0.01699f
C14477 VDD.n5475 Vbias 0.03902f
C14478 VDD.n5476 Vbias 0.03694f
C14479 VDD.n5477 Vbias 0.0216f
C14480 VDD.n5478 Vbias 0.01836f
C14481 VDD.t1089 Vbias 0.46278f
C14482 VDD.n5479 Vbias 0.03694f
C14483 VDD.n5480 Vbias 0.03694f
C14484 VDD.n5481 Vbias 0.06648f
C14485 VDD.n5482 Vbias 0.03639f
C14486 VDD.t280 Vbias 0.46278f
C14487 VDD.n5483 Vbias 0.03694f
C14488 VDD.n5484 Vbias 0.03694f
C14489 VDD.n5485 Vbias 0.0216f
C14490 VDD.n5486 Vbias 0.01836f
C14491 VDD.t1090 Vbias 0.017f
C14492 VDD.n5487 Vbias 0.01309f
C14493 VDD.n5488 Vbias 0.05322f
C14494 VDD.n5489 Vbias 0.01699f
C14495 VDD.n5490 Vbias 0.03902f
C14496 VDD.n5491 Vbias 0.03694f
C14497 VDD.n5492 Vbias 0.0216f
C14498 VDD.n5493 Vbias 0.01836f
C14499 VDD.n5494 Vbias 0.03639f
C14500 VDD.t365 Vbias 0.46278f
C14501 VDD.n5495 Vbias 0.03694f
C14502 VDD.n5496 Vbias 0.03694f
C14503 VDD.n5497 Vbias 0.0216f
C14504 VDD.n5498 Vbias 0.01836f
C14505 VDD.t841 Vbias 0.0169f
C14506 VDD.t965 Vbias 0.0169f
C14507 VDD.n5499 Vbias 0.07902f
C14508 VDD.t281 Vbias 0.0169f
C14509 VDD.t366 Vbias 0.0169f
C14510 VDD.n5500 Vbias 0.07902f
C14511 VDD.n5501 Vbias 0.03023f
C14512 VDD.n5502 Vbias 0.02305f
C14513 VDD.n5503 Vbias 0.03902f
C14514 VDD.n5504 Vbias 0.03694f
C14515 VDD.n5505 Vbias 0.0216f
C14516 VDD.n5506 Vbias 0.01836f
C14517 VDD.n5507 Vbias 0.03639f
C14518 VDD.t81 Vbias 0.46278f
C14519 VDD.n5508 Vbias 0.03694f
C14520 VDD.n5509 Vbias 0.03694f
C14521 VDD.n5510 Vbias 0.0216f
C14522 VDD.n5511 Vbias 0.01836f
C14523 VDD.n5512 Vbias 0.01914f
C14524 VDD.n5513 Vbias 0.03902f
C14525 VDD.n5514 Vbias 0.03694f
C14526 VDD.n5515 Vbias 0.0216f
C14527 VDD.n5516 Vbias 0.01836f
C14528 VDD.n5517 Vbias 0.03639f
C14529 VDD.t1002 Vbias 0.46278f
C14530 VDD.n5518 Vbias 0.03694f
C14531 VDD.n5519 Vbias 0.03694f
C14532 VDD.n5520 Vbias 0.0216f
C14533 VDD.n5521 Vbias 0.01836f
C14534 VDD.t82 Vbias 0.017f
C14535 VDD.t815 Vbias 0.017f
C14536 VDD.n5522 Vbias 0.09713f
C14537 VDD.n5523 Vbias 0.01699f
C14538 VDD.n5524 Vbias 0.03902f
C14539 VDD.n5525 Vbias 0.03694f
C14540 VDD.n5526 Vbias 0.0216f
C14541 VDD.n5527 Vbias 0.01836f
C14542 VDD.n5528 Vbias 0.03639f
C14543 VDD.t254 Vbias 0.46278f
C14544 VDD.n5529 Vbias 0.03694f
C14545 VDD.n5530 Vbias 0.03694f
C14546 VDD.n5531 Vbias 0.0216f
C14547 VDD.n5532 Vbias 0.01836f
C14548 VDD.t1003 Vbias 0.0169f
C14549 VDD.t825 Vbias 0.0169f
C14550 VDD.n5533 Vbias 0.07902f
C14551 VDD.t1047 Vbias 0.0169f
C14552 VDD.t255 Vbias 0.0169f
C14553 VDD.n5534 Vbias 0.07902f
C14554 VDD.n5535 Vbias 0.03023f
C14555 VDD.n5536 Vbias 0.02305f
C14556 VDD.n5537 Vbias 0.03902f
C14557 VDD.n5538 Vbias 0.03694f
C14558 VDD.n5539 Vbias 0.0216f
C14559 VDD.n5540 Vbias 0.01836f
C14560 VDD.n5541 Vbias 0.03639f
C14561 VDD.t33 Vbias 0.46278f
C14562 VDD.n5542 Vbias 0.03694f
C14563 VDD.n5543 Vbias 0.03694f
C14564 VDD.n5544 Vbias 0.0216f
C14565 VDD.n5545 Vbias 0.01836f
C14566 VDD.n5546 Vbias 0.01914f
C14567 VDD.n5547 Vbias 0.03902f
C14568 VDD.n5548 Vbias 0.03694f
C14569 VDD.n5549 Vbias 0.0216f
C14570 VDD.n5550 Vbias 0.01836f
C14571 VDD.t829 Vbias 0.54191f
C14572 VDD.n5551 Vbias 0.03694f
C14573 VDD.n5552 Vbias 0.03694f
C14574 VDD.n5553 Vbias 0.0216f
C14575 VDD.n5555 Vbias 0.45845f
C14576 VDD.n5556 Vbias 0.01999f
C14577 VDD.t789 Vbias 0.017f
C14578 VDD.t34 Vbias 0.017f
C14579 VDD.n5557 Vbias 0.09713f
C14580 VDD.t830 Vbias 0.017f
C14581 VDD.t312 Vbias 0.0169f
C14582 VDD.t185 Vbias 0.0169f
C14583 VDD.n5558 Vbias 0.07902f
C14584 VDD.t831 Vbias 0.0169f
C14585 VDD.t278 Vbias 0.0169f
C14586 VDD.n5559 Vbias 0.07902f
C14587 VDD.n5560 Vbias 0.03023f
C14588 VDD.n5561 Vbias 0.03902f
C14589 VDD.n5562 Vbias 0.03694f
C14590 VDD.n5563 Vbias 0.03902f
C14591 VDD.n5564 Vbias 0.03639f
C14592 VDD.n5565 Vbias 0.03639f
C14593 VDD.n5566 Vbias 0.50118f
C14594 VDD.n5567 Vbias 0.01836f
C14595 VDD.n5568 Vbias 0.01836f
C14596 VDD.n5569 Vbias 0.0216f
C14597 VDD.n5570 Vbias 0.03694f
C14598 VDD.n5571 Vbias 0.03639f
C14599 VDD.t184 Vbias 0.46278f
C14600 VDD.n5572 Vbias 0.03694f
C14601 VDD.n5573 Vbias 0.03694f
C14602 VDD.n5574 Vbias 0.0216f
C14603 VDD.n5575 Vbias 0.01836f
C14604 VDD.n5576 Vbias 0.02305f
C14605 VDD.n5577 Vbias 0.03902f
C14606 VDD.n5578 Vbias 0.03694f
C14607 VDD.n5579 Vbias 0.0216f
C14608 VDD.n5580 Vbias 0.01836f
C14609 VDD.n5581 Vbias 0.03639f
C14610 VDD.t103 Vbias 0.46278f
C14611 VDD.n5582 Vbias 0.03694f
C14612 VDD.n5583 Vbias 0.03694f
C14613 VDD.n5584 Vbias 0.0216f
C14614 VDD.n5585 Vbias 0.01836f
C14615 VDD.n5586 Vbias 0.01914f
C14616 VDD.n5587 Vbias 0.03902f
C14617 VDD.n5588 Vbias 0.03694f
C14618 VDD.n5589 Vbias 0.0216f
C14619 VDD.n5590 Vbias 0.01836f
C14620 VDD.n5591 Vbias 0.03639f
C14621 VDD.t855 Vbias 0.46278f
C14622 VDD.n5592 Vbias 0.03694f
C14623 VDD.n5593 Vbias 0.03694f
C14624 VDD.n5594 Vbias 0.0216f
C14625 VDD.n5595 Vbias 0.01836f
C14626 VDD.t104 Vbias 0.017f
C14627 VDD.t731 Vbias 0.017f
C14628 VDD.n5596 Vbias 0.09713f
C14629 VDD.n5597 Vbias 0.01699f
C14630 VDD.n5598 Vbias 0.03902f
C14631 VDD.n5599 Vbias 0.03694f
C14632 VDD.n5600 Vbias 0.0216f
C14633 VDD.n5601 Vbias 0.01836f
C14634 VDD.n5602 Vbias 0.03639f
C14635 VDD.t301 Vbias 0.46278f
C14636 VDD.n5603 Vbias 0.03694f
C14637 VDD.n5604 Vbias 0.03694f
C14638 VDD.n5605 Vbias 0.0216f
C14639 VDD.n5606 Vbias 0.01836f
C14640 VDD.t856 Vbias 0.0169f
C14641 VDD.t449 Vbias 0.0169f
C14642 VDD.n5607 Vbias 0.07902f
C14643 VDD.t857 Vbias 0.0169f
C14644 VDD.t302 Vbias 0.0169f
C14645 VDD.n5608 Vbias 0.07902f
C14646 VDD.n5609 Vbias 0.03023f
C14647 VDD.n5610 Vbias 0.01699f
C14648 VDD.n5611 Vbias 0.03902f
C14649 VDD.n5612 Vbias 0.03694f
C14650 VDD.n5613 Vbias 0.0216f
C14651 VDD.n5614 Vbias 0.01836f
C14652 VDD.t1054 Vbias 0.46278f
C14653 VDD.n5615 Vbias 0.03694f
C14654 VDD.n5616 Vbias 0.03694f
C14655 VDD.n5617 Vbias 0.06648f
C14656 VDD.n5618 Vbias 0.03639f
C14657 VDD.t303 Vbias 0.46278f
C14658 VDD.n5619 Vbias 0.03694f
C14659 VDD.n5620 Vbias 0.03694f
C14660 VDD.n5621 Vbias 0.0216f
C14661 VDD.n5622 Vbias 0.01836f
C14662 VDD.t1055 Vbias 0.017f
C14663 VDD.n5623 Vbias 0.01309f
C14664 VDD.n5624 Vbias 0.05322f
C14665 VDD.n5625 Vbias 0.01699f
C14666 VDD.n5626 Vbias 0.03902f
C14667 VDD.n5627 Vbias 0.03694f
C14668 VDD.n5628 Vbias 0.0216f
C14669 VDD.n5629 Vbias 0.01836f
C14670 VDD.n5630 Vbias 0.03639f
C14671 VDD.t548 Vbias 0.46278f
C14672 VDD.n5631 Vbias 0.03694f
C14673 VDD.n5632 Vbias 0.03694f
C14674 VDD.n5633 Vbias 0.0216f
C14675 VDD.n5634 Vbias 0.01836f
C14676 VDD.t304 Vbias 0.0169f
C14677 VDD.t549 Vbias 0.0169f
C14678 VDD.n5635 Vbias 0.07902f
C14679 VDD.t450 Vbias 0.0169f
C14680 VDD.t924 Vbias 0.0169f
C14681 VDD.n5636 Vbias 0.07902f
C14682 VDD.n5637 Vbias 0.03023f
C14683 VDD.n5638 Vbias 0.02305f
C14684 VDD.n5639 Vbias 0.03902f
C14685 VDD.n5640 Vbias 0.03694f
C14686 VDD.n5641 Vbias 0.0216f
C14687 VDD.n5642 Vbias 0.01836f
C14688 VDD.n5643 Vbias 0.03639f
C14689 VDD.t43 Vbias 0.46278f
C14690 VDD.n5644 Vbias 0.03694f
C14691 VDD.n5645 Vbias 0.03694f
C14692 VDD.n5646 Vbias 0.0216f
C14693 VDD.n5647 Vbias 0.01836f
C14694 VDD.n5648 Vbias 0.01914f
C14695 VDD.n5649 Vbias 0.03902f
C14696 VDD.n5650 Vbias 0.03694f
C14697 VDD.n5651 Vbias 0.0216f
C14698 VDD.n5652 Vbias 0.01836f
C14699 VDD.n5653 Vbias 0.03639f
C14700 VDD.t1028 Vbias 0.46278f
C14701 VDD.n5654 Vbias 0.03694f
C14702 VDD.n5655 Vbias 0.03694f
C14703 VDD.n5656 Vbias 0.0216f
C14704 VDD.n5657 Vbias 0.01836f
C14705 VDD.t44 Vbias 0.017f
C14706 VDD.t773 Vbias 0.017f
C14707 VDD.n5658 Vbias 0.09713f
C14708 VDD.n5659 Vbias 0.01699f
C14709 VDD.n5660 Vbias 0.03902f
C14710 VDD.n5661 Vbias 0.03694f
C14711 VDD.n5662 Vbias 0.0216f
C14712 VDD.n5663 Vbias 0.01836f
C14713 VDD.n5664 Vbias 0.03639f
C14714 VDD.t377 Vbias 0.46278f
C14715 VDD.n5665 Vbias 0.03694f
C14716 VDD.n5666 Vbias 0.03694f
C14717 VDD.n5667 Vbias 0.0216f
C14718 VDD.n5668 Vbias 0.01836f
C14719 VDD.t1029 Vbias 0.0169f
C14720 VDD.t378 Vbias 0.0169f
C14721 VDD.n5669 Vbias 0.07902f
C14722 VDD.t1070 Vbias 0.0169f
C14723 VDD.t624 Vbias 0.0169f
C14724 VDD.n5670 Vbias 0.07902f
C14725 VDD.n5671 Vbias 0.03023f
C14726 VDD.n5672 Vbias 0.02305f
C14727 VDD.n5673 Vbias 0.03902f
C14728 VDD.n5674 Vbias 0.03694f
C14729 VDD.n5675 Vbias 0.0216f
C14730 VDD.n5676 Vbias 0.01836f
C14731 VDD.n5677 Vbias 0.03639f
C14732 VDD.t53 Vbias 0.46278f
C14733 VDD.n5678 Vbias 0.03694f
C14734 VDD.n5679 Vbias 0.03694f
C14735 VDD.n5680 Vbias 0.0216f
C14736 VDD.n5681 Vbias 0.01836f
C14737 VDD.n5682 Vbias 0.01914f
C14738 VDD.n5683 Vbias 0.03902f
C14739 VDD.n5684 Vbias 0.03694f
C14740 VDD.n5685 Vbias 0.0216f
C14741 VDD.n5686 Vbias 0.01836f
C14742 VDD.t209 Vbias 0.54191f
C14743 VDD.n5687 Vbias 0.03694f
C14744 VDD.n5688 Vbias 0.03694f
C14745 VDD.n5689 Vbias 0.0216f
C14746 VDD.n5691 Vbias 0.45845f
C14747 VDD.n5692 Vbias 0.01999f
C14748 VDD.t807 Vbias 0.017f
C14749 VDD.t54 Vbias 0.017f
C14750 VDD.n5693 Vbias 0.09713f
C14751 VDD.t210 Vbias 0.017f
C14752 VDD.t997 Vbias 0.0169f
C14753 VDD.t570 Vbias 0.0169f
C14754 VDD.n5694 Vbias 0.07902f
C14755 VDD.t208 Vbias 0.0169f
C14756 VDD.t352 Vbias 0.0169f
C14757 VDD.n5695 Vbias 0.07902f
C14758 VDD.n5696 Vbias 0.03023f
C14759 VDD.n5697 Vbias 0.03902f
C14760 VDD.n5698 Vbias 0.03694f
C14761 VDD.n5699 Vbias 0.03902f
C14762 VDD.n5700 Vbias 0.03639f
C14763 VDD.n5701 Vbias 0.03639f
C14764 VDD.n5702 Vbias 0.50118f
C14765 VDD.n5703 Vbias 0.01836f
C14766 VDD.n5704 Vbias 0.01836f
C14767 VDD.n5705 Vbias 0.0216f
C14768 VDD.n5706 Vbias 0.03694f
C14769 VDD.n5707 Vbias 0.03639f
C14770 VDD.t351 Vbias 0.46278f
C14771 VDD.n5708 Vbias 0.03694f
C14772 VDD.n5709 Vbias 0.03694f
C14773 VDD.n5710 Vbias 0.0216f
C14774 VDD.n5711 Vbias 0.01836f
C14775 VDD.n5712 Vbias 0.02305f
C14776 VDD.n5713 Vbias 0.03902f
C14777 VDD.n5714 Vbias 0.03694f
C14778 VDD.n5715 Vbias 0.0216f
C14779 VDD.n5716 Vbias 0.01836f
C14780 VDD.n5717 Vbias 0.03639f
C14781 VDD.t25 Vbias 0.46278f
C14782 VDD.n5718 Vbias 0.03694f
C14783 VDD.n5719 Vbias 0.03694f
C14784 VDD.n5720 Vbias 0.0216f
C14785 VDD.n5721 Vbias 0.01836f
C14786 VDD.n5722 Vbias 0.01914f
C14787 VDD.n5723 Vbias 0.03902f
C14788 VDD.n5724 Vbias 0.03694f
C14789 VDD.n5725 Vbias 0.0216f
C14790 VDD.n5726 Vbias 0.01836f
C14791 VDD.n5727 Vbias 0.03639f
C14792 VDD.t529 Vbias 0.46278f
C14793 VDD.n5728 Vbias 0.03694f
C14794 VDD.n5729 Vbias 0.03694f
C14795 VDD.n5730 Vbias 0.0216f
C14796 VDD.n5731 Vbias 0.01836f
C14797 VDD.t26 Vbias 0.017f
C14798 VDD.t759 Vbias 0.017f
C14799 VDD.n5732 Vbias 0.09713f
C14800 VDD.n5733 Vbias 0.01699f
C14801 VDD.n5734 Vbias 0.03902f
C14802 VDD.n5735 Vbias 0.03694f
C14803 VDD.n5736 Vbias 0.0216f
C14804 VDD.n5737 Vbias 0.01836f
C14805 VDD.n5738 Vbias 0.03639f
C14806 VDD.t490 Vbias 0.46278f
C14807 VDD.n5739 Vbias 0.03694f
C14808 VDD.n5740 Vbias 0.03694f
C14809 VDD.n5741 Vbias 0.0216f
C14810 VDD.n5742 Vbias 0.01836f
C14811 VDD.t531 Vbias 0.0169f
C14812 VDD.t491 Vbias 0.0169f
C14813 VDD.n5743 Vbias 0.07902f
C14814 VDD.t530 Vbias 0.0169f
C14815 VDD.t500 Vbias 0.0169f
C14816 VDD.n5744 Vbias 0.07902f
C14817 VDD.n5745 Vbias 0.03023f
C14818 VDD.n5746 Vbias 0.01699f
C14819 VDD.n5747 Vbias 0.03902f
C14820 VDD.n5748 Vbias 0.03694f
C14821 VDD.n5749 Vbias 0.0216f
C14822 VDD.n5750 Vbias 0.01836f
C14823 VDD.t1079 Vbias 0.46278f
C14824 VDD.n5751 Vbias 0.03694f
C14825 VDD.n5752 Vbias 0.03694f
C14826 VDD.n5753 Vbias 0.06648f
C14827 VDD.n5754 Vbias 0.03639f
C14828 VDD.t501 Vbias 0.46278f
C14829 VDD.n5755 Vbias 0.03694f
C14830 VDD.n5756 Vbias 0.03694f
C14831 VDD.n5757 Vbias 0.0216f
C14832 VDD.n5758 Vbias 0.01836f
C14833 VDD.t1080 Vbias 0.017f
C14834 VDD.n5759 Vbias 0.01309f
C14835 VDD.n5760 Vbias 0.05322f
C14836 VDD.n5761 Vbias 0.01699f
C14837 VDD.n5762 Vbias 0.03902f
C14838 VDD.n5763 Vbias 0.03694f
C14839 VDD.n5764 Vbias 0.0216f
C14840 VDD.n5765 Vbias 0.01836f
C14841 VDD.n5766 Vbias 0.03639f
C14842 VDD.t299 Vbias 0.46278f
C14843 VDD.n5767 Vbias 0.03694f
C14844 VDD.n5768 Vbias 0.03694f
C14845 VDD.n5769 Vbias 0.0216f
C14846 VDD.n5770 Vbias 0.01836f
C14847 VDD.t502 Vbias 0.0169f
C14848 VDD.t333 Vbias 0.0169f
C14849 VDD.n5771 Vbias 0.07902f
C14850 VDD.t816 Vbias 0.0169f
C14851 VDD.t300 Vbias 0.0169f
C14852 VDD.n5772 Vbias 0.07902f
C14853 VDD.n5773 Vbias 0.03023f
C14854 VDD.n5774 Vbias 0.02305f
C14855 VDD.n5775 Vbias 0.03902f
C14856 VDD.n5776 Vbias 0.03694f
C14857 VDD.n5777 Vbias 0.0216f
C14858 VDD.n5778 Vbias 0.01836f
C14859 VDD.n5779 Vbias 0.03639f
C14860 VDD.t61 Vbias 0.46278f
C14861 VDD.n5780 Vbias 0.03694f
C14862 VDD.n5781 Vbias 0.03694f
C14863 VDD.n5782 Vbias 0.0216f
C14864 VDD.n5783 Vbias 0.01836f
C14865 VDD.n5784 Vbias 0.01914f
C14866 VDD.n5785 Vbias 0.03902f
C14867 VDD.n5786 Vbias 0.03694f
C14868 VDD.n5787 Vbias 0.0216f
C14869 VDD.n5788 Vbias 0.01836f
C14870 VDD.n5789 Vbias 0.03639f
C14871 VDD.t1056 Vbias 0.46278f
C14872 VDD.n5790 Vbias 0.03694f
C14873 VDD.n5791 Vbias 0.03694f
C14874 VDD.n5792 Vbias 0.0216f
C14875 VDD.n5793 Vbias 0.01836f
C14876 VDD.t62 Vbias 0.017f
C14877 VDD.t793 Vbias 0.017f
C14878 VDD.n5794 Vbias 0.09713f
C14879 VDD.n5795 Vbias 0.01699f
C14880 VDD.n5796 Vbias 0.03902f
C14881 VDD.n5797 Vbias 0.03694f
C14882 VDD.n5798 Vbias 0.0216f
C14883 VDD.n5799 Vbias 0.01836f
C14884 VDD.n5800 Vbias 0.03639f
C14885 VDD.t468 Vbias 0.46278f
C14886 VDD.n5801 Vbias 0.03694f
C14887 VDD.n5802 Vbias 0.03694f
C14888 VDD.n5803 Vbias 0.0216f
C14889 VDD.n5804 Vbias 0.01836f
C14890 VDD.t1057 Vbias 0.0169f
C14891 VDD.t469 Vbias 0.0169f
C14892 VDD.n5805 Vbias 0.07902f
C14893 VDD.t1088 Vbias 0.0169f
C14894 VDD.t611 Vbias 0.0169f
C14895 VDD.n5806 Vbias 0.07902f
C14896 VDD.n5807 Vbias 0.03023f
C14897 VDD.n5808 Vbias 0.02305f
C14898 VDD.n5809 Vbias 0.03902f
C14899 VDD.n5810 Vbias 0.03694f
C14900 VDD.n5811 Vbias 0.0216f
C14901 VDD.n5812 Vbias 0.01836f
C14902 VDD.n5813 Vbias 0.03639f
C14903 VDD.t107 Vbias 0.46278f
C14904 VDD.n5814 Vbias 0.03694f
C14905 VDD.n5815 Vbias 0.03694f
C14906 VDD.n5816 Vbias 0.0216f
C14907 VDD.n5817 Vbias 0.01836f
C14908 VDD.n5818 Vbias 0.01914f
C14909 VDD.n5819 Vbias 0.03902f
C14910 VDD.n5820 Vbias 0.03694f
C14911 VDD.n5821 Vbias 0.0216f
C14912 VDD.n5822 Vbias 0.01836f
C14913 VDD.t946 Vbias 0.54191f
C14914 VDD.n5823 Vbias 0.03694f
C14915 VDD.n5824 Vbias 0.03694f
C14916 VDD.n5825 Vbias 0.0216f
C14917 VDD.n5827 Vbias 0.45845f
C14918 VDD.n5828 Vbias 0.01999f
C14919 VDD.t761 Vbias 0.017f
C14920 VDD.t108 Vbias 0.017f
C14921 VDD.n5829 Vbias 0.09713f
C14922 VDD.t947 Vbias 0.017f
C14923 VDD.t918 Vbias 0.0169f
C14924 VDD.t707 Vbias 0.0169f
C14925 VDD.n5830 Vbias 0.07902f
C14926 VDD.t391 Vbias 0.0169f
C14927 VDD.t889 Vbias 0.0169f
C14928 VDD.n5831 Vbias 0.07902f
C14929 VDD.n5832 Vbias 0.03023f
C14930 VDD.n5833 Vbias 0.03902f
C14931 VDD.n5834 Vbias 0.03694f
C14932 VDD.n5835 Vbias 0.03902f
C14933 VDD.n5836 Vbias 0.03639f
C14934 VDD.n5837 Vbias 0.03639f
C14935 VDD.n5838 Vbias 0.50118f
C14936 VDD.n5839 Vbias 0.01836f
C14937 VDD.n5840 Vbias 0.01836f
C14938 VDD.n5841 Vbias 0.0216f
C14939 VDD.n5842 Vbias 0.03694f
C14940 VDD.n5843 Vbias 0.03639f
C14941 VDD.t706 Vbias 0.46278f
C14942 VDD.n5844 Vbias 0.03694f
C14943 VDD.n5845 Vbias 0.03694f
C14944 VDD.n5846 Vbias 0.0216f
C14945 VDD.n5847 Vbias 0.01836f
C14946 VDD.n5848 Vbias 0.02305f
C14947 VDD.n5849 Vbias 0.03902f
C14948 VDD.n5850 Vbias 0.03694f
C14949 VDD.n5851 Vbias 0.0216f
C14950 VDD.n5852 Vbias 0.01836f
C14951 VDD.n5853 Vbias 0.03639f
C14952 VDD.t121 Vbias 0.46278f
C14953 VDD.n5854 Vbias 0.03694f
C14954 VDD.n5855 Vbias 0.03694f
C14955 VDD.n5856 Vbias 0.0216f
C14956 VDD.n5857 Vbias 0.01836f
C14957 VDD.n5858 Vbias 0.01914f
C14958 VDD.n5859 Vbias 0.03902f
C14959 VDD.n5860 Vbias 0.03694f
C14960 VDD.n5861 Vbias 0.0216f
C14961 VDD.n5862 Vbias 0.01836f
C14962 VDD.n5863 Vbias 0.03639f
C14963 VDD.t297 Vbias 0.46278f
C14964 VDD.n5864 Vbias 0.03694f
C14965 VDD.n5865 Vbias 0.03694f
C14966 VDD.n5866 Vbias 0.0216f
C14967 VDD.n5867 Vbias 0.01836f
C14968 VDD.t779 Vbias 0.017f
C14969 VDD.t122 Vbias 0.017f
C14970 VDD.n5868 Vbias 0.09713f
C14971 VDD.n5869 Vbias 0.01699f
C14972 VDD.n5870 Vbias 0.03902f
C14973 VDD.n5871 Vbias 0.03694f
C14974 VDD.n5872 Vbias 0.0216f
C14975 VDD.n5873 Vbias 0.01836f
C14976 VDD.n5874 Vbias 0.03639f
C14977 VDD.t274 Vbias 0.46278f
C14978 VDD.n5875 Vbias 0.03694f
C14979 VDD.n5876 Vbias 0.03694f
C14980 VDD.n5877 Vbias 0.0216f
C14981 VDD.n5878 Vbias 0.01836f
C14982 VDD.t387 Vbias 0.0169f
C14983 VDD.t275 Vbias 0.0169f
C14984 VDD.n5879 Vbias 0.07902f
C14985 VDD.t298 Vbias 0.0169f
C14986 VDD.t951 Vbias 0.0169f
C14987 VDD.n5880 Vbias 0.07902f
C14988 VDD.n5881 Vbias 0.03023f
C14989 VDD.n5882 Vbias 0.01699f
C14990 VDD.n5883 Vbias 0.03902f
C14991 VDD.n5884 Vbias 0.03694f
C14992 VDD.n5885 Vbias 0.0216f
C14993 VDD.n5886 Vbias 0.01836f
C14994 VDD.t1024 Vbias 0.46278f
C14995 VDD.n5887 Vbias 0.03694f
C14996 VDD.n5888 Vbias 0.03694f
C14997 VDD.n5889 Vbias 0.06648f
C14998 VDD.n5890 Vbias 0.03639f
C14999 VDD.t276 Vbias 0.46278f
C15000 VDD.n5891 Vbias 0.03694f
C15001 VDD.n5892 Vbias 0.03694f
C15002 VDD.n5893 Vbias 0.0216f
C15003 VDD.n5894 Vbias 0.01836f
C15004 VDD.t1025 Vbias 0.017f
C15005 VDD.n5895 Vbias 0.01309f
C15006 VDD.n5896 Vbias 0.05322f
C15007 VDD.n5897 Vbias 0.01699f
C15008 VDD.n5898 Vbias 0.03902f
C15009 VDD.n5899 Vbias 0.03694f
C15010 VDD.n5900 Vbias 0.0216f
C15011 VDD.n5901 Vbias 0.01836f
C15012 VDD.n5902 Vbias 0.03639f
C15013 VDD.t219 Vbias 0.46278f
C15014 VDD.n5903 Vbias 0.03694f
C15015 VDD.n5904 Vbias 0.03694f
C15016 VDD.n5905 Vbias 0.0216f
C15017 VDD.n5906 Vbias 0.01836f
C15018 VDD.t952 Vbias 0.0169f
C15019 VDD.t220 Vbias 0.0169f
C15020 VDD.n5907 Vbias 0.07902f
C15021 VDD.t277 Vbias 0.0169f
C15022 VDD.t899 Vbias 0.0169f
C15023 VDD.n5908 Vbias 0.07902f
C15024 VDD.n5909 Vbias 0.03023f
C15025 VDD.n5910 Vbias 0.02305f
C15026 VDD.n5911 Vbias 0.03902f
C15027 VDD.n5912 Vbias 0.03694f
C15028 VDD.n5913 Vbias 0.0216f
C15029 VDD.n5914 Vbias 0.01836f
C15030 VDD.n5915 Vbias 0.03639f
C15031 VDD.t125 Vbias 0.46278f
C15032 VDD.n5916 Vbias 0.03694f
C15033 VDD.n5917 Vbias 0.03694f
C15034 VDD.n5918 Vbias 0.0216f
C15035 VDD.n5919 Vbias 0.01836f
C15036 VDD.n5920 Vbias 0.01914f
C15037 VDD.n5921 Vbias 0.03902f
C15038 VDD.n5922 Vbias 0.03694f
C15039 VDD.n5923 Vbias 0.0216f
C15040 VDD.n5924 Vbias 0.01836f
C15041 VDD.n5925 Vbias 0.03639f
C15042 VDD.t1000 Vbias 0.46278f
C15043 VDD.n5926 Vbias 0.03694f
C15044 VDD.n5927 Vbias 0.03694f
C15045 VDD.n5928 Vbias 0.0216f
C15046 VDD.n5929 Vbias 0.01836f
C15047 VDD.t781 Vbias 0.017f
C15048 VDD.t126 Vbias 0.017f
C15049 VDD.n5930 Vbias 0.09713f
C15050 VDD.n5931 Vbias 0.01699f
C15051 VDD.n5932 Vbias 0.03902f
C15052 VDD.n5933 Vbias 0.03694f
C15053 VDD.n5934 Vbias 0.0216f
C15054 VDD.n5935 Vbias 0.01836f
C15055 VDD.n5936 Vbias 0.03639f
C15056 VDD.t343 Vbias 0.46278f
C15057 VDD.n5937 Vbias 0.03694f
C15058 VDD.n5938 Vbias 0.03694f
C15059 VDD.n5939 Vbias 0.0216f
C15060 VDD.n5940 Vbias 0.01836f
C15061 VDD.t1001 Vbias 0.0169f
C15062 VDD.t344 Vbias 0.0169f
C15063 VDD.n5941 Vbias 0.07902f
C15064 VDD.t1044 Vbias 0.0169f
C15065 VDD.t563 Vbias 0.0169f
C15066 VDD.n5942 Vbias 0.07902f
C15067 VDD.n5943 Vbias 0.03023f
C15068 VDD.n5944 Vbias 0.02305f
C15069 VDD.n5945 Vbias 0.03902f
C15070 VDD.n5946 Vbias 0.03694f
C15071 VDD.n5947 Vbias 0.0216f
C15072 VDD.n5948 Vbias 0.01836f
C15073 VDD.n5949 Vbias 0.03639f
C15074 VDD.t85 Vbias 0.46278f
C15075 VDD.n5950 Vbias 0.03694f
C15076 VDD.n5951 Vbias 0.03694f
C15077 VDD.n5952 Vbias 0.0216f
C15078 VDD.n5953 Vbias 0.01836f
C15079 VDD.n5954 Vbias 0.01914f
C15080 VDD.n5955 Vbias 0.03902f
C15081 VDD.n5956 Vbias 0.03694f
C15082 VDD.n5957 Vbias 0.0216f
C15083 VDD.n5958 Vbias 0.01836f
C15084 VDD.t345 Vbias 0.54191f
C15085 VDD.n5959 Vbias 0.03694f
C15086 VDD.n5960 Vbias 0.03694f
C15087 VDD.n5961 Vbias 0.0216f
C15088 VDD.n5963 Vbias 0.45845f
C15089 VDD.n5964 Vbias 0.01999f
C15090 VDD.t86 Vbias 0.017f
C15091 VDD.t719 Vbias 0.017f
C15092 VDD.n5965 Vbias 0.09713f
C15093 VDD.t346 Vbias 0.017f
C15094 VDD.n5966 Vbias 0.05322f
C15095 VDD.n5967 Vbias 0.01309f
C15096 VDD.n5968 Vbias 0.06648f
C15097 VDD.n5969 Vbias 0.01999f
C15098 VDD.n5970 Vbias 0.03639f
C15099 VDD.n5971 Vbias 0.50118f
C15100 VDD.n5972 Vbias 0.01836f
C15101 VDD.n5973 Vbias 0.03639f
C15102 VDD.n5974 Vbias 0.50118f
C15103 VDD.n5975 Vbias 0.03639f
C15104 VDD.n5976 Vbias 0.03694f
C15105 VDD.n5977 Vbias 0.04583f
C15106 VDD.n5978 Vbias 0.03902f
C15107 VDD.n5979 Vbias 0.01836f
C15108 VDD.n5980 Vbias 0.03639f
C15109 VDD.n5981 Vbias 0.37318f
C15110 VDD.n5982 Vbias 0.01836f
C15111 VDD.n5983 Vbias 0.03639f
C15112 VDD.n5984 Vbias 0.37318f
C15113 VDD.n5985 Vbias 0.03639f
C15114 VDD.n5986 Vbias 0.03694f
C15115 VDD.n5987 Vbias 0.04583f
C15116 VDD.n5988 Vbias 0.03902f
C15117 VDD.n5989 Vbias 0.01836f
C15118 VDD.n5990 Vbias 0.03639f
C15119 VDD.n5991 Vbias 0.37318f
C15120 VDD.n5992 Vbias 0.01836f
C15121 VDD.n5993 Vbias 0.03639f
C15122 VDD.n5994 Vbias 0.37318f
C15123 VDD.n5995 Vbias 0.03639f
C15124 VDD.n5996 Vbias 0.03694f
C15125 VDD.n5997 Vbias 0.04583f
C15126 VDD.n5998 Vbias 0.03902f
C15127 VDD.n5999 Vbias 0.01836f
C15128 VDD.n6000 Vbias 0.03639f
C15129 VDD.n6001 Vbias 0.50118f
C15130 VDD.n6002 Vbias 0.01836f
C15131 VDD.n6003 Vbias 0.03639f
C15132 VDD.n6004 Vbias 0.50118f
C15133 VDD.n6005 Vbias 0.03639f
C15134 VDD.n6006 Vbias 0.03694f
C15135 VDD.n6007 Vbias 0.04583f
C15136 VDD.n6008 Vbias 0.03902f
C15137 VDD.n6009 Vbias 0.01836f
C15138 VDD.n6010 Vbias 0.03639f
C15139 VDD.n6011 Vbias 0.37318f
C15140 VDD.n6012 Vbias 0.01836f
C15141 VDD.n6013 Vbias 0.03639f
C15142 VDD.n6014 Vbias 0.37318f
C15143 VDD.n6015 Vbias 0.03639f
C15144 VDD.n6016 Vbias 0.03694f
C15145 VDD.n6017 Vbias 0.04583f
C15146 VDD.n6018 Vbias 0.03902f
C15147 VDD.n6019 Vbias 0.01836f
C15148 VDD.n6020 Vbias 0.03639f
C15149 VDD.n6021 Vbias 0.37318f
C15150 VDD.n6022 Vbias 0.01836f
C15151 VDD.n6023 Vbias 0.03639f
C15152 VDD.n6024 Vbias 0.37318f
C15153 VDD.n6025 Vbias 0.03639f
C15154 VDD.n6026 Vbias 0.03694f
C15155 VDD.n6027 Vbias 0.04583f
C15156 VDD.n6028 Vbias 0.03902f
C15157 VDD.n6029 Vbias 0.01836f
C15158 VDD.n6030 Vbias 0.03639f
C15159 VDD.n6031 Vbias 0.50118f
C15160 VDD.n6032 Vbias 0.50118f
C15161 VDD.n6033 Vbias 0.03639f
C15162 VDD.n6034 Vbias 0.01999f
C15163 VDD.n6035 Vbias 0.0216f
C15164 VDD.n6036 Vbias 0.01999f
C15165 VDD.n6037 Vbias 0.03639f
C15166 VDD.n6038 Vbias 0.50118f
C15167 VDD.n6039 Vbias 0.01836f
C15168 VDD.n6040 Vbias 0.03639f
C15169 VDD.n6041 Vbias 0.50118f
C15170 VDD.n6042 Vbias 0.03639f
C15171 VDD.n6043 Vbias 0.03694f
C15172 VDD.n6044 Vbias 0.04583f
C15173 VDD.n6045 Vbias 0.03902f
C15174 VDD.n6046 Vbias 0.01836f
C15175 VDD.n6047 Vbias 0.03639f
C15176 VDD.n6048 Vbias 0.37318f
C15177 VDD.n6049 Vbias 0.01836f
C15178 VDD.n6050 Vbias 0.03639f
C15179 VDD.n6051 Vbias 0.37318f
C15180 VDD.n6052 Vbias 0.03639f
C15181 VDD.n6053 Vbias 0.03694f
C15182 VDD.n6054 Vbias 0.04583f
C15183 VDD.n6055 Vbias 0.03902f
C15184 VDD.n6056 Vbias 0.01836f
C15185 VDD.n6057 Vbias 0.03639f
C15186 VDD.n6058 Vbias 0.50118f
C15187 VDD.n6059 Vbias 0.01836f
C15188 VDD.n6060 Vbias 0.03639f
C15189 VDD.n6061 Vbias 0.50118f
C15190 VDD.n6062 Vbias 0.03639f
C15191 VDD.n6063 Vbias 0.03694f
C15192 VDD.n6064 Vbias 0.04583f
C15193 VDD.n6065 Vbias 0.03902f
C15194 VDD.n6066 Vbias 0.01836f
C15195 VDD.n6067 Vbias 0.03639f
C15196 VDD.n6068 Vbias 0.37318f
C15197 VDD.n6069 Vbias 0.01836f
C15198 VDD.n6070 Vbias 0.03639f
C15199 VDD.n6071 Vbias 0.37318f
C15200 VDD.n6072 Vbias 0.03639f
C15201 VDD.n6073 Vbias 0.03694f
C15202 VDD.n6074 Vbias 0.04583f
C15203 VDD.n6075 Vbias 0.03902f
C15204 VDD.n6076 Vbias 0.01836f
C15205 VDD.n6077 Vbias 0.03639f
C15206 VDD.n6078 Vbias 0.37318f
C15207 VDD.n6079 Vbias 0.37318f
C15208 VDD.n6080 Vbias 0.03639f
C15209 VDD.n6081 Vbias 0.03639f
C15210 VDD.n6082 Vbias 0.01836f
C15211 VDD.n6083 Vbias 0.01836f
C15212 VDD.n6084 Vbias 0.0216f
C15213 VDD.n6085 Vbias 0.03694f
C15214 VDD.t390 Vbias 0.46278f
C15215 VDD.n6086 Vbias 0.03694f
C15216 VDD.n6087 Vbias 0.04583f
C15217 VDD.n6088 Vbias 0.074f
C15218 VDD.n6089 Vbias 0.05322f
C15219 VDD.n6090 Vbias 0.01309f
C15220 VDD.n6091 Vbias 0.06648f
C15221 VDD.n6092 Vbias 0.01999f
C15222 VDD.n6093 Vbias 0.03639f
C15223 VDD.n6094 Vbias 0.50118f
C15224 VDD.n6095 Vbias 0.01836f
C15225 VDD.n6096 Vbias 0.03639f
C15226 VDD.n6097 Vbias 0.50118f
C15227 VDD.n6098 Vbias 0.03639f
C15228 VDD.n6099 Vbias 0.03694f
C15229 VDD.n6100 Vbias 0.04583f
C15230 VDD.n6101 Vbias 0.03902f
C15231 VDD.n6102 Vbias 0.01836f
C15232 VDD.n6103 Vbias 0.03639f
C15233 VDD.n6104 Vbias 0.37318f
C15234 VDD.n6105 Vbias 0.01836f
C15235 VDD.n6106 Vbias 0.03639f
C15236 VDD.n6107 Vbias 0.37318f
C15237 VDD.n6108 Vbias 0.03639f
C15238 VDD.n6109 Vbias 0.03694f
C15239 VDD.n6110 Vbias 0.04583f
C15240 VDD.n6111 Vbias 0.03902f
C15241 VDD.n6112 Vbias 0.01836f
C15242 VDD.n6113 Vbias 0.03639f
C15243 VDD.n6114 Vbias 0.37318f
C15244 VDD.n6115 Vbias 0.01836f
C15245 VDD.n6116 Vbias 0.03639f
C15246 VDD.n6117 Vbias 0.37318f
C15247 VDD.n6118 Vbias 0.03639f
C15248 VDD.n6119 Vbias 0.03694f
C15249 VDD.n6120 Vbias 0.04583f
C15250 VDD.n6121 Vbias 0.03902f
C15251 VDD.n6122 Vbias 0.01836f
C15252 VDD.n6123 Vbias 0.03639f
C15253 VDD.n6124 Vbias 0.50118f
C15254 VDD.n6125 Vbias 0.01836f
C15255 VDD.n6126 Vbias 0.03639f
C15256 VDD.n6127 Vbias 0.50118f
C15257 VDD.n6128 Vbias 0.03639f
C15258 VDD.n6129 Vbias 0.03694f
C15259 VDD.n6130 Vbias 0.04583f
C15260 VDD.n6131 Vbias 0.03902f
C15261 VDD.n6132 Vbias 0.01836f
C15262 VDD.n6133 Vbias 0.03639f
C15263 VDD.n6134 Vbias 0.37318f
C15264 VDD.n6135 Vbias 0.01836f
C15265 VDD.n6136 Vbias 0.03639f
C15266 VDD.n6137 Vbias 0.37318f
C15267 VDD.n6138 Vbias 0.03639f
C15268 VDD.n6139 Vbias 0.03694f
C15269 VDD.n6140 Vbias 0.04583f
C15270 VDD.n6141 Vbias 0.03902f
C15271 VDD.n6142 Vbias 0.01836f
C15272 VDD.n6143 Vbias 0.03639f
C15273 VDD.n6144 Vbias 0.37318f
C15274 VDD.n6145 Vbias 0.01836f
C15275 VDD.n6146 Vbias 0.03639f
C15276 VDD.n6147 Vbias 0.37318f
C15277 VDD.n6148 Vbias 0.03639f
C15278 VDD.n6149 Vbias 0.03694f
C15279 VDD.n6150 Vbias 0.04583f
C15280 VDD.n6151 Vbias 0.03902f
C15281 VDD.n6152 Vbias 0.01836f
C15282 VDD.n6153 Vbias 0.03639f
C15283 VDD.n6154 Vbias 0.50118f
C15284 VDD.n6155 Vbias 0.50118f
C15285 VDD.n6156 Vbias 0.03639f
C15286 VDD.n6157 Vbias 0.01999f
C15287 VDD.n6158 Vbias 0.0216f
C15288 VDD.n6159 Vbias 0.01999f
C15289 VDD.n6160 Vbias 0.03639f
C15290 VDD.n6161 Vbias 0.50118f
C15291 VDD.n6162 Vbias 0.01836f
C15292 VDD.n6163 Vbias 0.03639f
C15293 VDD.n6164 Vbias 0.50118f
C15294 VDD.n6165 Vbias 0.03639f
C15295 VDD.n6166 Vbias 0.03694f
C15296 VDD.n6167 Vbias 0.04583f
C15297 VDD.n6168 Vbias 0.03902f
C15298 VDD.n6169 Vbias 0.01836f
C15299 VDD.n6170 Vbias 0.03639f
C15300 VDD.n6171 Vbias 0.37318f
C15301 VDD.n6172 Vbias 0.01836f
C15302 VDD.n6173 Vbias 0.03639f
C15303 VDD.n6174 Vbias 0.37318f
C15304 VDD.n6175 Vbias 0.03639f
C15305 VDD.n6176 Vbias 0.03694f
C15306 VDD.n6177 Vbias 0.04583f
C15307 VDD.n6178 Vbias 0.03902f
C15308 VDD.n6179 Vbias 0.01836f
C15309 VDD.n6180 Vbias 0.03639f
C15310 VDD.n6181 Vbias 0.50118f
C15311 VDD.n6182 Vbias 0.01836f
C15312 VDD.n6183 Vbias 0.03639f
C15313 VDD.n6184 Vbias 0.50118f
C15314 VDD.n6185 Vbias 0.03639f
C15315 VDD.n6186 Vbias 0.03694f
C15316 VDD.n6187 Vbias 0.04583f
C15317 VDD.n6188 Vbias 0.03902f
C15318 VDD.n6189 Vbias 0.01836f
C15319 VDD.n6190 Vbias 0.03639f
C15320 VDD.n6191 Vbias 0.37318f
C15321 VDD.n6192 Vbias 0.01836f
C15322 VDD.n6193 Vbias 0.03639f
C15323 VDD.n6194 Vbias 0.37318f
C15324 VDD.n6195 Vbias 0.03639f
C15325 VDD.n6196 Vbias 0.03694f
C15326 VDD.n6197 Vbias 0.04583f
C15327 VDD.n6198 Vbias 0.03902f
C15328 VDD.n6199 Vbias 0.01836f
C15329 VDD.n6200 Vbias 0.03639f
C15330 VDD.n6201 Vbias 0.37318f
C15331 VDD.n6202 Vbias 0.37318f
C15332 VDD.n6203 Vbias 0.03639f
C15333 VDD.n6204 Vbias 0.03639f
C15334 VDD.n6205 Vbias 0.01836f
C15335 VDD.n6206 Vbias 0.01836f
C15336 VDD.n6207 Vbias 0.0216f
C15337 VDD.n6208 Vbias 0.03694f
C15338 VDD.t207 Vbias 0.46278f
C15339 VDD.n6209 Vbias 0.03694f
C15340 VDD.n6210 Vbias 0.04583f
C15341 VDD.n6211 Vbias 0.074f
C15342 VDD.n6212 Vbias 0.05322f
C15343 VDD.n6213 Vbias 0.01309f
C15344 VDD.n6214 Vbias 0.06648f
C15345 VDD.n6215 Vbias 0.01999f
C15346 VDD.n6216 Vbias 0.03639f
C15347 VDD.n6217 Vbias 0.50118f
C15348 VDD.n6218 Vbias 0.01836f
C15349 VDD.n6219 Vbias 0.03639f
C15350 VDD.n6220 Vbias 0.50118f
C15351 VDD.n6221 Vbias 0.03639f
C15352 VDD.n6222 Vbias 0.03694f
C15353 VDD.n6223 Vbias 0.04583f
C15354 VDD.n6224 Vbias 0.03902f
C15355 VDD.n6225 Vbias 0.01836f
C15356 VDD.n6226 Vbias 0.03639f
C15357 VDD.n6227 Vbias 0.37318f
C15358 VDD.n6228 Vbias 0.01836f
C15359 VDD.n6229 Vbias 0.03639f
C15360 VDD.n6230 Vbias 0.37318f
C15361 VDD.n6231 Vbias 0.03639f
C15362 VDD.n6232 Vbias 0.03694f
C15363 VDD.n6233 Vbias 0.04583f
C15364 VDD.n6234 Vbias 0.03902f
C15365 VDD.n6235 Vbias 0.01836f
C15366 VDD.n6236 Vbias 0.03639f
C15367 VDD.n6237 Vbias 0.37318f
C15368 VDD.n6238 Vbias 0.01836f
C15369 VDD.n6239 Vbias 0.03639f
C15370 VDD.n6240 Vbias 0.37318f
C15371 VDD.n6241 Vbias 0.03639f
C15372 VDD.n6242 Vbias 0.03694f
C15373 VDD.n6243 Vbias 0.04583f
C15374 VDD.n6244 Vbias 0.03902f
C15375 VDD.n6245 Vbias 0.01836f
C15376 VDD.n6246 Vbias 0.03639f
C15377 VDD.n6247 Vbias 0.50118f
C15378 VDD.n6248 Vbias 0.01836f
C15379 VDD.n6249 Vbias 0.03639f
C15380 VDD.n6250 Vbias 0.50118f
C15381 VDD.n6251 Vbias 0.03639f
C15382 VDD.n6252 Vbias 0.03694f
C15383 VDD.n6253 Vbias 0.04583f
C15384 VDD.n6254 Vbias 0.03902f
C15385 VDD.n6255 Vbias 0.01836f
C15386 VDD.n6256 Vbias 0.03639f
C15387 VDD.n6257 Vbias 0.37318f
C15388 VDD.n6258 Vbias 0.01836f
C15389 VDD.n6259 Vbias 0.03639f
C15390 VDD.n6260 Vbias 0.37318f
C15391 VDD.n6261 Vbias 0.03639f
C15392 VDD.n6262 Vbias 0.03694f
C15393 VDD.n6263 Vbias 0.04583f
C15394 VDD.n6264 Vbias 0.03902f
C15395 VDD.n6265 Vbias 0.01836f
C15396 VDD.n6266 Vbias 0.03639f
C15397 VDD.n6267 Vbias 0.37318f
C15398 VDD.n6268 Vbias 0.01836f
C15399 VDD.n6269 Vbias 0.03639f
C15400 VDD.n6270 Vbias 0.37318f
C15401 VDD.n6271 Vbias 0.03639f
C15402 VDD.n6272 Vbias 0.03694f
C15403 VDD.n6273 Vbias 0.04583f
C15404 VDD.n6274 Vbias 0.03902f
C15405 VDD.n6275 Vbias 0.01836f
C15406 VDD.n6276 Vbias 0.03639f
C15407 VDD.n6277 Vbias 0.50118f
C15408 VDD.n6278 Vbias 0.50118f
C15409 VDD.n6279 Vbias 0.03639f
C15410 VDD.n6280 Vbias 0.01999f
C15411 VDD.n6281 Vbias 0.0216f
C15412 VDD.n6282 Vbias 0.01999f
C15413 VDD.n6283 Vbias 0.03639f
C15414 VDD.n6284 Vbias 0.50118f
C15415 VDD.n6285 Vbias 0.01836f
C15416 VDD.n6286 Vbias 0.03639f
C15417 VDD.n6287 Vbias 0.50118f
C15418 VDD.n6288 Vbias 0.03639f
C15419 VDD.n6289 Vbias 0.03694f
C15420 VDD.n6290 Vbias 0.04583f
C15421 VDD.n6291 Vbias 0.03902f
C15422 VDD.n6292 Vbias 0.01836f
C15423 VDD.n6293 Vbias 0.03639f
C15424 VDD.n6294 Vbias 0.37318f
C15425 VDD.n6295 Vbias 0.01836f
C15426 VDD.n6296 Vbias 0.03639f
C15427 VDD.n6297 Vbias 0.37318f
C15428 VDD.n6298 Vbias 0.03639f
C15429 VDD.n6299 Vbias 0.03694f
C15430 VDD.n6300 Vbias 0.04583f
C15431 VDD.n6301 Vbias 0.03902f
C15432 VDD.n6302 Vbias 0.01836f
C15433 VDD.n6303 Vbias 0.03639f
C15434 VDD.n6304 Vbias 0.50118f
C15435 VDD.n6305 Vbias 0.01836f
C15436 VDD.n6306 Vbias 0.03639f
C15437 VDD.n6307 Vbias 0.50118f
C15438 VDD.n6308 Vbias 0.03639f
C15439 VDD.n6309 Vbias 0.03694f
C15440 VDD.n6310 Vbias 0.04583f
C15441 VDD.n6311 Vbias 0.03902f
C15442 VDD.n6312 Vbias 0.01836f
C15443 VDD.n6313 Vbias 0.03639f
C15444 VDD.n6314 Vbias 0.37318f
C15445 VDD.n6315 Vbias 0.01836f
C15446 VDD.n6316 Vbias 0.03639f
C15447 VDD.n6317 Vbias 0.37318f
C15448 VDD.n6318 Vbias 0.03639f
C15449 VDD.n6319 Vbias 0.03694f
C15450 VDD.n6320 Vbias 0.04583f
C15451 VDD.n6321 Vbias 0.03902f
C15452 VDD.n6322 Vbias 0.01836f
C15453 VDD.n6323 Vbias 0.03639f
C15454 VDD.n6324 Vbias 0.37318f
C15455 VDD.n6325 Vbias 0.37318f
C15456 VDD.n6326 Vbias 0.03639f
C15457 VDD.n6327 Vbias 0.03639f
C15458 VDD.n6328 Vbias 0.01836f
C15459 VDD.n6329 Vbias 0.01836f
C15460 VDD.n6330 Vbias 0.0216f
C15461 VDD.n6331 Vbias 0.03694f
C15462 VDD.t311 Vbias 0.46278f
C15463 VDD.n6332 Vbias 0.03694f
C15464 VDD.n6333 Vbias 0.04583f
C15465 VDD.n6334 Vbias 0.074f
C15466 VDD.n6335 Vbias 0.05322f
C15467 VDD.n6336 Vbias 0.01309f
C15468 VDD.n6337 Vbias 0.06648f
C15469 VDD.n6338 Vbias 0.01999f
C15470 VDD.n6339 Vbias 0.03639f
C15471 VDD.n6340 Vbias 0.50118f
C15472 VDD.n6341 Vbias 0.01836f
C15473 VDD.n6342 Vbias 0.03639f
C15474 VDD.n6343 Vbias 0.50118f
C15475 VDD.n6344 Vbias 0.03639f
C15476 VDD.n6345 Vbias 0.03694f
C15477 VDD.n6346 Vbias 0.04583f
C15478 VDD.n6347 Vbias 0.03902f
C15479 VDD.n6348 Vbias 0.01836f
C15480 VDD.n6349 Vbias 0.03639f
C15481 VDD.n6350 Vbias 0.37318f
C15482 VDD.n6351 Vbias 0.01836f
C15483 VDD.n6352 Vbias 0.03639f
C15484 VDD.n6353 Vbias 0.37318f
C15485 VDD.n6354 Vbias 0.03639f
C15486 VDD.n6355 Vbias 0.03694f
C15487 VDD.n6356 Vbias 0.04583f
C15488 VDD.n6357 Vbias 0.03902f
C15489 VDD.n6358 Vbias 0.01836f
C15490 VDD.n6359 Vbias 0.03639f
C15491 VDD.n6360 Vbias 0.37318f
C15492 VDD.n6361 Vbias 0.01836f
C15493 VDD.n6362 Vbias 0.03639f
C15494 VDD.n6363 Vbias 0.37318f
C15495 VDD.n6364 Vbias 0.03639f
C15496 VDD.n6365 Vbias 0.03694f
C15497 VDD.n6366 Vbias 0.04583f
C15498 VDD.n6367 Vbias 0.03902f
C15499 VDD.n6368 Vbias 0.01836f
C15500 VDD.n6369 Vbias 0.03639f
C15501 VDD.n6370 Vbias 0.50118f
C15502 VDD.n6371 Vbias 0.01836f
C15503 VDD.n6372 Vbias 0.03639f
C15504 VDD.n6373 Vbias 0.50118f
C15505 VDD.n6374 Vbias 0.03639f
C15506 VDD.n6375 Vbias 0.03694f
C15507 VDD.n6376 Vbias 0.04583f
C15508 VDD.n6377 Vbias 0.03902f
C15509 VDD.n6378 Vbias 0.01836f
C15510 VDD.n6379 Vbias 0.03639f
C15511 VDD.n6380 Vbias 0.37318f
C15512 VDD.n6381 Vbias 0.01836f
C15513 VDD.n6382 Vbias 0.03639f
C15514 VDD.n6383 Vbias 0.37318f
C15515 VDD.n6384 Vbias 0.03639f
C15516 VDD.n6385 Vbias 0.03694f
C15517 VDD.n6386 Vbias 0.04583f
C15518 VDD.n6387 Vbias 0.03902f
C15519 VDD.n6388 Vbias 0.01836f
C15520 VDD.n6389 Vbias 0.03639f
C15521 VDD.n6390 Vbias 0.37318f
C15522 VDD.n6391 Vbias 0.01836f
C15523 VDD.n6392 Vbias 0.03639f
C15524 VDD.n6393 Vbias 0.37318f
C15525 VDD.n6394 Vbias 0.03639f
C15526 VDD.n6395 Vbias 0.03694f
C15527 VDD.n6396 Vbias 0.04583f
C15528 VDD.n6397 Vbias 0.03902f
C15529 VDD.n6398 Vbias 0.01836f
C15530 VDD.n6399 Vbias 0.03639f
C15531 VDD.n6400 Vbias 0.50118f
C15532 VDD.n6401 Vbias 0.50118f
C15533 VDD.n6402 Vbias 0.03639f
C15534 VDD.n6403 Vbias 0.01999f
C15535 VDD.n6404 Vbias 0.0216f
C15536 VDD.n6405 Vbias 0.01999f
C15537 VDD.n6406 Vbias 0.03639f
C15538 VDD.n6407 Vbias 0.50118f
C15539 VDD.n6408 Vbias 0.01836f
C15540 VDD.n6409 Vbias 0.03639f
C15541 VDD.n6410 Vbias 0.50118f
C15542 VDD.n6411 Vbias 0.03639f
C15543 VDD.n6412 Vbias 0.03694f
C15544 VDD.n6413 Vbias 0.04583f
C15545 VDD.n6414 Vbias 0.03902f
C15546 VDD.n6415 Vbias 0.01836f
C15547 VDD.n6416 Vbias 0.03639f
C15548 VDD.n6417 Vbias 0.37318f
C15549 VDD.n6418 Vbias 0.01836f
C15550 VDD.n6419 Vbias 0.03639f
C15551 VDD.n6420 Vbias 0.37318f
C15552 VDD.n6421 Vbias 0.03639f
C15553 VDD.n6422 Vbias 0.03694f
C15554 VDD.n6423 Vbias 0.04583f
C15555 VDD.n6424 Vbias 0.03902f
C15556 VDD.n6425 Vbias 0.01836f
C15557 VDD.n6426 Vbias 0.03639f
C15558 VDD.n6427 Vbias 0.50118f
C15559 VDD.n6428 Vbias 0.01836f
C15560 VDD.n6429 Vbias 0.03639f
C15561 VDD.n6430 Vbias 0.50118f
C15562 VDD.n6431 Vbias 0.03639f
C15563 VDD.n6432 Vbias 0.03694f
C15564 VDD.n6433 Vbias 0.04583f
C15565 VDD.n6434 Vbias 0.03902f
C15566 VDD.n6435 Vbias 0.01836f
C15567 VDD.n6436 Vbias 0.03639f
C15568 VDD.n6437 Vbias 0.37318f
C15569 VDD.n6438 Vbias 0.01836f
C15570 VDD.n6439 Vbias 0.03639f
C15571 VDD.n6440 Vbias 0.37318f
C15572 VDD.n6441 Vbias 0.03639f
C15573 VDD.n6442 Vbias 0.03694f
C15574 VDD.n6443 Vbias 0.04583f
C15575 VDD.n6444 Vbias 0.03902f
C15576 VDD.n6445 Vbias 0.01836f
C15577 VDD.n6446 Vbias 0.03639f
C15578 VDD.n6447 Vbias 0.37318f
C15579 VDD.n6448 Vbias 0.37318f
C15580 VDD.n6449 Vbias 0.03639f
C15581 VDD.n6450 Vbias 0.03639f
C15582 VDD.n6451 Vbias 0.01836f
C15583 VDD.n6452 Vbias 0.01836f
C15584 VDD.n6453 Vbias 0.0216f
C15585 VDD.n6454 Vbias 0.03694f
C15586 VDD.t658 Vbias 0.46278f
C15587 VDD.n6455 Vbias 0.03694f
C15588 VDD.n6456 Vbias 0.04583f
C15589 VDD.n6457 Vbias 0.074f
C15590 VDD.n6458 Vbias 0.05322f
C15591 VDD.n6459 Vbias 0.01309f
C15592 VDD.n6460 Vbias 0.06648f
C15593 VDD.n6461 Vbias 0.01999f
C15594 VDD.n6462 Vbias 0.03639f
C15595 VDD.n6463 Vbias 0.50118f
C15596 VDD.n6464 Vbias 0.01836f
C15597 VDD.n6465 Vbias 0.03639f
C15598 VDD.n6466 Vbias 0.50118f
C15599 VDD.n6467 Vbias 0.03639f
C15600 VDD.n6468 Vbias 0.03694f
C15601 VDD.n6469 Vbias 0.04583f
C15602 VDD.n6470 Vbias 0.03902f
C15603 VDD.n6471 Vbias 0.01836f
C15604 VDD.n6472 Vbias 0.03639f
C15605 VDD.n6473 Vbias 0.37318f
C15606 VDD.n6474 Vbias 0.01836f
C15607 VDD.n6475 Vbias 0.03639f
C15608 VDD.n6476 Vbias 0.37318f
C15609 VDD.n6477 Vbias 0.03639f
C15610 VDD.n6478 Vbias 0.03694f
C15611 VDD.n6479 Vbias 0.04583f
C15612 VDD.n6480 Vbias 0.03902f
C15613 VDD.n6481 Vbias 0.01836f
C15614 VDD.n6482 Vbias 0.03639f
C15615 VDD.n6483 Vbias 0.37318f
C15616 VDD.n6484 Vbias 0.01836f
C15617 VDD.n6485 Vbias 0.03639f
C15618 VDD.n6486 Vbias 0.37318f
C15619 VDD.n6487 Vbias 0.03639f
C15620 VDD.n6488 Vbias 0.03694f
C15621 VDD.n6489 Vbias 0.04583f
C15622 VDD.n6490 Vbias 0.03902f
C15623 VDD.n6491 Vbias 0.01836f
C15624 VDD.n6492 Vbias 0.03639f
C15625 VDD.n6493 Vbias 0.50118f
C15626 VDD.n6494 Vbias 0.01836f
C15627 VDD.n6495 Vbias 0.03639f
C15628 VDD.n6496 Vbias 0.50118f
C15629 VDD.n6497 Vbias 0.03639f
C15630 VDD.n6498 Vbias 0.03694f
C15631 VDD.n6499 Vbias 0.04583f
C15632 VDD.n6500 Vbias 0.03902f
C15633 VDD.n6501 Vbias 0.01836f
C15634 VDD.n6502 Vbias 0.03639f
C15635 VDD.n6503 Vbias 0.37318f
C15636 VDD.n6504 Vbias 0.01836f
C15637 VDD.n6505 Vbias 0.03639f
C15638 VDD.n6506 Vbias 0.37318f
C15639 VDD.n6507 Vbias 0.03639f
C15640 VDD.n6508 Vbias 0.03694f
C15641 VDD.n6509 Vbias 0.04583f
C15642 VDD.n6510 Vbias 0.03902f
C15643 VDD.n6511 Vbias 0.01836f
C15644 VDD.n6512 Vbias 0.03639f
C15645 VDD.n6513 Vbias 0.37318f
C15646 VDD.n6514 Vbias 0.01836f
C15647 VDD.n6515 Vbias 0.03639f
C15648 VDD.n6516 Vbias 0.37318f
C15649 VDD.n6517 Vbias 0.03639f
C15650 VDD.n6518 Vbias 0.03694f
C15651 VDD.n6519 Vbias 0.04583f
C15652 VDD.n6520 Vbias 0.03902f
C15653 VDD.n6521 Vbias 0.01836f
C15654 VDD.n6522 Vbias 0.03639f
C15655 VDD.n6523 Vbias 0.50118f
C15656 VDD.n6524 Vbias 0.50118f
C15657 VDD.n6525 Vbias 0.03639f
C15658 VDD.n6526 Vbias 0.01999f
C15659 VDD.n6527 Vbias 0.0216f
C15660 VDD.n6528 Vbias 0.01999f
C15661 VDD.n6529 Vbias 0.03639f
C15662 VDD.n6530 Vbias 0.50118f
C15663 VDD.n6531 Vbias 0.01836f
C15664 VDD.n6532 Vbias 0.03639f
C15665 VDD.n6533 Vbias 0.50118f
C15666 VDD.n6534 Vbias 0.03639f
C15667 VDD.n6535 Vbias 0.03694f
C15668 VDD.n6536 Vbias 0.04583f
C15669 VDD.n6537 Vbias 0.03902f
C15670 VDD.n6538 Vbias 0.01836f
C15671 VDD.n6539 Vbias 0.03639f
C15672 VDD.n6540 Vbias 0.37318f
C15673 VDD.n6541 Vbias 0.01836f
C15674 VDD.n6542 Vbias 0.03639f
C15675 VDD.n6543 Vbias 0.37318f
C15676 VDD.n6544 Vbias 0.03639f
C15677 VDD.n6545 Vbias 0.03694f
C15678 VDD.n6546 Vbias 0.04583f
C15679 VDD.n6547 Vbias 0.03902f
C15680 VDD.n6548 Vbias 0.01836f
C15681 VDD.n6549 Vbias 0.03639f
C15682 VDD.n6550 Vbias 0.50118f
C15683 VDD.n6551 Vbias 0.01836f
C15684 VDD.n6552 Vbias 0.03639f
C15685 VDD.n6553 Vbias 0.50118f
C15686 VDD.n6554 Vbias 0.03639f
C15687 VDD.n6555 Vbias 0.03694f
C15688 VDD.n6556 Vbias 0.04583f
C15689 VDD.n6557 Vbias 0.03902f
C15690 VDD.n6558 Vbias 0.01836f
C15691 VDD.n6559 Vbias 0.03639f
C15692 VDD.n6560 Vbias 0.37318f
C15693 VDD.n6561 Vbias 0.01836f
C15694 VDD.n6562 Vbias 0.03639f
C15695 VDD.n6563 Vbias 0.37318f
C15696 VDD.n6564 Vbias 0.03639f
C15697 VDD.n6565 Vbias 0.03694f
C15698 VDD.n6566 Vbias 0.04583f
C15699 VDD.n6567 Vbias 0.03902f
C15700 VDD.n6568 Vbias 0.01836f
C15701 VDD.n6569 Vbias 0.03639f
C15702 VDD.n6570 Vbias 0.37318f
C15703 VDD.n6571 Vbias 0.37318f
C15704 VDD.n6572 Vbias 0.03639f
C15705 VDD.n6573 Vbias 0.03639f
C15706 VDD.n6574 Vbias 0.01836f
C15707 VDD.n6575 Vbias 0.01836f
C15708 VDD.n6576 Vbias 0.0216f
C15709 VDD.n6577 Vbias 0.03694f
C15710 VDD.t151 Vbias 0.46278f
C15711 VDD.n6578 Vbias 0.03694f
C15712 VDD.n6579 Vbias 0.04583f
C15713 VDD.n6580 Vbias 0.074f
C15714 VDD.n6581 Vbias 0.05322f
C15715 VDD.n6582 Vbias 0.01309f
C15716 VDD.n6583 Vbias 0.06648f
C15717 VDD.n6584 Vbias 0.01999f
C15718 VDD.n6585 Vbias 0.03639f
C15719 VDD.n6586 Vbias 0.50118f
C15720 VDD.n6587 Vbias 0.01836f
C15721 VDD.n6588 Vbias 0.03639f
C15722 VDD.n6589 Vbias 0.50118f
C15723 VDD.n6590 Vbias 0.03639f
C15724 VDD.n6591 Vbias 0.03694f
C15725 VDD.n6592 Vbias 0.04583f
C15726 VDD.n6593 Vbias 0.03902f
C15727 VDD.n6594 Vbias 0.01836f
C15728 VDD.n6595 Vbias 0.03639f
C15729 VDD.n6596 Vbias 0.37318f
C15730 VDD.n6597 Vbias 0.01836f
C15731 VDD.n6598 Vbias 0.03639f
C15732 VDD.n6599 Vbias 0.37318f
C15733 VDD.n6600 Vbias 0.03639f
C15734 VDD.n6601 Vbias 0.03694f
C15735 VDD.n6602 Vbias 0.04583f
C15736 VDD.n6603 Vbias 0.03902f
C15737 VDD.n6604 Vbias 0.01836f
C15738 VDD.n6605 Vbias 0.03639f
C15739 VDD.n6606 Vbias 0.37318f
C15740 VDD.n6607 Vbias 0.01836f
C15741 VDD.n6608 Vbias 0.03639f
C15742 VDD.n6609 Vbias 0.37318f
C15743 VDD.n6610 Vbias 0.03639f
C15744 VDD.n6611 Vbias 0.03694f
C15745 VDD.n6612 Vbias 0.04583f
C15746 VDD.n6613 Vbias 0.03902f
C15747 VDD.n6614 Vbias 0.01836f
C15748 VDD.n6615 Vbias 0.03639f
C15749 VDD.n6616 Vbias 0.50118f
C15750 VDD.n6617 Vbias 0.01836f
C15751 VDD.n6618 Vbias 0.03639f
C15752 VDD.n6619 Vbias 0.50118f
C15753 VDD.n6620 Vbias 0.03639f
C15754 VDD.n6621 Vbias 0.03694f
C15755 VDD.n6622 Vbias 0.04583f
C15756 VDD.n6623 Vbias 0.03902f
C15757 VDD.n6624 Vbias 0.01836f
C15758 VDD.n6625 Vbias 0.03639f
C15759 VDD.n6626 Vbias 0.37318f
C15760 VDD.n6627 Vbias 0.01836f
C15761 VDD.n6628 Vbias 0.03639f
C15762 VDD.n6629 Vbias 0.37318f
C15763 VDD.n6630 Vbias 0.03639f
C15764 VDD.n6631 Vbias 0.03694f
C15765 VDD.n6632 Vbias 0.04583f
C15766 VDD.n6633 Vbias 0.03902f
C15767 VDD.n6634 Vbias 0.01836f
C15768 VDD.n6635 Vbias 0.03639f
C15769 VDD.n6636 Vbias 0.37318f
C15770 VDD.n6637 Vbias 0.01836f
C15771 VDD.n6638 Vbias 0.03639f
C15772 VDD.n6639 Vbias 0.37318f
C15773 VDD.n6640 Vbias 0.03639f
C15774 VDD.n6641 Vbias 0.03694f
C15775 VDD.n6642 Vbias 0.04583f
C15776 VDD.n6643 Vbias 0.03902f
C15777 VDD.n6644 Vbias 0.01836f
C15778 VDD.n6645 Vbias 0.03639f
C15779 VDD.n6646 Vbias 0.50118f
C15780 VDD.n6647 Vbias 0.50118f
C15781 VDD.n6648 Vbias 0.03639f
C15782 VDD.n6649 Vbias 0.01999f
C15783 VDD.n6650 Vbias 0.0216f
C15784 VDD.n6651 Vbias 0.01999f
C15785 VDD.n6652 Vbias 0.03639f
C15786 VDD.n6653 Vbias 0.50118f
C15787 VDD.n6654 Vbias 0.01836f
C15788 VDD.n6655 Vbias 0.03639f
C15789 VDD.n6656 Vbias 0.50118f
C15790 VDD.n6657 Vbias 0.03639f
C15791 VDD.n6658 Vbias 0.03694f
C15792 VDD.n6659 Vbias 0.04583f
C15793 VDD.n6660 Vbias 0.03902f
C15794 VDD.n6661 Vbias 0.01836f
C15795 VDD.n6662 Vbias 0.03639f
C15796 VDD.n6663 Vbias 0.37318f
C15797 VDD.n6664 Vbias 0.01836f
C15798 VDD.n6665 Vbias 0.03639f
C15799 VDD.n6666 Vbias 0.37318f
C15800 VDD.n6667 Vbias 0.03639f
C15801 VDD.n6668 Vbias 0.03694f
C15802 VDD.n6669 Vbias 0.04583f
C15803 VDD.n6670 Vbias 0.03902f
C15804 VDD.n6671 Vbias 0.01836f
C15805 VDD.n6672 Vbias 0.03639f
C15806 VDD.n6673 Vbias 0.50118f
C15807 VDD.n6674 Vbias 0.01836f
C15808 VDD.n6675 Vbias 0.03639f
C15809 VDD.n6676 Vbias 0.50118f
C15810 VDD.n6677 Vbias 0.03639f
C15811 VDD.n6678 Vbias 0.03694f
C15812 VDD.n6679 Vbias 0.04583f
C15813 VDD.n6680 Vbias 0.03902f
C15814 VDD.n6681 Vbias 0.01836f
C15815 VDD.n6682 Vbias 0.03639f
C15816 VDD.n6683 Vbias 0.37318f
C15817 VDD.n6684 Vbias 0.01836f
C15818 VDD.n6685 Vbias 0.03639f
C15819 VDD.n6686 Vbias 0.37318f
C15820 VDD.n6687 Vbias 0.03639f
C15821 VDD.n6688 Vbias 0.03694f
C15822 VDD.n6689 Vbias 0.04583f
C15823 VDD.n6690 Vbias 0.03902f
C15824 VDD.n6691 Vbias 0.01836f
C15825 VDD.n6692 Vbias 0.03639f
C15826 VDD.n6693 Vbias 0.37318f
C15827 VDD.n6694 Vbias 0.37318f
C15828 VDD.n6695 Vbias 0.03639f
C15829 VDD.n6696 Vbias 0.03639f
C15830 VDD.n6697 Vbias 0.01836f
C15831 VDD.n6698 Vbias 0.01836f
C15832 VDD.n6699 Vbias 0.0216f
C15833 VDD.n6700 Vbias 0.03694f
C15834 VDD.t862 Vbias 0.46278f
C15835 VDD.n6701 Vbias 0.03694f
C15836 VDD.n6702 Vbias 0.04583f
C15837 VDD.n6703 Vbias 0.074f
C15838 VDD.n6704 Vbias 0.05322f
C15839 VDD.n6705 Vbias 0.01309f
C15840 VDD.n6706 Vbias 0.06648f
C15841 VDD.n6707 Vbias 0.01999f
C15842 VDD.n6708 Vbias 0.03639f
C15843 VDD.n6709 Vbias 0.50118f
C15844 VDD.n6710 Vbias 0.01836f
C15845 VDD.n6711 Vbias 0.03639f
C15846 VDD.n6712 Vbias 0.50118f
C15847 VDD.n6713 Vbias 0.03639f
C15848 VDD.n6714 Vbias 0.03694f
C15849 VDD.n6715 Vbias 0.04583f
C15850 VDD.n6716 Vbias 0.03902f
C15851 VDD.n6717 Vbias 0.01836f
C15852 VDD.n6718 Vbias 0.03639f
C15853 VDD.n6719 Vbias 0.37318f
C15854 VDD.n6720 Vbias 0.01836f
C15855 VDD.n6721 Vbias 0.03639f
C15856 VDD.n6722 Vbias 0.37318f
C15857 VDD.n6723 Vbias 0.03639f
C15858 VDD.n6724 Vbias 0.03694f
C15859 VDD.n6725 Vbias 0.04583f
C15860 VDD.n6726 Vbias 0.03902f
C15861 VDD.n6727 Vbias 0.01836f
C15862 VDD.n6728 Vbias 0.03639f
C15863 VDD.n6729 Vbias 0.37318f
C15864 VDD.n6730 Vbias 0.01836f
C15865 VDD.n6731 Vbias 0.03639f
C15866 VDD.n6732 Vbias 0.37318f
C15867 VDD.n6733 Vbias 0.03639f
C15868 VDD.n6734 Vbias 0.03694f
C15869 VDD.n6735 Vbias 0.04583f
C15870 VDD.n6736 Vbias 0.03902f
C15871 VDD.n6737 Vbias 0.01836f
C15872 VDD.n6738 Vbias 0.03639f
C15873 VDD.n6739 Vbias 0.50118f
C15874 VDD.n6740 Vbias 0.01836f
C15875 VDD.n6741 Vbias 0.03639f
C15876 VDD.n6742 Vbias 0.50118f
C15877 VDD.n6743 Vbias 0.03639f
C15878 VDD.n6744 Vbias 0.03694f
C15879 VDD.n6745 Vbias 0.04583f
C15880 VDD.n6746 Vbias 0.03902f
C15881 VDD.n6747 Vbias 0.01836f
C15882 VDD.n6748 Vbias 0.03639f
C15883 VDD.n6749 Vbias 0.37318f
C15884 VDD.n6750 Vbias 0.01836f
C15885 VDD.n6751 Vbias 0.03639f
C15886 VDD.n6752 Vbias 0.37318f
C15887 VDD.n6753 Vbias 0.03639f
C15888 VDD.n6754 Vbias 0.03694f
C15889 VDD.n6755 Vbias 0.04583f
C15890 VDD.n6756 Vbias 0.03902f
C15891 VDD.n6757 Vbias 0.01836f
C15892 VDD.n6758 Vbias 0.03639f
C15893 VDD.n6759 Vbias 0.37318f
C15894 VDD.n6760 Vbias 0.01836f
C15895 VDD.n6761 Vbias 0.03639f
C15896 VDD.n6762 Vbias 0.37318f
C15897 VDD.n6763 Vbias 0.03639f
C15898 VDD.n6764 Vbias 0.03694f
C15899 VDD.n6765 Vbias 0.04583f
C15900 VDD.n6766 Vbias 0.03902f
C15901 VDD.n6767 Vbias 0.01836f
C15902 VDD.n6768 Vbias 0.03639f
C15903 VDD.n6769 Vbias 0.50118f
C15904 VDD.n6770 Vbias 0.50118f
C15905 VDD.n6771 Vbias 0.03639f
C15906 VDD.n6772 Vbias 0.01999f
C15907 VDD.n6773 Vbias 0.0216f
C15908 VDD.n6774 Vbias 0.01999f
C15909 VDD.n6775 Vbias 0.03639f
C15910 VDD.n6776 Vbias 0.50118f
C15911 VDD.n6777 Vbias 0.01836f
C15912 VDD.n6778 Vbias 0.03639f
C15913 VDD.n6779 Vbias 0.50118f
C15914 VDD.n6780 Vbias 0.03639f
C15915 VDD.n6781 Vbias 0.03694f
C15916 VDD.n6782 Vbias 0.04583f
C15917 VDD.n6783 Vbias 0.03902f
C15918 VDD.n6784 Vbias 0.01836f
C15919 VDD.n6785 Vbias 0.03639f
C15920 VDD.n6786 Vbias 0.37318f
C15921 VDD.n6787 Vbias 0.01836f
C15922 VDD.n6788 Vbias 0.03639f
C15923 VDD.n6789 Vbias 0.37318f
C15924 VDD.n6790 Vbias 0.03639f
C15925 VDD.n6791 Vbias 0.03694f
C15926 VDD.n6792 Vbias 0.04583f
C15927 VDD.n6793 Vbias 0.03902f
C15928 VDD.n6794 Vbias 0.01836f
C15929 VDD.n6795 Vbias 0.03639f
C15930 VDD.n6796 Vbias 0.50118f
C15931 VDD.n6797 Vbias 0.01836f
C15932 VDD.n6798 Vbias 0.03639f
C15933 VDD.n6799 Vbias 0.50118f
C15934 VDD.n6800 Vbias 0.03639f
C15935 VDD.n6801 Vbias 0.03694f
C15936 VDD.n6802 Vbias 0.04583f
C15937 VDD.n6803 Vbias 0.03902f
C15938 VDD.n6804 Vbias 0.01836f
C15939 VDD.n6805 Vbias 0.03639f
C15940 VDD.n6806 Vbias 0.37318f
C15941 VDD.n6807 Vbias 0.01836f
C15942 VDD.n6808 Vbias 0.03639f
C15943 VDD.n6809 Vbias 0.37318f
C15944 VDD.n6810 Vbias 0.03639f
C15945 VDD.n6811 Vbias 0.03694f
C15946 VDD.n6812 Vbias 0.04583f
C15947 VDD.n6813 Vbias 0.03902f
C15948 VDD.n6814 Vbias 0.01836f
C15949 VDD.n6815 Vbias 0.03639f
C15950 VDD.n6816 Vbias 0.37318f
C15951 VDD.n6817 Vbias 0.37318f
C15952 VDD.n6818 Vbias 0.03639f
C15953 VDD.n6819 Vbias 0.03639f
C15954 VDD.n6820 Vbias 0.01836f
C15955 VDD.n6821 Vbias 0.01836f
C15956 VDD.n6822 Vbias 0.0216f
C15957 VDD.n6823 Vbias 0.03694f
C15958 VDD.t937 Vbias 0.46278f
C15959 VDD.n6824 Vbias 0.03694f
C15960 VDD.n6825 Vbias 0.04583f
C15961 VDD.n6826 Vbias 0.05308f
C15962 VDD.n6827 Vbias 0.89624f
C15963 VDD.t410 Vbias 0.0169f
C15964 VDD.t1009 Vbias 0.0169f
C15965 VDD.n6829 Vbias 0.07902f
C15966 VDD.n6830 Vbias 0.0228f
C15967 VDD.n6831 Vbias 0.01999f
C15968 VDD.n6832 Vbias 0.01999f
C15969 VDD.n6833 Vbias 0.03639f
C15970 VDD.n6834 Vbias 0.03639f
C15971 VDD.t589 Vbias 0.24595f
C15972 VDD.n6835 Vbias 0.03694f
C15973 VDD.n6836 Vbias 0.03694f
C15974 VDD.t590 Vbias 0.017f
C15975 VDD.n6837 Vbias 0.07133f
C15976 VDD.n6838 Vbias 0.06984f
C15977 VDD.n6840 Vbias 0.26017f
C15978 VDD.n6841 Vbias 0.01999f
C15979 VDD.n6842 Vbias 0.0216f
C15980 VDD.n6843 Vbias 0.01999f
C15981 VDD.n6844 Vbias 0.03639f
C15982 VDD.n6845 Vbias 0.24422f
C15983 VDD.n6846 Vbias 0.24422f
C15984 VDD.t1008 Vbias 0.24595f
C15985 VDD.n6847 Vbias 0.03694f
C15986 VDD.n6848 Vbias 0.03694f
C15987 VDD.t368 Vbias 0.0169f
C15988 VDD.t871 Vbias 0.0169f
C15989 VDD.n6849 Vbias 0.07902f
C15990 VDD.n6850 Vbias 0.0228f
C15991 VDD.n6851 Vbias 0.01999f
C15992 VDD.n6852 Vbias 0.03694f
C15993 VDD.n6853 Vbias 0.0216f
C15994 VDD.n6854 Vbias 0.03694f
C15995 VDD.n6855 Vbias 0.26017f
C15996 VDD.t367 Vbias 0.24595f
C15997 VDD.t870 Vbias 0.24595f
C15998 VDD.n6857 Vbias 0.03694f
C15999 VDD.n6858 Vbias 0.03694f
C16000 VDD.t601 Vbias 0.017f
C16001 VDD.n6859 Vbias 0.05322f
C16002 VDD.n6860 Vbias 0.01999f
C16003 VDD.n6861 Vbias 0.03694f
C16004 VDD.n6862 Vbias 0.0216f
C16005 VDD.n6863 Vbias 0.03694f
C16006 VDD.n6864 Vbias 0.26017f
C16007 VDD.t600 Vbias 0.24595f
C16008 VDD.t958 Vbias 0.22551f
C16009 VDD.n6866 Vbias 0.03694f
C16010 VDD.n6867 Vbias 0.03694f
C16011 VDD.n6868 Vbias 0.06648f
C16012 VDD.t1040 Vbias 0.24595f
C16013 VDD.n6869 Vbias 0.03694f
C16014 VDD.n6870 Vbias 0.03694f
C16015 VDD.t959 Vbias 0.0169f
C16016 VDD.t1041 Vbias 0.0169f
C16017 VDD.n6871 Vbias 0.07902f
C16018 VDD.n6872 Vbias 0.01699f
C16019 VDD.n6873 Vbias 0.0228f
C16020 VDD.t583 Vbias 0.0169f
C16021 VDD.t906 Vbias 0.0169f
C16022 VDD.n6874 Vbias 0.07902f
C16023 VDD.n6875 Vbias 0.0228f
C16024 VDD.n6876 Vbias 0.01999f
C16025 VDD.n6877 Vbias 0.03694f
C16026 VDD.n6878 Vbias 0.0216f
C16027 VDD.n6879 Vbias 0.03694f
C16028 VDD.n6880 Vbias 0.26017f
C16029 VDD.t582 Vbias 0.24595f
C16030 VDD.t905 Vbias 0.24595f
C16031 VDD.n6882 Vbias 0.03694f
C16032 VDD.n6883 Vbias 0.03694f
C16033 VDD.t577 Vbias 0.017f
C16034 VDD.n6884 Vbias 0.05322f
C16035 VDD.n6885 Vbias 0.01999f
C16036 VDD.n6886 Vbias 0.03694f
C16037 VDD.n6887 Vbias 0.0216f
C16038 VDD.n6888 Vbias 0.03694f
C16039 VDD.n6889 Vbias 0.26017f
C16040 VDD.t576 Vbias 0.24595f
C16041 VDD.t620 Vbias 0.22551f
C16042 VDD.n6891 Vbias 0.03694f
C16043 VDD.n6892 Vbias 0.03694f
C16044 VDD.n6893 Vbias 0.06648f
C16045 VDD.t1012 Vbias 0.24595f
C16046 VDD.n6894 Vbias 0.03694f
C16047 VDD.n6895 Vbias 0.03694f
C16048 VDD.t621 Vbias 0.0169f
C16049 VDD.t1013 Vbias 0.0169f
C16050 VDD.n6896 Vbias 0.07902f
C16051 VDD.n6897 Vbias 0.01699f
C16052 VDD.n6898 Vbias 0.0228f
C16053 VDD.t358 Vbias 0.0169f
C16054 VDD.t879 Vbias 0.0169f
C16055 VDD.n6899 Vbias 0.07902f
C16056 VDD.n6900 Vbias 0.0228f
C16057 VDD.n6901 Vbias 0.01999f
C16058 VDD.n6902 Vbias 0.03694f
C16059 VDD.n6903 Vbias 0.0216f
C16060 VDD.n6904 Vbias 0.03694f
C16061 VDD.n6905 Vbias 0.26017f
C16062 VDD.t357 Vbias 0.24595f
C16063 VDD.t878 Vbias 0.24595f
C16064 VDD.n6907 Vbias 0.03694f
C16065 VDD.n6908 Vbias 0.03694f
C16066 VDD.t325 Vbias 0.017f
C16067 VDD.n6909 Vbias 0.05322f
C16068 VDD.n6910 Vbias 0.01999f
C16069 VDD.n6911 Vbias 0.03694f
C16070 VDD.n6912 Vbias 0.0216f
C16071 VDD.n6913 Vbias 0.03694f
C16072 VDD.n6914 Vbias 0.26017f
C16073 VDD.t324 Vbias 0.24595f
C16074 VDD.t339 Vbias 0.22551f
C16075 VDD.n6916 Vbias 0.03694f
C16076 VDD.n6917 Vbias 0.03694f
C16077 VDD.n6918 Vbias 0.06648f
C16078 VDD.t1036 Vbias 0.24595f
C16079 VDD.n6919 Vbias 0.03694f
C16080 VDD.n6920 Vbias 0.03694f
C16081 VDD.t340 Vbias 0.0169f
C16082 VDD.t1037 Vbias 0.0169f
C16083 VDD.n6921 Vbias 0.07902f
C16084 VDD.n6922 Vbias 0.01699f
C16085 VDD.n6923 Vbias 0.0228f
C16086 VDD.t330 Vbias 0.0169f
C16087 VDD.t695 Vbias 0.0169f
C16088 VDD.n6924 Vbias 0.07902f
C16089 VDD.n6925 Vbias 0.0228f
C16090 VDD.n6926 Vbias 0.01999f
C16091 VDD.n6927 Vbias 0.03694f
C16092 VDD.n6928 Vbias 0.0216f
C16093 VDD.n6929 Vbias 0.03694f
C16094 VDD.n6930 Vbias 0.26017f
C16095 VDD.t329 Vbias 0.24595f
C16096 VDD.t694 Vbias 0.24595f
C16097 VDD.n6932 Vbias 0.03694f
C16098 VDD.n6933 Vbias 0.03694f
C16099 VDD.n6934 Vbias 0.01699f
C16100 VDD.n6935 Vbias 0.06648f
C16101 VDD.n6937 Vbias 0.26017f
C16102 VDD.n6938 Vbias 0.01999f
C16103 VDD.n6939 Vbias 0.0216f
C16104 VDD.n6940 Vbias 0.01999f
C16105 VDD.n6941 Vbias 0.03639f
C16106 VDD.n6942 Vbias 0.18185f
C16107 VDD.n6943 Vbias 0.18185f
C16108 VDD.n6944 Vbias 0.03639f
C16109 VDD.n6945 Vbias 0.01999f
C16110 VDD.n6946 Vbias 0.06648f
C16111 VDD.n6947 Vbias 0.24997f
C16112 VDD.n6948 Vbias 0.01699f
C16113 VDD.n6949 Vbias 0.06648f
C16114 VDD.n6951 Vbias 0.26017f
C16115 VDD.n6952 Vbias 0.01999f
C16116 VDD.n6953 Vbias 0.0216f
C16117 VDD.n6954 Vbias 0.01999f
C16118 VDD.n6955 Vbias 0.03639f
C16119 VDD.n6956 Vbias 0.18185f
C16120 VDD.n6957 Vbias 0.18185f
C16121 VDD.n6958 Vbias 0.03639f
C16122 VDD.n6959 Vbias 0.01999f
C16123 VDD.n6960 Vbias 0.0216f
C16124 VDD.n6961 Vbias 0.01999f
C16125 VDD.n6962 Vbias 0.03639f
C16126 VDD.n6963 Vbias 0.24422f
C16127 VDD.n6964 Vbias 0.24422f
C16128 VDD.n6965 Vbias 0.03639f
C16129 VDD.n6966 Vbias 0.01999f
C16130 VDD.n6967 Vbias 0.06648f
C16131 VDD.n6968 Vbias 0.24606f
C16132 VDD.n6969 Vbias 0.01699f
C16133 VDD.n6970 Vbias 0.06648f
C16134 VDD.n6972 Vbias 0.26017f
C16135 VDD.n6973 Vbias 0.01999f
C16136 VDD.n6974 Vbias 0.0216f
C16137 VDD.n6975 Vbias 0.01999f
C16138 VDD.n6976 Vbias 0.03639f
C16139 VDD.n6977 Vbias 0.18185f
C16140 VDD.n6978 Vbias 0.18185f
C16141 VDD.n6979 Vbias 0.03639f
C16142 VDD.n6980 Vbias 0.01999f
C16143 VDD.n6981 Vbias 0.06648f
C16144 VDD.n6982 Vbias 0.24997f
C16145 VDD.n6983 Vbias 0.01699f
C16146 VDD.n6984 Vbias 0.06648f
C16147 VDD.n6986 Vbias 0.26017f
C16148 VDD.n6987 Vbias 0.01999f
C16149 VDD.n6988 Vbias 0.0216f
C16150 VDD.n6989 Vbias 0.01999f
C16151 VDD.n6990 Vbias 0.03639f
C16152 VDD.n6991 Vbias 0.18185f
C16153 VDD.n6992 Vbias 0.18185f
C16154 VDD.n6993 Vbias 0.03639f
C16155 VDD.n6994 Vbias 0.01999f
C16156 VDD.n6995 Vbias 0.0216f
C16157 VDD.n6996 Vbias 0.01999f
C16158 VDD.n6997 Vbias 0.03639f
C16159 VDD.n6998 Vbias 0.24422f
C16160 VDD.n6999 Vbias 0.24422f
C16161 VDD.n7000 Vbias 0.03639f
C16162 VDD.n7001 Vbias 0.01999f
C16163 VDD.n7002 Vbias 0.06648f
C16164 VDD.n7003 Vbias 0.24606f
C16165 VDD.n7004 Vbias 0.01699f
C16166 VDD.n7005 Vbias 0.06648f
C16167 VDD.n7007 Vbias 0.26017f
C16168 VDD.n7008 Vbias 0.01999f
C16169 VDD.n7009 Vbias 0.0216f
C16170 VDD.n7010 Vbias 0.01999f
C16171 VDD.n7011 Vbias 0.03639f
C16172 VDD.n7012 Vbias 0.18185f
C16173 VDD.n7013 Vbias 0.18185f
C16174 VDD.n7014 Vbias 0.03639f
C16175 VDD.n7015 Vbias 0.01999f
C16176 VDD.n7016 Vbias 0.06648f
C16177 VDD.n7017 Vbias 0.24997f
C16178 VDD.n7018 Vbias 0.01699f
C16179 VDD.n7019 Vbias 0.06648f
C16180 VDD.n7021 Vbias 0.26017f
C16181 VDD.n7022 Vbias 0.01999f
C16182 VDD.n7023 Vbias 0.0216f
C16183 VDD.n7024 Vbias 0.01999f
C16184 VDD.n7025 Vbias 0.03639f
C16185 VDD.n7026 Vbias 0.18185f
C16186 VDD.n7027 Vbias 0.18185f
C16187 VDD.n7028 Vbias 0.03639f
C16188 VDD.n7029 Vbias 0.01999f
C16189 VDD.n7030 Vbias 0.0216f
C16190 VDD.n7031 Vbias 0.01999f
C16191 VDD.n7032 Vbias 0.03639f
C16192 VDD.n7033 Vbias 0.24422f
C16193 VDD.n7034 Vbias 0.24422f
C16194 VDD.n7035 Vbias 0.03639f
C16195 VDD.n7036 Vbias 0.01999f
C16196 VDD.n7037 Vbias 0.06648f
C16197 VDD.n7038 Vbias 0.24606f
C16198 VDD.n7039 Vbias 0.01699f
C16199 VDD.n7040 Vbias 0.06648f
C16200 VDD.n7042 Vbias 0.26017f
C16201 VDD.n7043 Vbias 0.01999f
C16202 VDD.n7044 Vbias 0.0216f
C16203 VDD.n7045 Vbias 0.01999f
C16204 VDD.n7046 Vbias 0.03639f
C16205 VDD.n7047 Vbias 0.18185f
C16206 VDD.n7048 Vbias 0.18185f
C16207 VDD.n7049 Vbias 0.03639f
C16208 VDD.n7050 Vbias 0.01999f
C16209 VDD.n7051 Vbias 0.06648f
C16210 VDD.n7052 Vbias 0.24997f
C16211 VDD.n7053 Vbias 0.01699f
C16212 VDD.n7054 Vbias 0.06648f
C16213 VDD.n7056 Vbias 0.26017f
C16214 VDD.n7057 Vbias 0.01999f
C16215 VDD.n7058 Vbias 0.0216f
C16216 VDD.n7059 Vbias 0.01999f
C16217 VDD.n7060 Vbias 0.03639f
C16218 VDD.n7061 Vbias 0.18185f
C16219 VDD.n7062 Vbias 0.18185f
C16220 VDD.n7063 Vbias 0.0216f
C16221 VDD.n7064 Vbias 0.03694f
C16222 VDD.t409 Vbias 0.22551f
C16223 VDD.n7065 Vbias 0.03694f
C16224 VDD.n7066 Vbias 0.06648f
C16225 VDD.n7067 Vbias 0.01632f
C16226 VDD.n7068 Vbias 0.05591f
C16227 VDD.n7070 Vbias 1.55381f
C16228 VDD.n7071 Vbias 0.10375f
C16229 VDD.n7072 Vbias 0.01699f
C16230 VDD.n7073 Vbias 0.03902f
C16231 VDD.n7074 Vbias 0.03694f
C16232 VDD.n7075 Vbias 0.0216f
C16233 VDD.n7076 Vbias 0.01836f
C16234 VDD.n7077 Vbias 0.01836f
C16235 VDD.n7078 Vbias 0.03639f
C16236 VDD.n7079 Vbias 0.50118f
C16237 VDD.n7080 Vbias 0.03639f
C16238 VDD.n7081 Vbias 0.03694f
C16239 VDD.n7082 Vbias 0.04583f
C16240 VDD.n7083 Vbias 0.03902f
C16241 VDD.n7084 Vbias 0.01836f
C16242 VDD.n7085 Vbias 0.03639f
C16243 VDD.n7086 Vbias 0.37318f
C16244 VDD.n7087 Vbias 0.01836f
C16245 VDD.n7088 Vbias 0.03639f
C16246 VDD.n7089 Vbias 0.37318f
C16247 VDD.n7090 Vbias 0.03639f
C16248 VDD.n7091 Vbias 0.03694f
C16249 VDD.n7092 Vbias 0.04583f
C16250 VDD.n7093 Vbias 0.03902f
C16251 VDD.n7094 Vbias 0.01836f
C16252 VDD.n7095 Vbias 0.03639f
C16253 VDD.n7096 Vbias 0.37318f
C16254 VDD.n7097 Vbias 0.01836f
C16255 VDD.n7098 Vbias 0.03639f
C16256 VDD.n7099 Vbias 0.37318f
C16257 VDD.n7100 Vbias 0.03639f
C16258 VDD.n7101 Vbias 0.03694f
C16259 VDD.n7102 Vbias 0.04583f
C16260 VDD.n7103 Vbias 0.03902f
C16261 VDD.n7104 Vbias 0.01836f
C16262 VDD.n7105 Vbias 0.03639f
C16263 VDD.n7106 Vbias 0.50118f
C16264 VDD.n7107 Vbias 0.01836f
C16265 VDD.n7108 Vbias 0.03639f
C16266 VDD.n7109 Vbias 0.50118f
C16267 VDD.n7110 Vbias 0.03639f
C16268 VDD.n7111 Vbias 0.03694f
C16269 VDD.n7112 Vbias 0.04583f
C16270 VDD.n7113 Vbias 0.03902f
C16271 VDD.n7114 Vbias 0.01836f
C16272 VDD.n7115 Vbias 0.03639f
C16273 VDD.n7116 Vbias 0.37318f
C16274 VDD.n7117 Vbias 0.01836f
C16275 VDD.n7118 Vbias 0.03639f
C16276 VDD.n7119 Vbias 0.37318f
C16277 VDD.n7120 Vbias 0.03639f
C16278 VDD.n7121 Vbias 0.03694f
C16279 VDD.n7122 Vbias 0.04583f
C16280 VDD.n7123 Vbias 0.03902f
C16281 VDD.n7124 Vbias 0.01836f
C16282 VDD.n7125 Vbias 0.03639f
C16283 VDD.n7126 Vbias 0.50118f
C16284 VDD.n7127 Vbias 0.50118f
C16285 VDD.n7128 Vbias 0.03639f
C16286 VDD.n7129 Vbias 0.01999f
C16287 VDD.n7130 Vbias 0.0216f
C16288 VDD.n7131 Vbias 0.01999f
C16289 VDD.n7132 Vbias 0.03639f
C16290 VDD.n7133 Vbias 0.50118f
C16291 VDD.n7134 Vbias 0.50118f
C16292 VDD.n7135 Vbias 0.03639f
C16293 VDD.n7136 Vbias 0.03639f
C16294 VDD.n7137 Vbias 0.01836f
C16295 VDD.n7138 Vbias 0.01836f
C16296 VDD.n7139 Vbias 0.0216f
C16297 VDD.n7140 Vbias 0.03694f
C16298 VDD.t423 Vbias 0.46278f
C16299 VDD.n7141 Vbias 0.03694f
C16300 VDD.n7142 Vbias 0.04583f
C16301 VDD.n7143 Vbias 0.01699f
C16302 VDD.n7144 Vbias 0.03023f
C16303 VDD.n7145 Vbias 0.02225f
C16304 VDD.n7146 Vbias 0.04583f
C16305 VDD.n7147 Vbias 0.03902f
C16306 VDD.n7148 Vbias 0.01836f
C16307 VDD.n7149 Vbias 0.03639f
C16308 VDD.n7150 Vbias 0.37318f
C16309 VDD.n7151 Vbias 0.01836f
C16310 VDD.n7152 Vbias 0.03639f
C16311 VDD.n7153 Vbias 0.37318f
C16312 VDD.n7154 Vbias 0.03639f
C16313 VDD.n7155 Vbias 0.03694f
C16314 VDD.n7156 Vbias 0.04583f
C16315 VDD.n7157 Vbias 0.03902f
C16316 VDD.n7158 Vbias 0.01836f
C16317 VDD.n7159 Vbias 0.03639f
C16318 VDD.n7160 Vbias 0.50118f
C16319 VDD.n7161 Vbias 0.01836f
C16320 VDD.n7162 Vbias 0.03639f
C16321 VDD.n7163 Vbias 0.50118f
C16322 VDD.n7164 Vbias 0.03639f
C16323 VDD.n7165 Vbias 0.03694f
C16324 VDD.n7166 Vbias 0.04583f
C16325 VDD.n7167 Vbias 0.03902f
C16326 VDD.n7168 Vbias 0.01836f
C16327 VDD.n7169 Vbias 0.03639f
C16328 VDD.n7170 Vbias 0.37318f
C16329 VDD.n7171 Vbias 0.01836f
C16330 VDD.n7172 Vbias 0.03639f
C16331 VDD.n7173 Vbias 0.37318f
C16332 VDD.n7174 Vbias 0.03639f
C16333 VDD.n7175 Vbias 0.03694f
C16334 VDD.n7176 Vbias 0.04583f
C16335 VDD.n7177 Vbias 0.03902f
C16336 VDD.n7178 Vbias 0.01836f
C16337 VDD.n7179 Vbias 0.03639f
C16338 VDD.n7180 Vbias 0.37318f
C16339 VDD.n7181 Vbias 0.01836f
C16340 VDD.n7182 Vbias 0.03639f
C16341 VDD.n7183 Vbias 0.37318f
C16342 VDD.n7184 Vbias 0.03639f
C16343 VDD.n7185 Vbias 0.03694f
C16344 VDD.n7186 Vbias 0.04583f
C16345 VDD.n7187 Vbias 0.03902f
C16346 VDD.n7188 Vbias 0.01836f
C16347 VDD.n7189 Vbias 0.03639f
C16348 VDD.n7190 Vbias 0.50118f
C16349 VDD.n7191 Vbias 0.50118f
C16350 VDD.n7192 Vbias 0.03639f
C16351 VDD.n7193 Vbias 0.01999f
C16352 VDD.n7194 Vbias 0.06648f
C16353 VDD.n7195 Vbias 0.01309f
C16354 VDD.n7196 Vbias 0.05169f
C16355 VDD.n7197 Vbias 0.34538f
C16356 VDD.t851 Vbias 0.017f
C16357 VDD.n7198 Vbias 0.01999f
C16358 VDD.n7199 Vbias 0.03694f
C16359 VDD.n7200 Vbias 0.0216f
C16360 VDD.n7201 Vbias 0.03694f
C16361 VDD.n7202 Vbias 0.45845f
C16362 VDD.t850 Vbias 0.54191f
C16363 VDD.n7204 Vbias 0.03639f
C16364 VDD.t650 Vbias 0.46278f
C16365 VDD.n7205 Vbias 0.03694f
C16366 VDD.n7206 Vbias 0.03694f
C16367 VDD.n7207 Vbias 0.0216f
C16368 VDD.n7208 Vbias 0.01836f
C16369 VDD.t651 Vbias 0.017f
C16370 VDD.t1104 Vbias 0.017f
C16371 VDD.n7209 Vbias 0.09713f
C16372 VDD.n7210 Vbias 0.01914f
C16373 VDD.n7211 Vbias 0.03902f
C16374 VDD.n7212 Vbias 0.03694f
C16375 VDD.n7213 Vbias 0.0216f
C16376 VDD.n7214 Vbias 0.01836f
C16377 VDD.n7215 Vbias 0.03639f
C16378 VDD.t604 Vbias 0.46278f
C16379 VDD.n7216 Vbias 0.03694f
C16380 VDD.n7217 Vbias 0.03694f
C16381 VDD.n7218 Vbias 0.0216f
C16382 VDD.n7219 Vbias 0.01836f
C16383 VDD.n7220 Vbias 0.02305f
C16384 VDD.n7221 Vbias 0.03902f
C16385 VDD.n7222 Vbias 0.03694f
C16386 VDD.n7223 Vbias 0.0216f
C16387 VDD.n7224 Vbias 0.01836f
C16388 VDD.n7225 Vbias 0.03639f
C16389 VDD.t269 Vbias 0.46278f
C16390 VDD.n7226 Vbias 0.03694f
C16391 VDD.n7227 Vbias 0.03694f
C16392 VDD.n7228 Vbias 0.0216f
C16393 VDD.n7229 Vbias 0.01836f
C16394 VDD.t981 Vbias 0.0169f
C16395 VDD.t270 Vbias 0.0169f
C16396 VDD.n7230 Vbias 0.07902f
C16397 VDD.t605 Vbias 0.0169f
C16398 VDD.t273 Vbias 0.0169f
C16399 VDD.n7231 Vbias 0.07902f
C16400 VDD.n7232 Vbias 0.03023f
C16401 VDD.n7233 Vbias 0.01699f
C16402 VDD.n7234 Vbias 0.03902f
C16403 VDD.n7235 Vbias 0.03694f
C16404 VDD.n7236 Vbias 0.0216f
C16405 VDD.n7237 Vbias 0.01836f
C16406 VDD.n7238 Vbias 0.03639f
C16407 VDD.t985 Vbias 0.46278f
C16408 VDD.n7239 Vbias 0.03694f
C16409 VDD.n7240 Vbias 0.03694f
C16410 VDD.n7241 Vbias 0.0216f
C16411 VDD.n7242 Vbias 0.01836f
C16412 VDD.t1101 Vbias 0.017f
C16413 VDD.t986 Vbias 0.017f
C16414 VDD.n7243 Vbias 0.09713f
C16415 VDD.n7244 Vbias 0.01914f
C16416 VDD.n7245 Vbias 0.03902f
C16417 VDD.n7246 Vbias 0.03694f
C16418 VDD.n7247 Vbias 0.0216f
C16419 VDD.n7248 Vbias 0.01836f
C16420 VDD.n7249 Vbias 0.03639f
C16421 VDD.t309 Vbias 0.46278f
C16422 VDD.n7250 Vbias 0.03694f
C16423 VDD.n7251 Vbias 0.03694f
C16424 VDD.n7252 Vbias 0.0216f
C16425 VDD.n7253 Vbias 0.01836f
C16426 VDD.n7254 Vbias 0.02305f
C16427 VDD.n7255 Vbias 0.03902f
C16428 VDD.n7256 Vbias 0.03694f
C16429 VDD.n7257 Vbias 0.0216f
C16430 VDD.n7258 Vbias 0.01836f
C16431 VDD.n7259 Vbias 0.03639f
C16432 VDD.t873 Vbias 0.46278f
C16433 VDD.n7260 Vbias 0.03694f
C16434 VDD.n7261 Vbias 0.03694f
C16435 VDD.n7262 Vbias 0.0216f
C16436 VDD.n7263 Vbias 0.01836f
C16437 VDD.t669 Vbias 0.0169f
C16438 VDD.t874 Vbias 0.0169f
C16439 VDD.n7264 Vbias 0.07902f
C16440 VDD.t310 Vbias 0.0169f
C16441 VDD.t923 Vbias 0.0169f
C16442 VDD.n7265 Vbias 0.07902f
C16443 VDD.n7266 Vbias 0.03023f
C16444 VDD.n7267 Vbias 0.01699f
C16445 VDD.n7268 Vbias 0.03902f
C16446 VDD.n7269 Vbias 0.03694f
C16447 VDD.n7270 Vbias 0.0216f
C16448 VDD.n7271 Vbias 0.01836f
C16449 VDD.t271 Vbias 0.46278f
C16450 VDD.n7272 Vbias 0.03694f
C16451 VDD.n7273 Vbias 0.03694f
C16452 VDD.n7274 Vbias 0.06648f
C16453 VDD.n7275 Vbias 0.03639f
C16454 VDD.t375 Vbias 0.46278f
C16455 VDD.n7276 Vbias 0.03694f
C16456 VDD.n7277 Vbias 0.03694f
C16457 VDD.n7278 Vbias 0.0216f
C16458 VDD.n7279 Vbias 0.01836f
C16459 VDD.t272 Vbias 0.017f
C16460 VDD.n7280 Vbias 0.05322f
C16461 VDD.n7281 Vbias 0.01309f
C16462 VDD.n7282 Vbias 0.01699f
C16463 VDD.n7283 Vbias 0.03902f
C16464 VDD.n7284 Vbias 0.03694f
C16465 VDD.n7285 Vbias 0.0216f
C16466 VDD.n7286 Vbias 0.01836f
C16467 VDD.n7287 Vbias 0.03639f
C16468 VDD.t258 Vbias 0.46278f
C16469 VDD.n7288 Vbias 0.03694f
C16470 VDD.n7289 Vbias 0.03694f
C16471 VDD.n7290 Vbias 0.0216f
C16472 VDD.n7291 Vbias 0.01836f
C16473 VDD.t922 Vbias 0.0169f
C16474 VDD.t260 Vbias 0.0169f
C16475 VDD.n7292 Vbias 0.07902f
C16476 VDD.t376 Vbias 0.0169f
C16477 VDD.t259 Vbias 0.0169f
C16478 VDD.n7293 Vbias 0.07902f
C16479 VDD.n7294 Vbias 0.03023f
C16480 VDD.n7295 Vbias 0.01699f
C16481 VDD.n7296 Vbias 0.03902f
C16482 VDD.n7297 Vbias 0.03694f
C16483 VDD.n7298 Vbias 0.0216f
C16484 VDD.n7299 Vbias 0.01836f
C16485 VDD.n7300 Vbias 0.03639f
C16486 VDD.t331 Vbias 0.46278f
C16487 VDD.n7301 Vbias 0.03694f
C16488 VDD.n7302 Vbias 0.03694f
C16489 VDD.n7303 Vbias 0.0216f
C16490 VDD.n7304 Vbias 0.01836f
C16491 VDD.t332 Vbias 0.017f
C16492 VDD.t431 Vbias 0.017f
C16493 VDD.n7305 Vbias 0.09713f
C16494 VDD.n7306 Vbias 0.01914f
C16495 VDD.n7307 Vbias 0.03902f
C16496 VDD.n7308 Vbias 0.03694f
C16497 VDD.n7309 Vbias 0.0216f
C16498 VDD.n7310 Vbias 0.01836f
C16499 VDD.n7311 Vbias 0.03639f
C16500 VDD.t472 Vbias 0.46278f
C16501 VDD.n7312 Vbias 0.03694f
C16502 VDD.n7313 Vbias 0.03694f
C16503 VDD.n7314 Vbias 0.0216f
C16504 VDD.n7315 Vbias 0.01836f
C16505 VDD.n7316 Vbias 0.02305f
C16506 VDD.n7317 Vbias 0.03902f
C16507 VDD.n7318 Vbias 0.03694f
C16508 VDD.n7319 Vbias 0.0216f
C16509 VDD.n7320 Vbias 0.01836f
C16510 VDD.n7321 Vbias 0.03639f
C16511 VDD.t498 Vbias 0.46278f
C16512 VDD.n7322 Vbias 0.03694f
C16513 VDD.n7323 Vbias 0.03694f
C16514 VDD.n7324 Vbias 0.0216f
C16515 VDD.n7325 Vbias 0.01836f
C16516 VDD.t473 Vbias 0.0169f
C16517 VDD.t928 Vbias 0.0169f
C16518 VDD.n7326 Vbias 0.07902f
C16519 VDD.t489 Vbias 0.0169f
C16520 VDD.t499 Vbias 0.0169f
C16521 VDD.n7327 Vbias 0.07902f
C16522 VDD.n7328 Vbias 0.03023f
C16523 VDD.n7329 Vbias 0.01699f
C16524 VDD.n7330 Vbias 0.03902f
C16525 VDD.n7331 Vbias 0.03694f
C16526 VDD.n7332 Vbias 0.0216f
C16527 VDD.n7333 Vbias 0.01836f
C16528 VDD.n7334 Vbias 0.01836f
C16529 VDD.n7335 Vbias 0.03639f
C16530 VDD.n7336 Vbias 0.50118f
C16531 VDD.n7337 Vbias 0.03639f
C16532 VDD.n7338 Vbias 0.03694f
C16533 VDD.n7339 Vbias 0.04583f
C16534 VDD.n7340 Vbias 0.03902f
C16535 VDD.n7341 Vbias 0.01836f
C16536 VDD.n7342 Vbias 0.03639f
C16537 VDD.n7343 Vbias 0.37318f
C16538 VDD.n7344 Vbias 0.01836f
C16539 VDD.n7345 Vbias 0.03639f
C16540 VDD.n7346 Vbias 0.37318f
C16541 VDD.n7347 Vbias 0.03639f
C16542 VDD.n7348 Vbias 0.03694f
C16543 VDD.n7349 Vbias 0.04583f
C16544 VDD.n7350 Vbias 0.03902f
C16545 VDD.n7351 Vbias 0.01836f
C16546 VDD.n7352 Vbias 0.03639f
C16547 VDD.n7353 Vbias 0.37318f
C16548 VDD.n7354 Vbias 0.01836f
C16549 VDD.n7355 Vbias 0.03639f
C16550 VDD.n7356 Vbias 0.37318f
C16551 VDD.n7357 Vbias 0.03639f
C16552 VDD.n7358 Vbias 0.03694f
C16553 VDD.n7359 Vbias 0.04583f
C16554 VDD.n7360 Vbias 0.03902f
C16555 VDD.n7361 Vbias 0.01836f
C16556 VDD.n7362 Vbias 0.03639f
C16557 VDD.n7363 Vbias 0.50118f
C16558 VDD.n7364 Vbias 0.01836f
C16559 VDD.n7365 Vbias 0.03639f
C16560 VDD.n7366 Vbias 0.50118f
C16561 VDD.n7367 Vbias 0.03639f
C16562 VDD.n7368 Vbias 0.03694f
C16563 VDD.n7369 Vbias 0.04583f
C16564 VDD.n7370 Vbias 0.03902f
C16565 VDD.n7371 Vbias 0.01836f
C16566 VDD.n7372 Vbias 0.03639f
C16567 VDD.n7373 Vbias 0.37318f
C16568 VDD.n7374 Vbias 0.01836f
C16569 VDD.n7375 Vbias 0.03639f
C16570 VDD.n7376 Vbias 0.37318f
C16571 VDD.n7377 Vbias 0.03639f
C16572 VDD.n7378 Vbias 0.03694f
C16573 VDD.n7379 Vbias 0.04583f
C16574 VDD.n7380 Vbias 0.03902f
C16575 VDD.n7381 Vbias 0.01836f
C16576 VDD.n7382 Vbias 0.03639f
C16577 VDD.n7383 Vbias 0.50118f
C16578 VDD.n7384 Vbias 0.50118f
C16579 VDD.n7385 Vbias 0.03639f
C16580 VDD.n7386 Vbias 0.01999f
C16581 VDD.n7387 Vbias 0.0216f
C16582 VDD.n7388 Vbias 0.01999f
C16583 VDD.n7389 Vbias 0.03639f
C16584 VDD.n7390 Vbias 0.50118f
C16585 VDD.n7391 Vbias 0.01836f
C16586 VDD.n7392 Vbias 0.03639f
C16587 VDD.n7393 Vbias 0.50118f
C16588 VDD.n7394 Vbias 0.03639f
C16589 VDD.n7395 Vbias 0.03694f
C16590 VDD.n7396 Vbias 0.04583f
C16591 VDD.n7397 Vbias 0.03902f
C16592 VDD.n7398 Vbias 0.01836f
C16593 VDD.n7399 Vbias 0.03639f
C16594 VDD.n7400 Vbias 0.37318f
C16595 VDD.n7401 Vbias 0.01836f
C16596 VDD.n7402 Vbias 0.03639f
C16597 VDD.n7403 Vbias 0.37318f
C16598 VDD.n7404 Vbias 0.03639f
C16599 VDD.n7405 Vbias 0.03694f
C16600 VDD.n7406 Vbias 0.04583f
C16601 VDD.n7407 Vbias 0.03902f
C16602 VDD.n7408 Vbias 0.01836f
C16603 VDD.n7409 Vbias 0.03639f
C16604 VDD.n7410 Vbias 0.37318f
C16605 VDD.n7411 Vbias 0.01836f
C16606 VDD.n7412 Vbias 0.03639f
C16607 VDD.n7413 Vbias 0.37318f
C16608 VDD.n7414 Vbias 0.03639f
C16609 VDD.n7415 Vbias 0.03694f
C16610 VDD.n7416 Vbias 0.04583f
C16611 VDD.n7417 Vbias 0.03902f
C16612 VDD.n7418 Vbias 0.01836f
C16613 VDD.n7419 Vbias 0.03639f
C16614 VDD.n7420 Vbias 0.50118f
C16615 VDD.n7421 Vbias 0.01836f
C16616 VDD.n7422 Vbias 0.03639f
C16617 VDD.n7423 Vbias 0.50118f
C16618 VDD.n7424 Vbias 0.03639f
C16619 VDD.n7425 Vbias 0.03694f
C16620 VDD.n7426 Vbias 0.04583f
C16621 VDD.n7427 Vbias 0.03902f
C16622 VDD.n7428 Vbias 0.01836f
C16623 VDD.n7429 Vbias 0.03639f
C16624 VDD.n7430 Vbias 0.37318f
C16625 VDD.n7431 Vbias 0.01836f
C16626 VDD.n7432 Vbias 0.03639f
C16627 VDD.n7433 Vbias 0.37318f
C16628 VDD.n7434 Vbias 0.03639f
C16629 VDD.n7435 Vbias 0.03694f
C16630 VDD.n7436 Vbias 0.04583f
C16631 VDD.n7437 Vbias 0.03902f
C16632 VDD.n7438 Vbias 0.01836f
C16633 VDD.n7439 Vbias 0.03639f
C16634 VDD.n7440 Vbias 0.37318f
C16635 VDD.n7441 Vbias 0.01836f
C16636 VDD.n7442 Vbias 0.03639f
C16637 VDD.n7443 Vbias 0.37318f
C16638 VDD.n7444 Vbias 0.03639f
C16639 VDD.n7445 Vbias 0.03694f
C16640 VDD.n7446 Vbias 0.04583f
C16641 VDD.n7447 Vbias 0.03902f
C16642 VDD.n7448 Vbias 0.01836f
C16643 VDD.n7449 Vbias 0.03639f
C16644 VDD.n7450 Vbias 0.50118f
C16645 VDD.n7451 Vbias 0.50118f
C16646 VDD.n7452 Vbias 0.03639f
C16647 VDD.n7453 Vbias 0.01999f
C16648 VDD.n7454 Vbias 0.06648f
C16649 VDD.n7455 Vbias 0.01309f
C16650 VDD.n7456 Vbias 0.07184f
C16651 VDD.n7457 Vbias 0.65261f
C16652 VDD.n7458 Vbias 0.23842f
C16653 VDD.n7459 Vbias 0.07184f
C16654 VDD.n7460 Vbias 0.01309f
C16655 VDD.t397 Vbias 0.017f
C16656 VDD.t521 Vbias 0.017f
C16657 VDD.n7461 Vbias 0.02305f
C16658 VDD.n7462 Vbias 0.03902f
C16659 VDD.n7463 Vbias 0.03694f
C16660 VDD.n7464 Vbias 0.03902f
C16661 VDD.n7465 Vbias 0.03639f
C16662 VDD.n7466 Vbias 0.03639f
C16663 VDD.t943 Vbias 0.54191f
C16664 VDD.n7467 Vbias 0.03694f
C16665 VDD.n7468 Vbias 0.03694f
C16666 VDD.n7469 Vbias 0.0216f
C16667 VDD.n7471 Vbias 0.45845f
C16668 VDD.n7472 Vbias 0.01999f
C16669 VDD.n7473 Vbias 0.06648f
C16670 VDD.n7474 Vbias 0.01999f
C16671 VDD.n7475 Vbias 0.03639f
C16672 VDD.n7476 Vbias 0.50118f
C16673 VDD.n7477 Vbias 0.50118f
C16674 VDD.n7478 Vbias 0.01836f
C16675 VDD.n7479 Vbias 0.01836f
C16676 VDD.n7480 Vbias 0.0216f
C16677 VDD.n7481 Vbias 0.03694f
C16678 VDD.n7482 Vbias 0.03639f
C16679 VDD.t846 Vbias 0.46278f
C16680 VDD.n7483 Vbias 0.03694f
C16681 VDD.n7484 Vbias 0.03694f
C16682 VDD.n7485 Vbias 0.0216f
C16683 VDD.n7486 Vbias 0.01836f
C16684 VDD.n7487 Vbias 0.03902f
C16685 VDD.n7488 Vbias 0.03694f
C16686 VDD.n7489 Vbias 0.0216f
C16687 VDD.n7490 Vbias 0.01836f
C16688 VDD.n7491 Vbias 0.03639f
C16689 VDD.t146 Vbias 0.46278f
C16690 VDD.n7492 Vbias 0.03694f
C16691 VDD.n7493 Vbias 0.03694f
C16692 VDD.n7494 Vbias 0.0216f
C16693 VDD.n7495 Vbias 0.01836f
C16694 VDD.t847 Vbias 0.0169f
C16695 VDD.t147 Vbias 0.0169f
C16696 VDD.n7496 Vbias 0.07902f
C16697 VDD.t866 Vbias 0.0169f
C16698 VDD.t150 Vbias 0.0169f
C16699 VDD.n7497 Vbias 0.07902f
C16700 VDD.n7498 Vbias 0.03023f
C16701 VDD.n7499 Vbias 0.01699f
C16702 VDD.n7500 Vbias 0.03902f
C16703 VDD.n7501 Vbias 0.03694f
C16704 VDD.n7502 Vbias 0.0216f
C16705 VDD.n7503 Vbias 0.01836f
C16706 VDD.n7504 Vbias 0.03639f
C16707 VDD.t470 Vbias 0.46278f
C16708 VDD.n7505 Vbias 0.03694f
C16709 VDD.n7506 Vbias 0.03694f
C16710 VDD.n7507 Vbias 0.0216f
C16711 VDD.n7508 Vbias 0.01836f
C16712 VDD.t520 Vbias 0.017f
C16713 VDD.t471 Vbias 0.017f
C16714 VDD.n7509 Vbias 0.09713f
C16715 VDD.n7510 Vbias 0.01914f
C16716 VDD.n7511 Vbias 0.03902f
C16717 VDD.n7512 Vbias 0.03694f
C16718 VDD.n7513 Vbias 0.0216f
C16719 VDD.n7514 Vbias 0.01836f
C16720 VDD.n7515 Vbias 0.03639f
C16721 VDD.t712 Vbias 0.46278f
C16722 VDD.n7516 Vbias 0.03694f
C16723 VDD.n7517 Vbias 0.03694f
C16724 VDD.n7518 Vbias 0.0216f
C16725 VDD.n7519 Vbias 0.01836f
C16726 VDD.n7520 Vbias 0.02305f
C16727 VDD.n7521 Vbias 0.03902f
C16728 VDD.n7522 Vbias 0.03694f
C16729 VDD.n7523 Vbias 0.0216f
C16730 VDD.n7524 Vbias 0.01836f
C16731 VDD.n7525 Vbias 0.03639f
C16732 VDD.t553 Vbias 0.46278f
C16733 VDD.n7526 Vbias 0.03694f
C16734 VDD.n7527 Vbias 0.03694f
C16735 VDD.n7528 Vbias 0.0216f
C16736 VDD.n7529 Vbias 0.01836f
C16737 VDD.t900 Vbias 0.0169f
C16738 VDD.t554 Vbias 0.0169f
C16739 VDD.n7530 Vbias 0.07902f
C16740 VDD.t713 Vbias 0.0169f
C16741 VDD.t950 Vbias 0.0169f
C16742 VDD.n7531 Vbias 0.07902f
C16743 VDD.n7532 Vbias 0.03023f
C16744 VDD.n7533 Vbias 0.01699f
C16745 VDD.n7534 Vbias 0.03902f
C16746 VDD.n7535 Vbias 0.03694f
C16747 VDD.n7536 Vbias 0.0216f
C16748 VDD.n7537 Vbias 0.01836f
C16749 VDD.t148 Vbias 0.46278f
C16750 VDD.n7538 Vbias 0.03694f
C16751 VDD.n7539 Vbias 0.03694f
C16752 VDD.n7540 Vbias 0.06648f
C16753 VDD.n7541 Vbias 0.03639f
C16754 VDD.t555 Vbias 0.46278f
C16755 VDD.n7542 Vbias 0.03694f
C16756 VDD.n7543 Vbias 0.03694f
C16757 VDD.n7544 Vbias 0.0216f
C16758 VDD.n7545 Vbias 0.01836f
C16759 VDD.t149 Vbias 0.017f
C16760 VDD.n7546 Vbias 0.05322f
C16761 VDD.n7547 Vbias 0.01309f
C16762 VDD.n7548 Vbias 0.01699f
C16763 VDD.n7549 Vbias 0.03902f
C16764 VDD.n7550 Vbias 0.03694f
C16765 VDD.n7551 Vbias 0.0216f
C16766 VDD.n7552 Vbias 0.01836f
C16767 VDD.n7553 Vbias 0.03639f
C16768 VDD.t890 Vbias 0.46278f
C16769 VDD.n7554 Vbias 0.03694f
C16770 VDD.n7555 Vbias 0.03694f
C16771 VDD.n7556 Vbias 0.0216f
C16772 VDD.n7557 Vbias 0.01836f
C16773 VDD.t949 Vbias 0.0169f
C16774 VDD.t891 Vbias 0.0169f
C16775 VDD.n7558 Vbias 0.07902f
C16776 VDD.t556 Vbias 0.0169f
C16777 VDD.t892 Vbias 0.0169f
C16778 VDD.n7559 Vbias 0.07902f
C16779 VDD.n7560 Vbias 0.03023f
C16780 VDD.n7561 Vbias 0.01699f
C16781 VDD.n7562 Vbias 0.03902f
C16782 VDD.n7563 Vbias 0.03694f
C16783 VDD.n7564 Vbias 0.0216f
C16784 VDD.n7565 Vbias 0.01836f
C16785 VDD.n7566 Vbias 0.03639f
C16786 VDD.t194 Vbias 0.46278f
C16787 VDD.n7567 Vbias 0.03694f
C16788 VDD.n7568 Vbias 0.03694f
C16789 VDD.n7569 Vbias 0.0216f
C16790 VDD.n7570 Vbias 0.01836f
C16791 VDD.t359 Vbias 0.017f
C16792 VDD.t195 Vbias 0.017f
C16793 VDD.n7571 Vbias 0.09713f
C16794 VDD.n7572 Vbias 0.01914f
C16795 VDD.n7573 Vbias 0.03902f
C16796 VDD.n7574 Vbias 0.03694f
C16797 VDD.n7575 Vbias 0.0216f
C16798 VDD.n7576 Vbias 0.01836f
C16799 VDD.n7577 Vbias 0.03639f
C16800 VDD.t662 Vbias 0.46278f
C16801 VDD.n7578 Vbias 0.03694f
C16802 VDD.n7579 Vbias 0.03694f
C16803 VDD.n7580 Vbias 0.0216f
C16804 VDD.n7581 Vbias 0.01836f
C16805 VDD.n7582 Vbias 0.02305f
C16806 VDD.n7583 Vbias 0.03902f
C16807 VDD.n7584 Vbias 0.03694f
C16808 VDD.n7585 Vbias 0.0216f
C16809 VDD.n7586 Vbias 0.01836f
C16810 VDD.n7587 Vbias 0.03639f
C16811 VDD.t157 Vbias 0.46278f
C16812 VDD.n7588 Vbias 0.03694f
C16813 VDD.n7589 Vbias 0.03694f
C16814 VDD.n7590 Vbias 0.0216f
C16815 VDD.n7591 Vbias 0.01836f
C16816 VDD.t663 Vbias 0.0169f
C16817 VDD.t915 Vbias 0.0169f
C16818 VDD.n7592 Vbias 0.07902f
C16819 VDD.t893 Vbias 0.0169f
C16820 VDD.t158 Vbias 0.0169f
C16821 VDD.n7593 Vbias 0.07902f
C16822 VDD.n7594 Vbias 0.03023f
C16823 VDD.n7595 Vbias 0.01699f
C16824 VDD.n7596 Vbias 0.03902f
C16825 VDD.n7597 Vbias 0.03694f
C16826 VDD.n7598 Vbias 0.0216f
C16827 VDD.n7599 Vbias 0.01836f
C16828 VDD.n7600 Vbias 0.01836f
C16829 VDD.n7601 Vbias 0.03639f
C16830 VDD.n7602 Vbias 0.50118f
C16831 VDD.n7603 Vbias 0.03639f
C16832 VDD.n7604 Vbias 0.03694f
C16833 VDD.n7605 Vbias 0.04583f
C16834 VDD.n7606 Vbias 0.03902f
C16835 VDD.n7607 Vbias 0.01836f
C16836 VDD.n7608 Vbias 0.03639f
C16837 VDD.n7609 Vbias 0.37318f
C16838 VDD.n7610 Vbias 0.01836f
C16839 VDD.n7611 Vbias 0.03639f
C16840 VDD.n7612 Vbias 0.37318f
C16841 VDD.n7613 Vbias 0.03639f
C16842 VDD.n7614 Vbias 0.03694f
C16843 VDD.n7615 Vbias 0.04583f
C16844 VDD.n7616 Vbias 0.03902f
C16845 VDD.n7617 Vbias 0.01836f
C16846 VDD.n7618 Vbias 0.03639f
C16847 VDD.n7619 Vbias 0.37318f
C16848 VDD.n7620 Vbias 0.01836f
C16849 VDD.n7621 Vbias 0.03639f
C16850 VDD.n7622 Vbias 0.37318f
C16851 VDD.n7623 Vbias 0.03639f
C16852 VDD.n7624 Vbias 0.03694f
C16853 VDD.n7625 Vbias 0.04583f
C16854 VDD.n7626 Vbias 0.03902f
C16855 VDD.n7627 Vbias 0.01836f
C16856 VDD.n7628 Vbias 0.03639f
C16857 VDD.n7629 Vbias 0.50118f
C16858 VDD.n7630 Vbias 0.01836f
C16859 VDD.n7631 Vbias 0.03639f
C16860 VDD.n7632 Vbias 0.50118f
C16861 VDD.n7633 Vbias 0.03639f
C16862 VDD.n7634 Vbias 0.03694f
C16863 VDD.n7635 Vbias 0.04583f
C16864 VDD.n7636 Vbias 0.03902f
C16865 VDD.n7637 Vbias 0.01836f
C16866 VDD.n7638 Vbias 0.03639f
C16867 VDD.n7639 Vbias 0.37318f
C16868 VDD.n7640 Vbias 0.01836f
C16869 VDD.n7641 Vbias 0.03639f
C16870 VDD.n7642 Vbias 0.37318f
C16871 VDD.n7643 Vbias 0.03639f
C16872 VDD.n7644 Vbias 0.03694f
C16873 VDD.n7645 Vbias 0.04583f
C16874 VDD.n7646 Vbias 0.03902f
C16875 VDD.n7647 Vbias 0.01836f
C16876 VDD.n7648 Vbias 0.03639f
C16877 VDD.n7649 Vbias 0.50118f
C16878 VDD.n7650 Vbias 0.50118f
C16879 VDD.n7651 Vbias 0.03639f
C16880 VDD.n7652 Vbias 0.01999f
C16881 VDD.n7653 Vbias 0.0216f
C16882 VDD.n7654 Vbias 0.01999f
C16883 VDD.n7655 Vbias 0.03639f
C16884 VDD.n7656 Vbias 0.50118f
C16885 VDD.n7657 Vbias 0.01836f
C16886 VDD.n7658 Vbias 0.03639f
C16887 VDD.n7659 Vbias 0.50118f
C16888 VDD.n7660 Vbias 0.03639f
C16889 VDD.n7661 Vbias 0.03694f
C16890 VDD.n7662 Vbias 0.04583f
C16891 VDD.n7663 Vbias 0.03902f
C16892 VDD.n7664 Vbias 0.01836f
C16893 VDD.n7665 Vbias 0.03639f
C16894 VDD.n7666 Vbias 0.37318f
C16895 VDD.n7667 Vbias 0.01836f
C16896 VDD.n7668 Vbias 0.03639f
C16897 VDD.n7669 Vbias 0.37318f
C16898 VDD.n7670 Vbias 0.03639f
C16899 VDD.n7671 Vbias 0.03694f
C16900 VDD.n7672 Vbias 0.04583f
C16901 VDD.n7673 Vbias 0.03902f
C16902 VDD.n7674 Vbias 0.01836f
C16903 VDD.n7675 Vbias 0.03639f
C16904 VDD.n7676 Vbias 0.37318f
C16905 VDD.n7677 Vbias 0.01836f
C16906 VDD.n7678 Vbias 0.03639f
C16907 VDD.n7679 Vbias 0.37318f
C16908 VDD.n7680 Vbias 0.03639f
C16909 VDD.n7681 Vbias 0.03694f
C16910 VDD.n7682 Vbias 0.04583f
C16911 VDD.n7683 Vbias 0.03902f
C16912 VDD.n7684 Vbias 0.01836f
C16913 VDD.n7685 Vbias 0.03639f
C16914 VDD.n7686 Vbias 0.50118f
C16915 VDD.n7687 Vbias 0.01836f
C16916 VDD.n7688 Vbias 0.03639f
C16917 VDD.n7689 Vbias 0.50118f
C16918 VDD.n7690 Vbias 0.03639f
C16919 VDD.n7691 Vbias 0.03694f
C16920 VDD.n7692 Vbias 0.04583f
C16921 VDD.n7693 Vbias 0.03902f
C16922 VDD.n7694 Vbias 0.01836f
C16923 VDD.n7695 Vbias 0.03639f
C16924 VDD.n7696 Vbias 0.37318f
C16925 VDD.n7697 Vbias 0.01836f
C16926 VDD.n7698 Vbias 0.03639f
C16927 VDD.n7699 Vbias 0.37318f
C16928 VDD.n7700 Vbias 0.03639f
C16929 VDD.n7701 Vbias 0.03694f
C16930 VDD.n7702 Vbias 0.04583f
C16931 VDD.n7703 Vbias 0.03902f
C16932 VDD.n7704 Vbias 0.01836f
C16933 VDD.n7705 Vbias 0.03639f
C16934 VDD.n7706 Vbias 0.37318f
C16935 VDD.n7707 Vbias 0.37318f
C16936 VDD.n7708 Vbias 0.03639f
C16937 VDD.n7709 Vbias 0.03639f
C16938 VDD.n7710 Vbias 0.01836f
C16939 VDD.n7711 Vbias 0.01836f
C16940 VDD.n7712 Vbias 0.0216f
C16941 VDD.n7713 Vbias 0.03694f
C16942 VDD.t396 Vbias 0.46278f
C16943 VDD.n7714 Vbias 0.03694f
C16944 VDD.n7715 Vbias 0.04583f
C16945 VDD.n7716 Vbias 0.01914f
C16946 VDD.n7717 Vbias 0.09713f
C16947 Nand_Gate_4.A.t10 Vbias 0.27993f
C16948 Nand_Gate_4.A.n0 Vbias 0.08177f
C16949 Nand_Gate_4.A.n1 Vbias 0.03548f
C16950 Nand_Gate_4.A.n2 Vbias 0.15601f
C16951 Nand_Gate_4.A.t4 Vbias 0.1302f
C16952 Nand_Gate_4.A.n3 Vbias 0.04085f
C16953 Nand_Gate_4.A.t1 Vbias 0.03651f
C16954 Nand_Gate_4.A.n4 Vbias 0.159f
C16955 Nand_Gate_4.A.n5 Vbias 0.03942f
C16956 Nand_Gate_4.A.t5 Vbias 0.27994f
C16957 Nand_Gate_4.A.n6 Vbias 0.27511f
C16958 Nand_Gate_4.A.n7 Vbias 0.03007f
C16959 Nand_Gate_4.A.t11 Vbias 0.14554f
C16960 Nand_Gate_4.A.n8 Vbias 0.04192f
C16961 Nand_Gate_4.A.n9 Vbias 0.01797f
C16962 Nand_Gate_4.A.n10 Vbias 0.03367f
C16963 Nand_Gate_4.A.n11 Vbias 0.04236f
C16964 Nand_Gate_4.A.t9 Vbias 0.27994f
C16965 Nand_Gate_4.A.n12 Vbias 0.27511f
C16966 Nand_Gate_4.A.n13 Vbias 0.03007f
C16967 Nand_Gate_4.A.t7 Vbias 0.14554f
C16968 Nand_Gate_4.A.n14 Vbias 0.04192f
C16969 Nand_Gate_4.A.n15 Vbias 0.01797f
C16970 Nand_Gate_4.A.n16 Vbias 0.03367f
C16971 Nand_Gate_4.A.n18 Vbias 0.12656f
C16972 Nand_Gate_4.A.n19 Vbias 0.03459f
C16973 Nand_Gate_4.A.n20 Vbias 0.09204f
C16974 Nand_Gate_4.A.t8 Vbias 0.14555f
C16975 Nand_Gate_4.A.n21 Vbias 0.14257f
C16976 Nand_Gate_4.A.n22 Vbias 0.03007f
C16977 Nand_Gate_4.A.t6 Vbias 0.27993f
C16978 Nand_Gate_4.A.n23 Vbias 0.08177f
C16979 Nand_Gate_4.A.n24 Vbias 0.02035f
C16980 Nand_Gate_4.A.n25 Vbias 0.0296f
C16981 Nand_Gate_4.A.n26 Vbias 0.14551f
C16982 Nand_Gate_4.A.n27 Vbias 0.25531f
C16983 Nand_Gate_4.A.n28 Vbias 0.15873f
C16984 Nand_Gate_4.A.n29 Vbias 0.34318f
C16985 Nand_Gate_4.A.n31 Vbias 0.04546f
C16986 Nand_Gate_4.A.n32 Vbias 0.02608f
C16987 Nand_Gate_4.A.t0 Vbias 0.03876f
C16988 Nand_Gate_4.A.t3 Vbias 0.03797f
C16989 Nand_Gate_4.A.n33 Vbias 0.21593f
C16990 Nand_Gate_4.A.n34 Vbias 0.07184f
C16991 Nand_Gate_4.A.t2 Vbias 0.03797f
C16992 Nand_Gate_4.A.n35 Vbias 0.05849f
C16993 Nand_Gate_4.A.n36 Vbias 0.10356f
C16994 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t3 Vbias 0.07037f
C16995 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n0 Vbias 0.16004f
C16996 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n1 Vbias 0.07725f
C16997 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t5 Vbias 0.2799f
C16998 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n2 Vbias 0.27418f
C16999 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n3 Vbias 0.05783f
C17000 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t4 Vbias 0.53832f
C17001 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n4 Vbias 0.15726f
C17002 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n5 Vbias 0.03913f
C17003 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n6 Vbias 0.05692f
C17004 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n7 Vbias 0.14585f
C17005 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n8 Vbias 0.14585f
C17006 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n9 Vbias 0.07581f
C17007 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t2 Vbias 0.07318f
C17008 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t0 Vbias 0.07454f
C17009 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.t1 Vbias 0.07302f
C17010 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n10 Vbias 0.41525f
C17011 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n11 Vbias 0.23391f
C17012 RingCounter_0.D_FlipFlop_8.3-input-nand_1.Vout.n12 Vbias 0.22303f
C17013 CLK.t64 Vbias 0.34775f
C17014 CLK.n0 Vbias 0.36055f
C17015 CLK.n1 Vbias 0.03901f
C17016 CLK.n2 Vbias 0.05208f
C17017 CLK.t95 Vbias 0.16006f
C17018 CLK.n3 Vbias 0.13494f
C17019 CLK.n4 Vbias 0.04584f
C17020 CLK.t86 Vbias 0.34774f
C17021 CLK.t33 Vbias 0.1808f
C17022 CLK.n5 Vbias 0.19066f
C17023 CLK.t82 Vbias 0.34774f
C17024 CLK.n6 Vbias 0.30782f
C17025 CLK.n7 Vbias 0.30867f
C17026 CLK.n8 Vbias 0.19316f
C17027 CLK.t42 Vbias 0.16007f
C17028 CLK.n9 Vbias 0.01795f
C17029 CLK.n10 Vbias 0.04351f
C17030 CLK.n11 Vbias 0.46223f
C17031 CLK.t46 Vbias 0.34775f
C17032 CLK.n12 Vbias 0.36055f
C17033 CLK.n13 Vbias 0.03901f
C17034 CLK.n14 Vbias 0.05208f
C17035 CLK.t27 Vbias 0.16006f
C17036 CLK.n15 Vbias 0.13494f
C17037 CLK.n16 Vbias 0.04584f
C17038 CLK.t79 Vbias 0.34774f
C17039 CLK.t57 Vbias 0.1808f
C17040 CLK.n17 Vbias 0.19066f
C17041 CLK.t7 Vbias 0.34774f
C17042 CLK.n18 Vbias 0.30782f
C17043 CLK.n19 Vbias 0.30867f
C17044 CLK.n20 Vbias 0.19316f
C17045 CLK.t113 Vbias 0.16007f
C17046 CLK.n21 Vbias 0.01795f
C17047 CLK.n22 Vbias 0.04351f
C17048 CLK.n23 Vbias 0.161f
C17049 CLK.t9 Vbias 0.34775f
C17050 CLK.n24 Vbias 0.36055f
C17051 CLK.n25 Vbias 0.03901f
C17052 CLK.n26 Vbias 0.05208f
C17053 CLK.t117 Vbias 0.16006f
C17054 CLK.n27 Vbias 0.13494f
C17055 CLK.n28 Vbias 0.04584f
C17056 CLK.t36 Vbias 0.34774f
C17057 CLK.t88 Vbias 0.1808f
C17058 CLK.n29 Vbias 0.19066f
C17059 CLK.t73 Vbias 0.34774f
C17060 CLK.n30 Vbias 0.30782f
C17061 CLK.n31 Vbias 0.30867f
C17062 CLK.n32 Vbias 0.19316f
C17063 CLK.t70 Vbias 0.16007f
C17064 CLK.n33 Vbias 0.01795f
C17065 CLK.n34 Vbias 0.04351f
C17066 CLK.n35 Vbias 0.74111f
C17067 CLK.t71 Vbias 0.34775f
C17068 CLK.n36 Vbias 0.36055f
C17069 CLK.n37 Vbias 0.03901f
C17070 CLK.n38 Vbias 0.05208f
C17071 CLK.t54 Vbias 0.16006f
C17072 CLK.n39 Vbias 0.13494f
C17073 CLK.n40 Vbias 0.04584f
C17074 CLK.t112 Vbias 0.34774f
C17075 CLK.t28 Vbias 0.1808f
C17076 CLK.n41 Vbias 0.19066f
C17077 CLK.t101 Vbias 0.34774f
C17078 CLK.n42 Vbias 0.30782f
C17079 CLK.n43 Vbias 0.30867f
C17080 CLK.n44 Vbias 0.19316f
C17081 CLK.t19 Vbias 0.16007f
C17082 CLK.n45 Vbias 0.01795f
C17083 CLK.n46 Vbias 0.04351f
C17084 CLK.n48 Vbias 2.31789f
C17085 CLK.t99 Vbias 0.34775f
C17086 CLK.n49 Vbias 0.36055f
C17087 CLK.n50 Vbias 0.03901f
C17088 CLK.n51 Vbias 0.05208f
C17089 CLK.t84 Vbias 0.16006f
C17090 CLK.n52 Vbias 0.13494f
C17091 CLK.n53 Vbias 0.04584f
C17092 CLK.t14 Vbias 0.34774f
C17093 CLK.t55 Vbias 0.1808f
C17094 CLK.n54 Vbias 0.19066f
C17095 CLK.t4 Vbias 0.34774f
C17096 CLK.n55 Vbias 0.30782f
C17097 CLK.n56 Vbias 0.30867f
C17098 CLK.n57 Vbias 0.19316f
C17099 CLK.t38 Vbias 0.16007f
C17100 CLK.n58 Vbias 0.01795f
C17101 CLK.n59 Vbias 0.04351f
C17102 CLK.n61 Vbias 2.02899f
C17103 CLK.t41 Vbias 0.34775f
C17104 CLK.n62 Vbias 0.36055f
C17105 CLK.n63 Vbias 0.03901f
C17106 CLK.n64 Vbias 0.05208f
C17107 CLK.t114 Vbias 0.16006f
C17108 CLK.n65 Vbias 0.13494f
C17109 CLK.n66 Vbias 0.04584f
C17110 CLK.t76 Vbias 0.34774f
C17111 CLK.t11 Vbias 0.1808f
C17112 CLK.n67 Vbias 0.19066f
C17113 CLK.t66 Vbias 0.34774f
C17114 CLK.n68 Vbias 0.30782f
C17115 CLK.n69 Vbias 0.30867f
C17116 CLK.n70 Vbias 0.19316f
C17117 CLK.t63 Vbias 0.16007f
C17118 CLK.n71 Vbias 0.01795f
C17119 CLK.n72 Vbias 0.04351f
C17120 CLK.n74 Vbias 2.02899f
C17121 CLK.t65 Vbias 0.34775f
C17122 CLK.n75 Vbias 0.36055f
C17123 CLK.n76 Vbias 0.03901f
C17124 CLK.n77 Vbias 0.05208f
C17125 CLK.t51 Vbias 0.16006f
C17126 CLK.n78 Vbias 0.13494f
C17127 CLK.n79 Vbias 0.04584f
C17128 CLK.t109 Vbias 0.34774f
C17129 CLK.t25 Vbias 0.1808f
C17130 CLK.n80 Vbias 0.19066f
C17131 CLK.t92 Vbias 0.34774f
C17132 CLK.n81 Vbias 0.30782f
C17133 CLK.n82 Vbias 0.30867f
C17134 CLK.n83 Vbias 0.19316f
C17135 CLK.t16 Vbias 0.16007f
C17136 CLK.n84 Vbias 0.01795f
C17137 CLK.n85 Vbias 0.04351f
C17138 CLK.n87 Vbias 2.02899f
C17139 CLK.t91 Vbias 0.34775f
C17140 CLK.n88 Vbias 0.36055f
C17141 CLK.n89 Vbias 0.03901f
C17142 CLK.n90 Vbias 0.05208f
C17143 CLK.t80 Vbias 0.16006f
C17144 CLK.n91 Vbias 0.13494f
C17145 CLK.n92 Vbias 0.04584f
C17146 CLK.t12 Vbias 0.34774f
C17147 CLK.t52 Vbias 0.1808f
C17148 CLK.n93 Vbias 0.19066f
C17149 CLK.t32 Vbias 0.34774f
C17150 CLK.n94 Vbias 0.30782f
C17151 CLK.n95 Vbias 0.30867f
C17152 CLK.n96 Vbias 0.19316f
C17153 CLK.t30 Vbias 0.16007f
C17154 CLK.n97 Vbias 0.01795f
C17155 CLK.n98 Vbias 0.04351f
C17156 CLK.n100 Vbias 2.02899f
C17157 CLK.t20 Vbias 0.34775f
C17158 CLK.n101 Vbias 0.36055f
C17159 CLK.n102 Vbias 0.03901f
C17160 CLK.n103 Vbias 0.05208f
C17161 CLK.t13 Vbias 0.16006f
C17162 CLK.n104 Vbias 0.13494f
C17163 CLK.n105 Vbias 0.04584f
C17164 CLK.t50 Vbias 0.34774f
C17165 CLK.t31 Vbias 0.1808f
C17166 CLK.n106 Vbias 0.19066f
C17167 CLK.t104 Vbias 0.34774f
C17168 CLK.n107 Vbias 0.30782f
C17169 CLK.n108 Vbias 0.30867f
C17170 CLK.n109 Vbias 0.19316f
C17171 CLK.t83 Vbias 0.16007f
C17172 CLK.n110 Vbias 0.01795f
C17173 CLK.n111 Vbias 0.04351f
C17174 CLK.n113 Vbias 1.6993f
C17175 CLK.n114 Vbias 1.33849f
C17176 CLK.n115 Vbias 3.26289f
C17177 CLK.t77 Vbias 0.1808f
C17178 CLK.t3 Vbias 0.34774f
C17179 CLK.n116 Vbias 0.10158f
C17180 CLK.n117 Vbias 0.04344f
C17181 CLK.n118 Vbias 0.08021f
C17182 CLK.n119 Vbias 1.49061f
C17183 CLK.t105 Vbias 0.1808f
C17184 CLK.t21 Vbias 0.34774f
C17185 CLK.n120 Vbias 0.10158f
C17186 CLK.n121 Vbias 0.04344f
C17187 CLK.n122 Vbias 0.08021f
C17188 CLK.n123 Vbias 0.04177f
C17189 CLK.n124 Vbias 2.2385f
C17190 CLK.t18 Vbias 0.1808f
C17191 CLK.n125 Vbias 0.19316f
C17192 CLK.t49 Vbias 0.34774f
C17193 CLK.n126 Vbias 0.78151f
C17194 CLK.n127 Vbias 1.66232f
C17195 CLK.t44 Vbias 0.1808f
C17196 CLK.n128 Vbias 0.19316f
C17197 CLK.t81 Vbias 0.34774f
C17198 CLK.n129 Vbias 0.1094f
C17199 CLK.n130 Vbias 2.33217f
C17200 CLK.t87 Vbias 0.1808f
C17201 CLK.n131 Vbias 0.19316f
C17202 CLK.t48 Vbias 0.34774f
C17203 CLK.n132 Vbias 0.1094f
C17204 CLK.n133 Vbias 1.80643f
C17205 CLK.t34 Vbias 0.1808f
C17206 CLK.n134 Vbias 0.19316f
C17207 CLK.t43 Vbias 0.34774f
C17208 CLK.n135 Vbias 1.30135f
C17209 CLK.n136 Vbias 4.44918f
C17210 CLK.n137 Vbias 4.34264f
C17211 CLK.t74 Vbias 0.1808f
C17212 CLK.t115 Vbias 0.34774f
C17213 CLK.n138 Vbias 0.10158f
C17214 CLK.n139 Vbias 0.04344f
C17215 CLK.n140 Vbias 0.08021f
C17216 CLK.n141 Vbias 0.04177f
C17217 CLK.n142 Vbias 2.54051f
C17218 CLK.t110 Vbias 0.1808f
C17219 CLK.t61 Vbias 0.34774f
C17220 CLK.n143 Vbias 0.10158f
C17221 CLK.n144 Vbias 0.04344f
C17222 CLK.n145 Vbias 0.08021f
C17223 CLK.n146 Vbias 0.04177f
C17224 CLK.n147 Vbias 1.63439f
C17225 CLK.n148 Vbias 3.26269f
C17226 CLK.n149 Vbias 1.09574f
C17227 CLK.n150 Vbias 0.6418f
C17228 CLK.t68 Vbias 0.34775f
C17229 CLK.n151 Vbias 0.36055f
C17230 CLK.n152 Vbias 0.03901f
C17231 CLK.n153 Vbias 0.05208f
C17232 CLK.t102 Vbias 0.16006f
C17233 CLK.n154 Vbias 0.13494f
C17234 CLK.n155 Vbias 0.04584f
C17235 CLK.t90 Vbias 0.34774f
C17236 CLK.t17 Vbias 0.1808f
C17237 CLK.n156 Vbias 0.19066f
C17238 CLK.t106 Vbias 0.34774f
C17239 CLK.n157 Vbias 0.30782f
C17240 CLK.n158 Vbias 0.30867f
C17241 CLK.n159 Vbias 0.19316f
C17242 CLK.t45 Vbias 0.16007f
C17243 CLK.n160 Vbias 0.01795f
C17244 CLK.n161 Vbias 0.04351f
C17245 CLK.n162 Vbias 0.74111f
C17246 CLK.t96 Vbias 0.34775f
C17247 CLK.n163 Vbias 0.36055f
C17248 CLK.n164 Vbias 0.03901f
C17249 CLK.n165 Vbias 0.05208f
C17250 CLK.t5 Vbias 0.16006f
C17251 CLK.n166 Vbias 0.13494f
C17252 CLK.n167 Vbias 0.04584f
C17253 CLK.t0 Vbias 0.34774f
C17254 CLK.t78 Vbias 0.1808f
C17255 CLK.n168 Vbias 0.19066f
C17256 CLK.t10 Vbias 0.34774f
C17257 CLK.n169 Vbias 0.30782f
C17258 CLK.n170 Vbias 0.30867f
C17259 CLK.n171 Vbias 0.19316f
C17260 CLK.t69 Vbias 0.16007f
C17261 CLK.n172 Vbias 0.01795f
C17262 CLK.n173 Vbias 0.04351f
C17263 CLK.n175 Vbias 2.31789f
C17264 CLK.t35 Vbias 0.34775f
C17265 CLK.n176 Vbias 0.36055f
C17266 CLK.n177 Vbias 0.03901f
C17267 CLK.n178 Vbias 0.05208f
C17268 CLK.t22 Vbias 0.16006f
C17269 CLK.n179 Vbias 0.13494f
C17270 CLK.n180 Vbias 0.04584f
C17271 CLK.t56 Vbias 0.34774f
C17272 CLK.t111 Vbias 0.1808f
C17273 CLK.n181 Vbias 0.19066f
C17274 CLK.t24 Vbias 0.34774f
C17275 CLK.n182 Vbias 0.30782f
C17276 CLK.n183 Vbias 0.30867f
C17277 CLK.n184 Vbias 0.19316f
C17278 CLK.t97 Vbias 0.16007f
C17279 CLK.n185 Vbias 0.01795f
C17280 CLK.n186 Vbias 0.04351f
C17281 CLK.n188 Vbias 2.02899f
C17282 CLK.t60 Vbias 0.34775f
C17283 CLK.n189 Vbias 0.36055f
C17284 CLK.n190 Vbias 0.03901f
C17285 CLK.n191 Vbias 0.05208f
C17286 CLK.t93 Vbias 0.16006f
C17287 CLK.n192 Vbias 0.13494f
C17288 CLK.n193 Vbias 0.04584f
C17289 CLK.t85 Vbias 0.34774f
C17290 CLK.t47 Vbias 0.1808f
C17291 CLK.n194 Vbias 0.19066f
C17292 CLK.t103 Vbias 0.34774f
C17293 CLK.n195 Vbias 0.30782f
C17294 CLK.n196 Vbias 0.30867f
C17295 CLK.n197 Vbias 0.19316f
C17296 CLK.t37 Vbias 0.16007f
C17297 CLK.n198 Vbias 0.01795f
C17298 CLK.n199 Vbias 0.04351f
C17299 CLK.n201 Vbias 2.02899f
C17300 CLK.t89 Vbias 0.34775f
C17301 CLK.n202 Vbias 0.36055f
C17302 CLK.n203 Vbias 0.03901f
C17303 CLK.n204 Vbias 0.05208f
C17304 CLK.t2 Vbias 0.16006f
C17305 CLK.n205 Vbias 0.13494f
C17306 CLK.n206 Vbias 0.04584f
C17307 CLK.t116 Vbias 0.34774f
C17308 CLK.t75 Vbias 0.1808f
C17309 CLK.n207 Vbias 0.19066f
C17310 CLK.t6 Vbias 0.34774f
C17311 CLK.n208 Vbias 0.30782f
C17312 CLK.n209 Vbias 0.30867f
C17313 CLK.n210 Vbias 0.19316f
C17314 CLK.t62 Vbias 0.16007f
C17315 CLK.n211 Vbias 0.01795f
C17316 CLK.n212 Vbias 0.04351f
C17317 CLK.n214 Vbias 2.02899f
C17318 CLK.t29 Vbias 0.34775f
C17319 CLK.n215 Vbias 0.36055f
C17320 CLK.n216 Vbias 0.03901f
C17321 CLK.n217 Vbias 0.05208f
C17322 CLK.t59 Vbias 0.16006f
C17323 CLK.n218 Vbias 0.13494f
C17324 CLK.n219 Vbias 0.04584f
C17325 CLK.t53 Vbias 0.34774f
C17326 CLK.t108 Vbias 0.1808f
C17327 CLK.n220 Vbias 0.19066f
C17328 CLK.t67 Vbias 0.34774f
C17329 CLK.n221 Vbias 0.30782f
C17330 CLK.n222 Vbias 0.30867f
C17331 CLK.n223 Vbias 0.19316f
C17332 CLK.t15 Vbias 0.16007f
C17333 CLK.n224 Vbias 0.01795f
C17334 CLK.n225 Vbias 0.04351f
C17335 CLK.n227 Vbias 2.02899f
C17336 CLK.t98 Vbias 0.34775f
C17337 CLK.n228 Vbias 0.36055f
C17338 CLK.n229 Vbias 0.03901f
C17339 CLK.n230 Vbias 0.05208f
C17340 CLK.t8 Vbias 0.16006f
C17341 CLK.n231 Vbias 0.13494f
C17342 CLK.n232 Vbias 0.04584f
C17343 CLK.t1 Vbias 0.34774f
C17344 CLK.t26 Vbias 0.1808f
C17345 CLK.n233 Vbias 0.19066f
C17346 CLK.t94 Vbias 0.34774f
C17347 CLK.n234 Vbias 0.30782f
C17348 CLK.n235 Vbias 0.30867f
C17349 CLK.n236 Vbias 0.19316f
C17350 CLK.t72 Vbias 0.16007f
C17351 CLK.n237 Vbias 0.01795f
C17352 CLK.n238 Vbias 0.04351f
C17353 CLK.n240 Vbias 2.02899f
C17354 CLK.t40 Vbias 0.34775f
C17355 CLK.n241 Vbias 0.36055f
C17356 CLK.n242 Vbias 0.03901f
C17357 CLK.n243 Vbias 0.05208f
C17358 CLK.t23 Vbias 0.16006f
C17359 CLK.n244 Vbias 0.13494f
C17360 CLK.n245 Vbias 0.04584f
C17361 CLK.t58 Vbias 0.34774f
C17362 CLK.t39 Vbias 0.1808f
C17363 CLK.n246 Vbias 0.19066f
C17364 CLK.t107 Vbias 0.34774f
C17365 CLK.n247 Vbias 0.30782f
C17366 CLK.n248 Vbias 0.30867f
C17367 CLK.n249 Vbias 0.19316f
C17368 CLK.t100 Vbias 0.16007f
C17369 CLK.n250 Vbias 0.01795f
C17370 CLK.n251 Vbias 0.04351f
C17371 CLK.n253 Vbias 1.01773f
C17372 CLK.n254 Vbias 0.30418f
C17373 EN.t16 Vbias 0.26445f
C17374 EN.n0 Vbias 0.07618f
C17375 EN.n1 Vbias 0.02029f
C17376 EN.n2 Vbias 0.03162f
C17377 EN.t54 Vbias 0.50863f
C17378 EN.n3 Vbias 0.14859f
C17379 EN.n4 Vbias 0.06447f
C17380 EN.n5 Vbias 0.28347f
C17381 EN.t98 Vbias 0.23655f
C17382 EN.n6 Vbias 0.13574f
C17383 EN.n7 Vbias 0.42089f
C17384 EN.t74 Vbias 0.50866f
C17385 EN.n8 Vbias 0.51224f
C17386 EN.n9 Vbias 0.05464f
C17387 EN.t38 Vbias 0.26445f
C17388 EN.n10 Vbias 0.07618f
C17389 EN.n11 Vbias 0.02029f
C17390 EN.n12 Vbias 0.03162f
C17391 EN.n14 Vbias 0.81908f
C17392 EN.n15 Vbias 0.31544f
C17393 EN.n16 Vbias 0.05464f
C17394 EN.n17 Vbias 2.28323f
C17395 EN.t86 Vbias 0.50866f
C17396 EN.n18 Vbias 0.51224f
C17397 EN.n19 Vbias 0.05464f
C17398 EN.t106 Vbias 0.26445f
C17399 EN.n20 Vbias 0.07618f
C17400 EN.n21 Vbias 0.02029f
C17401 EN.n22 Vbias 0.03162f
C17402 EN.n23 Vbias 0.31544f
C17403 EN.t8 Vbias 0.50866f
C17404 EN.n24 Vbias 0.51224f
C17405 EN.n25 Vbias 0.05464f
C17406 EN.t29 Vbias 0.26445f
C17407 EN.n26 Vbias 0.07618f
C17408 EN.n27 Vbias 0.02029f
C17409 EN.n28 Vbias 0.03162f
C17410 EN.n30 Vbias 0.70253f
C17411 EN.t65 Vbias 0.50863f
C17412 EN.n31 Vbias 0.14859f
C17413 EN.n32 Vbias 0.06447f
C17414 EN.n33 Vbias 0.28347f
C17415 EN.t81 Vbias 0.23655f
C17416 EN.n34 Vbias 0.13574f
C17417 EN.n35 Vbias 0.3113f
C17418 EN.n36 Vbias 0.38457f
C17419 EN.t7 Vbias 0.50866f
C17420 EN.n37 Vbias 0.51224f
C17421 EN.n38 Vbias 0.05464f
C17422 EN.t26 Vbias 0.26445f
C17423 EN.n39 Vbias 0.07618f
C17424 EN.n40 Vbias 0.02029f
C17425 EN.n41 Vbias 0.03162f
C17426 EN.n42 Vbias 0.31544f
C17427 EN.t64 Vbias 0.50866f
C17428 EN.n43 Vbias 0.51224f
C17429 EN.n44 Vbias 0.05464f
C17430 EN.t49 Vbias 0.26445f
C17431 EN.n45 Vbias 0.07618f
C17432 EN.n46 Vbias 0.02029f
C17433 EN.n47 Vbias 0.03162f
C17434 EN.n49 Vbias 0.70253f
C17435 EN.t84 Vbias 0.50863f
C17436 EN.n50 Vbias 0.14859f
C17437 EN.n51 Vbias 0.06447f
C17438 EN.n52 Vbias 0.28347f
C17439 EN.t40 Vbias 0.23655f
C17440 EN.n53 Vbias 0.13574f
C17441 EN.n54 Vbias 0.3113f
C17442 EN.n55 Vbias 0.38457f
C17443 EN.n56 Vbias 2.21237f
C17444 EN.n57 Vbias 5.01882f
C17445 EN.t41 Vbias 0.50866f
C17446 EN.n58 Vbias 0.52738f
C17447 EN.n59 Vbias 0.05705f
C17448 EN.n60 Vbias 0.07618f
C17449 EN.t56 Vbias 0.23758f
C17450 EN.n61 Vbias 0.47754f
C17451 EN.n62 Vbias 0.13574f
C17452 EN.t61 Vbias 0.26446f
C17453 EN.n63 Vbias 0.2467f
C17454 EN.n64 Vbias 0.05464f
C17455 EN.t87 Vbias 0.50863f
C17456 EN.n65 Vbias 0.14859f
C17457 EN.n66 Vbias 0.04933f
C17458 EN.n67 Vbias 0.08333f
C17459 EN.n68 Vbias 0.31544f
C17460 EN.t6 Vbias 0.26446f
C17461 EN.n69 Vbias 0.2467f
C17462 EN.n70 Vbias 0.05464f
C17463 EN.t43 Vbias 0.50863f
C17464 EN.n71 Vbias 0.14859f
C17465 EN.n72 Vbias 0.04933f
C17466 EN.n73 Vbias 0.08333f
C17467 EN.n75 Vbias 0.80102f
C17468 EN.n76 Vbias 2.60416f
C17469 EN.n77 Vbias 2.39848f
C17470 EN.n78 Vbias 4.41011f
C17471 EN.n79 Vbias 7.03069f
C17472 EN.n80 Vbias 1.6489f
C17473 EN.n81 Vbias 2.28323f
C17474 EN.t27 Vbias 0.50866f
C17475 EN.n82 Vbias 0.51224f
C17476 EN.n83 Vbias 0.05464f
C17477 EN.t45 Vbias 0.26445f
C17478 EN.n84 Vbias 0.07618f
C17479 EN.n85 Vbias 0.02029f
C17480 EN.n86 Vbias 0.03162f
C17481 EN.n87 Vbias 0.31544f
C17482 EN.t83 Vbias 0.50866f
C17483 EN.n88 Vbias 0.51224f
C17484 EN.n89 Vbias 0.05464f
C17485 EN.t66 Vbias 0.26445f
C17486 EN.n90 Vbias 0.07618f
C17487 EN.n91 Vbias 0.02029f
C17488 EN.n92 Vbias 0.03162f
C17489 EN.n94 Vbias 0.70253f
C17490 EN.t102 Vbias 0.50863f
C17491 EN.n95 Vbias 0.14859f
C17492 EN.n96 Vbias 0.06447f
C17493 EN.n97 Vbias 0.28347f
C17494 EN.t60 Vbias 0.23655f
C17495 EN.n98 Vbias 0.13574f
C17496 EN.n99 Vbias 0.3113f
C17497 EN.n100 Vbias 0.38457f
C17498 EN.t11 Vbias 0.26445f
C17499 EN.n101 Vbias 0.07618f
C17500 EN.n102 Vbias 0.02029f
C17501 EN.n103 Vbias 0.03162f
C17502 EN.t70 Vbias 0.50863f
C17503 EN.n104 Vbias 0.14859f
C17504 EN.n105 Vbias 0.06447f
C17505 EN.n106 Vbias 0.28347f
C17506 EN.t35 Vbias 0.23655f
C17507 EN.n107 Vbias 0.13574f
C17508 EN.n108 Vbias 0.42089f
C17509 EN.t22 Vbias 0.50866f
C17510 EN.n109 Vbias 0.51224f
C17511 EN.n110 Vbias 0.05464f
C17512 EN.t18 Vbias 0.26445f
C17513 EN.n111 Vbias 0.07618f
C17514 EN.n112 Vbias 0.02029f
C17515 EN.n113 Vbias 0.03162f
C17516 EN.n115 Vbias 0.81908f
C17517 EN.n116 Vbias 0.31544f
C17518 EN.n117 Vbias 0.05464f
C17519 EN.n118 Vbias 0.51224f
C17520 EN.t19 Vbias 0.45736f
C17521 EN.n119 Vbias 2.28323f
C17522 EN.t4 Vbias 0.50866f
C17523 EN.n120 Vbias 0.51224f
C17524 EN.n121 Vbias 0.05464f
C17525 EN.t25 Vbias 0.26445f
C17526 EN.n122 Vbias 0.07618f
C17527 EN.n123 Vbias 0.02029f
C17528 EN.n124 Vbias 0.03162f
C17529 EN.n125 Vbias 0.31544f
C17530 EN.t0 Vbias 0.50866f
C17531 EN.n126 Vbias 0.51224f
C17532 EN.n127 Vbias 0.05464f
C17533 EN.t89 Vbias 0.26445f
C17534 EN.n128 Vbias 0.07618f
C17535 EN.n129 Vbias 0.02029f
C17536 EN.n130 Vbias 0.03162f
C17537 EN.n132 Vbias 0.70253f
C17538 EN.t32 Vbias 0.50863f
C17539 EN.n133 Vbias 0.14859f
C17540 EN.n134 Vbias 0.06447f
C17541 EN.n135 Vbias 0.28347f
C17542 EN.t77 Vbias 0.23655f
C17543 EN.n136 Vbias 0.13574f
C17544 EN.n137 Vbias 0.3113f
C17545 EN.n138 Vbias 0.38457f
C17546 EN.t12 Vbias 0.26446f
C17547 EN.n139 Vbias 0.2467f
C17548 EN.n140 Vbias 0.05464f
C17549 EN.t95 Vbias 0.50863f
C17550 EN.n141 Vbias 0.14859f
C17551 EN.n142 Vbias 0.04933f
C17552 EN.n143 Vbias 0.08333f
C17553 EN.n144 Vbias 0.31544f
C17554 EN.t10 Vbias 0.26446f
C17555 EN.n145 Vbias 0.2467f
C17556 EN.n146 Vbias 0.05464f
C17557 EN.t62 Vbias 0.50863f
C17558 EN.n147 Vbias 0.14859f
C17559 EN.n148 Vbias 0.04933f
C17560 EN.n149 Vbias 0.08333f
C17561 EN.n151 Vbias 0.70253f
C17562 EN.t20 Vbias 0.50866f
C17563 EN.n152 Vbias 0.52738f
C17564 EN.n153 Vbias 0.05705f
C17565 EN.n154 Vbias 0.07618f
C17566 EN.t42 Vbias 0.23758f
C17567 EN.n155 Vbias 0.47754f
C17568 EN.n156 Vbias 0.13574f
C17569 EN.n157 Vbias 0.24515f
C17570 EN.t93 Vbias 0.26445f
C17571 EN.n158 Vbias 0.07618f
C17572 EN.n159 Vbias 0.02029f
C17573 EN.n160 Vbias 0.03162f
C17574 EN.t3 Vbias 0.50863f
C17575 EN.n161 Vbias 0.14859f
C17576 EN.n162 Vbias 0.06447f
C17577 EN.n163 Vbias 0.28347f
C17578 EN.t37 Vbias 0.23655f
C17579 EN.n164 Vbias 0.13574f
C17580 EN.n165 Vbias 0.42089f
C17581 EN.t107 Vbias 0.50866f
C17582 EN.n166 Vbias 0.51224f
C17583 EN.n167 Vbias 0.05464f
C17584 EN.t101 Vbias 0.26445f
C17585 EN.n168 Vbias 0.07618f
C17586 EN.n169 Vbias 0.02029f
C17587 EN.n170 Vbias 0.03162f
C17588 EN.n172 Vbias 0.81908f
C17589 EN.n173 Vbias 0.31544f
C17590 EN.n174 Vbias 0.05464f
C17591 EN.n175 Vbias 0.51224f
C17592 EN.t73 Vbias 0.45736f
C17593 EN.t94 Vbias 0.26445f
C17594 EN.n176 Vbias 0.07618f
C17595 EN.n177 Vbias 0.02029f
C17596 EN.n178 Vbias 0.03162f
C17597 EN.t59 Vbias 0.50863f
C17598 EN.n179 Vbias 0.14859f
C17599 EN.n180 Vbias 0.06447f
C17600 EN.n181 Vbias 0.28347f
C17601 EN.t13 Vbias 0.23655f
C17602 EN.n182 Vbias 0.13574f
C17603 EN.n183 Vbias 0.42089f
C17604 EN.t57 Vbias 0.50866f
C17605 EN.n184 Vbias 0.51224f
C17606 EN.n185 Vbias 0.05464f
C17607 EN.t50 Vbias 0.26445f
C17608 EN.n186 Vbias 0.07618f
C17609 EN.n187 Vbias 0.02029f
C17610 EN.n188 Vbias 0.03162f
C17611 EN.n190 Vbias 0.81908f
C17612 EN.n191 Vbias 0.31544f
C17613 EN.n192 Vbias 0.05464f
C17614 EN.n193 Vbias 0.51224f
C17615 EN.t1 Vbias 0.8262f
C17616 EN.n194 Vbias 3.30704f
C17617 EN.n195 Vbias 4.64174f
C17618 EN.n196 Vbias 5.73599f
C17619 EN.t85 Vbias 0.50866f
C17620 EN.n197 Vbias 0.51224f
C17621 EN.n198 Vbias 0.05464f
C17622 EN.t104 Vbias 0.26445f
C17623 EN.n199 Vbias 0.07618f
C17624 EN.n200 Vbias 0.02029f
C17625 EN.n201 Vbias 0.03162f
C17626 EN.n202 Vbias 0.31544f
C17627 EN.t58 Vbias 0.50866f
C17628 EN.n203 Vbias 0.51224f
C17629 EN.n204 Vbias 0.05464f
C17630 EN.t71 Vbias 0.26445f
C17631 EN.n205 Vbias 0.07618f
C17632 EN.n206 Vbias 0.02029f
C17633 EN.n207 Vbias 0.03162f
C17634 EN.n209 Vbias 0.70253f
C17635 EN.t2 Vbias 0.50863f
C17636 EN.n210 Vbias 0.14859f
C17637 EN.n211 Vbias 0.06447f
C17638 EN.n212 Vbias 0.28347f
C17639 EN.t21 Vbias 0.23655f
C17640 EN.n213 Vbias 0.13574f
C17641 EN.n214 Vbias 0.3113f
C17642 EN.n215 Vbias 0.38457f
C17643 EN.t15 Vbias 0.26445f
C17644 EN.n216 Vbias 0.07618f
C17645 EN.n217 Vbias 0.02029f
C17646 EN.n218 Vbias 0.03162f
C17647 EN.t33 Vbias 0.50863f
C17648 EN.n219 Vbias 0.14859f
C17649 EN.n220 Vbias 0.06447f
C17650 EN.n221 Vbias 0.28347f
C17651 EN.t88 Vbias 0.23655f
C17652 EN.n222 Vbias 0.13574f
C17653 EN.n223 Vbias 0.42089f
C17654 EN.t28 Vbias 0.50866f
C17655 EN.n224 Vbias 0.51224f
C17656 EN.n225 Vbias 0.05464f
C17657 EN.t23 Vbias 0.26445f
C17658 EN.n226 Vbias 0.07618f
C17659 EN.n227 Vbias 0.02029f
C17660 EN.n228 Vbias 0.03162f
C17661 EN.n230 Vbias 0.81908f
C17662 EN.n231 Vbias 0.31544f
C17663 EN.n232 Vbias 0.05464f
C17664 EN.n233 Vbias 0.51224f
C17665 EN.t91 Vbias 0.45736f
C17666 EN.n234 Vbias 4.64174f
C17667 EN.n235 Vbias 5.02091f
C17668 EN.n236 Vbias 2.40127f
C17669 EN.n237 Vbias 2.28323f
C17670 EN.n238 Vbias 5.02091f
C17671 EN.t72 Vbias 0.26445f
C17672 EN.n239 Vbias 0.07618f
C17673 EN.n240 Vbias 0.02029f
C17674 EN.n241 Vbias 0.03162f
C17675 EN.t52 Vbias 0.50863f
C17676 EN.n242 Vbias 0.14859f
C17677 EN.n243 Vbias 0.06447f
C17678 EN.n244 Vbias 0.28347f
C17679 EN.t9 Vbias 0.23655f
C17680 EN.n245 Vbias 0.13574f
C17681 EN.n246 Vbias 0.42089f
C17682 EN.t82 Vbias 0.50866f
C17683 EN.n247 Vbias 0.51224f
C17684 EN.n248 Vbias 0.05464f
C17685 EN.t47 Vbias 0.26445f
C17686 EN.n249 Vbias 0.07618f
C17687 EN.n250 Vbias 0.02029f
C17688 EN.n251 Vbias 0.03162f
C17689 EN.n253 Vbias 0.81908f
C17690 EN.n254 Vbias 0.31544f
C17691 EN.n255 Vbias 0.05464f
C17692 EN.n256 Vbias 0.51224f
C17693 EN.t48 Vbias 0.45736f
C17694 EN.n257 Vbias 4.64174f
C17695 EN.n258 Vbias 2.28323f
C17696 EN.t63 Vbias 0.50866f
C17697 EN.n259 Vbias 0.51224f
C17698 EN.n260 Vbias 0.05464f
C17699 EN.t80 Vbias 0.26445f
C17700 EN.n261 Vbias 0.07618f
C17701 EN.n262 Vbias 0.02029f
C17702 EN.n263 Vbias 0.03162f
C17703 EN.n264 Vbias 0.31544f
C17704 EN.t31 Vbias 0.50866f
C17705 EN.n265 Vbias 0.51224f
C17706 EN.n266 Vbias 0.05464f
C17707 EN.t46 Vbias 0.26445f
C17708 EN.n267 Vbias 0.07618f
C17709 EN.n268 Vbias 0.02029f
C17710 EN.n269 Vbias 0.03162f
C17711 EN.n271 Vbias 0.70253f
C17712 EN.t51 Vbias 0.50863f
C17713 EN.n272 Vbias 0.14859f
C17714 EN.n273 Vbias 0.06447f
C17715 EN.n274 Vbias 0.28347f
C17716 EN.t96 Vbias 0.23655f
C17717 EN.n275 Vbias 0.13574f
C17718 EN.n276 Vbias 0.3113f
C17719 EN.n277 Vbias 0.38457f
C17720 EN.n278 Vbias 5.02091f
C17721 EN.t90 Vbias 0.26445f
C17722 EN.n279 Vbias 0.07618f
C17723 EN.n280 Vbias 0.02029f
C17724 EN.n281 Vbias 0.03162f
C17725 EN.t103 Vbias 0.50863f
C17726 EN.n282 Vbias 0.14859f
C17727 EN.n283 Vbias 0.06447f
C17728 EN.n284 Vbias 0.28347f
C17729 EN.t36 Vbias 0.23655f
C17730 EN.n285 Vbias 0.13574f
C17731 EN.n286 Vbias 0.42089f
C17732 EN.t99 Vbias 0.50866f
C17733 EN.n287 Vbias 0.51224f
C17734 EN.n288 Vbias 0.05464f
C17735 EN.t97 Vbias 0.26445f
C17736 EN.n289 Vbias 0.07618f
C17737 EN.n290 Vbias 0.02029f
C17738 EN.n291 Vbias 0.03162f
C17739 EN.n293 Vbias 0.81908f
C17740 EN.n294 Vbias 0.31544f
C17741 EN.n295 Vbias 0.05464f
C17742 EN.n296 Vbias 0.51224f
C17743 EN.t69 Vbias 0.45736f
C17744 EN.n297 Vbias 4.64174f
C17745 EN.n298 Vbias 2.28323f
C17746 EN.n299 Vbias 2.28323f
C17747 EN.n300 Vbias 4.64174f
C17748 EN.n301 Vbias 5.02091f
C17749 EN.n302 Vbias 2.28323f
C17750 EN.t68 Vbias 0.50866f
C17751 EN.n303 Vbias 0.51224f
C17752 EN.n304 Vbias 0.05464f
C17753 EN.t55 Vbias 0.26445f
C17754 EN.n305 Vbias 0.07618f
C17755 EN.n306 Vbias 0.02029f
C17756 EN.n307 Vbias 0.03162f
C17757 EN.n308 Vbias 0.31544f
C17758 EN.t100 Vbias 0.50866f
C17759 EN.n309 Vbias 0.51224f
C17760 EN.n310 Vbias 0.05464f
C17761 EN.t17 Vbias 0.26445f
C17762 EN.n311 Vbias 0.07618f
C17763 EN.n312 Vbias 0.02029f
C17764 EN.n313 Vbias 0.03162f
C17765 EN.n315 Vbias 0.70253f
C17766 EN.t24 Vbias 0.50863f
C17767 EN.n316 Vbias 0.14859f
C17768 EN.n317 Vbias 0.06447f
C17769 EN.n318 Vbias 0.28347f
C17770 EN.t76 Vbias 0.23655f
C17771 EN.n319 Vbias 0.13574f
C17772 EN.n320 Vbias 0.3113f
C17773 EN.n321 Vbias 0.38457f
C17774 EN.t67 Vbias 0.26445f
C17775 EN.n322 Vbias 0.07618f
C17776 EN.n323 Vbias 0.02029f
C17777 EN.n324 Vbias 0.03162f
C17778 EN.t5 Vbias 0.50863f
C17779 EN.n325 Vbias 0.14859f
C17780 EN.n326 Vbias 0.06447f
C17781 EN.n327 Vbias 0.28347f
C17782 EN.t39 Vbias 0.23655f
C17783 EN.n328 Vbias 0.13574f
C17784 EN.n329 Vbias 0.42089f
C17785 EN.t78 Vbias 0.50866f
C17786 EN.n330 Vbias 0.51224f
C17787 EN.n331 Vbias 0.05464f
C17788 EN.t92 Vbias 0.26445f
C17789 EN.n332 Vbias 0.07618f
C17790 EN.n333 Vbias 0.02029f
C17791 EN.n334 Vbias 0.03162f
C17792 EN.n336 Vbias 0.81908f
C17793 EN.n337 Vbias 0.31544f
C17794 EN.n338 Vbias 0.05464f
C17795 EN.n339 Vbias 0.51224f
C17796 EN.t44 Vbias 0.45736f
C17797 EN.n340 Vbias 4.64174f
C17798 EN.n341 Vbias 5.02091f
C17799 EN.n342 Vbias 2.28323f
C17800 EN.n343 Vbias 2.40127f
C17801 EN.n344 Vbias 5.02091f
C17802 EN.t75 Vbias 0.26445f
C17803 EN.n345 Vbias 0.07618f
C17804 EN.n346 Vbias 0.02029f
C17805 EN.n347 Vbias 0.03162f
C17806 EN.t34 Vbias 0.50863f
C17807 EN.n348 Vbias 0.14859f
C17808 EN.n349 Vbias 0.06447f
C17809 EN.n350 Vbias 0.28347f
C17810 EN.t79 Vbias 0.23655f
C17811 EN.n351 Vbias 0.13574f
C17812 EN.n352 Vbias 0.42089f
C17813 EN.t30 Vbias 0.50866f
C17814 EN.n353 Vbias 0.51224f
C17815 EN.n354 Vbias 0.05464f
C17816 EN.t14 Vbias 0.26445f
C17817 EN.n355 Vbias 0.07618f
C17818 EN.n356 Vbias 0.02029f
C17819 EN.n357 Vbias 0.03162f
C17820 EN.n359 Vbias 0.81908f
C17821 EN.n360 Vbias 0.31544f
C17822 EN.n361 Vbias 0.05464f
C17823 EN.n362 Vbias 0.51224f
C17824 EN.t53 Vbias 0.45736f
C17825 EN.n363 Vbias 4.64174f
C17826 EN.n364 Vbias 2.40127f
C17827 EN.n365 Vbias 1.269f
C17828 EN.t105 Vbias 0.45736f
C17829 EN.n366 Vbias 0.51224f
C17830 CDAC8_0.switch_7.Z.t3 Vbias 0.03153f
C17831 CDAC8_0.switch_7.Z.t1 Vbias 0.03153f
C17832 CDAC8_0.switch_7.Z.n0 Vbias 0.11392f
C17833 CDAC8_0.switch_7.Z.n1 Vbias 0.2622f
C17834 CDAC8_0.switch_7.Z.t0 Vbias 0.0331f
C17835 CDAC8_0.switch_7.Z.n2 Vbias 2.15483f
C17836 CDAC8_0.switch_7.Z.n3 Vbias 0.71553f
C17837 CDAC8_0.switch_7.Z.t71 Vbias 5.57036f
C17838 CDAC8_0.switch_7.Z.n4 Vbias 1.29163f
C17839 CDAC8_0.switch_7.Z.n5 Vbias 0.84016f
C17840 CDAC8_0.switch_7.Z.t14 Vbias 5.57036f
C17841 CDAC8_0.switch_7.Z.n6 Vbias 1.29163f
C17842 CDAC8_0.switch_7.Z.t62 Vbias 5.57036f
C17843 CDAC8_0.switch_7.Z.n7 Vbias 1.29163f
C17844 CDAC8_0.switch_7.Z.n8 Vbias 0.71553f
C17845 CDAC8_0.switch_7.Z.n9 Vbias 1.0317f
C17846 CDAC8_0.switch_7.Z.t68 Vbias 5.57036f
C17847 CDAC8_0.switch_7.Z.n10 Vbias 1.29163f
C17848 CDAC8_0.switch_7.Z.t121 Vbias 5.57036f
C17849 CDAC8_0.switch_7.Z.n11 Vbias 1.29163f
C17850 CDAC8_0.switch_7.Z.t51 Vbias 5.57036f
C17851 CDAC8_0.switch_7.Z.n12 Vbias 1.29163f
C17852 CDAC8_0.switch_7.Z.n13 Vbias 1.0317f
C17853 CDAC8_0.switch_7.Z.t103 Vbias 5.57036f
C17854 CDAC8_0.switch_7.Z.n14 Vbias 1.29163f
C17855 CDAC8_0.switch_7.Z.n15 Vbias 1.0317f
C17856 CDAC8_0.switch_7.Z.t106 Vbias 5.57036f
C17857 CDAC8_0.switch_7.Z.n16 Vbias 1.43387f
C17858 CDAC8_0.switch_7.Z.t81 Vbias 5.57036f
C17859 CDAC8_0.switch_7.Z.n17 Vbias 1.63982f
C17860 CDAC8_0.switch_7.Z.n18 Vbias 1.0317f
C17861 CDAC8_0.switch_7.Z.t57 Vbias 5.57036f
C17862 CDAC8_0.switch_7.Z.n19 Vbias 1.29163f
C17863 CDAC8_0.switch_7.Z.n20 Vbias 0.84016f
C17864 CDAC8_0.switch_7.Z.t17 Vbias 5.57036f
C17865 CDAC8_0.switch_7.Z.n21 Vbias 1.29163f
C17866 CDAC8_0.switch_7.Z.n22 Vbias 0.84016f
C17867 CDAC8_0.switch_7.Z.t12 Vbias 5.57036f
C17868 CDAC8_0.switch_7.Z.n23 Vbias 1.29163f
C17869 CDAC8_0.switch_7.Z.n24 Vbias 0.84016f
C17870 CDAC8_0.switch_7.Z.t125 Vbias 5.57036f
C17871 CDAC8_0.switch_7.Z.n25 Vbias 1.29163f
C17872 CDAC8_0.switch_7.Z.n26 Vbias 0.84016f
C17873 CDAC8_0.switch_7.Z.t117 Vbias 5.65115f
C17874 CDAC8_0.switch_7.Z.t98 Vbias 5.65115f
C17875 CDAC8_0.switch_7.Z.t58 Vbias 5.57036f
C17876 CDAC8_0.switch_7.Z.n27 Vbias 1.29163f
C17877 CDAC8_0.switch_7.Z.n28 Vbias 1.0317f
C17878 CDAC8_0.switch_7.Z.t39 Vbias 5.57036f
C17879 CDAC8_0.switch_7.Z.n29 Vbias 1.29163f
C17880 CDAC8_0.switch_7.Z.n30 Vbias 1.0317f
C17881 CDAC8_0.switch_7.Z.t113 Vbias 5.57036f
C17882 CDAC8_0.switch_7.Z.n31 Vbias 1.29163f
C17883 CDAC8_0.switch_7.Z.n32 Vbias 1.0317f
C17884 CDAC8_0.switch_7.Z.t120 Vbias 5.57036f
C17885 CDAC8_0.switch_7.Z.n33 Vbias 1.29163f
C17886 CDAC8_0.switch_7.Z.n34 Vbias 1.0317f
C17887 CDAC8_0.switch_7.Z.t92 Vbias 5.57036f
C17888 CDAC8_0.switch_7.Z.n35 Vbias 1.29163f
C17889 CDAC8_0.switch_7.Z.n36 Vbias 2.08292f
C17890 CDAC8_0.switch_7.Z.t36 Vbias 5.65115f
C17891 CDAC8_0.switch_7.Z.n37 Vbias 0.60915f
C17892 CDAC8_0.switch_7.Z.t100 Vbias 5.57036f
C17893 CDAC8_0.switch_7.Z.n38 Vbias 1.29163f
C17894 CDAC8_0.switch_7.Z.n39 Vbias 0.60915f
C17895 CDAC8_0.switch_7.Z.t48 Vbias 5.57036f
C17896 CDAC8_0.switch_7.Z.n40 Vbias 1.29163f
C17897 CDAC8_0.switch_7.Z.n41 Vbias 0.60915f
C17898 CDAC8_0.switch_7.Z.t54 Vbias 5.57036f
C17899 CDAC8_0.switch_7.Z.n42 Vbias 1.29163f
C17900 CDAC8_0.switch_7.Z.n43 Vbias 0.60915f
C17901 CDAC8_0.switch_7.Z.t29 Vbias 5.57036f
C17902 CDAC8_0.switch_7.Z.n44 Vbias 1.29163f
C17903 CDAC8_0.switch_7.Z.n45 Vbias 1.66037f
C17904 CDAC8_0.switch_7.Z.n46 Vbias 0.84016f
C17905 CDAC8_0.switch_7.Z.t129 Vbias 5.65115f
C17906 CDAC8_0.switch_7.Z.n47 Vbias 2.08292f
C17907 CDAC8_0.switch_7.Z.n48 Vbias 0.84016f
C17908 CDAC8_0.switch_7.Z.n49 Vbias 1.66037f
C17909 CDAC8_0.switch_7.Z.t111 Vbias 5.57036f
C17910 CDAC8_0.switch_7.Z.n50 Vbias 1.29163f
C17911 CDAC8_0.switch_7.Z.n51 Vbias 0.60915f
C17912 CDAC8_0.switch_7.Z.n52 Vbias 0.84016f
C17913 CDAC8_0.switch_7.Z.n53 Vbias 1.0317f
C17914 CDAC8_0.switch_7.Z.t23 Vbias 5.57036f
C17915 CDAC8_0.switch_7.Z.n54 Vbias 1.29163f
C17916 CDAC8_0.switch_7.Z.n55 Vbias 1.0317f
C17917 CDAC8_0.switch_7.Z.n56 Vbias 0.84016f
C17918 CDAC8_0.switch_7.Z.n57 Vbias 0.60915f
C17919 CDAC8_0.switch_7.Z.t5 Vbias 5.57036f
C17920 CDAC8_0.switch_7.Z.n58 Vbias 1.29163f
C17921 CDAC8_0.switch_7.Z.n59 Vbias 0.60915f
C17922 CDAC8_0.switch_7.Z.n60 Vbias 0.84016f
C17923 CDAC8_0.switch_7.Z.n61 Vbias 1.0317f
C17924 CDAC8_0.switch_7.Z.t66 Vbias 5.57036f
C17925 CDAC8_0.switch_7.Z.n62 Vbias 1.29163f
C17926 CDAC8_0.switch_7.Z.t85 Vbias 5.57036f
C17927 CDAC8_0.switch_7.Z.n63 Vbias 1.29163f
C17928 CDAC8_0.switch_7.Z.n64 Vbias 1.0317f
C17929 CDAC8_0.switch_7.Z.n65 Vbias 0.84016f
C17930 CDAC8_0.switch_7.Z.n66 Vbias 0.60915f
C17931 CDAC8_0.switch_7.Z.t74 Vbias 5.57036f
C17932 CDAC8_0.switch_7.Z.n67 Vbias 1.29163f
C17933 CDAC8_0.switch_7.Z.n68 Vbias 0.60915f
C17934 CDAC8_0.switch_7.Z.n69 Vbias 0.84016f
C17935 CDAC8_0.switch_7.Z.n70 Vbias 0.84016f
C17936 CDAC8_0.switch_7.Z.n71 Vbias 0.60915f
C17937 CDAC8_0.switch_7.Z.t114 Vbias 5.57036f
C17938 CDAC8_0.switch_7.Z.n72 Vbias 1.29163f
C17939 CDAC8_0.switch_7.Z.n73 Vbias 0.60915f
C17940 CDAC8_0.switch_7.Z.n74 Vbias 0.87809f
C17941 CDAC8_0.switch_7.Z.n75 Vbias 1.0317f
C17942 CDAC8_0.switch_7.Z.t97 Vbias 5.57036f
C17943 CDAC8_0.switch_7.Z.n76 Vbias 1.29163f
C17944 CDAC8_0.switch_7.Z.n77 Vbias 0.60915f
C17945 CDAC8_0.switch_7.Z.t91 Vbias 5.57036f
C17946 CDAC8_0.switch_7.Z.n78 Vbias 1.29163f
C17947 CDAC8_0.switch_7.Z.t42 Vbias 5.57036f
C17948 CDAC8_0.switch_7.Z.n79 Vbias 1.29163f
C17949 CDAC8_0.switch_7.Z.n80 Vbias 0.84016f
C17950 CDAC8_0.switch_7.Z.t35 Vbias 5.57036f
C17951 CDAC8_0.switch_7.Z.n81 Vbias 1.29163f
C17952 CDAC8_0.switch_7.Z.t46 Vbias 5.57036f
C17953 CDAC8_0.switch_7.Z.n82 Vbias 1.29163f
C17954 CDAC8_0.switch_7.Z.n83 Vbias 0.84016f
C17955 CDAC8_0.switch_7.Z.t55 Vbias 5.57036f
C17956 CDAC8_0.switch_7.Z.n84 Vbias 1.29163f
C17957 CDAC8_0.switch_7.Z.n85 Vbias 0.84016f
C17958 CDAC8_0.switch_7.Z.t122 Vbias 5.57036f
C17959 CDAC8_0.switch_7.Z.n86 Vbias 1.29163f
C17960 CDAC8_0.switch_7.Z.n87 Vbias 0.84016f
C17961 CDAC8_0.switch_7.Z.t104 Vbias 5.57036f
C17962 CDAC8_0.switch_7.Z.n88 Vbias 1.29163f
C17963 CDAC8_0.switch_7.Z.n89 Vbias 0.84016f
C17964 CDAC8_0.switch_7.Z.t9 Vbias 5.79939f
C17965 CDAC8_0.switch_7.Z.n90 Vbias 0.71553f
C17966 CDAC8_0.switch_7.Z.t15 Vbias 5.57036f
C17967 CDAC8_0.switch_7.Z.n91 Vbias 1.29163f
C17968 CDAC8_0.switch_7.Z.n92 Vbias 0.84016f
C17969 CDAC8_0.switch_7.Z.t59 Vbias 5.57036f
C17970 CDAC8_0.switch_7.Z.n93 Vbias 1.29163f
C17971 CDAC8_0.switch_7.Z.t72 Vbias 5.57036f
C17972 CDAC8_0.switch_7.Z.n94 Vbias 1.29163f
C17973 CDAC8_0.switch_7.Z.n95 Vbias 0.84016f
C17974 CDAC8_0.switch_7.Z.t31 Vbias 5.57036f
C17975 CDAC8_0.switch_7.Z.n96 Vbias 1.29163f
C17976 CDAC8_0.switch_7.Z.n97 Vbias 0.84016f
C17977 CDAC8_0.switch_7.Z.t24 Vbias 5.57036f
C17978 CDAC8_0.switch_7.Z.n98 Vbias 1.29163f
C17979 CDAC8_0.switch_7.Z.n99 Vbias 0.84016f
C17980 CDAC8_0.switch_7.Z.t79 Vbias 5.57036f
C17981 CDAC8_0.switch_7.Z.n100 Vbias 1.29163f
C17982 CDAC8_0.switch_7.Z.n101 Vbias 0.84016f
C17983 CDAC8_0.switch_7.Z.t40 Vbias 5.79939f
C17984 CDAC8_0.switch_7.Z.t19 Vbias 5.79939f
C17985 CDAC8_0.switch_7.Z.n102 Vbias 2.24911f
C17986 CDAC8_0.switch_7.Z.t47 Vbias 5.57036f
C17987 CDAC8_0.switch_7.Z.n103 Vbias 1.29163f
C17988 CDAC8_0.switch_7.Z.t126 Vbias 5.57036f
C17989 CDAC8_0.switch_7.Z.n104 Vbias 1.29163f
C17990 CDAC8_0.switch_7.Z.n105 Vbias 1.0317f
C17991 CDAC8_0.switch_7.Z.t130 Vbias 5.57036f
C17992 CDAC8_0.switch_7.Z.n106 Vbias 1.29163f
C17993 CDAC8_0.switch_7.Z.n107 Vbias 1.0317f
C17994 CDAC8_0.switch_7.Z.t73 Vbias 5.57036f
C17995 CDAC8_0.switch_7.Z.n108 Vbias 1.29163f
C17996 CDAC8_0.switch_7.Z.n109 Vbias 1.0317f
C17997 CDAC8_0.switch_7.Z.t56 Vbias 5.57036f
C17998 CDAC8_0.switch_7.Z.n110 Vbias 1.29163f
C17999 CDAC8_0.switch_7.Z.n111 Vbias 1.0317f
C18000 CDAC8_0.switch_7.Z.t60 Vbias 5.57036f
C18001 CDAC8_0.switch_7.Z.n112 Vbias 1.29163f
C18002 CDAC8_0.switch_7.Z.n113 Vbias 1.0317f
C18003 CDAC8_0.switch_7.Z.t41 Vbias 5.57036f
C18004 CDAC8_0.switch_7.Z.n114 Vbias 1.29163f
C18005 CDAC8_0.switch_7.Z.n115 Vbias 1.0317f
C18006 CDAC8_0.switch_7.Z.t7 Vbias 5.57036f
C18007 CDAC8_0.switch_7.Z.n116 Vbias 1.29163f
C18008 CDAC8_0.switch_7.Z.t110 Vbias 5.57036f
C18009 CDAC8_0.switch_7.Z.n117 Vbias 1.29163f
C18010 CDAC8_0.switch_7.Z.n118 Vbias 1.0317f
C18011 CDAC8_0.switch_7.Z.t27 Vbias 5.57036f
C18012 CDAC8_0.switch_7.Z.n119 Vbias 1.29163f
C18013 CDAC8_0.switch_7.Z.t116 Vbias 5.57036f
C18014 CDAC8_0.switch_7.Z.n120 Vbias 1.29163f
C18015 CDAC8_0.switch_7.Z.n121 Vbias 1.0317f
C18016 CDAC8_0.switch_7.Z.n122 Vbias 0.71553f
C18017 CDAC8_0.switch_7.Z.t115 Vbias 5.57036f
C18018 CDAC8_0.switch_7.Z.n123 Vbias 1.29163f
C18019 CDAC8_0.switch_7.Z.n124 Vbias 0.84016f
C18020 CDAC8_0.switch_7.Z.t32 Vbias 5.57036f
C18021 CDAC8_0.switch_7.Z.n125 Vbias 1.29163f
C18022 CDAC8_0.switch_7.Z.n126 Vbias 0.84016f
C18023 CDAC8_0.switch_7.Z.t45 Vbias 5.57036f
C18024 CDAC8_0.switch_7.Z.n127 Vbias 1.29163f
C18025 CDAC8_0.switch_7.Z.n128 Vbias 0.84016f
C18026 CDAC8_0.switch_7.Z.t112 Vbias 5.57036f
C18027 CDAC8_0.switch_7.Z.n129 Vbias 1.29163f
C18028 CDAC8_0.switch_7.Z.n130 Vbias 0.84016f
C18029 CDAC8_0.switch_7.Z.t25 Vbias 5.57036f
C18030 CDAC8_0.switch_7.Z.n131 Vbias 1.29163f
C18031 CDAC8_0.switch_7.Z.n132 Vbias 0.84016f
C18032 CDAC8_0.switch_7.Z.t90 Vbias 5.65115f
C18033 CDAC8_0.switch_7.Z.t8 Vbias 5.65115f
C18034 CDAC8_0.switch_7.Z.t88 Vbias 5.57036f
C18035 CDAC8_0.switch_7.Z.n133 Vbias 1.29163f
C18036 CDAC8_0.switch_7.Z.n134 Vbias 1.0317f
C18037 CDAC8_0.switch_7.Z.t96 Vbias 5.57036f
C18038 CDAC8_0.switch_7.Z.n135 Vbias 1.29163f
C18039 CDAC8_0.switch_7.Z.n136 Vbias 1.0317f
C18040 CDAC8_0.switch_7.Z.t75 Vbias 5.57036f
C18041 CDAC8_0.switch_7.Z.n137 Vbias 1.29163f
C18042 CDAC8_0.switch_7.Z.n138 Vbias 1.0317f
C18043 CDAC8_0.switch_7.Z.t26 Vbias 5.57036f
C18044 CDAC8_0.switch_7.Z.n139 Vbias 1.29163f
C18045 CDAC8_0.switch_7.Z.n140 Vbias 1.0317f
C18046 CDAC8_0.switch_7.Z.t33 Vbias 5.57036f
C18047 CDAC8_0.switch_7.Z.n141 Vbias 1.29163f
C18048 CDAC8_0.switch_7.Z.n142 Vbias 1.0317f
C18049 CDAC8_0.switch_7.Z.t4 Vbias 5.57036f
C18050 CDAC8_0.switch_7.Z.n143 Vbias 1.29163f
C18051 CDAC8_0.switch_7.Z.n144 Vbias 2.08292f
C18052 CDAC8_0.switch_7.Z.t70 Vbias 5.65115f
C18053 CDAC8_0.switch_7.Z.n145 Vbias 0.60915f
C18054 CDAC8_0.switch_7.Z.t34 Vbias 5.57036f
C18055 CDAC8_0.switch_7.Z.n146 Vbias 1.29163f
C18056 CDAC8_0.switch_7.Z.n147 Vbias 0.60915f
C18057 CDAC8_0.switch_7.Z.t13 Vbias 5.57036f
C18058 CDAC8_0.switch_7.Z.n148 Vbias 1.29163f
C18059 CDAC8_0.switch_7.Z.n149 Vbias 0.60915f
C18060 CDAC8_0.switch_7.Z.t87 Vbias 5.57036f
C18061 CDAC8_0.switch_7.Z.n150 Vbias 1.29163f
C18062 CDAC8_0.switch_7.Z.n151 Vbias 0.60915f
C18063 CDAC8_0.switch_7.Z.t93 Vbias 5.57036f
C18064 CDAC8_0.switch_7.Z.n152 Vbias 1.29163f
C18065 CDAC8_0.switch_7.Z.n153 Vbias 0.60915f
C18066 CDAC8_0.switch_7.Z.t67 Vbias 5.57036f
C18067 CDAC8_0.switch_7.Z.n154 Vbias 1.29163f
C18068 CDAC8_0.switch_7.Z.n155 Vbias 1.66037f
C18069 CDAC8_0.switch_7.Z.n156 Vbias 0.84016f
C18070 CDAC8_0.switch_7.Z.t30 Vbias 5.65115f
C18071 CDAC8_0.switch_7.Z.n157 Vbias 1.66037f
C18072 CDAC8_0.switch_7.Z.n158 Vbias 0.84016f
C18073 CDAC8_0.switch_7.Z.n159 Vbias 2.08292f
C18074 CDAC8_0.switch_7.Z.t86 Vbias 5.57036f
C18075 CDAC8_0.switch_7.Z.n160 Vbias 1.29163f
C18076 CDAC8_0.switch_7.Z.n161 Vbias 1.0317f
C18077 CDAC8_0.switch_7.Z.n162 Vbias 0.84016f
C18078 CDAC8_0.switch_7.Z.n163 Vbias 0.60915f
C18079 CDAC8_0.switch_7.Z.t50 Vbias 5.57036f
C18080 CDAC8_0.switch_7.Z.n164 Vbias 1.29163f
C18081 CDAC8_0.switch_7.Z.n165 Vbias 0.60915f
C18082 CDAC8_0.switch_7.Z.n166 Vbias 0.84016f
C18083 CDAC8_0.switch_7.Z.n167 Vbias 1.0317f
C18084 CDAC8_0.switch_7.Z.t107 Vbias 5.57036f
C18085 CDAC8_0.switch_7.Z.n168 Vbias 1.29163f
C18086 CDAC8_0.switch_7.Z.n169 Vbias 1.0317f
C18087 CDAC8_0.switch_7.Z.n170 Vbias 0.84016f
C18088 CDAC8_0.switch_7.Z.n171 Vbias 0.60915f
C18089 CDAC8_0.switch_7.Z.t95 Vbias 5.57036f
C18090 CDAC8_0.switch_7.Z.n172 Vbias 1.29163f
C18091 CDAC8_0.switch_7.Z.n173 Vbias 0.60915f
C18092 CDAC8_0.switch_7.Z.n174 Vbias 0.84016f
C18093 CDAC8_0.switch_7.Z.n175 Vbias 1.0317f
C18094 CDAC8_0.switch_7.Z.t49 Vbias 5.57036f
C18095 CDAC8_0.switch_7.Z.n176 Vbias 1.29163f
C18096 CDAC8_0.switch_7.Z.t44 Vbias 5.57036f
C18097 CDAC8_0.switch_7.Z.n177 Vbias 1.29163f
C18098 CDAC8_0.switch_7.Z.n178 Vbias 1.0317f
C18099 CDAC8_0.switch_7.Z.n179 Vbias 0.84016f
C18100 CDAC8_0.switch_7.Z.n180 Vbias 0.60915f
C18101 CDAC8_0.switch_7.Z.t108 Vbias 5.57036f
C18102 CDAC8_0.switch_7.Z.n181 Vbias 1.29163f
C18103 CDAC8_0.switch_7.Z.n182 Vbias 0.60915f
C18104 CDAC8_0.switch_7.Z.n183 Vbias 0.84016f
C18105 CDAC8_0.switch_7.Z.n184 Vbias 0.84016f
C18106 CDAC8_0.switch_7.Z.n185 Vbias 0.60915f
C18107 CDAC8_0.switch_7.Z.t53 Vbias 5.57036f
C18108 CDAC8_0.switch_7.Z.n186 Vbias 1.29163f
C18109 CDAC8_0.switch_7.Z.n187 Vbias 0.60915f
C18110 CDAC8_0.switch_7.Z.n188 Vbias 0.84016f
C18111 CDAC8_0.switch_7.Z.t69 Vbias 5.57036f
C18112 CDAC8_0.switch_7.Z.n189 Vbias 1.17533f
C18113 CDAC8_0.switch_7.Z.t65 Vbias 5.57036f
C18114 CDAC8_0.switch_7.Z.n190 Vbias 1.29163f
C18115 CDAC8_0.switch_7.Z.n191 Vbias 1.0317f
C18116 CDAC8_0.switch_7.Z.n192 Vbias 0.84016f
C18117 CDAC8_0.switch_7.Z.n193 Vbias 0.60915f
C18118 CDAC8_0.switch_7.Z.t131 Vbias 5.57036f
C18119 CDAC8_0.switch_7.Z.n194 Vbias 1.29163f
C18120 CDAC8_0.switch_7.Z.n195 Vbias 0.60915f
C18121 CDAC8_0.switch_7.Z.n196 Vbias 0.84016f
C18122 CDAC8_0.switch_7.Z.n197 Vbias 0.84016f
C18123 CDAC8_0.switch_7.Z.n198 Vbias 0.60915f
C18124 CDAC8_0.switch_7.Z.t102 Vbias 5.57036f
C18125 CDAC8_0.switch_7.Z.n199 Vbias 1.29163f
C18126 CDAC8_0.switch_7.Z.n200 Vbias 0.60915f
C18127 CDAC8_0.switch_7.Z.t124 Vbias 5.57036f
C18128 CDAC8_0.switch_7.Z.n201 Vbias 1.29163f
C18129 CDAC8_0.switch_7.Z.n202 Vbias 0.60915f
C18130 CDAC8_0.switch_7.Z.t119 Vbias 5.57036f
C18131 CDAC8_0.switch_7.Z.n203 Vbias 1.29163f
C18132 CDAC8_0.switch_7.Z.n204 Vbias 0.60915f
C18133 CDAC8_0.switch_7.Z.t11 Vbias 5.57036f
C18134 CDAC8_0.switch_7.Z.n205 Vbias 1.29163f
C18135 CDAC8_0.switch_7.Z.n206 Vbias 0.60915f
C18136 CDAC8_0.switch_7.Z.t63 Vbias 5.57036f
C18137 CDAC8_0.switch_7.Z.n207 Vbias 1.29163f
C18138 CDAC8_0.switch_7.Z.n208 Vbias 0.60915f
C18139 CDAC8_0.switch_7.Z.t61 Vbias 5.57036f
C18140 CDAC8_0.switch_7.Z.n209 Vbias 1.29163f
C18141 CDAC8_0.switch_7.Z.t80 Vbias 5.79939f
C18142 CDAC8_0.switch_7.Z.n210 Vbias 1.82656f
C18143 CDAC8_0.switch_7.Z.n211 Vbias 0.84016f
C18144 CDAC8_0.switch_7.Z.t101 Vbias 5.79939f
C18145 CDAC8_0.switch_7.Z.n212 Vbias 2.24911f
C18146 CDAC8_0.switch_7.Z.n213 Vbias 0.84016f
C18147 CDAC8_0.switch_7.Z.n214 Vbias 1.82656f
C18148 CDAC8_0.switch_7.Z.t18 Vbias 5.57036f
C18149 CDAC8_0.switch_7.Z.n215 Vbias 1.29163f
C18150 CDAC8_0.switch_7.Z.n216 Vbias 0.60915f
C18151 CDAC8_0.switch_7.Z.n217 Vbias 0.84016f
C18152 CDAC8_0.switch_7.Z.n218 Vbias 1.0317f
C18153 CDAC8_0.switch_7.Z.t83 Vbias 5.57036f
C18154 CDAC8_0.switch_7.Z.n219 Vbias 1.29163f
C18155 CDAC8_0.switch_7.Z.n220 Vbias 1.0317f
C18156 CDAC8_0.switch_7.Z.n221 Vbias 0.84016f
C18157 CDAC8_0.switch_7.Z.n222 Vbias 0.60915f
C18158 CDAC8_0.switch_7.Z.t94 Vbias 5.57036f
C18159 CDAC8_0.switch_7.Z.n223 Vbias 1.29163f
C18160 CDAC8_0.switch_7.Z.n224 Vbias 0.60915f
C18161 CDAC8_0.switch_7.Z.n225 Vbias 0.84016f
C18162 CDAC8_0.switch_7.Z.n226 Vbias 1.0317f
C18163 CDAC8_0.switch_7.Z.t10 Vbias 5.57036f
C18164 CDAC8_0.switch_7.Z.n227 Vbias 1.29163f
C18165 CDAC8_0.switch_7.Z.n228 Vbias 1.0317f
C18166 CDAC8_0.switch_7.Z.n229 Vbias 0.84016f
C18167 CDAC8_0.switch_7.Z.n230 Vbias 0.60915f
C18168 CDAC8_0.switch_7.Z.t78 Vbias 5.57036f
C18169 CDAC8_0.switch_7.Z.n231 Vbias 1.29163f
C18170 CDAC8_0.switch_7.Z.n232 Vbias 0.60915f
C18171 CDAC8_0.switch_7.Z.n233 Vbias 0.84016f
C18172 CDAC8_0.switch_7.Z.n234 Vbias 1.0317f
C18173 CDAC8_0.switch_7.Z.t123 Vbias 5.57036f
C18174 CDAC8_0.switch_7.Z.n235 Vbias 1.17533f
C18175 CDAC8_0.switch_7.Z.n236 Vbias 3.78864f
C18176 CDAC8_0.switch_7.Z.n237 Vbias 3.78864f
C18177 CDAC8_0.switch_7.Z.t128 Vbias 5.57036f
C18178 CDAC8_0.switch_7.Z.n238 Vbias 1.17533f
C18179 CDAC8_0.switch_7.Z.n239 Vbias 1.0317f
C18180 CDAC8_0.switch_7.Z.t21 Vbias 5.57036f
C18181 CDAC8_0.switch_7.Z.n240 Vbias 1.29163f
C18182 CDAC8_0.switch_7.Z.n241 Vbias 1.0317f
C18183 CDAC8_0.switch_7.Z.t16 Vbias 5.57036f
C18184 CDAC8_0.switch_7.Z.n242 Vbias 1.29163f
C18185 CDAC8_0.switch_7.Z.n243 Vbias 1.0317f
C18186 CDAC8_0.switch_7.Z.t38 Vbias 5.57036f
C18187 CDAC8_0.switch_7.Z.n244 Vbias 1.29163f
C18188 CDAC8_0.switch_7.Z.n245 Vbias 1.0317f
C18189 CDAC8_0.switch_7.Z.t89 Vbias 5.57036f
C18190 CDAC8_0.switch_7.Z.n246 Vbias 1.29163f
C18191 CDAC8_0.switch_7.Z.n247 Vbias 1.0317f
C18192 CDAC8_0.switch_7.Z.t84 Vbias 5.57036f
C18193 CDAC8_0.switch_7.Z.n248 Vbias 1.29163f
C18194 CDAC8_0.switch_7.Z.t105 Vbias 5.79939f
C18195 CDAC8_0.switch_7.Z.n249 Vbias 2.24911f
C18196 CDAC8_0.switch_7.Z.n250 Vbias 0.60915f
C18197 CDAC8_0.switch_7.Z.t82 Vbias 5.57036f
C18198 CDAC8_0.switch_7.Z.n251 Vbias 1.29163f
C18199 CDAC8_0.switch_7.Z.n252 Vbias 0.60915f
C18200 CDAC8_0.switch_7.Z.t77 Vbias 5.57036f
C18201 CDAC8_0.switch_7.Z.n253 Vbias 1.29163f
C18202 CDAC8_0.switch_7.Z.n254 Vbias 0.60915f
C18203 CDAC8_0.switch_7.Z.t99 Vbias 5.57036f
C18204 CDAC8_0.switch_7.Z.n255 Vbias 1.29163f
C18205 CDAC8_0.switch_7.Z.n256 Vbias 0.60915f
C18206 CDAC8_0.switch_7.Z.t28 Vbias 5.57036f
C18207 CDAC8_0.switch_7.Z.n257 Vbias 1.29163f
C18208 CDAC8_0.switch_7.Z.n258 Vbias 0.60915f
C18209 CDAC8_0.switch_7.Z.t22 Vbias 5.57036f
C18210 CDAC8_0.switch_7.Z.n259 Vbias 1.29163f
C18211 CDAC8_0.switch_7.Z.t43 Vbias 5.79939f
C18212 CDAC8_0.switch_7.Z.n260 Vbias 1.82656f
C18213 CDAC8_0.switch_7.Z.n261 Vbias 0.84016f
C18214 CDAC8_0.switch_7.Z.t127 Vbias 5.79939f
C18215 CDAC8_0.switch_7.Z.n262 Vbias 1.82656f
C18216 CDAC8_0.switch_7.Z.n263 Vbias 0.84016f
C18217 CDAC8_0.switch_7.Z.n264 Vbias 2.24911f
C18218 CDAC8_0.switch_7.Z.t118 Vbias 5.57036f
C18219 CDAC8_0.switch_7.Z.n265 Vbias 1.29163f
C18220 CDAC8_0.switch_7.Z.n266 Vbias 1.0317f
C18221 CDAC8_0.switch_7.Z.n267 Vbias 0.84016f
C18222 CDAC8_0.switch_7.Z.n268 Vbias 0.60915f
C18223 CDAC8_0.switch_7.Z.t109 Vbias 5.57036f
C18224 CDAC8_0.switch_7.Z.n269 Vbias 1.29163f
C18225 CDAC8_0.switch_7.Z.n270 Vbias 0.60915f
C18226 CDAC8_0.switch_7.Z.n271 Vbias 0.84016f
C18227 CDAC8_0.switch_7.Z.n272 Vbias 1.0317f
C18228 CDAC8_0.switch_7.Z.t64 Vbias 5.57036f
C18229 CDAC8_0.switch_7.Z.n273 Vbias 1.29163f
C18230 CDAC8_0.switch_7.Z.n274 Vbias 1.0317f
C18231 CDAC8_0.switch_7.Z.n275 Vbias 0.84016f
C18232 CDAC8_0.switch_7.Z.n276 Vbias 0.60915f
C18233 CDAC8_0.switch_7.Z.t37 Vbias 5.57036f
C18234 CDAC8_0.switch_7.Z.n277 Vbias 1.29163f
C18235 CDAC8_0.switch_7.Z.n278 Vbias 0.60915f
C18236 CDAC8_0.switch_7.Z.n279 Vbias 0.84016f
C18237 CDAC8_0.switch_7.Z.n280 Vbias 1.0317f
C18238 CDAC8_0.switch_7.Z.t52 Vbias 5.57036f
C18239 CDAC8_0.switch_7.Z.n281 Vbias 1.29163f
C18240 CDAC8_0.switch_7.Z.n282 Vbias 1.0317f
C18241 CDAC8_0.switch_7.Z.n283 Vbias 0.84016f
C18242 CDAC8_0.switch_7.Z.n284 Vbias 0.60915f
C18243 CDAC8_0.switch_7.Z.t20 Vbias 5.57036f
C18244 CDAC8_0.switch_7.Z.n285 Vbias 1.29163f
C18245 CDAC8_0.switch_7.Z.n286 Vbias 0.60915f
C18246 CDAC8_0.switch_7.Z.n287 Vbias 0.84016f
C18247 CDAC8_0.switch_7.Z.n288 Vbias 0.84016f
C18248 CDAC8_0.switch_7.Z.n289 Vbias 0.60915f
C18249 CDAC8_0.switch_7.Z.t6 Vbias 5.57036f
C18250 CDAC8_0.switch_7.Z.n290 Vbias 1.29163f
C18251 CDAC8_0.switch_7.Z.n291 Vbias 0.60915f
C18252 CDAC8_0.switch_7.Z.n292 Vbias 0.84016f
C18253 CDAC8_0.switch_7.Z.n293 Vbias 1.0317f
C18254 CDAC8_0.switch_7.Z.t76 Vbias 5.57036f
C18255 CDAC8_0.switch_7.Z.n294 Vbias 1.17533f
C18256 CDAC8_0.switch_7.Z.n295 Vbias 2.11553f
C18257 CDAC8_0.switch_7.Z.n296 Vbias 3.35902f
C18258 CDAC8_0.switch_7.Z.n297 Vbias 0.13266f
C18259 CDAC8_0.switch_7.Z.t2 Vbias 0.03308f
.ends

