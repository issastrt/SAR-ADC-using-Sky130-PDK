magic
tech sky130A
magscale 1 2
timestamp 1755875457
<< metal1 >>
rect 11040 40339 97170 40385
rect 19709 39536 19773 39542
rect 19709 39484 19715 39536
rect 19767 39484 19773 39536
rect 19709 39478 19773 39484
rect 22508 39536 22572 39542
rect 22508 39484 22514 39536
rect 22566 39484 22572 39536
rect 22508 39478 22572 39484
rect 30749 39536 30813 39542
rect 30749 39484 30755 39536
rect 30807 39484 30813 39536
rect 30749 39478 30813 39484
rect 33548 39536 33612 39542
rect 33548 39484 33554 39536
rect 33606 39484 33612 39536
rect 33548 39478 33612 39484
rect 41789 39536 41853 39542
rect 41789 39484 41795 39536
rect 41847 39484 41853 39536
rect 41789 39478 41853 39484
rect 44588 39536 44652 39542
rect 44588 39484 44594 39536
rect 44646 39484 44652 39536
rect 44588 39478 44652 39484
rect 52829 39536 52893 39542
rect 52829 39484 52835 39536
rect 52887 39484 52893 39536
rect 52829 39478 52893 39484
rect 55628 39536 55692 39542
rect 55628 39484 55634 39536
rect 55686 39484 55692 39536
rect 55628 39478 55692 39484
rect 63869 39536 63933 39542
rect 63869 39484 63875 39536
rect 63927 39484 63933 39536
rect 63869 39478 63933 39484
rect 66668 39536 66732 39542
rect 66668 39484 66674 39536
rect 66726 39484 66732 39536
rect 66668 39478 66732 39484
rect 74909 39536 74973 39542
rect 74909 39484 74915 39536
rect 74967 39484 74973 39536
rect 74909 39478 74973 39484
rect 77708 39536 77772 39542
rect 77708 39484 77714 39536
rect 77766 39484 77772 39536
rect 77708 39478 77772 39484
rect 85949 39536 86013 39542
rect 85949 39484 85955 39536
rect 86007 39484 86013 39536
rect 85949 39478 86013 39484
rect 88748 39536 88812 39542
rect 88748 39484 88754 39536
rect 88806 39484 88812 39536
rect 88748 39478 88812 39484
rect 87549 38606 87613 38612
rect 87549 38603 87555 38606
rect 11128 38557 87555 38603
rect 87549 38554 87555 38557
rect 87607 38603 87613 38606
rect 87607 38557 97170 38603
rect 87607 38554 87613 38557
rect 87549 38548 87613 38554
rect 96766 37050 96830 37056
rect 96766 36998 96772 37050
rect 96824 36998 96830 37050
rect 96766 36992 96830 36998
rect 86765 36824 86829 36830
rect 86765 36821 86771 36824
rect 11040 36775 86771 36821
rect 86765 36772 86771 36775
rect 86823 36821 86829 36824
rect 86823 36775 97170 36821
rect 86823 36772 86829 36775
rect 86765 36766 86829 36772
rect 86765 3613 86829 3619
rect 86765 3610 86771 3613
rect 88 3564 86771 3610
rect 86765 3561 86771 3564
rect 86823 3610 86829 3613
rect 86823 3564 97198 3610
rect 86823 3561 86829 3564
rect 86765 3555 86829 3561
rect 1656 3387 1720 3393
rect 1656 3335 1662 3387
rect 1714 3335 1720 3387
rect 1656 3329 1720 3335
rect 12696 3387 12760 3393
rect 12696 3335 12702 3387
rect 12754 3335 12760 3387
rect 12696 3329 12760 3335
rect 23736 3387 23800 3393
rect 23736 3335 23742 3387
rect 23794 3335 23800 3387
rect 23736 3329 23800 3335
rect 34776 3387 34840 3393
rect 34776 3335 34782 3387
rect 34834 3335 34840 3387
rect 34776 3329 34840 3335
rect 45816 3387 45880 3393
rect 45816 3335 45822 3387
rect 45874 3335 45880 3387
rect 45816 3329 45880 3335
rect 56856 3387 56920 3393
rect 56856 3335 56862 3387
rect 56914 3335 56920 3387
rect 56856 3329 56920 3335
rect 67896 3387 67960 3393
rect 67896 3335 67902 3387
rect 67954 3335 67960 3387
rect 67896 3329 67960 3335
rect 78936 3387 79000 3393
rect 78936 3335 78942 3387
rect 78994 3335 79000 3387
rect 78936 3329 79000 3335
rect 89976 3387 90040 3393
rect 89976 3335 89982 3387
rect 90034 3335 90040 3387
rect 89976 3329 90040 3335
rect 96766 3387 96830 3393
rect 96766 3335 96772 3387
rect 96824 3335 96830 3387
rect 96766 3329 96830 3335
rect 8446 2761 8510 2767
rect 8446 2709 8452 2761
rect 8504 2709 8510 2761
rect 8446 2703 8510 2709
rect 11245 2761 11309 2767
rect 11245 2709 11251 2761
rect 11303 2709 11309 2761
rect 11245 2703 11309 2709
rect 19486 2761 19550 2767
rect 19486 2709 19492 2761
rect 19544 2709 19550 2761
rect 19486 2703 19550 2709
rect 22285 2761 22349 2767
rect 22285 2709 22291 2761
rect 22343 2709 22349 2761
rect 22285 2703 22349 2709
rect 30526 2761 30590 2767
rect 30526 2709 30532 2761
rect 30584 2709 30590 2761
rect 30526 2703 30590 2709
rect 33325 2761 33389 2767
rect 33325 2709 33331 2761
rect 33383 2709 33389 2761
rect 33325 2703 33389 2709
rect 41566 2761 41630 2767
rect 41566 2709 41572 2761
rect 41624 2709 41630 2761
rect 41566 2703 41630 2709
rect 44365 2761 44429 2767
rect 44365 2709 44371 2761
rect 44423 2709 44429 2761
rect 44365 2703 44429 2709
rect 52606 2761 52670 2767
rect 52606 2709 52612 2761
rect 52664 2709 52670 2761
rect 52606 2703 52670 2709
rect 55405 2761 55469 2767
rect 55405 2709 55411 2761
rect 55463 2709 55469 2761
rect 55405 2703 55469 2709
rect 63646 2761 63710 2767
rect 63646 2709 63652 2761
rect 63704 2709 63710 2761
rect 63646 2703 63710 2709
rect 66445 2761 66509 2767
rect 66445 2709 66451 2761
rect 66503 2709 66509 2761
rect 66445 2703 66509 2709
rect 74686 2761 74750 2767
rect 74686 2709 74692 2761
rect 74744 2709 74750 2761
rect 74686 2703 74750 2709
rect 77485 2761 77549 2767
rect 77485 2709 77491 2761
rect 77543 2709 77549 2761
rect 77485 2703 77549 2709
rect 85726 2761 85790 2767
rect 85726 2709 85732 2761
rect 85784 2709 85790 2761
rect 85726 2703 85790 2709
rect 88525 2761 88589 2767
rect 88525 2709 88531 2761
rect 88583 2709 88589 2761
rect 88525 2703 88589 2709
rect 5730 1831 5794 1837
rect 5730 1828 5736 1831
rect 88 1782 5736 1828
rect 5730 1779 5736 1782
rect 5788 1828 5794 1831
rect 16770 1831 16834 1837
rect 16770 1828 16776 1831
rect 5788 1782 16776 1828
rect 5788 1779 5794 1782
rect 5730 1773 5794 1779
rect 16770 1779 16776 1782
rect 16828 1828 16834 1831
rect 27810 1831 27874 1837
rect 27810 1828 27816 1831
rect 16828 1782 27816 1828
rect 16828 1779 16834 1782
rect 16770 1773 16834 1779
rect 27810 1779 27816 1782
rect 27868 1828 27874 1831
rect 38850 1831 38914 1837
rect 38850 1828 38856 1831
rect 27868 1782 38856 1828
rect 27868 1779 27874 1782
rect 27810 1773 27874 1779
rect 38850 1779 38856 1782
rect 38908 1828 38914 1831
rect 49890 1831 49954 1837
rect 49890 1828 49896 1831
rect 38908 1782 49896 1828
rect 38908 1779 38914 1782
rect 38850 1773 38914 1779
rect 49890 1779 49896 1782
rect 49948 1828 49954 1831
rect 60930 1831 60994 1837
rect 60930 1828 60936 1831
rect 49948 1782 60936 1828
rect 49948 1779 49954 1782
rect 49890 1773 49954 1779
rect 60930 1779 60936 1782
rect 60988 1828 60994 1831
rect 71970 1831 72034 1837
rect 71970 1828 71976 1831
rect 60988 1782 71976 1828
rect 60988 1779 60994 1782
rect 60930 1773 60994 1779
rect 71970 1779 71976 1782
rect 72028 1828 72034 1831
rect 83010 1831 83074 1837
rect 83010 1828 83016 1831
rect 72028 1782 83016 1828
rect 72028 1779 72034 1782
rect 71970 1773 72034 1779
rect 83010 1779 83016 1782
rect 83068 1828 83074 1831
rect 87549 1831 87613 1837
rect 87549 1828 87555 1831
rect 83068 1782 87555 1828
rect 83068 1779 83074 1782
rect 83010 1773 83074 1779
rect 87549 1779 87555 1782
rect 87607 1828 87613 1831
rect 94050 1831 94114 1837
rect 94050 1828 94056 1831
rect 87607 1782 94056 1828
rect 87607 1779 87613 1782
rect 87549 1773 87613 1779
rect 94050 1779 94056 1782
rect 94108 1828 94114 1831
rect 94108 1782 97170 1828
rect 94108 1779 94114 1782
rect 94050 1773 94114 1779
rect 5730 1575 5794 1581
rect 5730 1523 5736 1575
rect 5788 1523 5794 1575
rect 5730 1517 5794 1523
rect 16770 1575 16834 1581
rect 16770 1523 16776 1575
rect 16828 1523 16834 1575
rect 16770 1517 16834 1523
rect 27810 1575 27874 1581
rect 27810 1523 27816 1575
rect 27868 1523 27874 1575
rect 27810 1517 27874 1523
rect 38850 1575 38914 1581
rect 38850 1523 38856 1575
rect 38908 1523 38914 1575
rect 38850 1517 38914 1523
rect 49890 1575 49954 1581
rect 49890 1523 49896 1575
rect 49948 1523 49954 1575
rect 49890 1517 49954 1523
rect 60930 1575 60994 1581
rect 60930 1523 60936 1575
rect 60988 1523 60994 1575
rect 60930 1517 60994 1523
rect 71970 1575 72034 1581
rect 71970 1523 71976 1575
rect 72028 1523 72034 1575
rect 71970 1517 72034 1523
rect 83010 1575 83074 1581
rect 83010 1523 83016 1575
rect 83068 1523 83074 1575
rect 83010 1517 83074 1523
rect 94050 1575 94114 1581
rect 94050 1523 94056 1575
rect 94108 1523 94114 1575
rect 94050 1517 94114 1523
rect 88 0 97198 46
<< via1 >>
rect 19715 39484 19767 39536
rect 22514 39484 22566 39536
rect 30755 39484 30807 39536
rect 33554 39484 33606 39536
rect 41795 39484 41847 39536
rect 44594 39484 44646 39536
rect 52835 39484 52887 39536
rect 55634 39484 55686 39536
rect 63875 39484 63927 39536
rect 66674 39484 66726 39536
rect 74915 39484 74967 39536
rect 77714 39484 77766 39536
rect 85955 39484 86007 39536
rect 88754 39484 88806 39536
rect 87555 38554 87607 38606
rect 96772 36998 96824 37050
rect 86771 36772 86823 36824
rect 86771 3561 86823 3613
rect 1662 3335 1714 3387
rect 12702 3335 12754 3387
rect 23742 3335 23794 3387
rect 34782 3335 34834 3387
rect 45822 3335 45874 3387
rect 56862 3335 56914 3387
rect 67902 3335 67954 3387
rect 78942 3335 78994 3387
rect 89982 3335 90034 3387
rect 96772 3335 96824 3387
rect 8452 2709 8504 2761
rect 11251 2709 11303 2761
rect 19492 2709 19544 2761
rect 22291 2709 22343 2761
rect 30532 2709 30584 2761
rect 33331 2709 33383 2761
rect 41572 2709 41624 2761
rect 44371 2709 44423 2761
rect 52612 2709 52664 2761
rect 55411 2709 55463 2761
rect 63652 2709 63704 2761
rect 66451 2709 66503 2761
rect 74692 2709 74744 2761
rect 77491 2709 77543 2761
rect 85732 2709 85784 2761
rect 88531 2709 88583 2761
rect 5736 1779 5788 1831
rect 16776 1779 16828 1831
rect 27816 1779 27868 1831
rect 38856 1779 38908 1831
rect 49896 1779 49948 1831
rect 60936 1779 60988 1831
rect 71976 1779 72028 1831
rect 83016 1779 83068 1831
rect 87555 1779 87607 1831
rect 94056 1779 94108 1831
rect 5736 1523 5788 1575
rect 16776 1523 16828 1575
rect 27816 1523 27868 1575
rect 38856 1523 38908 1575
rect 49896 1523 49948 1575
rect 60936 1523 60988 1575
rect 71976 1523 72028 1575
rect 83016 1523 83068 1575
rect 94056 1523 94108 1575
<< metal2 >>
rect 322 39538 396 39547
rect 322 39482 331 39538
rect 387 39533 396 39538
rect 19709 39536 19773 39542
rect 387 39487 11523 39533
rect 387 39482 396 39487
rect 322 39473 396 39482
rect 19709 39484 19715 39536
rect 19767 39533 19773 39536
rect 22508 39536 22572 39542
rect 22508 39533 22514 39536
rect 19767 39487 22514 39533
rect 19767 39484 19773 39487
rect 19709 39478 19773 39484
rect 22508 39484 22514 39487
rect 22566 39484 22572 39536
rect 22508 39478 22572 39484
rect 30749 39536 30813 39542
rect 30749 39484 30755 39536
rect 30807 39533 30813 39536
rect 33548 39536 33612 39542
rect 33548 39533 33554 39536
rect 30807 39487 33554 39533
rect 30807 39484 30813 39487
rect 30749 39478 30813 39484
rect 33548 39484 33554 39487
rect 33606 39484 33612 39536
rect 33548 39478 33612 39484
rect 41789 39536 41853 39542
rect 41789 39484 41795 39536
rect 41847 39533 41853 39536
rect 44588 39536 44652 39542
rect 44588 39533 44594 39536
rect 41847 39487 44594 39533
rect 41847 39484 41853 39487
rect 41789 39478 41853 39484
rect 44588 39484 44594 39487
rect 44646 39484 44652 39536
rect 44588 39478 44652 39484
rect 52829 39536 52893 39542
rect 52829 39484 52835 39536
rect 52887 39533 52893 39536
rect 55628 39536 55692 39542
rect 55628 39533 55634 39536
rect 52887 39487 55634 39533
rect 52887 39484 52893 39487
rect 52829 39478 52893 39484
rect 55628 39484 55634 39487
rect 55686 39484 55692 39536
rect 55628 39478 55692 39484
rect 63869 39536 63933 39542
rect 63869 39484 63875 39536
rect 63927 39533 63933 39536
rect 66668 39536 66732 39542
rect 66668 39533 66674 39536
rect 63927 39487 66674 39533
rect 63927 39484 63933 39487
rect 63869 39478 63933 39484
rect 66668 39484 66674 39487
rect 66726 39484 66732 39536
rect 66668 39478 66732 39484
rect 74909 39536 74973 39542
rect 74909 39484 74915 39536
rect 74967 39533 74973 39536
rect 77708 39536 77772 39542
rect 77708 39533 77714 39536
rect 74967 39487 77714 39533
rect 74967 39484 74973 39487
rect 74909 39478 74973 39484
rect 77708 39484 77714 39487
rect 77766 39484 77772 39536
rect 77708 39478 77772 39484
rect 85949 39536 86013 39542
rect 85949 39484 85955 39536
rect 86007 39533 86013 39536
rect 88748 39536 88812 39542
rect 88748 39533 88754 39536
rect 86007 39487 88754 39533
rect 86007 39484 86013 39487
rect 85949 39478 86013 39484
rect 88748 39484 88754 39487
rect 88806 39484 88812 39536
rect 88748 39478 88812 39484
rect 16765 39418 16839 39427
rect 16765 39362 16774 39418
rect 16830 39362 16839 39418
rect 16765 39353 16839 39362
rect 23731 39418 23805 39427
rect 23731 39362 23740 39418
rect 23796 39362 23805 39418
rect 23731 39353 23805 39362
rect 34771 39418 34845 39427
rect 34771 39362 34780 39418
rect 34836 39362 34845 39418
rect 34771 39353 34845 39362
rect 45811 39418 45885 39427
rect 45811 39362 45820 39418
rect 45876 39362 45885 39418
rect 45811 39353 45885 39362
rect 56851 39418 56925 39427
rect 56851 39362 56860 39418
rect 56916 39362 56925 39418
rect 56851 39353 56925 39362
rect 67891 39418 67965 39427
rect 67891 39362 67900 39418
rect 67956 39362 67965 39418
rect 67891 39353 67965 39362
rect 78931 39418 79005 39427
rect 78931 39362 78940 39418
rect 78996 39362 79005 39418
rect 78931 39353 79005 39362
rect 89971 39418 90045 39427
rect 89971 39362 89980 39418
rect 90036 39362 90045 39418
rect 89971 39353 90045 39362
rect 87544 38608 87618 38617
rect 87544 38552 87553 38608
rect 87609 38552 87618 38608
rect 87544 38543 87618 38552
rect 12691 37798 12765 37807
rect 12691 37742 12700 37798
rect 12756 37742 12765 37798
rect 12691 37733 12765 37742
rect 27805 37798 27879 37807
rect 27805 37742 27814 37798
rect 27870 37742 27879 37798
rect 27805 37733 27879 37742
rect 38845 37798 38919 37807
rect 38845 37742 38854 37798
rect 38910 37742 38919 37798
rect 38845 37733 38919 37742
rect 49885 37798 49959 37807
rect 49885 37742 49894 37798
rect 49950 37742 49959 37798
rect 49885 37733 49959 37742
rect 60925 37798 60999 37807
rect 60925 37742 60934 37798
rect 60990 37742 60999 37798
rect 60925 37733 60999 37742
rect 71965 37798 72039 37807
rect 71965 37742 71974 37798
rect 72030 37742 72039 37798
rect 71965 37733 72039 37742
rect 83005 37798 83079 37807
rect 83005 37742 83014 37798
rect 83070 37742 83079 37798
rect 83005 37733 83079 37742
rect 94045 37798 94119 37807
rect 94045 37742 94054 37798
rect 94110 37742 94119 37798
rect 94045 37733 94119 37742
rect 96761 37052 96835 37061
rect 96761 36996 96770 37052
rect 96826 36996 96835 37052
rect 96761 36987 96835 36996
rect 86760 36826 86834 36835
rect 86760 36770 86769 36826
rect 86825 36770 86834 36826
rect 86760 36761 86834 36770
rect 16765 36734 16839 36743
rect 16765 36678 16774 36734
rect 16830 36729 16839 36734
rect 27805 36734 27879 36743
rect 27805 36729 27814 36734
rect 16830 36683 27814 36729
rect 16830 36678 16839 36683
rect 16765 36669 16839 36678
rect 27805 36678 27814 36683
rect 27870 36729 27879 36734
rect 38845 36734 38919 36743
rect 38845 36729 38854 36734
rect 27870 36683 38854 36729
rect 27870 36678 27879 36683
rect 27805 36669 27879 36678
rect 38845 36678 38854 36683
rect 38910 36729 38919 36734
rect 49885 36734 49959 36743
rect 49885 36729 49894 36734
rect 38910 36683 49894 36729
rect 38910 36678 38919 36683
rect 38845 36669 38919 36678
rect 49885 36678 49894 36683
rect 49950 36729 49959 36734
rect 60925 36734 60999 36743
rect 60925 36729 60934 36734
rect 49950 36683 60934 36729
rect 49950 36678 49959 36683
rect 49885 36669 49959 36678
rect 60925 36678 60934 36683
rect 60990 36729 60999 36734
rect 71965 36734 72039 36743
rect 71965 36729 71974 36734
rect 60990 36683 71974 36729
rect 60990 36678 60999 36683
rect 60925 36669 60999 36678
rect 71965 36678 71974 36683
rect 72030 36729 72039 36734
rect 83005 36734 83079 36743
rect 83005 36729 83014 36734
rect 72030 36683 83014 36729
rect 72030 36678 72039 36683
rect 71965 36669 72039 36678
rect 83005 36678 83014 36683
rect 83070 36729 83079 36734
rect 94045 36734 94119 36743
rect 94045 36729 94054 36734
rect 83070 36683 94054 36729
rect 83070 36678 83079 36683
rect 83005 36669 83079 36678
rect 94045 36678 94054 36683
rect 94110 36678 94119 36734
rect 94045 36669 94119 36678
rect 12691 36642 12765 36651
rect 12691 36586 12700 36642
rect 12756 36637 12765 36642
rect 23731 36642 23805 36651
rect 23731 36637 23740 36642
rect 12756 36591 23740 36637
rect 12756 36586 12765 36591
rect 12691 36577 12765 36586
rect 23731 36586 23740 36591
rect 23796 36637 23805 36642
rect 34771 36642 34845 36651
rect 34771 36637 34780 36642
rect 23796 36591 34780 36637
rect 23796 36586 23805 36591
rect 23731 36577 23805 36586
rect 34771 36586 34780 36591
rect 34836 36637 34845 36642
rect 45811 36642 45885 36651
rect 45811 36637 45820 36642
rect 34836 36591 45820 36637
rect 34836 36586 34845 36591
rect 34771 36577 34845 36586
rect 45811 36586 45820 36591
rect 45876 36637 45885 36642
rect 56851 36642 56925 36651
rect 56851 36637 56860 36642
rect 45876 36591 56860 36637
rect 45876 36586 45885 36591
rect 45811 36577 45885 36586
rect 56851 36586 56860 36591
rect 56916 36637 56925 36642
rect 67891 36642 67965 36651
rect 67891 36637 67900 36642
rect 56916 36591 67900 36637
rect 56916 36586 56925 36591
rect 56851 36577 56925 36586
rect 67891 36586 67900 36591
rect 67956 36637 67965 36642
rect 78931 36642 79005 36651
rect 78931 36637 78940 36642
rect 67956 36591 78940 36637
rect 67956 36586 67965 36591
rect 67891 36577 67965 36586
rect 78931 36586 78940 36591
rect 78996 36637 79005 36642
rect 89971 36642 90045 36651
rect 89971 36637 89980 36642
rect 78996 36591 89980 36637
rect 78996 36586 79005 36591
rect 78931 36577 79005 36586
rect 89971 36586 89980 36591
rect 90036 36586 90045 36642
rect 89971 36577 90045 36586
rect 1651 3799 1725 3808
rect 1651 3743 1660 3799
rect 1716 3794 1725 3799
rect 12691 3799 12765 3808
rect 12691 3794 12700 3799
rect 1716 3748 12700 3794
rect 1716 3743 1725 3748
rect 1651 3734 1725 3743
rect 12691 3743 12700 3748
rect 12756 3794 12765 3799
rect 23731 3799 23805 3808
rect 23731 3794 23740 3799
rect 12756 3748 23740 3794
rect 12756 3743 12765 3748
rect 12691 3734 12765 3743
rect 23731 3743 23740 3748
rect 23796 3794 23805 3799
rect 34771 3799 34845 3808
rect 34771 3794 34780 3799
rect 23796 3748 34780 3794
rect 23796 3743 23805 3748
rect 23731 3734 23805 3743
rect 34771 3743 34780 3748
rect 34836 3794 34845 3799
rect 45811 3799 45885 3808
rect 45811 3794 45820 3799
rect 34836 3748 45820 3794
rect 34836 3743 34845 3748
rect 34771 3734 34845 3743
rect 45811 3743 45820 3748
rect 45876 3794 45885 3799
rect 56851 3799 56925 3808
rect 56851 3794 56860 3799
rect 45876 3748 56860 3794
rect 45876 3743 45885 3748
rect 45811 3734 45885 3743
rect 56851 3743 56860 3748
rect 56916 3794 56925 3799
rect 67891 3799 67965 3808
rect 67891 3794 67900 3799
rect 56916 3748 67900 3794
rect 56916 3743 56925 3748
rect 56851 3734 56925 3743
rect 67891 3743 67900 3748
rect 67956 3794 67965 3799
rect 78931 3799 79005 3808
rect 78931 3794 78940 3799
rect 67956 3748 78940 3794
rect 67956 3743 67965 3748
rect 67891 3734 67965 3743
rect 78931 3743 78940 3748
rect 78996 3794 79005 3799
rect 89971 3799 90045 3808
rect 89971 3794 89980 3799
rect 78996 3748 89980 3794
rect 78996 3743 79005 3748
rect 78931 3734 79005 3743
rect 89971 3743 89980 3748
rect 90036 3743 90045 3799
rect 89971 3734 90045 3743
rect 5725 3707 5799 3716
rect 5725 3651 5734 3707
rect 5790 3702 5799 3707
rect 16765 3707 16839 3716
rect 16765 3702 16774 3707
rect 5790 3656 16774 3702
rect 5790 3651 5799 3656
rect 5725 3642 5799 3651
rect 16765 3651 16774 3656
rect 16830 3702 16839 3707
rect 27805 3707 27879 3716
rect 27805 3702 27814 3707
rect 16830 3656 27814 3702
rect 16830 3651 16839 3656
rect 16765 3642 16839 3651
rect 27805 3651 27814 3656
rect 27870 3702 27879 3707
rect 38845 3707 38919 3716
rect 38845 3702 38854 3707
rect 27870 3656 38854 3702
rect 27870 3651 27879 3656
rect 27805 3642 27879 3651
rect 38845 3651 38854 3656
rect 38910 3702 38919 3707
rect 49885 3707 49959 3716
rect 49885 3702 49894 3707
rect 38910 3656 49894 3702
rect 38910 3651 38919 3656
rect 38845 3642 38919 3651
rect 49885 3651 49894 3656
rect 49950 3702 49959 3707
rect 60925 3707 60999 3716
rect 60925 3702 60934 3707
rect 49950 3656 60934 3702
rect 49950 3651 49959 3656
rect 49885 3642 49959 3651
rect 60925 3651 60934 3656
rect 60990 3702 60999 3707
rect 71965 3707 72039 3716
rect 71965 3702 71974 3707
rect 60990 3656 71974 3702
rect 60990 3651 60999 3656
rect 60925 3642 60999 3651
rect 71965 3651 71974 3656
rect 72030 3702 72039 3707
rect 83005 3707 83079 3716
rect 83005 3702 83014 3707
rect 72030 3656 83014 3702
rect 72030 3651 72039 3656
rect 71965 3642 72039 3651
rect 83005 3651 83014 3656
rect 83070 3702 83079 3707
rect 94045 3707 94119 3716
rect 94045 3702 94054 3707
rect 83070 3656 94054 3702
rect 83070 3651 83079 3656
rect 83005 3642 83079 3651
rect 94045 3651 94054 3656
rect 94110 3651 94119 3707
rect 94045 3642 94119 3651
rect 86760 3615 86834 3624
rect 86760 3559 86769 3615
rect 86825 3559 86834 3615
rect 86760 3550 86834 3559
rect 1651 3389 1725 3398
rect 1651 3333 1660 3389
rect 1716 3333 1725 3389
rect 1651 3324 1725 3333
rect 12691 3389 12765 3398
rect 12691 3333 12700 3389
rect 12756 3333 12765 3389
rect 12691 3324 12765 3333
rect 23731 3389 23805 3398
rect 23731 3333 23740 3389
rect 23796 3333 23805 3389
rect 23731 3324 23805 3333
rect 34771 3389 34845 3398
rect 34771 3333 34780 3389
rect 34836 3333 34845 3389
rect 34771 3324 34845 3333
rect 45811 3389 45885 3398
rect 45811 3333 45820 3389
rect 45876 3333 45885 3389
rect 45811 3324 45885 3333
rect 56851 3389 56925 3398
rect 56851 3333 56860 3389
rect 56916 3333 56925 3389
rect 56851 3324 56925 3333
rect 67891 3389 67965 3398
rect 67891 3333 67900 3389
rect 67956 3333 67965 3389
rect 67891 3324 67965 3333
rect 78931 3389 79005 3398
rect 78931 3333 78940 3389
rect 78996 3333 79005 3389
rect 78931 3324 79005 3333
rect 89971 3389 90045 3398
rect 89971 3333 89980 3389
rect 90036 3333 90045 3389
rect 89971 3324 90045 3333
rect 96761 3389 96835 3398
rect 96761 3333 96770 3389
rect 96826 3333 96835 3389
rect 96761 3324 96835 3333
rect 8446 2761 8510 2767
rect 8446 2709 8452 2761
rect 8504 2758 8510 2761
rect 11245 2761 11309 2767
rect 11245 2758 11251 2761
rect 8504 2712 11251 2758
rect 8504 2709 8510 2712
rect 8446 2703 8510 2709
rect 11245 2709 11251 2712
rect 11303 2709 11309 2761
rect 11245 2703 11309 2709
rect 19486 2761 19550 2767
rect 19486 2709 19492 2761
rect 19544 2758 19550 2761
rect 22285 2761 22349 2767
rect 22285 2758 22291 2761
rect 19544 2712 22291 2758
rect 19544 2709 19550 2712
rect 19486 2703 19550 2709
rect 22285 2709 22291 2712
rect 22343 2709 22349 2761
rect 22285 2703 22349 2709
rect 30526 2761 30590 2767
rect 30526 2709 30532 2761
rect 30584 2758 30590 2761
rect 33325 2761 33389 2767
rect 33325 2758 33331 2761
rect 30584 2712 33331 2758
rect 30584 2709 30590 2712
rect 30526 2703 30590 2709
rect 33325 2709 33331 2712
rect 33383 2709 33389 2761
rect 33325 2703 33389 2709
rect 41566 2761 41630 2767
rect 41566 2709 41572 2761
rect 41624 2758 41630 2761
rect 44365 2761 44429 2767
rect 44365 2758 44371 2761
rect 41624 2712 44371 2758
rect 41624 2709 41630 2712
rect 41566 2703 41630 2709
rect 44365 2709 44371 2712
rect 44423 2709 44429 2761
rect 44365 2703 44429 2709
rect 52606 2761 52670 2767
rect 52606 2709 52612 2761
rect 52664 2758 52670 2761
rect 55405 2761 55469 2767
rect 55405 2758 55411 2761
rect 52664 2712 55411 2758
rect 52664 2709 52670 2712
rect 52606 2703 52670 2709
rect 55405 2709 55411 2712
rect 55463 2709 55469 2761
rect 55405 2703 55469 2709
rect 63646 2761 63710 2767
rect 63646 2709 63652 2761
rect 63704 2758 63710 2761
rect 66445 2761 66509 2767
rect 66445 2758 66451 2761
rect 63704 2712 66451 2758
rect 63704 2709 63710 2712
rect 63646 2703 63710 2709
rect 66445 2709 66451 2712
rect 66503 2709 66509 2761
rect 66445 2703 66509 2709
rect 74686 2761 74750 2767
rect 74686 2709 74692 2761
rect 74744 2758 74750 2761
rect 77485 2761 77549 2767
rect 77485 2758 77491 2761
rect 74744 2712 77491 2758
rect 74744 2709 74750 2712
rect 74686 2703 74750 2709
rect 77485 2709 77491 2712
rect 77543 2709 77549 2761
rect 77485 2703 77549 2709
rect 85726 2761 85790 2767
rect 85726 2709 85732 2761
rect 85784 2758 85790 2761
rect 88525 2761 88589 2767
rect 88525 2758 88531 2761
rect 85784 2712 88531 2758
rect 85784 2709 85790 2712
rect 85726 2703 85790 2709
rect 88525 2709 88531 2712
rect 88583 2709 88589 2761
rect 88525 2703 88589 2709
rect 5725 1833 5799 1842
rect 5725 1777 5734 1833
rect 5790 1777 5799 1833
rect 5725 1768 5799 1777
rect 16765 1833 16839 1842
rect 16765 1777 16774 1833
rect 16830 1777 16839 1833
rect 16765 1768 16839 1777
rect 27805 1833 27879 1842
rect 27805 1777 27814 1833
rect 27870 1777 27879 1833
rect 27805 1768 27879 1777
rect 38845 1833 38919 1842
rect 38845 1777 38854 1833
rect 38910 1777 38919 1833
rect 38845 1768 38919 1777
rect 49885 1833 49959 1842
rect 49885 1777 49894 1833
rect 49950 1777 49959 1833
rect 49885 1768 49959 1777
rect 60925 1833 60999 1842
rect 60925 1777 60934 1833
rect 60990 1777 60999 1833
rect 60925 1768 60999 1777
rect 71965 1833 72039 1842
rect 71965 1777 71974 1833
rect 72030 1777 72039 1833
rect 71965 1768 72039 1777
rect 83005 1833 83079 1842
rect 83005 1777 83014 1833
rect 83070 1777 83079 1833
rect 83005 1768 83079 1777
rect 87544 1833 87618 1842
rect 87544 1777 87553 1833
rect 87609 1777 87618 1833
rect 87544 1768 87618 1777
rect 94045 1833 94119 1842
rect 94045 1777 94054 1833
rect 94110 1777 94119 1833
rect 94045 1768 94119 1777
rect 5725 1577 5799 1586
rect 5725 1521 5734 1577
rect 5790 1521 5799 1577
rect 5725 1512 5799 1521
rect 16765 1577 16839 1586
rect 16765 1521 16774 1577
rect 16830 1521 16839 1577
rect 16765 1512 16839 1521
rect 27805 1577 27879 1586
rect 27805 1521 27814 1577
rect 27870 1521 27879 1577
rect 27805 1512 27879 1521
rect 38845 1577 38919 1586
rect 38845 1521 38854 1577
rect 38910 1521 38919 1577
rect 38845 1512 38919 1521
rect 49885 1577 49959 1586
rect 49885 1521 49894 1577
rect 49950 1521 49959 1577
rect 49885 1512 49959 1521
rect 60925 1577 60999 1586
rect 60925 1521 60934 1577
rect 60990 1521 60999 1577
rect 60925 1512 60999 1521
rect 71965 1577 72039 1586
rect 71965 1521 71974 1577
rect 72030 1521 72039 1577
rect 71965 1512 72039 1521
rect 83005 1577 83079 1586
rect 83005 1521 83014 1577
rect 83070 1521 83079 1577
rect 83005 1512 83079 1521
rect 94045 1577 94119 1586
rect 94045 1521 94054 1577
rect 94110 1521 94119 1577
rect 94045 1512 94119 1521
<< via2 >>
rect 331 39482 387 39538
rect 16774 39362 16830 39418
rect 23740 39362 23796 39418
rect 34780 39362 34836 39418
rect 45820 39362 45876 39418
rect 56860 39362 56916 39418
rect 67900 39362 67956 39418
rect 78940 39362 78996 39418
rect 89980 39362 90036 39418
rect 87553 38606 87609 38608
rect 87553 38554 87555 38606
rect 87555 38554 87607 38606
rect 87607 38554 87609 38606
rect 87553 38552 87609 38554
rect 12700 37742 12756 37798
rect 27814 37742 27870 37798
rect 38854 37742 38910 37798
rect 49894 37742 49950 37798
rect 60934 37742 60990 37798
rect 71974 37742 72030 37798
rect 83014 37742 83070 37798
rect 94054 37742 94110 37798
rect 96770 37050 96826 37052
rect 96770 36998 96772 37050
rect 96772 36998 96824 37050
rect 96824 36998 96826 37050
rect 96770 36996 96826 36998
rect 86769 36824 86825 36826
rect 86769 36772 86771 36824
rect 86771 36772 86823 36824
rect 86823 36772 86825 36824
rect 86769 36770 86825 36772
rect 16774 36678 16830 36734
rect 27814 36678 27870 36734
rect 38854 36678 38910 36734
rect 49894 36678 49950 36734
rect 60934 36678 60990 36734
rect 71974 36678 72030 36734
rect 83014 36678 83070 36734
rect 94054 36678 94110 36734
rect 12700 36586 12756 36642
rect 23740 36586 23796 36642
rect 34780 36586 34836 36642
rect 45820 36586 45876 36642
rect 56860 36586 56916 36642
rect 67900 36586 67956 36642
rect 78940 36586 78996 36642
rect 89980 36586 90036 36642
rect 1660 3743 1716 3799
rect 12700 3743 12756 3799
rect 23740 3743 23796 3799
rect 34780 3743 34836 3799
rect 45820 3743 45876 3799
rect 56860 3743 56916 3799
rect 67900 3743 67956 3799
rect 78940 3743 78996 3799
rect 89980 3743 90036 3799
rect 5734 3651 5790 3707
rect 16774 3651 16830 3707
rect 27814 3651 27870 3707
rect 38854 3651 38910 3707
rect 49894 3651 49950 3707
rect 60934 3651 60990 3707
rect 71974 3651 72030 3707
rect 83014 3651 83070 3707
rect 94054 3651 94110 3707
rect 86769 3613 86825 3615
rect 86769 3561 86771 3613
rect 86771 3561 86823 3613
rect 86823 3561 86825 3613
rect 86769 3559 86825 3561
rect 1660 3387 1716 3389
rect 1660 3335 1662 3387
rect 1662 3335 1714 3387
rect 1714 3335 1716 3387
rect 1660 3333 1716 3335
rect 12700 3387 12756 3389
rect 12700 3335 12702 3387
rect 12702 3335 12754 3387
rect 12754 3335 12756 3387
rect 12700 3333 12756 3335
rect 23740 3387 23796 3389
rect 23740 3335 23742 3387
rect 23742 3335 23794 3387
rect 23794 3335 23796 3387
rect 23740 3333 23796 3335
rect 34780 3387 34836 3389
rect 34780 3335 34782 3387
rect 34782 3335 34834 3387
rect 34834 3335 34836 3387
rect 34780 3333 34836 3335
rect 45820 3387 45876 3389
rect 45820 3335 45822 3387
rect 45822 3335 45874 3387
rect 45874 3335 45876 3387
rect 45820 3333 45876 3335
rect 56860 3387 56916 3389
rect 56860 3335 56862 3387
rect 56862 3335 56914 3387
rect 56914 3335 56916 3387
rect 56860 3333 56916 3335
rect 67900 3387 67956 3389
rect 67900 3335 67902 3387
rect 67902 3335 67954 3387
rect 67954 3335 67956 3387
rect 67900 3333 67956 3335
rect 78940 3387 78996 3389
rect 78940 3335 78942 3387
rect 78942 3335 78994 3387
rect 78994 3335 78996 3387
rect 78940 3333 78996 3335
rect 89980 3387 90036 3389
rect 89980 3335 89982 3387
rect 89982 3335 90034 3387
rect 90034 3335 90036 3387
rect 89980 3333 90036 3335
rect 96770 3387 96826 3389
rect 96770 3335 96772 3387
rect 96772 3335 96824 3387
rect 96824 3335 96826 3387
rect 96770 3333 96826 3335
rect 5734 1831 5790 1833
rect 5734 1779 5736 1831
rect 5736 1779 5788 1831
rect 5788 1779 5790 1831
rect 5734 1777 5790 1779
rect 16774 1831 16830 1833
rect 16774 1779 16776 1831
rect 16776 1779 16828 1831
rect 16828 1779 16830 1831
rect 16774 1777 16830 1779
rect 27814 1831 27870 1833
rect 27814 1779 27816 1831
rect 27816 1779 27868 1831
rect 27868 1779 27870 1831
rect 27814 1777 27870 1779
rect 38854 1831 38910 1833
rect 38854 1779 38856 1831
rect 38856 1779 38908 1831
rect 38908 1779 38910 1831
rect 38854 1777 38910 1779
rect 49894 1831 49950 1833
rect 49894 1779 49896 1831
rect 49896 1779 49948 1831
rect 49948 1779 49950 1831
rect 49894 1777 49950 1779
rect 60934 1831 60990 1833
rect 60934 1779 60936 1831
rect 60936 1779 60988 1831
rect 60988 1779 60990 1831
rect 60934 1777 60990 1779
rect 71974 1831 72030 1833
rect 71974 1779 71976 1831
rect 71976 1779 72028 1831
rect 72028 1779 72030 1831
rect 71974 1777 72030 1779
rect 83014 1831 83070 1833
rect 83014 1779 83016 1831
rect 83016 1779 83068 1831
rect 83068 1779 83070 1831
rect 83014 1777 83070 1779
rect 87553 1831 87609 1833
rect 87553 1779 87555 1831
rect 87555 1779 87607 1831
rect 87607 1779 87609 1831
rect 87553 1777 87609 1779
rect 94054 1831 94110 1833
rect 94054 1779 94056 1831
rect 94056 1779 94108 1831
rect 94108 1779 94110 1831
rect 94054 1777 94110 1779
rect 5734 1575 5790 1577
rect 5734 1523 5736 1575
rect 5736 1523 5788 1575
rect 5788 1523 5790 1575
rect 5734 1521 5790 1523
rect 16774 1575 16830 1577
rect 16774 1523 16776 1575
rect 16776 1523 16828 1575
rect 16828 1523 16830 1575
rect 16774 1521 16830 1523
rect 27814 1575 27870 1577
rect 27814 1523 27816 1575
rect 27816 1523 27868 1575
rect 27868 1523 27870 1575
rect 27814 1521 27870 1523
rect 38854 1575 38910 1577
rect 38854 1523 38856 1575
rect 38856 1523 38908 1575
rect 38908 1523 38910 1575
rect 38854 1521 38910 1523
rect 49894 1575 49950 1577
rect 49894 1523 49896 1575
rect 49896 1523 49948 1575
rect 49948 1523 49950 1575
rect 49894 1521 49950 1523
rect 60934 1575 60990 1577
rect 60934 1523 60936 1575
rect 60936 1523 60988 1575
rect 60988 1523 60990 1575
rect 60934 1521 60990 1523
rect 71974 1575 72030 1577
rect 71974 1523 71976 1575
rect 71976 1523 72028 1575
rect 72028 1523 72030 1575
rect 71974 1521 72030 1523
rect 83014 1575 83070 1577
rect 83014 1523 83016 1575
rect 83016 1523 83068 1575
rect 83068 1523 83070 1575
rect 83014 1521 83070 1523
rect 94054 1575 94110 1577
rect 94054 1523 94056 1575
rect 94056 1523 94108 1575
rect 94108 1523 94110 1575
rect 94054 1521 94110 1523
<< metal3 >>
rect 326 39538 392 39543
rect 326 39482 331 39538
rect 387 39482 392 39538
rect 326 39477 392 39482
rect 329 1577 389 39477
rect 16769 39418 16835 39423
rect 16769 39362 16774 39418
rect 16830 39362 16835 39418
rect 16769 39357 16835 39362
rect 23735 39418 23801 39423
rect 23735 39362 23740 39418
rect 23796 39362 23801 39418
rect 23735 39357 23801 39362
rect 34775 39418 34841 39423
rect 34775 39362 34780 39418
rect 34836 39362 34841 39418
rect 34775 39357 34841 39362
rect 45815 39418 45881 39423
rect 45815 39362 45820 39418
rect 45876 39362 45881 39418
rect 45815 39357 45881 39362
rect 56855 39418 56921 39423
rect 56855 39362 56860 39418
rect 56916 39362 56921 39418
rect 56855 39357 56921 39362
rect 67895 39418 67961 39423
rect 67895 39362 67900 39418
rect 67956 39362 67961 39418
rect 67895 39357 67961 39362
rect 78935 39418 79001 39423
rect 78935 39362 78940 39418
rect 78996 39362 79001 39418
rect 78935 39357 79001 39362
rect 89975 39418 90041 39423
rect 89975 39362 89980 39418
rect 90036 39362 90041 39418
rect 89975 39357 90041 39362
rect 13434 38612 13510 38618
rect 13434 38548 13440 38612
rect 13504 38548 13510 38612
rect 13434 38542 13510 38548
rect 12695 37798 12761 37803
rect 12695 37742 12700 37798
rect 12756 37742 12761 37798
rect 12695 37737 12761 37742
rect 12698 36647 12758 37737
rect 16772 36739 16832 39357
rect 16769 36734 16835 36739
rect 16769 36678 16774 36734
rect 16830 36678 16835 36734
rect 16769 36673 16835 36678
rect 12695 36642 12761 36647
rect 12695 36586 12700 36642
rect 12756 36586 12761 36642
rect 12695 36581 12761 36586
rect 12698 3804 12758 36581
rect 1655 3799 1721 3804
rect 1655 3743 1660 3799
rect 1716 3743 1721 3799
rect 1655 3738 1721 3743
rect 12695 3799 12761 3804
rect 12695 3743 12700 3799
rect 12756 3743 12761 3799
rect 12695 3738 12761 3743
rect 1658 3394 1718 3738
rect 5729 3707 5795 3712
rect 5729 3651 5734 3707
rect 5790 3651 5795 3707
rect 5729 3646 5795 3651
rect 1655 3389 1721 3394
rect 1655 3333 1660 3389
rect 1716 3333 1721 3389
rect 1655 3328 1721 3333
rect 5732 1838 5792 3646
rect 12698 3394 12758 3738
rect 16772 3712 16832 36673
rect 23738 36647 23798 39357
rect 24474 38612 24550 38618
rect 24474 38548 24480 38612
rect 24544 38548 24550 38612
rect 24474 38542 24550 38548
rect 27809 37798 27875 37803
rect 27809 37742 27814 37798
rect 27870 37742 27875 37798
rect 27809 37737 27875 37742
rect 27812 36739 27872 37737
rect 27809 36734 27875 36739
rect 27809 36678 27814 36734
rect 27870 36678 27875 36734
rect 27809 36673 27875 36678
rect 23735 36642 23801 36647
rect 23735 36586 23740 36642
rect 23796 36586 23801 36642
rect 23735 36581 23801 36586
rect 23738 3804 23798 36581
rect 23735 3799 23801 3804
rect 23735 3743 23740 3799
rect 23796 3743 23801 3799
rect 23735 3738 23801 3743
rect 16769 3707 16835 3712
rect 16769 3651 16774 3707
rect 16830 3651 16835 3707
rect 16769 3646 16835 3651
rect 12695 3389 12761 3394
rect 12695 3333 12700 3389
rect 12756 3333 12761 3389
rect 12695 3328 12761 3333
rect 5729 1833 5795 1838
rect 5729 1777 5734 1833
rect 5790 1777 5795 1833
rect 5729 1772 5795 1777
rect 6468 1837 6544 1843
rect 16772 1838 16832 3646
rect 23738 3394 23798 3738
rect 27812 3712 27872 36673
rect 34778 36647 34838 39357
rect 35514 38612 35590 38618
rect 35514 38548 35520 38612
rect 35584 38548 35590 38612
rect 35514 38542 35590 38548
rect 38849 37798 38915 37803
rect 38849 37742 38854 37798
rect 38910 37742 38915 37798
rect 38849 37737 38915 37742
rect 38852 36739 38912 37737
rect 38849 36734 38915 36739
rect 38849 36678 38854 36734
rect 38910 36678 38915 36734
rect 38849 36673 38915 36678
rect 34775 36642 34841 36647
rect 34775 36586 34780 36642
rect 34836 36586 34841 36642
rect 34775 36581 34841 36586
rect 34778 3804 34838 36581
rect 34775 3799 34841 3804
rect 34775 3743 34780 3799
rect 34836 3743 34841 3799
rect 34775 3738 34841 3743
rect 27809 3707 27875 3712
rect 27809 3651 27814 3707
rect 27870 3651 27875 3707
rect 27809 3646 27875 3651
rect 23735 3389 23801 3394
rect 23735 3333 23740 3389
rect 23796 3333 23801 3389
rect 23735 3328 23801 3333
rect 6468 1773 6474 1837
rect 6538 1773 6544 1837
rect 5732 1582 5792 1772
rect 6468 1767 6544 1773
rect 16769 1833 16835 1838
rect 16769 1777 16774 1833
rect 16830 1777 16835 1833
rect 16769 1772 16835 1777
rect 17508 1837 17584 1843
rect 27812 1838 27872 3646
rect 34778 3394 34838 3738
rect 38852 3712 38912 36673
rect 45818 36647 45878 39357
rect 46554 38612 46630 38618
rect 46554 38548 46560 38612
rect 46624 38548 46630 38612
rect 46554 38542 46630 38548
rect 49889 37798 49955 37803
rect 49889 37742 49894 37798
rect 49950 37742 49955 37798
rect 49889 37737 49955 37742
rect 49892 36739 49952 37737
rect 49889 36734 49955 36739
rect 49889 36678 49894 36734
rect 49950 36678 49955 36734
rect 49889 36673 49955 36678
rect 45815 36642 45881 36647
rect 45815 36586 45820 36642
rect 45876 36586 45881 36642
rect 45815 36581 45881 36586
rect 45818 3804 45878 36581
rect 45815 3799 45881 3804
rect 45815 3743 45820 3799
rect 45876 3743 45881 3799
rect 45815 3738 45881 3743
rect 38849 3707 38915 3712
rect 38849 3651 38854 3707
rect 38910 3651 38915 3707
rect 38849 3646 38915 3651
rect 34775 3389 34841 3394
rect 34775 3333 34780 3389
rect 34836 3333 34841 3389
rect 34775 3328 34841 3333
rect 17508 1773 17514 1837
rect 17578 1773 17584 1837
rect 16772 1582 16832 1772
rect 17508 1767 17584 1773
rect 27809 1833 27875 1838
rect 27809 1777 27814 1833
rect 27870 1777 27875 1833
rect 27809 1772 27875 1777
rect 28548 1837 28624 1843
rect 38852 1838 38912 3646
rect 45818 3394 45878 3738
rect 49892 3712 49952 36673
rect 56858 36647 56918 39357
rect 57594 38612 57670 38618
rect 57594 38548 57600 38612
rect 57664 38548 57670 38612
rect 57594 38542 57670 38548
rect 60929 37798 60995 37803
rect 60929 37742 60934 37798
rect 60990 37742 60995 37798
rect 60929 37737 60995 37742
rect 60932 36739 60992 37737
rect 60929 36734 60995 36739
rect 60929 36678 60934 36734
rect 60990 36678 60995 36734
rect 60929 36673 60995 36678
rect 56855 36642 56921 36647
rect 56855 36586 56860 36642
rect 56916 36586 56921 36642
rect 56855 36581 56921 36586
rect 56858 3804 56918 36581
rect 56855 3799 56921 3804
rect 56855 3743 56860 3799
rect 56916 3743 56921 3799
rect 56855 3738 56921 3743
rect 49889 3707 49955 3712
rect 49889 3651 49894 3707
rect 49950 3651 49955 3707
rect 49889 3646 49955 3651
rect 45815 3389 45881 3394
rect 45815 3333 45820 3389
rect 45876 3333 45881 3389
rect 45815 3328 45881 3333
rect 28548 1773 28554 1837
rect 28618 1773 28624 1837
rect 27812 1582 27872 1772
rect 28548 1767 28624 1773
rect 38849 1833 38915 1838
rect 38849 1777 38854 1833
rect 38910 1777 38915 1833
rect 38849 1772 38915 1777
rect 39588 1837 39664 1843
rect 49892 1838 49952 3646
rect 56858 3394 56918 3738
rect 60932 3712 60992 36673
rect 67898 36647 67958 39357
rect 68634 38612 68710 38618
rect 68634 38548 68640 38612
rect 68704 38548 68710 38612
rect 68634 38542 68710 38548
rect 71969 37798 72035 37803
rect 71969 37742 71974 37798
rect 72030 37742 72035 37798
rect 71969 37737 72035 37742
rect 71972 36739 72032 37737
rect 71969 36734 72035 36739
rect 71969 36678 71974 36734
rect 72030 36678 72035 36734
rect 71969 36673 72035 36678
rect 67895 36642 67961 36647
rect 67895 36586 67900 36642
rect 67956 36586 67961 36642
rect 67895 36581 67961 36586
rect 67898 3804 67958 36581
rect 67895 3799 67961 3804
rect 67895 3743 67900 3799
rect 67956 3743 67961 3799
rect 67895 3738 67961 3743
rect 60929 3707 60995 3712
rect 60929 3651 60934 3707
rect 60990 3651 60995 3707
rect 60929 3646 60995 3651
rect 56855 3389 56921 3394
rect 56855 3333 56860 3389
rect 56916 3333 56921 3389
rect 56855 3328 56921 3333
rect 39588 1773 39594 1837
rect 39658 1773 39664 1837
rect 38852 1582 38912 1772
rect 39588 1767 39664 1773
rect 49889 1833 49955 1838
rect 49889 1777 49894 1833
rect 49950 1777 49955 1833
rect 49889 1772 49955 1777
rect 50628 1837 50704 1843
rect 60932 1838 60992 3646
rect 67898 3394 67958 3738
rect 71972 3712 72032 36673
rect 78938 36647 78998 39357
rect 79674 38612 79750 38618
rect 79674 38548 79680 38612
rect 79744 38548 79750 38612
rect 79674 38542 79750 38548
rect 87124 38612 87200 38618
rect 87124 38548 87130 38612
rect 87194 38548 87200 38612
rect 87124 38542 87200 38548
rect 87548 38608 87614 38613
rect 87548 38552 87553 38608
rect 87609 38552 87614 38608
rect 87548 38547 87614 38552
rect 83009 37798 83075 37803
rect 83009 37742 83014 37798
rect 83070 37742 83075 37798
rect 83009 37737 83075 37742
rect 83012 36739 83072 37737
rect 86764 36826 86830 36831
rect 86764 36770 86769 36826
rect 86825 36770 86830 36826
rect 86764 36765 86830 36770
rect 83009 36734 83075 36739
rect 83009 36678 83014 36734
rect 83070 36678 83075 36734
rect 83009 36673 83075 36678
rect 78935 36642 79001 36647
rect 78935 36586 78940 36642
rect 78996 36586 79001 36642
rect 78935 36581 79001 36586
rect 78938 3804 78998 36581
rect 78935 3799 79001 3804
rect 78935 3743 78940 3799
rect 78996 3743 79001 3799
rect 78935 3738 79001 3743
rect 71969 3707 72035 3712
rect 71969 3651 71974 3707
rect 72030 3651 72035 3707
rect 71969 3646 72035 3651
rect 67895 3389 67961 3394
rect 67895 3333 67900 3389
rect 67956 3333 67961 3389
rect 67895 3328 67961 3333
rect 50628 1773 50634 1837
rect 50698 1773 50704 1837
rect 49892 1582 49952 1772
rect 50628 1767 50704 1773
rect 60929 1833 60995 1838
rect 60929 1777 60934 1833
rect 60990 1777 60995 1833
rect 60929 1772 60995 1777
rect 61668 1837 61744 1843
rect 71972 1838 72032 3646
rect 78938 3394 78998 3738
rect 83012 3712 83072 36673
rect 83009 3707 83075 3712
rect 83009 3651 83014 3707
rect 83070 3651 83075 3707
rect 83009 3646 83075 3651
rect 78935 3389 79001 3394
rect 78935 3333 78940 3389
rect 78996 3333 79001 3389
rect 78935 3328 79001 3333
rect 61668 1773 61674 1837
rect 61738 1773 61744 1837
rect 60932 1582 60992 1772
rect 61668 1767 61744 1773
rect 71969 1833 72035 1838
rect 71969 1777 71974 1833
rect 72030 1777 72035 1833
rect 71969 1772 72035 1777
rect 72708 1837 72784 1843
rect 83012 1838 83072 3646
rect 86767 3620 86827 36765
rect 86764 3615 86830 3620
rect 86764 3559 86769 3615
rect 86825 3559 86830 3615
rect 86764 3554 86830 3559
rect 87132 1843 87192 38542
rect 72708 1773 72714 1837
rect 72778 1773 72784 1837
rect 71972 1582 72032 1772
rect 72708 1767 72784 1773
rect 83009 1833 83075 1838
rect 83009 1777 83014 1833
rect 83070 1777 83075 1833
rect 83009 1772 83075 1777
rect 83748 1837 83824 1843
rect 83748 1773 83754 1837
rect 83818 1773 83824 1837
rect 83012 1582 83072 1772
rect 83748 1767 83824 1773
rect 87124 1837 87200 1843
rect 87551 1838 87611 38547
rect 89978 36647 90038 39357
rect 90714 38612 90790 38618
rect 90714 38548 90720 38612
rect 90784 38548 90790 38612
rect 90714 38542 90790 38548
rect 94049 37798 94115 37803
rect 94049 37742 94054 37798
rect 94110 37742 94115 37798
rect 94049 37737 94115 37742
rect 94052 36739 94112 37737
rect 96765 37052 96831 37057
rect 96765 36996 96770 37052
rect 96826 36996 96831 37052
rect 96765 36991 96831 36996
rect 94049 36734 94115 36739
rect 94049 36678 94054 36734
rect 94110 36678 94115 36734
rect 94049 36673 94115 36678
rect 89975 36642 90041 36647
rect 89975 36586 89980 36642
rect 90036 36586 90041 36642
rect 89975 36581 90041 36586
rect 89978 3804 90038 36581
rect 89975 3799 90041 3804
rect 89975 3743 89980 3799
rect 90036 3743 90041 3799
rect 89975 3738 90041 3743
rect 89978 3394 90038 3738
rect 94052 3712 94112 36673
rect 94049 3707 94115 3712
rect 94049 3651 94054 3707
rect 94110 3651 94115 3707
rect 94049 3646 94115 3651
rect 89975 3389 90041 3394
rect 89975 3333 89980 3389
rect 90036 3333 90041 3389
rect 89975 3328 90041 3333
rect 94052 1838 94112 3646
rect 96768 3394 96828 36991
rect 96765 3389 96831 3394
rect 96765 3333 96770 3389
rect 96826 3333 96831 3389
rect 96765 3328 96831 3333
rect 87124 1773 87130 1837
rect 87194 1773 87200 1837
rect 87124 1767 87200 1773
rect 87548 1833 87614 1838
rect 87548 1777 87553 1833
rect 87609 1777 87614 1833
rect 87548 1772 87614 1777
rect 94049 1833 94115 1838
rect 94049 1777 94054 1833
rect 94110 1777 94115 1833
rect 94049 1772 94115 1777
rect 94788 1837 94864 1843
rect 94788 1773 94794 1837
rect 94858 1773 94864 1837
rect 94052 1582 94112 1772
rect 94788 1767 94864 1773
rect 5729 1577 5795 1582
rect 5729 1521 5734 1577
rect 5790 1521 5795 1577
rect 5729 1516 5795 1521
rect 16769 1577 16835 1582
rect 16769 1521 16774 1577
rect 16830 1521 16835 1577
rect 16769 1516 16835 1521
rect 27809 1577 27875 1582
rect 27809 1521 27814 1577
rect 27870 1521 27875 1577
rect 27809 1516 27875 1521
rect 38849 1577 38915 1582
rect 38849 1521 38854 1577
rect 38910 1521 38915 1577
rect 38849 1516 38915 1521
rect 49889 1577 49955 1582
rect 49889 1521 49894 1577
rect 49950 1521 49955 1577
rect 49889 1516 49955 1521
rect 60929 1577 60995 1582
rect 60929 1521 60934 1577
rect 60990 1521 60995 1577
rect 60929 1516 60995 1521
rect 71969 1577 72035 1582
rect 71969 1521 71974 1577
rect 72030 1521 72035 1577
rect 71969 1516 72035 1521
rect 83009 1577 83075 1582
rect 83009 1521 83014 1577
rect 83070 1521 83075 1577
rect 83009 1516 83075 1521
rect 94049 1577 94115 1582
rect 94049 1521 94054 1577
rect 94110 1521 94115 1577
rect 94049 1516 94115 1521
rect 97205 51 97265 3559
<< via3 >>
rect 13440 38548 13504 38612
rect 24480 38548 24544 38612
rect 35520 38548 35584 38612
rect 6474 1773 6538 1837
rect 46560 38548 46624 38612
rect 17514 1773 17578 1837
rect 57600 38548 57664 38612
rect 28554 1773 28618 1837
rect 68640 38548 68704 38612
rect 39594 1773 39658 1837
rect 79680 38548 79744 38612
rect 87130 38548 87194 38612
rect 50634 1773 50698 1837
rect 61674 1773 61738 1837
rect 72714 1773 72778 1837
rect 83754 1773 83818 1837
rect 90720 38548 90784 38612
rect 87130 1773 87194 1837
rect 94794 1773 94858 1837
<< metal4 >>
rect 13439 38612 13505 38613
rect 13439 38548 13440 38612
rect 13504 38610 13505 38612
rect 24479 38612 24545 38613
rect 24479 38610 24480 38612
rect 13504 38550 24480 38610
rect 13504 38548 13505 38550
rect 13439 38547 13505 38548
rect 24479 38548 24480 38550
rect 24544 38610 24545 38612
rect 35519 38612 35585 38613
rect 35519 38610 35520 38612
rect 24544 38550 35520 38610
rect 24544 38548 24545 38550
rect 24479 38547 24545 38548
rect 35519 38548 35520 38550
rect 35584 38610 35585 38612
rect 46559 38612 46625 38613
rect 46559 38610 46560 38612
rect 35584 38550 46560 38610
rect 35584 38548 35585 38550
rect 35519 38547 35585 38548
rect 46559 38548 46560 38550
rect 46624 38610 46625 38612
rect 57599 38612 57665 38613
rect 57599 38610 57600 38612
rect 46624 38550 57600 38610
rect 46624 38548 46625 38550
rect 46559 38547 46625 38548
rect 57599 38548 57600 38550
rect 57664 38610 57665 38612
rect 68639 38612 68705 38613
rect 68639 38610 68640 38612
rect 57664 38550 68640 38610
rect 57664 38548 57665 38550
rect 57599 38547 57665 38548
rect 68639 38548 68640 38550
rect 68704 38610 68705 38612
rect 79679 38612 79745 38613
rect 79679 38610 79680 38612
rect 68704 38550 79680 38610
rect 68704 38548 68705 38550
rect 68639 38547 68705 38548
rect 79679 38548 79680 38550
rect 79744 38610 79745 38612
rect 87129 38612 87195 38613
rect 87129 38610 87130 38612
rect 79744 38550 87130 38610
rect 79744 38548 79745 38550
rect 79679 38547 79745 38548
rect 87129 38548 87130 38550
rect 87194 38610 87195 38612
rect 90719 38612 90785 38613
rect 90719 38610 90720 38612
rect 87194 38550 90720 38610
rect 87194 38548 87195 38550
rect 87129 38547 87195 38548
rect 90719 38548 90720 38550
rect 90784 38548 90785 38612
rect 90719 38547 90785 38548
rect 6473 1837 6539 1838
rect 6473 1773 6474 1837
rect 6538 1835 6539 1837
rect 17513 1837 17579 1838
rect 17513 1835 17514 1837
rect 6538 1775 17514 1835
rect 6538 1773 6539 1775
rect 6473 1772 6539 1773
rect 17513 1773 17514 1775
rect 17578 1835 17579 1837
rect 28553 1837 28619 1838
rect 28553 1835 28554 1837
rect 17578 1775 28554 1835
rect 17578 1773 17579 1775
rect 17513 1772 17579 1773
rect 28553 1773 28554 1775
rect 28618 1835 28619 1837
rect 39593 1837 39659 1838
rect 39593 1835 39594 1837
rect 28618 1775 39594 1835
rect 28618 1773 28619 1775
rect 28553 1772 28619 1773
rect 39593 1773 39594 1775
rect 39658 1835 39659 1837
rect 50633 1837 50699 1838
rect 50633 1835 50634 1837
rect 39658 1775 50634 1835
rect 39658 1773 39659 1775
rect 39593 1772 39659 1773
rect 50633 1773 50634 1775
rect 50698 1835 50699 1837
rect 61673 1837 61739 1838
rect 61673 1835 61674 1837
rect 50698 1775 61674 1835
rect 50698 1773 50699 1775
rect 50633 1772 50699 1773
rect 61673 1773 61674 1775
rect 61738 1835 61739 1837
rect 72713 1837 72779 1838
rect 72713 1835 72714 1837
rect 61738 1775 72714 1835
rect 61738 1773 61739 1775
rect 61673 1772 61739 1773
rect 72713 1773 72714 1775
rect 72778 1835 72779 1837
rect 83753 1837 83819 1838
rect 83753 1835 83754 1837
rect 72778 1775 83754 1835
rect 72778 1773 72779 1775
rect 72713 1772 72779 1773
rect 83753 1773 83754 1775
rect 83818 1835 83819 1837
rect 87129 1837 87195 1838
rect 87129 1835 87130 1837
rect 83818 1775 87130 1835
rect 83818 1773 83819 1775
rect 83753 1772 83819 1773
rect 87129 1773 87130 1775
rect 87194 1835 87195 1837
rect 94793 1837 94859 1838
rect 94793 1835 94794 1837
rect 87194 1775 94794 1835
rect 87194 1773 87195 1775
rect 87129 1772 87195 1773
rect 94793 1773 94794 1775
rect 94858 1773 94859 1837
rect 94793 1772 94859 1773
use D_FlipFlop  D_FlipFlop_1
timestamp 1755875389
transform 1 0 22168 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1755875389
transform 1 0 33208 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1755875389
transform 1 0 44248 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1755875389
transform 1 0 55288 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1755875389
transform 1 0 66328 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1755875389
transform 1 0 88408 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1755875389
transform 1 0 77368 0 1 38557
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_8
timestamp 1755875389
transform -1 0 19890 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_9
timestamp 1755875389
transform -1 0 86130 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_10
timestamp 1755875389
transform -1 0 97170 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_11
timestamp 1755875389
transform -1 0 75090 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_12
timestamp 1755875389
transform -1 0 64050 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_13
timestamp 1755875389
transform -1 0 53010 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_14
timestamp 1755875389
transform -1 0 41970 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_15
timestamp 1755875389
transform -1 0 30930 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_16
timestamp 1755875389
transform -1 0 8850 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_17
timestamp 1755875389
transform 1 0 11128 0 1 38557
box -102 -1796 8762 1842
<< labels >>
flabel metal3 96768 3389 96828 33240 0 FreeSans 160 0 0 0 Q7
port 7 nsew
flabel metal2 85784 2712 88531 2758 0 FreeSans 160 0 0 0 Q8
port 8 nsew
flabel metal2 74744 2712 77491 2758 0 FreeSans 160 0 0 0 Q9
port 9 nsew
flabel metal2 63704 2712 66451 2758 0 FreeSans 160 0 0 0 Q10
port 10 nsew
flabel metal2 52664 2712 55411 2758 0 FreeSans 160 0 0 0 Q11
port 11 nsew
flabel metal2 41624 2712 44371 2758 0 FreeSans 160 0 0 0 Q12
port 12 nsew
flabel metal2 30590 2712 33331 2758 0 FreeSans 160 0 0 0 Q13
port 13 nsew
flabel metal2 19544 2712 22291 2758 0 FreeSans 160 0 0 0 Q14
port 14 nsew
flabel metal2 8504 2712 11251 2758 0 FreeSans 160 0 0 0 Q15
port 15 nsew
flabel metal2 78996 3748 89980 3794 0 FreeSans 160 0 0 0 EN
port 16 nsew
flabel metal2 83070 3656 94054 3702 0 FreeSans 160 0 0 0 VDD
port 17 nsew
flabel metal3 97205 51 97265 3559 0 FreeSans 160 90 0 0 GND
port 20 nsew
flabel metal4 83818 1775 87130 1835 0 FreeSans 160 0 0 0 CLK
port 21 nsew
flabel metal2 19767 39487 22514 39533 0 FreeSans 160 0 0 0 Q0
port 0 nsew
flabel metal2 30807 39487 33554 39533 0 FreeSans 160 0 0 0 Q1
port 1 nsew
flabel metal2 41847 39487 44594 39533 0 FreeSans 160 0 0 0 Q2
port 2 nsew
flabel metal2 52887 39487 55634 39533 0 FreeSans 160 0 0 0 Q3
port 3 nsew
flabel metal2 63927 39487 66674 39533 0 FreeSans 160 0 0 0 Q4
port 4 nsew
flabel metal2 74967 39487 77714 39533 0 FreeSans 160 0 0 0 Q5
port 5 nsew
flabel metal2 86007 39487 88754 39533 0 FreeSans 160 0 0 0 Q6
port 6 nsew
<< end >>
