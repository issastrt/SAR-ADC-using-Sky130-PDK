** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_04-36-38/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.4870588235 8.5u 0.4870588235 8.500001u 0.488823529375 17u 0.488823529375 17.000001u 0.49058823525 25.5u
+ 0.49058823525 25.500001u 0.492352941125 34u 0.492352941125 34.000001u 0.494117647 42.5u 0.494117647 42.500001u 0.54352941175 51u 0.54352941175
+ 51.000001u 0.545294117625 59.5u 0.545294117625 59.500001u 0.5470588235 68u 0.5470588235 68.000001u 0.548823529375 76.5u 0.548823529375
+ 76.500001u 0.6 85u 0.6 85.000001u 0.601764705875 93.5u 0.601764705875 93.500001u 0.60352941175 102u 0.60352941175 102.000001u 0.605294117625
+ 110.5u 0.605294117625 110.500001u 0.656470588125 119u 0.656470588125 119.000001u 0.658235294 127.5u 0.658235294 127.500001u 0.66 136u
+ 0.66 136.000001u 0.661764705875 144.5u 0.661764705875 144.500001u 0.712941176375 153u 0.712941176375 153.000001u 0.71470588225 161.5u
+ 0.71470588225 161.500001u 0.716470588125 170u 0.716470588125 170.000001u 0.718235294 178.5u 0.718235294 178.500001u 0.769411764625 187u
+ 0.769411764625 187.000001u 0.7711764705 195.5u 0.7711764705 195.500001u 0.772941176375 204u 0.772941176375 204.000001u 0.77470588225 212.5u
+ 0.77470588225 212.500001u 0.776470588125 221u 0.776470588125 221.000001u 0.825882352875 229.5u 0.825882352875 229.500001u 0.82764705875 238u
+ 0.82764705875 238.000001u 0.829411764625 246.5u 0.829411764625 246.500001u 0.8311764705 255u 0.8311764705 255.000001u 0.882352941125 263.5u
+ 0.882352941125 263.500001u 0.884117647 272u 0.884117647 272.000001u 0.885882352875 280.5u 0.885882352875)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=125
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 280.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-13_04-36-38/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
