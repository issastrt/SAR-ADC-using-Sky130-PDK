magic
tech sky130A
timestamp 1753016136
<< pwell >>
rect -186 -201 186 201
<< mvnmos >>
rect -72 -72 72 72
<< mvndiff >>
rect -101 66 -72 72
rect -101 -66 -95 66
rect -78 -66 -72 66
rect -101 -72 -72 -66
rect 72 66 101 72
rect 72 -66 78 66
rect 95 -66 101 66
rect 72 -72 101 -66
<< mvndiffc >>
rect -95 -66 -78 66
rect 78 -66 95 66
<< mvpsubdiff >>
rect -168 177 168 183
rect -168 160 -114 177
rect 114 160 168 177
rect -168 154 168 160
rect -168 129 -139 154
rect -168 -129 -162 129
rect -145 -129 -139 129
rect 139 129 168 154
rect -168 -154 -139 -129
rect 139 -129 145 129
rect 162 -129 168 129
rect 139 -154 168 -129
rect -168 -160 168 -154
rect -168 -177 -114 -160
rect 114 -177 168 -160
rect -168 -183 168 -177
<< mvpsubdiffcont >>
rect -114 160 114 177
rect -162 -129 -145 129
rect 145 -129 162 129
rect -114 -177 114 -160
<< poly >>
rect -72 108 72 116
rect -72 91 -64 108
rect 64 91 72 108
rect -72 72 72 91
rect -72 -91 72 -72
rect -72 -108 -64 -91
rect 64 -108 72 -91
rect -72 -116 72 -108
<< polycont >>
rect -64 91 64 108
rect -64 -108 64 -91
<< locali >>
rect -162 160 -114 177
rect 114 160 162 177
rect -162 129 -145 160
rect 145 129 162 160
rect -72 91 -64 108
rect 64 91 72 108
rect -95 66 -78 74
rect -95 -74 -78 -66
rect 78 66 95 74
rect 78 -74 95 -66
rect -72 -108 -64 -91
rect 64 -108 72 -91
rect -162 -160 -145 -129
rect 145 -160 162 -129
rect -162 -177 -114 -160
rect 114 -177 162 -160
<< viali >>
rect -64 91 64 108
rect -95 -66 -78 66
rect 78 -66 95 66
rect -64 -108 64 -91
<< metal1 >>
rect -70 108 70 111
rect -70 91 -64 108
rect 64 91 70 108
rect -70 88 70 91
rect -98 66 -75 72
rect -98 -66 -95 66
rect -78 -66 -75 66
rect -98 -72 -75 -66
rect 75 66 98 72
rect 75 -66 78 66
rect 95 -66 98 66
rect 75 -72 98 -66
rect -70 -91 70 -88
rect -70 -108 -64 -91
rect 64 -108 70 -91
rect -70 -111 70 -108
<< properties >>
string FIXED_BBOX -153 -168 153 168
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.44 l 1.44 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
