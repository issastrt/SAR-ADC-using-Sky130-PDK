** sch_path: /home/issa/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-07_20-22-19/parameters/offset_error/run_2/offset_error.sch
**.subckt offset_error
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VVin Vin GND PWL(0u 0 8.5u 0 8.500001u 0.001 17u 0.001 17.000001u 0.002 25.5u 0.002 25.500001u 0.003 34u 0.003 34.000001u 0.004
+ 42.5u 0.004 42.500001u 0.005 51u 0.005 51.000001u 0.006 59.5u 0.006 59.500001u 0.007 68u 0.007 68.000001u 0.008 76.5u 0.008 76.500001u
+ 0.009 85u 0.009 85.000001u 0.010 93.5u 0.010 93.500001u 0.011 102u 0.011 102.000001u 0.012 110.5u 0.012 110.500001u 0.013 119u 0.013
+ 119.000001u 0.014 127.5u 0.014 127.500001u 0.015 136u 0.015)
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
R1 net1 GND 0.01 m=1
**** begin user architecture code

.control
tran 0.5u 136u uic
set wr_singlescale
wrdata /home/issa/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-07_20-22-19/parameters/offset_error/run_2/offset_error_2.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)
quit
.endc



* CACE gensim simulation file offset_error_2
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/issa/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice ss

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
