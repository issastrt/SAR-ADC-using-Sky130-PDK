** sch_path: /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_21-12-20/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.139411764125 8.5u 0.139411764125 8.500001u 0.141176470000 17u 0.141176470000 17.000001u 0.142941175875 25.5u
+ 0.142941175875 25.500001u 0.144705881750 34u 0.144705881750 34.000001u 0.146470587625 42.5u 0.146470587625 42.500001u 0.148235293500 51u
+ 0.148235293500 51.000001u 0.149999999375 59.5u 0.149999999375 59.500001u 0.151764705250 68u 0.151764705250 68.000001u 0.153529411125 76.5u
+ 0.153529411125 76.500001u 0.155294117000 85u 0.155294117000 85.000001u 0.157058822875 93.5u 0.157058822875 93.500001u 0.158823528750 102u
+ 0.158823528750 102.000001u 0.160588234625 110.5u 0.160588234625 110.500001u 0.162352940500 119u 0.162352940500 119.000001u 0.164117646375 127.5u
+ 0.164117646375 127.500001u 0.165882352250 136u 0.165882352250 136.000001u 0.167647058125 144.5u 0.167647058125 144.500001u 0.169411764000 153u
+ 0.169411764000 153.000001u 0.171176469875 161.5u 0.171176469875 161.500001u 0.172941175750 170u 0.172941175750 170.000001u 0.174705881625 178.5u
+ 0.174705881625 178.500001u 0.176470587500 187u 0.176470587500 187.000001u 0.178235293375 195.5u 0.178235293375 195.500001u 0.179999999250 204u
+ 0.179999999250 204.000001u 0.181764705125 212.5u 0.181764705125 212.500001u 0.183529411000 221u 0.183529411000 221.000001u 0.185294116875 229.5u
+ 0.185294116875 229.500001u 0.187058822750 238u 0.187058822750 238.000001u 0.188823528625 246.5u 0.188823528625 246.500001u 0.190588234500 255u
+ 0.190588234500 255.000001u 0.192352940375 263.5u 0.192352940375 263.500001u 0.194117646250 272u 0.194117646250 272.000001u 0.195882352125 280.5u
+ 0.195882352125 280.500001u 0.197647058000 289u 0.197647058000 289.000001u 0.199411763875 297.5u 0.199411763875 297.500001u 0.201176469750 306u
+ 0.201176469750 306.000001u 0.202941175625 314.5u 0.202941175625 314.500001u 0.204705881500 323u 0.204705881500 323.000001u 0.206470587375 331.5u
+ 0.206470587375 331.500001u 0.208235293250 340u 0.208235293250 340.000001u 0.210000000125 348.5u 0.210000000125 348.500001u 0.211764706000 357u
+ 0.211764706000 357.000001u 0.213529411875 365.5u 0.213529411875 365.500001u 0.215294117750 374u 0.215294117750 374.000001u 0.217058823625 382.5u
+ 0.217058823625 382.500001u 0.218823529500 391u 0.218823529500 391.000001u 0.220588235375 399.5u 0.220588235375 399.500001u 0.222352941250 408u
+ 0.222352941250 408.000001u 0.224117647125 416.5u 0.224117647125 416.500001u 0.225882353000 425u 0.225882353000 425.000001u 0.227647058875 433.5u
+ 0.227647058875 433.500001u 0.229411764750 442u 0.229411764750 442.000001u 0.231176470625 450.5u 0.231176470625 450.500001u 0.232941176500 459u
+ 0.232941176500 459.000001u 0.234705882375 467.5u 0.234705882375 467.500001u 0.236470588250 476u 0.236470588250 476.000001u 0.238235294125 484.5u
+ 0.238235294125 484.500001u 0.240000000000 493u 0.240000000000 493.000001u 0.241764705875 501.5u 0.241764705875 501.500001u 0.243529411750 510u
+ 0.243529411750 510.000001u 0.245294117625 518.5u 0.245294117625 518.500001u 0.247058823500 527u 0.247058823500 527.000001u 0.248823529375 535.5u
+ 0.248823529375 535.500001u 0.250588235250 544u 0.250588235250 544.000001u 0.252352941125 552.5u 0.252352941125 552.500001u 0.254117647000 561u
+ 0.254117647000 561.000001u 0.255882352875 569.5u 0.255882352875 569.500001u 0.257647058750 578u 0.257647058750 578.000001u 0.259411764625 586.5u
+ 0.259411764625 586.500001u 0.261176470500 595u 0.261176470500 595.000001u 0.262941176375 603.5u 0.262941176375 603.500001u 0.264705882250 612u
+ 0.264705882250 612.000001u 0.266470588125 620.5u 0.266470588125 620.500001u 0.268235294000 629u 0.268235294000 629.000001u 0.270000000000 637.5u
+ 0.270000000000 637.500001u 0.271764705875 646u 0.271764705875 646.000001u 0.273529411750 654.5u 0.273529411750 654.500001u 0.275294117625 663u
+ 0.275294117625 663.000001u 0.277058823500 671.5u 0.277058823500 671.500001u 0.278823529375 680u 0.278823529375)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/madra/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 680u uic
  wrdata /home/madra/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_21-12-20/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
