magic
tech sky130A
magscale 1 2
timestamp 1757233891
<< nwell >>
rect -2503 49987 -2429 50061
rect 6259 49987 6333 50061
rect 15021 49987 15095 50061
rect 23783 49987 23857 50061
rect 32545 49987 32619 50061
rect 41307 49987 41381 50061
rect 12794 46139 12868 46213
rect 16738 46139 16812 46213
rect 20682 46139 20756 46213
rect 24626 46139 24700 46213
rect 28570 46139 28644 46213
rect 32514 46139 32588 46213
rect 36458 46139 36532 46213
<< mvnsubdiff >>
rect -2436 49995 -2429 50061
rect 6326 49995 6333 50061
rect 15088 49995 15095 50061
rect 23850 49995 23857 50061
rect 32612 49995 32619 50061
rect 41374 49995 41381 50061
<< metal1 >>
rect 50604 55861 50668 55867
rect 50604 55809 50610 55861
rect 50662 55809 50668 55861
rect 50604 55803 50668 55809
rect -12804 53576 -12740 53582
rect -12804 53524 -12798 53576
rect -12746 53573 -12740 53576
rect 57650 53576 57714 53582
rect 57650 53573 57656 53576
rect -12746 53527 57656 53573
rect -12746 53524 -12740 53527
rect -12804 53518 -12740 53524
rect 57650 53524 57656 53527
rect 57708 53524 57714 53576
rect 57650 53518 57714 53524
rect -7180 53320 -7116 53326
rect -7180 53318 -7174 53320
rect -7185 53272 -7174 53318
rect -7180 53268 -7174 53272
rect -7122 53318 -7116 53320
rect -6566 53320 -6502 53326
rect -6566 53318 -6560 53320
rect -7122 53272 -7111 53318
rect -6571 53272 -6560 53318
rect -7122 53268 -7116 53272
rect -7180 53262 -7116 53268
rect -6566 53268 -6560 53272
rect -6508 53318 -6502 53320
rect 1582 53320 1646 53326
rect 1582 53318 1588 53320
rect -6508 53272 -6497 53318
rect 1577 53272 1588 53318
rect -6508 53268 -6502 53272
rect -6566 53262 -6502 53268
rect 1582 53268 1588 53272
rect 1640 53318 1646 53320
rect 2196 53320 2260 53326
rect 2196 53318 2202 53320
rect 1640 53272 1651 53318
rect 2191 53272 2202 53318
rect 1640 53268 1646 53272
rect 1582 53262 1646 53268
rect 2196 53268 2202 53272
rect 2254 53318 2260 53320
rect 10344 53320 10408 53326
rect 10344 53318 10350 53320
rect 2254 53272 2265 53318
rect 10339 53272 10350 53318
rect 2254 53268 2260 53272
rect 2196 53262 2260 53268
rect 10344 53268 10350 53272
rect 10402 53318 10408 53320
rect 10958 53320 11022 53326
rect 10958 53318 10964 53320
rect 10402 53272 10413 53318
rect 10953 53272 10964 53318
rect 10402 53268 10408 53272
rect 10344 53262 10408 53268
rect 10958 53268 10964 53272
rect 11016 53318 11022 53320
rect 19106 53320 19170 53326
rect 19106 53318 19112 53320
rect 11016 53272 11027 53318
rect 19101 53272 19112 53318
rect 11016 53268 11022 53272
rect 10958 53262 11022 53268
rect 19106 53268 19112 53272
rect 19164 53318 19170 53320
rect 19720 53320 19784 53326
rect 19720 53318 19726 53320
rect 19164 53272 19175 53318
rect 19715 53272 19726 53318
rect 19164 53268 19170 53272
rect 19106 53262 19170 53268
rect 19720 53268 19726 53272
rect 19778 53318 19784 53320
rect 27868 53320 27932 53326
rect 27868 53318 27874 53320
rect 19778 53272 19789 53318
rect 27863 53272 27874 53318
rect 19778 53268 19784 53272
rect 19720 53262 19784 53268
rect 27868 53268 27874 53272
rect 27926 53318 27932 53320
rect 28482 53320 28546 53326
rect 28482 53318 28488 53320
rect 27926 53272 27937 53318
rect 28477 53272 28488 53318
rect 27926 53268 27932 53272
rect 27868 53262 27932 53268
rect 28482 53268 28488 53272
rect 28540 53318 28546 53320
rect 36630 53320 36694 53326
rect 36630 53318 36636 53320
rect 28540 53272 28551 53318
rect 36625 53272 36636 53318
rect 28540 53268 28546 53272
rect 28482 53262 28546 53268
rect 36630 53268 36636 53272
rect 36688 53318 36694 53320
rect 37244 53320 37308 53326
rect 37244 53318 37250 53320
rect 36688 53272 36699 53318
rect 37239 53272 37250 53318
rect 36688 53268 36694 53272
rect 36630 53262 36694 53268
rect 37244 53268 37250 53272
rect 37302 53318 37308 53320
rect 45392 53320 45456 53326
rect 45392 53318 45398 53320
rect 37302 53272 37313 53318
rect 45387 53272 45398 53318
rect 37302 53268 37308 53272
rect 37244 53262 37308 53268
rect 45392 53268 45398 53272
rect 45450 53318 45456 53320
rect 46006 53320 46070 53326
rect 46006 53318 46012 53320
rect 45450 53272 45461 53318
rect 46001 53272 46012 53318
rect 45450 53268 45456 53272
rect 45392 53262 45456 53268
rect 46006 53268 46012 53272
rect 46064 53318 46070 53320
rect 54154 53320 54218 53326
rect 54154 53318 54160 53320
rect 46064 53272 46075 53318
rect 54149 53272 54160 53318
rect 46064 53268 46070 53272
rect 46006 53262 46070 53268
rect 54154 53268 54160 53272
rect 54212 53318 54218 53320
rect 54768 53319 54832 53325
rect 54212 53272 54223 53318
rect 54212 53268 54218 53272
rect 54154 53262 54218 53268
rect 54768 53267 54774 53319
rect 54826 53267 54832 53319
rect 54768 53261 54832 53267
rect -11319 52904 -11255 52910
rect -11319 52852 -11313 52904
rect -11261 52852 -11255 52904
rect -11319 52846 -11255 52852
rect -2557 52904 -2493 52910
rect -2557 52852 -2551 52904
rect -2499 52852 -2493 52904
rect -2557 52846 -2493 52852
rect 6205 52904 6269 52910
rect 6205 52852 6211 52904
rect 6263 52852 6269 52904
rect 6205 52846 6269 52852
rect 14967 52904 15031 52910
rect 14967 52852 14973 52904
rect 15025 52852 15031 52904
rect 14967 52846 15031 52852
rect 23729 52904 23793 52910
rect 23729 52852 23735 52904
rect 23787 52852 23793 52904
rect 23729 52846 23793 52852
rect 32491 52904 32555 52910
rect 32491 52852 32497 52904
rect 32549 52852 32555 52904
rect 32491 52846 32555 52852
rect 41253 52904 41317 52910
rect 41253 52852 41259 52904
rect 41311 52852 41317 52904
rect 41253 52846 41317 52852
rect 50015 52904 50079 52910
rect 50015 52852 50021 52904
rect 50073 52852 50079 52904
rect 50015 52846 50079 52852
rect -11933 52646 -11869 52652
rect -11933 52594 -11927 52646
rect -11875 52594 -11869 52646
rect -11933 52588 -11869 52594
rect -7403 52646 -7339 52652
rect -7403 52594 -7397 52646
rect -7345 52594 -7339 52646
rect -7403 52588 -7339 52594
rect -3171 52646 -3107 52652
rect -3171 52594 -3165 52646
rect -3113 52594 -3107 52646
rect -3171 52588 -3107 52594
rect 1359 52646 1423 52652
rect 1359 52594 1365 52646
rect 1417 52594 1423 52646
rect 1359 52588 1423 52594
rect 5591 52646 5655 52652
rect 5591 52594 5597 52646
rect 5649 52594 5655 52646
rect 5591 52588 5655 52594
rect 10121 52646 10185 52652
rect 10121 52594 10127 52646
rect 10179 52594 10185 52646
rect 10121 52588 10185 52594
rect 14353 52646 14417 52652
rect 14353 52594 14359 52646
rect 14411 52594 14417 52646
rect 14353 52588 14417 52594
rect 18883 52646 18947 52652
rect 18883 52594 18889 52646
rect 18941 52594 18947 52646
rect 18883 52588 18947 52594
rect 23115 52646 23179 52652
rect 23115 52594 23121 52646
rect 23173 52594 23179 52646
rect 23115 52588 23179 52594
rect 27645 52646 27709 52652
rect 27645 52594 27651 52646
rect 27703 52594 27709 52646
rect 27645 52588 27709 52594
rect 31877 52646 31941 52652
rect 31877 52594 31883 52646
rect 31935 52594 31941 52646
rect 31877 52588 31941 52594
rect 36407 52646 36471 52652
rect 36407 52594 36413 52646
rect 36465 52594 36471 52646
rect 36407 52588 36471 52594
rect 40639 52646 40703 52652
rect 40639 52594 40645 52646
rect 40697 52594 40703 52646
rect 40639 52588 40703 52594
rect 45169 52646 45233 52652
rect 45169 52594 45175 52646
rect 45227 52594 45233 52646
rect 45169 52588 45233 52594
rect 49401 52646 49465 52652
rect 49401 52594 49407 52646
rect 49459 52594 49465 52646
rect 49401 52588 49465 52594
rect 53931 52646 53995 52652
rect 53931 52594 53937 52646
rect 53989 52594 53995 52646
rect 53931 52588 53995 52594
rect -1581 52346 -1535 52351
rect 7181 52346 7227 52351
rect 15943 52346 15989 52351
rect 24705 52346 24751 52351
rect 33467 52346 33513 52351
rect 42229 52346 42275 52351
rect 50991 52346 51037 52351
rect -10352 52340 -10288 52346
rect -10352 52288 -10346 52340
rect -10294 52288 -10288 52340
rect -1590 52340 -1526 52346
rect -1590 52337 -1584 52340
rect -10352 52282 -10288 52288
rect -1595 52288 -1584 52337
rect -1532 52288 -1526 52340
rect 7172 52340 7236 52346
rect 7172 52337 7178 52340
rect -1595 52282 -1526 52288
rect 7167 52288 7178 52337
rect 7230 52288 7236 52340
rect 15934 52340 15998 52346
rect 15934 52337 15940 52340
rect 7167 52282 7236 52288
rect 15929 52288 15940 52337
rect 15992 52288 15998 52340
rect 24696 52340 24760 52346
rect 24696 52337 24702 52340
rect 15929 52282 15998 52288
rect 24691 52288 24702 52337
rect 24754 52288 24760 52340
rect 33458 52340 33522 52346
rect 33458 52337 33464 52340
rect 24691 52282 24760 52288
rect 33453 52288 33464 52337
rect 33516 52288 33522 52340
rect 42220 52340 42284 52346
rect 42220 52337 42226 52340
rect 33453 52282 33522 52288
rect 42215 52288 42226 52337
rect 42278 52288 42284 52340
rect 50982 52340 51046 52346
rect 50982 52337 50988 52340
rect 42215 52282 42284 52288
rect 50987 52288 50988 52337
rect 51040 52288 51046 52340
rect 50987 52282 51046 52288
rect -1595 52049 -1585 52282
rect 7167 52049 7177 52282
rect 15929 52049 15939 52282
rect 24691 52049 24701 52282
rect 33453 52049 33463 52282
rect 42215 52049 42225 52282
rect -12944 51760 57572 51791
rect -12946 51754 57574 51760
rect -12946 51702 -12940 51754
rect -12888 51702 57516 51754
rect 57568 51702 57574 51754
rect -12946 51696 57574 51702
rect -12944 51665 57572 51696
rect -10352 51488 -10288 51494
rect -10352 51436 -10346 51488
rect -10294 51436 -10288 51488
rect -1590 51488 -1526 51494
rect -1590 51485 -1584 51488
rect -1595 51439 -1584 51485
rect -10352 51430 -10288 51436
rect -1590 51436 -1584 51439
rect -1532 51485 -1526 51488
rect 7172 51488 7236 51494
rect 7172 51485 7178 51488
rect -1532 51439 -1521 51485
rect 7167 51439 7178 51485
rect -1532 51436 -1526 51439
rect -1590 51430 -1526 51436
rect 7172 51436 7178 51439
rect 7230 51485 7236 51488
rect 15934 51488 15998 51494
rect 15934 51485 15940 51488
rect 7230 51439 7241 51485
rect 15929 51439 15940 51485
rect 7230 51436 7236 51439
rect 7172 51430 7236 51436
rect 15934 51436 15940 51439
rect 15992 51485 15998 51488
rect 24696 51488 24760 51494
rect 24696 51485 24702 51488
rect 15992 51439 16003 51485
rect 24691 51439 24702 51485
rect 15992 51436 15998 51439
rect 15934 51430 15998 51436
rect 24696 51436 24702 51439
rect 24754 51485 24760 51488
rect 33458 51488 33522 51494
rect 33458 51485 33464 51488
rect 24754 51439 24765 51485
rect 33453 51439 33464 51485
rect 24754 51436 24760 51439
rect 24696 51430 24760 51436
rect 33458 51436 33464 51439
rect 33516 51485 33522 51488
rect 42220 51488 42284 51494
rect 42220 51485 42226 51488
rect 33516 51439 33527 51485
rect 42215 51439 42226 51485
rect 33516 51436 33522 51439
rect 33458 51430 33522 51436
rect 42220 51436 42226 51439
rect 42278 51485 42284 51488
rect 50982 51488 51046 51494
rect 50982 51485 50988 51488
rect 42278 51439 42289 51485
rect 50977 51439 50988 51485
rect 42278 51436 42284 51439
rect 42220 51430 42284 51436
rect 50982 51436 50988 51439
rect 51040 51485 51046 51488
rect 51040 51439 51051 51485
rect 51040 51436 51046 51439
rect 50982 51430 51046 51436
rect -12324 50954 -12260 50960
rect -12324 50902 -12318 50954
rect -12266 50902 -12260 50954
rect -12324 50896 -12260 50902
rect -3562 50954 -3498 50960
rect -3562 50902 -3556 50954
rect -3504 50902 -3498 50954
rect -3562 50896 -3498 50902
rect 5200 50954 5264 50960
rect 5200 50902 5206 50954
rect 5258 50902 5264 50954
rect 5200 50896 5264 50902
rect 13962 50954 14026 50960
rect 13962 50902 13968 50954
rect 14020 50902 14026 50954
rect 13962 50896 14026 50902
rect 22724 50954 22788 50960
rect 22724 50902 22730 50954
rect 22782 50902 22788 50954
rect 22724 50896 22788 50902
rect 31486 50954 31550 50960
rect 31486 50902 31492 50954
rect 31544 50902 31550 50954
rect 31486 50896 31550 50902
rect 40248 50954 40312 50960
rect 40248 50902 40254 50954
rect 40306 50902 40312 50954
rect 40248 50896 40312 50902
rect 49010 50954 49019 50960
rect 49065 50954 49074 50960
rect 49010 50902 49016 50954
rect 49068 50902 49074 50954
rect 49010 50896 49019 50902
rect 49065 50896 49074 50902
rect 49010 50188 49074 50194
rect 49010 50136 49016 50188
rect 49068 50136 49074 50188
rect 49010 50130 49074 50136
rect -12804 49932 -12740 49938
rect -12804 49880 -12798 49932
rect -12746 49929 -12740 49932
rect 57650 49932 57714 49938
rect 57650 49929 57656 49932
rect -12746 49883 -12664 49929
rect 57432 49883 57656 49929
rect -12746 49880 -12740 49883
rect -12804 49874 -12740 49880
rect 57650 49880 57656 49883
rect 57708 49880 57714 49932
rect 57650 49874 57714 49880
rect 51726 49676 51790 49682
rect 51726 49624 51732 49676
rect 51784 49624 51790 49676
rect 51726 49618 51790 49624
rect 57510 48150 57574 48156
rect 57510 48147 57516 48150
rect 57432 48101 57516 48147
rect 57510 48098 57516 48101
rect 57568 48098 57574 48150
rect 57510 48092 57574 48098
rect -12804 47012 -12740 47018
rect -12804 46960 -12798 47012
rect -12746 47009 -12740 47012
rect 50235 47012 50299 47018
rect 50235 47009 50241 47012
rect -12746 46963 7640 47009
rect 37174 46963 50241 47009
rect -12746 46960 -12740 46963
rect -12804 46954 -12740 46960
rect 50235 46960 50241 46963
rect 50293 47009 50299 47012
rect 55667 47012 55731 47018
rect 55667 47009 55673 47012
rect 50293 46963 55673 47009
rect 50293 46960 50299 46963
rect 50235 46954 50299 46960
rect 55667 46960 55673 46963
rect 55725 47009 55731 47012
rect 57650 47012 57714 47018
rect 57650 47009 57656 47012
rect 55725 46963 57656 47009
rect 55725 46960 55731 46963
rect 55667 46954 55731 46960
rect 57650 46960 57656 46963
rect 57708 46960 57714 47012
rect 57650 46954 57714 46960
rect 8855 46202 8919 46208
rect 8855 46150 8861 46202
rect 8913 46150 8919 46202
rect 12799 46202 12863 46208
rect 12799 46199 12805 46202
rect 12794 46153 12805 46199
rect 8855 46144 8919 46150
rect 12799 46150 12805 46153
rect 12857 46199 12863 46202
rect 16743 46202 16807 46208
rect 16743 46199 16749 46202
rect 12857 46153 12868 46199
rect 16738 46153 16749 46199
rect 12857 46150 12863 46153
rect 12799 46144 12863 46150
rect 16743 46150 16749 46153
rect 16801 46199 16807 46202
rect 20687 46202 20751 46208
rect 20687 46199 20693 46202
rect 16801 46153 16812 46199
rect 20682 46153 20693 46199
rect 16801 46150 16807 46153
rect 16743 46144 16807 46150
rect 20687 46150 20693 46153
rect 20745 46199 20751 46202
rect 24631 46202 24695 46208
rect 24631 46199 24637 46202
rect 20745 46153 20756 46199
rect 24626 46153 24637 46199
rect 20745 46150 20751 46153
rect 20687 46144 20751 46150
rect 24631 46150 24637 46153
rect 24689 46199 24695 46202
rect 28575 46202 28639 46208
rect 28575 46199 28581 46202
rect 24689 46153 24700 46199
rect 28570 46153 28581 46199
rect 24689 46150 24695 46153
rect 24631 46144 24695 46150
rect 28575 46150 28581 46153
rect 28633 46199 28639 46202
rect 32519 46202 32583 46208
rect 32519 46199 32525 46202
rect 28633 46153 28644 46199
rect 32514 46153 32525 46199
rect 28633 46150 28639 46153
rect 28575 46144 28639 46150
rect 32519 46150 32525 46153
rect 32577 46199 32583 46202
rect 36463 46202 36527 46208
rect 36463 46199 36469 46202
rect 32577 46153 32588 46199
rect 36458 46153 36469 46199
rect 32577 46150 32583 46153
rect 32519 46144 32583 46150
rect 36463 46150 36469 46153
rect 36521 46199 36527 46202
rect 36521 46153 36532 46199
rect 36521 46150 36527 46153
rect 36463 46144 36527 46150
rect -12946 45230 -12882 45236
rect -12946 45178 -12940 45230
rect -12888 45227 -12882 45230
rect 57510 45230 57574 45236
rect 57510 45227 57516 45230
rect -12888 45181 1445 45227
rect 42366 45181 57516 45227
rect -12888 45178 -12882 45181
rect -12946 45172 -12882 45178
rect 57510 45178 57516 45181
rect 57568 45178 57574 45230
rect 57510 45172 57574 45178
rect 55667 42090 55731 42096
rect 55667 42038 55673 42090
rect 55725 42038 55731 42090
rect 55667 42032 55731 42038
rect 50235 41563 50241 41615
rect 50293 41563 50299 41615
rect 50226 10356 55345 10402
<< via1 >>
rect 50610 55809 50662 55861
rect -12798 53524 -12746 53576
rect 57656 53524 57708 53576
rect -7174 53268 -7122 53320
rect -6560 53268 -6508 53320
rect 1588 53268 1640 53320
rect 2202 53268 2254 53320
rect 10350 53268 10402 53320
rect 10964 53268 11016 53320
rect 19112 53268 19164 53320
rect 19726 53268 19778 53320
rect 27874 53268 27926 53320
rect 28488 53268 28540 53320
rect 36636 53268 36688 53320
rect 37250 53268 37302 53320
rect 45398 53268 45450 53320
rect 46012 53268 46064 53320
rect 54160 53268 54212 53320
rect 54774 53267 54826 53319
rect -11313 52852 -11261 52904
rect -2551 52852 -2499 52904
rect 6211 52852 6263 52904
rect 14973 52852 15025 52904
rect 23735 52852 23787 52904
rect 32497 52852 32549 52904
rect 41259 52852 41311 52904
rect 50021 52852 50073 52904
rect -11927 52594 -11875 52646
rect -7397 52594 -7345 52646
rect -3165 52594 -3113 52646
rect 1365 52594 1417 52646
rect 5597 52594 5649 52646
rect 10127 52594 10179 52646
rect 14359 52594 14411 52646
rect 18889 52594 18941 52646
rect 23121 52594 23173 52646
rect 27651 52594 27703 52646
rect 31883 52594 31935 52646
rect 36413 52594 36465 52646
rect 40645 52594 40697 52646
rect 45175 52594 45227 52646
rect 49407 52594 49459 52646
rect 53937 52594 53989 52646
rect -10346 52288 -10294 52340
rect -1584 52288 -1532 52340
rect 7178 52288 7230 52340
rect 15940 52288 15992 52340
rect 24702 52288 24754 52340
rect 33464 52288 33516 52340
rect 42226 52288 42278 52340
rect 50988 52288 51040 52340
rect -12940 51702 -12888 51754
rect 57516 51702 57568 51754
rect -10346 51436 -10294 51488
rect -1584 51436 -1532 51488
rect 7178 51436 7230 51488
rect 15940 51436 15992 51488
rect 24702 51436 24754 51488
rect 33464 51436 33516 51488
rect 42226 51436 42278 51488
rect 50988 51436 51040 51488
rect -12318 50902 -12266 50954
rect -3556 50902 -3504 50954
rect 5206 50902 5258 50954
rect 13968 50902 14020 50954
rect 22730 50902 22782 50954
rect 31492 50902 31544 50954
rect 40254 50902 40306 50954
rect 49016 50902 49068 50954
rect 49016 50136 49068 50188
rect -12798 49880 -12746 49932
rect 57656 49880 57708 49932
rect 51732 49624 51784 49676
rect 57516 48098 57568 48150
rect -12798 46960 -12746 47012
rect 50241 46960 50293 47012
rect 55673 46960 55725 47012
rect 57656 46960 57708 47012
rect 8861 46150 8913 46202
rect 12805 46150 12857 46202
rect 16749 46150 16801 46202
rect 20693 46150 20745 46202
rect 24637 46150 24689 46202
rect 28581 46150 28633 46202
rect 32525 46150 32577 46202
rect 36469 46150 36521 46202
rect -12940 45178 -12888 45230
rect 57516 45178 57568 45230
rect 55673 42038 55725 42090
rect 50241 41563 50293 41615
<< metal2 >>
rect 51944 61738 52018 61747
rect 51944 61682 51953 61738
rect 52009 61733 52018 61738
rect 57645 61738 57719 61747
rect 57645 61733 57654 61738
rect 52009 61687 57654 61733
rect 52009 61682 52018 61687
rect 51944 61673 52018 61682
rect 57645 61682 57654 61687
rect 57710 61682 57719 61738
rect 57645 61673 57719 61682
rect -12809 61589 -12735 61598
rect -12809 61533 -12800 61589
rect -12744 61584 -12735 61589
rect -7291 61589 -7217 61598
rect -7291 61584 -7282 61589
rect -12744 61538 -7282 61584
rect -12744 61533 -12735 61538
rect -12809 61524 -12735 61533
rect -7291 61533 -7282 61538
rect -7226 61533 -7217 61589
rect -7291 61524 -7217 61533
rect 50599 55863 50673 55872
rect 50599 55807 50608 55863
rect 50664 55807 50673 55863
rect 50599 55798 50673 55807
rect -12809 53578 -12735 53587
rect -12809 53522 -12800 53578
rect -12744 53522 -12735 53578
rect -12809 53513 -12735 53522
rect 57645 53576 57719 53587
rect 57645 53524 57656 53576
rect 57708 53524 57719 53576
rect 57645 53513 57719 53524
rect -7185 53322 -7111 53331
rect -7185 53266 -7176 53322
rect -7120 53266 -7111 53322
rect -7185 53257 -7111 53266
rect -6571 53322 -6497 53331
rect -6571 53266 -6562 53322
rect -6506 53266 -6497 53322
rect -6571 53257 -6497 53266
rect 1577 53322 1651 53331
rect 1577 53266 1586 53322
rect 1642 53266 1651 53322
rect 1577 53257 1651 53266
rect 2191 53322 2265 53331
rect 2191 53266 2200 53322
rect 2256 53266 2265 53322
rect 2191 53257 2265 53266
rect 10339 53322 10413 53331
rect 10339 53266 10348 53322
rect 10404 53266 10413 53322
rect 10339 53257 10413 53266
rect 10953 53322 11027 53331
rect 10953 53266 10962 53322
rect 11018 53266 11027 53322
rect 10953 53257 11027 53266
rect 19101 53322 19175 53331
rect 19101 53266 19110 53322
rect 19166 53266 19175 53322
rect 19101 53257 19175 53266
rect 19715 53322 19789 53331
rect 19715 53266 19724 53322
rect 19780 53266 19789 53322
rect 19715 53257 19789 53266
rect 27863 53322 27937 53331
rect 27863 53266 27872 53322
rect 27928 53266 27937 53322
rect 27863 53257 27937 53266
rect 28477 53322 28551 53331
rect 28477 53266 28486 53322
rect 28542 53266 28551 53322
rect 28477 53257 28551 53266
rect 36625 53322 36699 53331
rect 36625 53266 36634 53322
rect 36690 53266 36699 53322
rect 36625 53257 36699 53266
rect 37239 53322 37313 53331
rect 37239 53266 37248 53322
rect 37304 53266 37313 53322
rect 37239 53257 37313 53266
rect 45387 53322 45461 53331
rect 45387 53266 45396 53322
rect 45452 53266 45461 53322
rect 45387 53257 45461 53266
rect 46001 53322 46075 53331
rect 46001 53266 46010 53322
rect 46066 53266 46075 53322
rect 46001 53257 46075 53266
rect 54149 53322 54223 53331
rect 54149 53266 54158 53322
rect 54214 53266 54223 53322
rect 54149 53257 54223 53266
rect 54763 53321 54837 53330
rect 54763 53265 54772 53321
rect 54828 53265 54837 53321
rect 54763 53256 54837 53265
rect -11319 52904 -11255 52910
rect -11319 52901 -11313 52904
rect -11355 52855 -11313 52901
rect -11319 52852 -11313 52855
rect -11261 52901 -11255 52904
rect -2557 52904 -2493 52910
rect -2557 52901 -2551 52904
rect -11261 52855 -2551 52901
rect -11261 52852 -11255 52855
rect -11319 52846 -11255 52852
rect -2557 52852 -2551 52855
rect -2499 52901 -2493 52904
rect 6205 52904 6269 52910
rect 6205 52901 6211 52904
rect -2499 52855 6211 52901
rect -2499 52852 -2493 52855
rect -2557 52846 -2493 52852
rect 6205 52852 6211 52855
rect 6263 52901 6269 52904
rect 14967 52904 15031 52910
rect 14967 52901 14973 52904
rect 6263 52855 14973 52901
rect 6263 52852 6269 52855
rect 6205 52846 6269 52852
rect 14967 52852 14973 52855
rect 15025 52901 15031 52904
rect 19343 52906 19417 52915
rect 19343 52901 19352 52906
rect 15025 52855 19352 52901
rect 15025 52852 15031 52855
rect 14967 52846 15031 52852
rect 19343 52850 19352 52855
rect 19408 52901 19417 52906
rect 23729 52904 23793 52910
rect 23729 52901 23735 52904
rect 19408 52855 23735 52901
rect 19408 52850 19417 52855
rect 19343 52841 19417 52850
rect 23729 52852 23735 52855
rect 23787 52901 23793 52904
rect 32491 52904 32555 52910
rect 32491 52901 32497 52904
rect 23787 52855 32497 52901
rect 23787 52852 23793 52855
rect 23729 52846 23793 52852
rect 32491 52852 32497 52855
rect 32549 52901 32555 52904
rect 41253 52904 41317 52910
rect 41253 52901 41259 52904
rect 32549 52855 41259 52901
rect 32549 52852 32555 52855
rect 32491 52846 32555 52852
rect 41253 52852 41259 52855
rect 41311 52901 41317 52904
rect 50015 52904 50079 52910
rect 50015 52901 50021 52904
rect 41311 52855 50021 52901
rect 41311 52852 41317 52855
rect 41253 52846 41317 52852
rect 50015 52852 50021 52855
rect 50073 52901 50079 52904
rect 50073 52855 50115 52901
rect 50073 52852 50079 52855
rect 50015 52846 50079 52852
rect -11933 52646 -11869 52652
rect -11933 52594 -11927 52646
rect -11875 52643 -11869 52646
rect -7403 52646 -7339 52652
rect -7403 52643 -7397 52646
rect -11875 52597 -7397 52643
rect -11875 52594 -11869 52597
rect -11933 52588 -11869 52594
rect -7403 52594 -7397 52597
rect -7345 52594 -7339 52646
rect -7403 52588 -7339 52594
rect -3171 52646 -3107 52652
rect -3171 52594 -3165 52646
rect -3113 52643 -3107 52646
rect 1359 52646 1423 52652
rect 1359 52643 1365 52646
rect -3113 52597 1365 52643
rect -3113 52594 -3107 52597
rect -3171 52588 -3107 52594
rect 1359 52594 1365 52597
rect 1417 52594 1423 52646
rect 1359 52588 1423 52594
rect 5591 52646 5655 52652
rect 5591 52594 5597 52646
rect 5649 52643 5655 52646
rect 10121 52646 10185 52652
rect 10121 52643 10127 52646
rect 5649 52597 10127 52643
rect 5649 52594 5655 52597
rect 5591 52588 5655 52594
rect 10121 52594 10127 52597
rect 10179 52594 10185 52646
rect 10121 52588 10185 52594
rect 14353 52646 14417 52652
rect 14353 52594 14359 52646
rect 14411 52643 14417 52646
rect 18883 52646 18947 52652
rect 18883 52643 18889 52646
rect 14411 52597 18889 52643
rect 14411 52594 14417 52597
rect 14353 52588 14417 52594
rect 18883 52594 18889 52597
rect 18941 52594 18947 52646
rect 18883 52588 18947 52594
rect 23115 52646 23179 52652
rect 23115 52594 23121 52646
rect 23173 52643 23179 52646
rect 27645 52646 27709 52652
rect 27645 52643 27651 52646
rect 23173 52597 27651 52643
rect 23173 52594 23179 52597
rect 23115 52588 23179 52594
rect 27645 52594 27651 52597
rect 27703 52594 27709 52646
rect 27645 52588 27709 52594
rect 31877 52646 31941 52652
rect 31877 52594 31883 52646
rect 31935 52643 31941 52646
rect 36407 52646 36471 52652
rect 36407 52643 36413 52646
rect 31935 52597 36413 52643
rect 31935 52594 31941 52597
rect 31877 52588 31941 52594
rect 36407 52594 36413 52597
rect 36465 52594 36471 52646
rect 36407 52588 36471 52594
rect 40639 52646 40703 52652
rect 40639 52594 40645 52646
rect 40697 52643 40703 52646
rect 45169 52646 45233 52652
rect 45169 52643 45175 52646
rect 40697 52597 45175 52643
rect 40697 52594 40703 52597
rect 40639 52588 40703 52594
rect 45169 52594 45175 52597
rect 45227 52594 45233 52646
rect 45169 52588 45233 52594
rect 49401 52646 49465 52652
rect 49401 52594 49407 52646
rect 49459 52643 49465 52646
rect 53931 52646 53995 52652
rect 53931 52643 53937 52646
rect 49459 52597 53937 52643
rect 49459 52594 49465 52597
rect 49401 52588 49465 52594
rect 53931 52594 53937 52597
rect 53989 52594 53995 52646
rect 53931 52588 53995 52594
rect -10357 52342 -10283 52351
rect -10357 52286 -10348 52342
rect -10292 52286 -10283 52342
rect -10357 52277 -10283 52286
rect -1595 52342 -1521 52351
rect -1595 52286 -1586 52342
rect -1530 52286 -1521 52342
rect -1595 52277 -1521 52286
rect 7167 52342 7241 52351
rect 7167 52286 7176 52342
rect 7232 52286 7241 52342
rect 7167 52277 7241 52286
rect 15929 52342 16003 52351
rect 15929 52286 15938 52342
rect 15994 52286 16003 52342
rect 15929 52277 16003 52286
rect 24691 52342 24765 52351
rect 24691 52286 24700 52342
rect 24756 52286 24765 52342
rect 24691 52277 24765 52286
rect 33453 52342 33527 52351
rect 33453 52286 33462 52342
rect 33518 52286 33527 52342
rect 33453 52277 33527 52286
rect 42215 52342 42289 52351
rect 42215 52286 42224 52342
rect 42280 52286 42289 52342
rect 42215 52277 42289 52286
rect 50977 52342 51051 52351
rect 50977 52286 50986 52342
rect 51042 52286 51051 52342
rect 50977 52277 51051 52286
rect -12951 51756 -12877 51765
rect -12951 51700 -12942 51756
rect -12886 51700 -12877 51756
rect -12951 51691 -12877 51700
rect 57505 51756 57579 51765
rect 57505 51700 57514 51756
rect 57570 51700 57579 51756
rect 57505 51691 57579 51700
rect -10357 51490 -10283 51499
rect -10357 51434 -10348 51490
rect -10292 51434 -10283 51490
rect -10357 51425 -10283 51434
rect -1595 51490 -1521 51499
rect -1595 51434 -1586 51490
rect -1530 51434 -1521 51490
rect -1595 51425 -1521 51434
rect 7167 51490 7241 51499
rect 7167 51434 7176 51490
rect 7232 51434 7241 51490
rect 7167 51425 7241 51434
rect 15929 51490 16003 51499
rect 15929 51434 15938 51490
rect 15994 51434 16003 51490
rect 15929 51425 16003 51434
rect 24691 51490 24765 51499
rect 24691 51434 24700 51490
rect 24756 51434 24765 51490
rect 24691 51425 24765 51434
rect 33453 51490 33527 51499
rect 33453 51434 33462 51490
rect 33518 51434 33527 51490
rect 33453 51425 33527 51434
rect 42215 51490 42289 51499
rect 42215 51434 42224 51490
rect 42280 51434 42289 51490
rect 42215 51425 42289 51434
rect 50977 51490 51051 51499
rect 50977 51434 50986 51490
rect 51042 51434 51051 51490
rect 50977 51425 51051 51434
rect -12324 50954 -12260 50960
rect -12324 50951 -12318 50954
rect -12432 50905 -12318 50951
rect -12324 50902 -12318 50905
rect -12266 50951 -12260 50954
rect -3562 50954 -3498 50960
rect -3562 50951 -3556 50954
rect -12266 50905 -3556 50951
rect -12266 50902 -12260 50905
rect -12324 50896 -12260 50902
rect -3562 50902 -3556 50905
rect -3504 50951 -3498 50954
rect 5200 50954 5264 50960
rect 5200 50951 5206 50954
rect -3504 50905 5206 50951
rect -3504 50902 -3498 50905
rect -3562 50896 -3498 50902
rect 5200 50902 5206 50905
rect 5258 50951 5264 50954
rect 13962 50954 14026 50960
rect 13962 50951 13968 50954
rect 5258 50905 13968 50951
rect 5258 50902 5264 50905
rect 5200 50896 5264 50902
rect 13962 50902 13968 50905
rect 14020 50951 14026 50954
rect 22724 50954 22788 50960
rect 22724 50951 22730 50954
rect 14020 50905 22730 50951
rect 14020 50902 14026 50905
rect 13962 50896 14026 50902
rect 22724 50902 22730 50905
rect 22782 50951 22788 50954
rect 31486 50954 31550 50960
rect 31486 50951 31492 50954
rect 22782 50905 31492 50951
rect 22782 50902 22788 50905
rect 22724 50896 22788 50902
rect 31486 50902 31492 50905
rect 31544 50951 31550 50954
rect 40248 50954 40312 50960
rect 40248 50951 40254 50954
rect 31544 50905 40254 50951
rect 31544 50902 31550 50905
rect 31486 50896 31550 50902
rect 40248 50902 40254 50905
rect 40306 50951 40312 50954
rect 49010 50954 49074 50960
rect 49010 50951 49016 50954
rect 40306 50905 49016 50951
rect 40306 50902 40312 50905
rect 40248 50896 40312 50902
rect 49010 50902 49016 50905
rect 49068 50951 49074 50954
rect 49068 50905 49182 50951
rect 49068 50902 49074 50905
rect 49010 50896 49074 50902
rect 49005 50190 49079 50199
rect 49005 50134 49014 50190
rect 49070 50134 49079 50190
rect 49005 50125 49079 50134
rect -11265 50052 -11191 50061
rect -11265 49996 -11256 50052
rect -11200 50047 -11191 50052
rect -2503 50052 -2429 50061
rect -2503 50047 -2494 50052
rect -11200 50001 -2494 50047
rect -11200 49996 -11191 50001
rect -11265 49987 -11191 49996
rect -2503 49996 -2494 50001
rect -2438 50047 -2429 50052
rect 6259 50052 6333 50061
rect 6259 50047 6268 50052
rect -2438 50001 6268 50047
rect -2438 49996 -2429 50001
rect -2503 49987 -2429 49996
rect 6259 49996 6268 50001
rect 6324 50047 6333 50052
rect 15021 50052 15095 50061
rect 15021 50047 15030 50052
rect 6324 50001 15030 50047
rect 6324 49996 6333 50001
rect 6259 49987 6333 49996
rect 15021 49996 15030 50001
rect 15086 50047 15095 50052
rect 23783 50052 23857 50061
rect 23783 50047 23792 50052
rect 15086 50001 23792 50047
rect 15086 49996 15095 50001
rect 15021 49987 15095 49996
rect 23783 49996 23792 50001
rect 23848 50047 23857 50052
rect 32545 50052 32619 50061
rect 32545 50047 32554 50052
rect 23848 50001 32554 50047
rect 23848 49996 23857 50001
rect 23783 49987 23857 49996
rect 32545 49996 32554 50001
rect 32610 50047 32619 50052
rect 41307 50052 41381 50061
rect 41307 50047 41316 50052
rect 32610 50001 41316 50047
rect 32610 49996 32619 50001
rect 32545 49987 32619 49996
rect 41307 49996 41316 50001
rect 41372 50047 41381 50052
rect 49920 50052 49994 50061
rect 49920 50047 49929 50052
rect 41372 50001 49929 50047
rect 41372 49996 41381 50001
rect 41307 49987 41381 49996
rect 49920 49996 49929 50001
rect 49985 50047 49994 50052
rect 49985 50001 50087 50047
rect 49985 49996 49994 50001
rect 49920 49987 49994 49996
rect -12809 49934 -12735 49943
rect -12809 49878 -12800 49934
rect -12744 49878 -12735 49934
rect -12809 49869 -12735 49878
rect 57645 49932 57719 49943
rect 57645 49880 57656 49932
rect 57708 49880 57719 49932
rect 57645 49869 57719 49880
rect 51721 49678 51795 49687
rect 51721 49622 51730 49678
rect 51786 49622 51795 49678
rect 51721 49613 51795 49622
rect 57505 48152 57579 48161
rect 57505 48096 57514 48152
rect 57570 48096 57579 48152
rect 57505 48087 57579 48096
rect -12809 47014 -12735 47023
rect -12809 46958 -12800 47014
rect -12744 46958 -12735 47014
rect -12809 46949 -12735 46958
rect 50230 47014 50304 47023
rect 50230 46958 50239 47014
rect 50295 46958 50304 47014
rect 50230 46949 50304 46958
rect 55662 47014 55736 47023
rect 55662 46958 55671 47014
rect 55727 46958 55736 47014
rect 55662 46949 55736 46958
rect 57645 47014 57719 47023
rect 57645 46958 57654 47014
rect 57710 46958 57719 47014
rect 57645 46949 57719 46958
rect 8850 46204 8924 46213
rect 8850 46148 8859 46204
rect 8915 46148 8924 46204
rect 8850 46139 8924 46148
rect 12794 46204 12868 46213
rect 12794 46148 12803 46204
rect 12859 46148 12868 46204
rect 12794 46139 12868 46148
rect 16738 46204 16812 46213
rect 16738 46148 16747 46204
rect 16803 46148 16812 46204
rect 16738 46139 16812 46148
rect 20682 46204 20756 46213
rect 20682 46148 20691 46204
rect 20747 46148 20756 46204
rect 20682 46139 20756 46148
rect 24626 46204 24700 46213
rect 24626 46148 24635 46204
rect 24691 46148 24700 46204
rect 24626 46139 24700 46148
rect 28570 46204 28644 46213
rect 28570 46148 28579 46204
rect 28635 46148 28644 46204
rect 28570 46139 28644 46148
rect 32514 46204 32588 46213
rect 32514 46148 32523 46204
rect 32579 46148 32588 46204
rect 32514 46139 32588 46148
rect 36458 46204 36532 46213
rect 36458 46148 36467 46204
rect 36523 46148 36532 46204
rect 36458 46139 36532 46148
rect -12951 45232 -12877 45241
rect -12951 45176 -12942 45232
rect -12886 45176 -12877 45232
rect -12951 45167 -12877 45176
rect 57505 45232 57579 45241
rect 57505 45176 57514 45232
rect 57570 45176 57579 45232
rect 57505 45167 57579 45176
rect 55662 42092 55736 42101
rect 55662 42036 55671 42092
rect 55727 42036 55736 42092
rect 55662 42027 55736 42036
rect 50237 41619 50297 41628
rect 50237 41550 50297 41559
rect 49005 29325 49079 29334
rect 49005 29269 49014 29325
rect 49070 29320 49079 29325
rect 49070 29274 50070 29320
rect 49070 29269 49079 29274
rect 49005 29260 49079 29269
<< via2 >>
rect 51953 61682 52009 61738
rect 57654 61682 57710 61738
rect -12800 61533 -12744 61589
rect -7282 61533 -7226 61589
rect 50608 55861 50664 55863
rect 50608 55809 50610 55861
rect 50610 55809 50662 55861
rect 50662 55809 50664 55861
rect 50608 55807 50664 55809
rect -12800 53576 -12744 53578
rect -12800 53524 -12798 53576
rect -12798 53524 -12746 53576
rect -12746 53524 -12744 53576
rect -12800 53522 -12744 53524
rect -7176 53320 -7120 53322
rect -7176 53268 -7174 53320
rect -7174 53268 -7122 53320
rect -7122 53268 -7120 53320
rect -7176 53266 -7120 53268
rect -6562 53320 -6506 53322
rect -6562 53268 -6560 53320
rect -6560 53268 -6508 53320
rect -6508 53268 -6506 53320
rect -6562 53266 -6506 53268
rect 1586 53320 1642 53322
rect 1586 53268 1588 53320
rect 1588 53268 1640 53320
rect 1640 53268 1642 53320
rect 1586 53266 1642 53268
rect 2200 53320 2256 53322
rect 2200 53268 2202 53320
rect 2202 53268 2254 53320
rect 2254 53268 2256 53320
rect 2200 53266 2256 53268
rect 10348 53320 10404 53322
rect 10348 53268 10350 53320
rect 10350 53268 10402 53320
rect 10402 53268 10404 53320
rect 10348 53266 10404 53268
rect 10962 53320 11018 53322
rect 10962 53268 10964 53320
rect 10964 53268 11016 53320
rect 11016 53268 11018 53320
rect 10962 53266 11018 53268
rect 19110 53320 19166 53322
rect 19110 53268 19112 53320
rect 19112 53268 19164 53320
rect 19164 53268 19166 53320
rect 19110 53266 19166 53268
rect 19724 53320 19780 53322
rect 19724 53268 19726 53320
rect 19726 53268 19778 53320
rect 19778 53268 19780 53320
rect 19724 53266 19780 53268
rect 27872 53320 27928 53322
rect 27872 53268 27874 53320
rect 27874 53268 27926 53320
rect 27926 53268 27928 53320
rect 27872 53266 27928 53268
rect 28486 53320 28542 53322
rect 28486 53268 28488 53320
rect 28488 53268 28540 53320
rect 28540 53268 28542 53320
rect 28486 53266 28542 53268
rect 36634 53320 36690 53322
rect 36634 53268 36636 53320
rect 36636 53268 36688 53320
rect 36688 53268 36690 53320
rect 36634 53266 36690 53268
rect 37248 53320 37304 53322
rect 37248 53268 37250 53320
rect 37250 53268 37302 53320
rect 37302 53268 37304 53320
rect 37248 53266 37304 53268
rect 45396 53320 45452 53322
rect 45396 53268 45398 53320
rect 45398 53268 45450 53320
rect 45450 53268 45452 53320
rect 45396 53266 45452 53268
rect 46010 53320 46066 53322
rect 46010 53268 46012 53320
rect 46012 53268 46064 53320
rect 46064 53268 46066 53320
rect 46010 53266 46066 53268
rect 54158 53320 54214 53322
rect 54158 53268 54160 53320
rect 54160 53268 54212 53320
rect 54212 53268 54214 53320
rect 54158 53266 54214 53268
rect 54772 53319 54828 53321
rect 54772 53267 54774 53319
rect 54774 53267 54826 53319
rect 54826 53267 54828 53319
rect 54772 53265 54828 53267
rect 19352 52850 19408 52906
rect -10348 52340 -10292 52342
rect -10348 52288 -10346 52340
rect -10346 52288 -10294 52340
rect -10294 52288 -10292 52340
rect -10348 52286 -10292 52288
rect -1586 52340 -1530 52342
rect -1586 52288 -1584 52340
rect -1584 52288 -1532 52340
rect -1532 52288 -1530 52340
rect -1586 52286 -1530 52288
rect 7176 52340 7232 52342
rect 7176 52288 7178 52340
rect 7178 52288 7230 52340
rect 7230 52288 7232 52340
rect 7176 52286 7232 52288
rect 15938 52340 15994 52342
rect 15938 52288 15940 52340
rect 15940 52288 15992 52340
rect 15992 52288 15994 52340
rect 15938 52286 15994 52288
rect 24700 52340 24756 52342
rect 24700 52288 24702 52340
rect 24702 52288 24754 52340
rect 24754 52288 24756 52340
rect 24700 52286 24756 52288
rect 33462 52340 33518 52342
rect 33462 52288 33464 52340
rect 33464 52288 33516 52340
rect 33516 52288 33518 52340
rect 33462 52286 33518 52288
rect 42224 52340 42280 52342
rect 42224 52288 42226 52340
rect 42226 52288 42278 52340
rect 42278 52288 42280 52340
rect 42224 52286 42280 52288
rect 50986 52340 51042 52342
rect 50986 52288 50988 52340
rect 50988 52288 51040 52340
rect 51040 52288 51042 52340
rect 50986 52286 51042 52288
rect -12942 51754 -12886 51756
rect -12942 51702 -12940 51754
rect -12940 51702 -12888 51754
rect -12888 51702 -12886 51754
rect -12942 51700 -12886 51702
rect 57514 51754 57570 51756
rect 57514 51702 57516 51754
rect 57516 51702 57568 51754
rect 57568 51702 57570 51754
rect 57514 51700 57570 51702
rect -10348 51488 -10292 51490
rect -10348 51436 -10346 51488
rect -10346 51436 -10294 51488
rect -10294 51436 -10292 51488
rect -10348 51434 -10292 51436
rect -1586 51488 -1530 51490
rect -1586 51436 -1584 51488
rect -1584 51436 -1532 51488
rect -1532 51436 -1530 51488
rect -1586 51434 -1530 51436
rect 7176 51488 7232 51490
rect 7176 51436 7178 51488
rect 7178 51436 7230 51488
rect 7230 51436 7232 51488
rect 7176 51434 7232 51436
rect 15938 51488 15994 51490
rect 15938 51436 15940 51488
rect 15940 51436 15992 51488
rect 15992 51436 15994 51488
rect 15938 51434 15994 51436
rect 24700 51488 24756 51490
rect 24700 51436 24702 51488
rect 24702 51436 24754 51488
rect 24754 51436 24756 51488
rect 24700 51434 24756 51436
rect 33462 51488 33518 51490
rect 33462 51436 33464 51488
rect 33464 51436 33516 51488
rect 33516 51436 33518 51488
rect 33462 51434 33518 51436
rect 42224 51488 42280 51490
rect 42224 51436 42226 51488
rect 42226 51436 42278 51488
rect 42278 51436 42280 51488
rect 42224 51434 42280 51436
rect 50986 51488 51042 51490
rect 50986 51436 50988 51488
rect 50988 51436 51040 51488
rect 51040 51436 51042 51488
rect 50986 51434 51042 51436
rect 49014 50188 49070 50190
rect 49014 50136 49016 50188
rect 49016 50136 49068 50188
rect 49068 50136 49070 50188
rect 49014 50134 49070 50136
rect -11256 49996 -11200 50052
rect -2494 49996 -2438 50052
rect 6268 49996 6324 50052
rect 15030 49996 15086 50052
rect 23792 49996 23848 50052
rect 32554 49996 32610 50052
rect 41316 49996 41372 50052
rect 49929 49996 49985 50052
rect -12800 49932 -12744 49934
rect -12800 49880 -12798 49932
rect -12798 49880 -12746 49932
rect -12746 49880 -12744 49932
rect -12800 49878 -12744 49880
rect 51730 49676 51786 49678
rect 51730 49624 51732 49676
rect 51732 49624 51784 49676
rect 51784 49624 51786 49676
rect 51730 49622 51786 49624
rect 57514 48150 57570 48152
rect 57514 48098 57516 48150
rect 57516 48098 57568 48150
rect 57568 48098 57570 48150
rect 57514 48096 57570 48098
rect -12800 47012 -12744 47014
rect -12800 46960 -12798 47012
rect -12798 46960 -12746 47012
rect -12746 46960 -12744 47012
rect -12800 46958 -12744 46960
rect 50239 47012 50295 47014
rect 50239 46960 50241 47012
rect 50241 46960 50293 47012
rect 50293 46960 50295 47012
rect 50239 46958 50295 46960
rect 55671 47012 55727 47014
rect 55671 46960 55673 47012
rect 55673 46960 55725 47012
rect 55725 46960 55727 47012
rect 55671 46958 55727 46960
rect 57654 47012 57710 47014
rect 57654 46960 57656 47012
rect 57656 46960 57708 47012
rect 57708 46960 57710 47012
rect 57654 46958 57710 46960
rect 8859 46202 8915 46204
rect 8859 46150 8861 46202
rect 8861 46150 8913 46202
rect 8913 46150 8915 46202
rect 8859 46148 8915 46150
rect 12803 46202 12859 46204
rect 12803 46150 12805 46202
rect 12805 46150 12857 46202
rect 12857 46150 12859 46202
rect 12803 46148 12859 46150
rect 16747 46202 16803 46204
rect 16747 46150 16749 46202
rect 16749 46150 16801 46202
rect 16801 46150 16803 46202
rect 16747 46148 16803 46150
rect 20691 46202 20747 46204
rect 20691 46150 20693 46202
rect 20693 46150 20745 46202
rect 20745 46150 20747 46202
rect 20691 46148 20747 46150
rect 24635 46202 24691 46204
rect 24635 46150 24637 46202
rect 24637 46150 24689 46202
rect 24689 46150 24691 46202
rect 24635 46148 24691 46150
rect 28579 46202 28635 46204
rect 28579 46150 28581 46202
rect 28581 46150 28633 46202
rect 28633 46150 28635 46202
rect 28579 46148 28635 46150
rect 32523 46202 32579 46204
rect 32523 46150 32525 46202
rect 32525 46150 32577 46202
rect 32577 46150 32579 46202
rect 32523 46148 32579 46150
rect 36467 46202 36523 46204
rect 36467 46150 36469 46202
rect 36469 46150 36521 46202
rect 36521 46150 36523 46202
rect 36467 46148 36523 46150
rect -12942 45230 -12886 45232
rect -12942 45178 -12940 45230
rect -12940 45178 -12888 45230
rect -12888 45178 -12886 45230
rect -12942 45176 -12886 45178
rect 57514 45230 57570 45232
rect 57514 45178 57516 45230
rect 57516 45178 57568 45230
rect 57568 45178 57570 45230
rect 57514 45176 57570 45178
rect 55671 42090 55727 42092
rect 55671 42038 55673 42090
rect 55673 42038 55725 42090
rect 55725 42038 55727 42090
rect 55671 42036 55727 42038
rect 50237 41615 50297 41619
rect 50237 41563 50241 41615
rect 50241 41563 50293 41615
rect 50293 41563 50297 41615
rect 50237 41559 50297 41563
rect 49014 29269 49070 29325
<< metal3 >>
rect -6944 62908 -1886 62968
rect 52642 62908 57572 62968
rect -12944 51761 -12884 62908
rect 51948 61740 52014 61743
rect -6421 61680 47040 61740
rect 47100 61680 48171 61740
rect 51669 61738 52014 61740
rect 51669 61682 51953 61738
rect 52009 61682 52014 61738
rect 51669 61680 52014 61682
rect 51948 61677 52014 61680
rect -12805 61589 -12739 61594
rect -12805 61533 -12800 61589
rect -12744 61533 -12739 61589
rect -12805 61528 -12739 61533
rect -7287 61591 -7221 61594
rect -7287 61589 -6974 61591
rect -7287 61533 -7282 61589
rect -7226 61533 -6974 61589
rect -7287 61531 -6974 61533
rect -7287 61528 -7221 61531
rect -12802 53583 -12742 61528
rect -6421 60623 47040 60683
rect 47100 60623 51181 60683
rect -4548 54476 -2183 54536
rect -984 54476 1381 54536
rect 2580 54476 4945 54536
rect 6144 54476 8509 54536
rect 9708 54476 12073 54536
rect 13272 54476 15637 54536
rect 16836 54476 19201 54536
rect -3396 53837 -3336 54476
rect -6572 53831 -6496 53837
rect -6572 53767 -6566 53831
rect -6502 53767 -6496 53831
rect -6572 53761 -6496 53767
rect -3404 53831 -3328 53837
rect -3404 53767 -3398 53831
rect -3334 53767 -3328 53831
rect -3404 53761 -3328 53767
rect -2653 53831 -2577 53837
rect -2653 53767 -2647 53831
rect -2583 53767 -2577 53831
rect -2653 53761 -2577 53767
rect -11415 53703 -11339 53709
rect -11415 53639 -11409 53703
rect -11345 53639 -11339 53703
rect -11415 53633 -11339 53639
rect -7186 53703 -7110 53709
rect -7186 53639 -7180 53703
rect -7116 53639 -7110 53703
rect -7186 53633 -7110 53639
rect -12805 53578 -12739 53583
rect -12805 53522 -12800 53578
rect -12744 53522 -12739 53578
rect -12805 53517 -12739 53522
rect -12947 51756 -12881 51761
rect -12947 51700 -12942 51756
rect -12886 51700 -12881 51756
rect -12947 51695 -12881 51700
rect -12944 45237 -12884 51695
rect -12802 49939 -12742 53517
rect -11407 50688 -11347 53633
rect -7178 53327 -7118 53633
rect -6564 53327 -6504 53761
rect -7181 53322 -7115 53327
rect -7181 53266 -7176 53322
rect -7120 53266 -7115 53322
rect -7181 53261 -7115 53266
rect -6567 53322 -6501 53327
rect -6567 53266 -6562 53322
rect -6506 53266 -6501 53322
rect -6567 53261 -6501 53266
rect -10353 52342 -10287 52347
rect -10353 52286 -10348 52342
rect -10292 52286 -10287 52342
rect -10353 52281 -10287 52286
rect -10350 51495 -10290 52281
rect -10353 51490 -10287 51495
rect -10353 51434 -10348 51490
rect -10292 51434 -10287 51490
rect -10353 51429 -10287 51434
rect -2645 50687 -2585 53761
rect 168 53709 228 54476
rect 1584 53837 1644 53846
rect 1576 53831 1652 53837
rect 1576 53767 1582 53831
rect 1646 53767 1652 53831
rect 1576 53761 1652 53767
rect 160 53703 236 53709
rect 160 53639 166 53703
rect 230 53639 236 53703
rect 160 53633 236 53639
rect 1584 53327 1644 53761
rect 3732 53709 3792 54476
rect 7296 53837 7356 54476
rect 7288 53831 7364 53837
rect 7288 53767 7294 53831
rect 7358 53767 7364 53831
rect 7288 53761 7364 53767
rect 2190 53703 2266 53709
rect 2190 53639 2196 53703
rect 2260 53639 2266 53703
rect 2190 53633 2266 53639
rect 3724 53703 3800 53709
rect 3724 53639 3730 53703
rect 3794 53639 3800 53703
rect 3724 53633 3800 53639
rect 6109 53703 6185 53709
rect 6109 53639 6115 53703
rect 6179 53639 6185 53703
rect 6109 53633 6185 53639
rect 10338 53703 10414 53709
rect 10338 53639 10344 53703
rect 10408 53639 10414 53703
rect 10338 53633 10414 53639
rect 2198 53327 2258 53633
rect 1581 53322 1647 53327
rect 1581 53266 1586 53322
rect 1642 53266 1647 53322
rect 1581 53261 1647 53266
rect 2195 53322 2261 53327
rect 2195 53266 2200 53322
rect 2256 53266 2261 53322
rect 2195 53261 2261 53266
rect -1591 52342 -1525 52347
rect -1591 52286 -1586 52342
rect -1530 52286 -1525 52342
rect -1591 52281 -1525 52286
rect -1588 51495 -1528 52281
rect -1591 51490 -1525 51495
rect -1591 51434 -1586 51490
rect -1530 51434 -1525 51490
rect -1591 51429 -1525 51434
rect 6117 50688 6177 53633
rect 10346 53327 10406 53633
rect 10960 53327 11020 54476
rect 14424 53709 14484 54476
rect 17988 53837 18048 54476
rect 17980 53831 18056 53837
rect 17980 53767 17986 53831
rect 18050 53767 18056 53831
rect 17980 53761 18056 53767
rect 14416 53703 14492 53709
rect 14416 53639 14422 53703
rect 14486 53639 14492 53703
rect 14416 53633 14492 53639
rect 14871 53703 14947 53709
rect 14871 53639 14877 53703
rect 14941 53639 14947 53703
rect 14871 53633 14947 53639
rect 19100 53703 19176 53709
rect 19100 53639 19106 53703
rect 19170 53639 19176 53703
rect 19100 53633 19176 53639
rect 10343 53322 10409 53327
rect 10343 53266 10348 53322
rect 10404 53266 10409 53322
rect 10343 53261 10409 53266
rect 10957 53322 11023 53327
rect 10957 53266 10962 53322
rect 11018 53266 11023 53322
rect 10957 53261 11023 53266
rect 7171 52342 7237 52347
rect 7171 52286 7176 52342
rect 7232 52286 7237 52342
rect 7171 52281 7237 52286
rect 7174 51495 7234 52281
rect 7171 51490 7237 51495
rect 7171 51434 7176 51490
rect 7232 51434 7237 51490
rect 7171 51429 7237 51434
rect 14879 50688 14939 53633
rect 19108 53327 19168 53633
rect 19105 53322 19171 53327
rect 19105 53266 19110 53322
rect 19166 53266 19171 53322
rect 19105 53261 19171 53266
rect 19350 52911 19410 60623
rect 28680 54536 28740 54655
rect 50064 54536 50124 56231
rect 50603 55865 50669 55868
rect 50603 55863 51788 55865
rect 50603 55807 50608 55863
rect 50664 55807 51788 55863
rect 50603 55805 51788 55807
rect 50603 55802 50669 55805
rect 20400 54476 22765 54536
rect 23964 54476 26329 54536
rect 27528 54476 29893 54536
rect 31092 54476 33457 54536
rect 34656 54476 37021 54536
rect 38220 54476 40585 54536
rect 41784 54476 44149 54536
rect 45348 54476 47713 54536
rect 48912 54476 51277 54536
rect 19714 53831 19790 53837
rect 19714 53767 19720 53831
rect 19784 53767 19790 53831
rect 19714 53761 19790 53767
rect 19722 53327 19782 53761
rect 21552 53709 21612 54476
rect 25116 53837 25176 54476
rect 25108 53831 25184 53837
rect 25108 53767 25114 53831
rect 25178 53767 25184 53831
rect 25108 53761 25184 53767
rect 28476 53831 28552 53837
rect 28476 53767 28482 53831
rect 28546 53767 28552 53831
rect 28476 53761 28552 53767
rect 27870 53709 27930 53720
rect 21544 53703 21620 53709
rect 21544 53639 21550 53703
rect 21614 53639 21620 53703
rect 21544 53633 21620 53639
rect 23633 53703 23709 53709
rect 23633 53639 23639 53703
rect 23703 53639 23709 53703
rect 23633 53633 23709 53639
rect 27862 53703 27938 53709
rect 27862 53639 27868 53703
rect 27932 53639 27938 53703
rect 27862 53633 27938 53639
rect 19719 53322 19785 53327
rect 19719 53266 19724 53322
rect 19780 53266 19785 53322
rect 19719 53261 19785 53266
rect 19347 52906 19413 52911
rect 19347 52850 19352 52906
rect 19408 52850 19413 52906
rect 19347 52845 19413 52850
rect 15933 52342 15999 52347
rect 15933 52286 15938 52342
rect 15994 52286 15999 52342
rect 15933 52281 15999 52286
rect 15936 51495 15996 52281
rect 15933 51490 15999 51495
rect 15933 51434 15938 51490
rect 15994 51434 15999 51490
rect 15933 51429 15999 51434
rect 23641 50688 23701 53633
rect 27870 53327 27930 53633
rect 28484 53327 28544 53761
rect 28680 53709 28740 54476
rect 32244 53837 32304 54476
rect 32236 53831 32312 53837
rect 32236 53767 32242 53831
rect 32306 53767 32312 53831
rect 32236 53761 32312 53767
rect 35808 53709 35868 54476
rect 39372 53837 39432 54476
rect 37238 53831 37314 53837
rect 37238 53767 37244 53831
rect 37308 53767 37314 53831
rect 37238 53761 37314 53767
rect 39364 53831 39440 53837
rect 39364 53767 39370 53831
rect 39434 53767 39440 53831
rect 39364 53761 39440 53767
rect 28672 53703 28748 53709
rect 28672 53639 28678 53703
rect 28742 53639 28748 53703
rect 28672 53633 28748 53639
rect 32395 53703 32471 53709
rect 32395 53639 32401 53703
rect 32465 53639 32471 53703
rect 32395 53633 32471 53639
rect 35800 53703 35876 53709
rect 35800 53639 35806 53703
rect 35870 53639 35876 53703
rect 35800 53633 35876 53639
rect 36624 53703 36700 53709
rect 36624 53639 36630 53703
rect 36694 53639 36700 53703
rect 36624 53633 36700 53639
rect 27867 53322 27933 53327
rect 27867 53266 27872 53322
rect 27928 53266 27933 53322
rect 27867 53261 27933 53266
rect 28481 53322 28547 53327
rect 28481 53266 28486 53322
rect 28542 53266 28547 53322
rect 28481 53261 28547 53266
rect 24695 52342 24761 52347
rect 24695 52286 24700 52342
rect 24756 52286 24761 52342
rect 24695 52281 24761 52286
rect 24698 51495 24758 52281
rect 24695 51490 24761 51495
rect 24695 51434 24700 51490
rect 24756 51434 24761 51490
rect 24695 51429 24761 51434
rect 32403 50688 32463 53633
rect 36632 53327 36692 53633
rect 37246 53327 37306 53761
rect 42936 53709 42996 54476
rect 46500 53837 46560 54476
rect 46000 53831 46076 53837
rect 46000 53767 46006 53831
rect 46070 53767 46076 53831
rect 46000 53761 46076 53767
rect 46492 53831 46568 53837
rect 46492 53767 46498 53831
rect 46562 53767 46568 53831
rect 46492 53761 46568 53767
rect 41157 53703 41233 53709
rect 41157 53639 41163 53703
rect 41227 53639 41233 53703
rect 41157 53633 41233 53639
rect 42928 53703 43004 53709
rect 42928 53639 42934 53703
rect 42998 53639 43004 53703
rect 42928 53633 43004 53639
rect 45386 53703 45462 53709
rect 45386 53639 45392 53703
rect 45456 53639 45462 53703
rect 45386 53633 45462 53639
rect 36629 53322 36695 53327
rect 36629 53266 36634 53322
rect 36690 53266 36695 53322
rect 36629 53261 36695 53266
rect 37243 53322 37309 53327
rect 37243 53266 37248 53322
rect 37304 53266 37309 53322
rect 37243 53261 37309 53266
rect 33457 52342 33523 52347
rect 33457 52286 33462 52342
rect 33518 52286 33523 52342
rect 33457 52281 33523 52286
rect 33460 51495 33520 52281
rect 33457 51490 33523 51495
rect 33457 51434 33462 51490
rect 33518 51434 33523 51490
rect 33457 51429 33523 51434
rect 41165 50688 41225 53633
rect 45394 53327 45454 53633
rect 46008 53327 46068 53761
rect 50064 53709 50124 54476
rect 49919 53703 49995 53709
rect 49919 53639 49925 53703
rect 49989 53639 49995 53703
rect 49919 53633 49995 53639
rect 50056 53703 50132 53709
rect 50056 53639 50062 53703
rect 50126 53639 50132 53703
rect 50056 53633 50132 53639
rect 45391 53322 45457 53327
rect 45391 53266 45396 53322
rect 45452 53266 45457 53322
rect 45391 53261 45457 53266
rect 46005 53322 46071 53327
rect 46005 53266 46010 53322
rect 46066 53266 46071 53322
rect 46005 53261 46071 53266
rect 45394 53064 45454 53261
rect 46008 53064 46068 53261
rect 42219 52342 42285 52347
rect 42219 52286 42224 52342
rect 42280 52286 42285 52342
rect 42219 52281 42285 52286
rect 42222 51495 42282 52281
rect 42219 51490 42285 51495
rect 42219 51434 42224 51490
rect 42280 51434 42285 51490
rect 42219 51429 42285 51434
rect 49927 50688 49987 53633
rect 50981 52342 51047 52347
rect 50981 52286 50986 52342
rect 51042 52286 51047 52342
rect 50981 52281 51047 52286
rect 50984 51495 51044 52281
rect 50981 51490 51047 51495
rect 50981 51434 50986 51490
rect 51042 51434 51047 51490
rect 50981 51429 51047 51434
rect 49009 50190 49075 50195
rect 49009 50134 49014 50190
rect 49070 50134 49075 50190
rect 49009 50129 49075 50134
rect 6266 50057 6326 50061
rect 15028 50057 15088 50061
rect 23790 50057 23850 50061
rect 32552 50057 32612 50061
rect 41314 50057 41374 50061
rect -11261 50052 -11195 50057
rect -11261 49996 -11256 50052
rect -11200 49996 -11195 50052
rect -11261 49991 -11195 49996
rect -2499 49991 -2496 50057
rect -2436 49991 -2433 50057
rect 6263 50052 6329 50057
rect 6263 49996 6268 50052
rect 6324 49996 6329 50052
rect 6263 49991 6329 49996
rect 15025 50052 15091 50057
rect 15025 49996 15030 50052
rect 15086 49996 15091 50052
rect 15025 49991 15091 49996
rect 23787 50052 23853 50057
rect 23787 49996 23792 50052
rect 23848 49996 23853 50052
rect 23787 49991 23853 49996
rect 32549 50052 32615 50057
rect 32549 49996 32554 50052
rect 32610 49996 32615 50052
rect 32549 49991 32615 49996
rect 41311 50052 41377 50057
rect 41311 49996 41316 50052
rect 41372 49996 41377 50052
rect 41311 49991 41377 49996
rect 6266 49987 6326 49991
rect 15028 49987 15088 49991
rect 23790 49987 23850 49991
rect 32552 49987 32612 49991
rect 41314 49987 41374 49991
rect -12805 49934 -12739 49939
rect -12805 49878 -12800 49934
rect -12744 49878 -12739 49934
rect -12805 49873 -12739 49878
rect -12802 47019 -12742 49873
rect -4203 47145 -4143 49678
rect 4559 47273 4619 49678
rect 13321 47401 13381 49678
rect 22083 47529 22143 49678
rect 28569 47779 28645 47785
rect 28569 47715 28575 47779
rect 28639 47715 28645 47779
rect 28569 47709 28645 47715
rect 24625 47651 24701 47657
rect 24625 47587 24631 47651
rect 24695 47587 24701 47651
rect 24625 47581 24701 47587
rect 20681 47523 20757 47529
rect 20681 47459 20687 47523
rect 20751 47459 20757 47523
rect 20681 47453 20757 47459
rect 22075 47523 22151 47529
rect 22075 47459 22081 47523
rect 22145 47459 22151 47523
rect 22075 47453 22151 47459
rect 13313 47395 13389 47401
rect 13313 47331 13319 47395
rect 13383 47331 13389 47395
rect 13313 47325 13389 47331
rect 16737 47395 16813 47401
rect 16737 47331 16743 47395
rect 16807 47331 16813 47395
rect 16737 47325 16813 47331
rect 4551 47267 4627 47273
rect 4551 47203 4557 47267
rect 4621 47203 4627 47267
rect 4551 47197 4627 47203
rect 12793 47267 12869 47273
rect 12793 47203 12799 47267
rect 12863 47203 12869 47267
rect 12793 47197 12869 47203
rect -4211 47139 -4135 47145
rect -4211 47075 -4205 47139
rect -4141 47075 -4135 47139
rect -4211 47069 -4135 47075
rect 8849 47139 8925 47145
rect 8849 47075 8855 47139
rect 8919 47075 8925 47139
rect 8849 47069 8925 47075
rect -12805 47014 -12739 47019
rect -12805 46958 -12800 47014
rect -12744 46958 -12739 47014
rect -12805 46953 -12739 46958
rect 8857 46209 8917 47069
rect 12801 46209 12861 47197
rect 16745 46209 16805 47325
rect 20689 46209 20749 47453
rect 24633 46209 24693 47581
rect 28577 46209 28637 47709
rect 30845 47657 30905 49678
rect 36457 48035 36533 48041
rect 36457 47971 36463 48035
rect 36527 47971 36533 48035
rect 36457 47965 36533 47971
rect 32513 47907 32589 47913
rect 32513 47843 32519 47907
rect 32583 47843 32589 47907
rect 32513 47837 32589 47843
rect 30837 47651 30913 47657
rect 30837 47587 30843 47651
rect 30907 47587 30913 47651
rect 30837 47581 30913 47587
rect 32521 46209 32581 47837
rect 36465 46209 36525 47965
rect 39607 47785 39667 49678
rect 48369 47913 48429 49678
rect 48361 47907 48437 47913
rect 48361 47843 48367 47907
rect 48431 47843 48437 47907
rect 48361 47837 48437 47843
rect 39599 47779 39675 47785
rect 39599 47715 39605 47779
rect 39669 47715 39675 47779
rect 39599 47709 39675 47715
rect 8854 46204 8920 46209
rect 8854 46148 8859 46204
rect 8915 46148 8920 46204
rect 8854 46143 8920 46148
rect 12798 46204 12864 46209
rect 12798 46148 12803 46204
rect 12859 46148 12864 46204
rect 12798 46143 12864 46148
rect 16742 46204 16808 46209
rect 16742 46148 16747 46204
rect 16803 46148 16808 46204
rect 16742 46143 16808 46148
rect 20686 46204 20752 46209
rect 20686 46148 20691 46204
rect 20747 46148 20752 46204
rect 20686 46143 20752 46148
rect 24630 46204 24696 46209
rect 24630 46148 24635 46204
rect 24691 46148 24696 46204
rect 24630 46143 24696 46148
rect 28574 46204 28640 46209
rect 28574 46148 28579 46204
rect 28635 46148 28640 46204
rect 28574 46143 28640 46148
rect 32518 46204 32584 46209
rect 32518 46148 32523 46204
rect 32579 46148 32584 46204
rect 32518 46143 32584 46148
rect 36462 46204 36528 46209
rect 36462 46148 36467 46204
rect 36523 46148 36528 46204
rect 36462 46143 36528 46148
rect -12947 45232 -12881 45237
rect -12947 45176 -12942 45232
rect -12886 45176 -12881 45232
rect -12947 45171 -12881 45176
rect 49012 29330 49072 50129
rect 49924 50052 49990 50057
rect 49924 49996 49929 50052
rect 49985 49996 49990 50052
rect 49924 49991 49990 49996
rect 51728 49683 51788 55805
rect 54762 53831 54838 53837
rect 54762 53767 54768 53831
rect 54832 53767 54838 53831
rect 54762 53761 54838 53767
rect 54148 53703 54224 53709
rect 54148 53639 54154 53703
rect 54218 53639 54224 53703
rect 54148 53633 54224 53639
rect 54156 53327 54216 53633
rect 54153 53322 54219 53327
rect 54770 53326 54830 53761
rect 54153 53266 54158 53322
rect 54214 53266 54219 53322
rect 54153 53261 54219 53266
rect 54767 53321 54833 53326
rect 54767 53265 54772 53321
rect 54828 53265 54833 53321
rect 54767 53260 54833 53265
rect 57512 51761 57572 62908
rect 57649 61738 57715 61743
rect 57649 61682 57654 61738
rect 57710 61682 57715 61738
rect 57649 61677 57715 61682
rect 57652 53583 57712 61677
rect 57649 53517 57715 53583
rect 57509 51756 57575 51761
rect 57509 51700 57514 51756
rect 57570 51700 57575 51756
rect 57509 51695 57575 51700
rect 51725 49678 51791 49683
rect 51725 49622 51730 49678
rect 51786 49622 51791 49678
rect 51725 49617 51791 49622
rect 57131 48041 57191 49678
rect 57512 48157 57572 51695
rect 57652 49939 57712 53517
rect 57649 49873 57715 49939
rect 57509 48152 57575 48157
rect 57509 48096 57514 48152
rect 57570 48096 57575 48152
rect 57509 48091 57575 48096
rect 57123 48035 57199 48041
rect 57123 47971 57129 48035
rect 57193 47971 57199 48035
rect 57123 47965 57199 47971
rect 50234 47014 50300 47019
rect 50234 46958 50239 47014
rect 50295 46958 50300 47014
rect 50234 46953 50300 46958
rect 55666 47014 55732 47019
rect 55666 46958 55671 47014
rect 55727 46958 55732 47014
rect 55666 46953 55732 46958
rect 50237 41624 50297 46953
rect 55669 42097 55729 46953
rect 57512 45237 57572 48091
rect 57652 47019 57712 49873
rect 57649 47014 57715 47019
rect 57649 46958 57654 47014
rect 57710 46958 57715 47014
rect 57649 46953 57715 46958
rect 57509 45232 57575 45237
rect 57509 45176 57514 45232
rect 57570 45176 57575 45232
rect 57509 45171 57575 45176
rect 55666 42092 55732 42097
rect 55666 42036 55671 42092
rect 55727 42036 55732 42092
rect 55666 42031 55732 42036
rect 50232 41619 50302 41624
rect 50232 41559 50237 41619
rect 50297 41559 50302 41619
rect 50232 41554 50302 41559
rect 49009 29325 49075 29330
rect 49009 29269 49014 29325
rect 49070 29269 49075 29325
rect 49009 29264 49075 29269
rect 41580 26826 41656 26832
rect 41580 26762 41586 26826
rect 41650 26824 41656 26826
rect 48674 26826 48750 26832
rect 48674 26824 48680 26826
rect 41650 26764 48680 26824
rect 41650 26762 41656 26764
rect 41580 26756 41656 26762
rect 48674 26762 48680 26764
rect 48744 26762 48750 26826
rect 48674 26756 48750 26762
rect 52220 26826 52296 26832
rect 52220 26762 52226 26826
rect 52290 26762 52296 26826
rect 52220 26756 52296 26762
rect 52228 24771 52288 26756
<< via3 >>
rect -6566 53767 -6502 53831
rect -3398 53767 -3334 53831
rect -2647 53767 -2583 53831
rect -11409 53639 -11345 53703
rect -7180 53639 -7116 53703
rect 1582 53767 1646 53831
rect 166 53639 230 53703
rect 7294 53767 7358 53831
rect 2196 53639 2260 53703
rect 3730 53639 3794 53703
rect 6115 53639 6179 53703
rect 10344 53639 10408 53703
rect 17986 53767 18050 53831
rect 14422 53639 14486 53703
rect 14877 53639 14941 53703
rect 19106 53639 19170 53703
rect 19720 53767 19784 53831
rect 25114 53767 25178 53831
rect 28482 53767 28546 53831
rect 21550 53639 21614 53703
rect 23639 53639 23703 53703
rect 27868 53639 27932 53703
rect 32242 53767 32306 53831
rect 37244 53767 37308 53831
rect 39370 53767 39434 53831
rect 28678 53639 28742 53703
rect 32401 53639 32465 53703
rect 35806 53639 35870 53703
rect 36630 53639 36694 53703
rect 46006 53767 46070 53831
rect 46498 53767 46562 53831
rect 41163 53639 41227 53703
rect 42934 53639 42998 53703
rect 45392 53639 45456 53703
rect 49925 53639 49989 53703
rect 50062 53639 50126 53703
rect 28575 47715 28639 47779
rect 24631 47587 24695 47651
rect 20687 47459 20751 47523
rect 22081 47459 22145 47523
rect 13319 47331 13383 47395
rect 16743 47331 16807 47395
rect 4557 47203 4621 47267
rect 12799 47203 12863 47267
rect -4205 47075 -4141 47139
rect 8855 47075 8919 47139
rect 36463 47971 36527 48035
rect 32519 47843 32583 47907
rect 30843 47587 30907 47651
rect 48367 47843 48431 47907
rect 39605 47715 39669 47779
rect 54768 53767 54832 53831
rect 54154 53639 54218 53703
rect 57129 47971 57193 48035
rect 41586 26762 41650 26826
rect 48680 26762 48744 26826
rect 52226 26762 52290 26826
<< metal4 >>
rect -6567 53831 -6501 53832
rect -6567 53767 -6566 53831
rect -6502 53829 -6501 53831
rect -3399 53831 -3333 53832
rect -3399 53829 -3398 53831
rect -6502 53769 -3398 53829
rect -6502 53767 -6501 53769
rect -6567 53766 -6501 53767
rect -3399 53767 -3398 53769
rect -3334 53767 -3333 53831
rect -3399 53766 -3333 53767
rect -2648 53831 -2582 53832
rect -2648 53767 -2647 53831
rect -2583 53829 -2582 53831
rect 1581 53831 1647 53832
rect 1581 53829 1582 53831
rect -2583 53769 1582 53829
rect -2583 53767 -2582 53769
rect -2648 53766 -2582 53767
rect 1581 53767 1582 53769
rect 1646 53829 1647 53831
rect 7293 53831 7359 53832
rect 7293 53829 7294 53831
rect 1646 53769 7294 53829
rect 1646 53767 1647 53769
rect 1581 53766 1647 53767
rect 7293 53767 7294 53769
rect 7358 53767 7359 53831
rect 7293 53766 7359 53767
rect 17985 53831 18051 53832
rect 17985 53767 17986 53831
rect 18050 53829 18051 53831
rect 19719 53831 19785 53832
rect 19719 53829 19720 53831
rect 18050 53769 19720 53829
rect 18050 53767 18051 53769
rect 17985 53766 18051 53767
rect 19719 53767 19720 53769
rect 19784 53767 19785 53831
rect 19719 53766 19785 53767
rect 25113 53831 25179 53832
rect 25113 53767 25114 53831
rect 25178 53829 25179 53831
rect 28481 53831 28547 53832
rect 28481 53829 28482 53831
rect 25178 53769 28482 53829
rect 25178 53767 25179 53769
rect 25113 53766 25179 53767
rect 28481 53767 28482 53769
rect 28546 53767 28547 53831
rect 28481 53766 28547 53767
rect 32241 53831 32307 53832
rect 32241 53767 32242 53831
rect 32306 53829 32307 53831
rect 37243 53831 37309 53832
rect 37243 53829 37244 53831
rect 32306 53769 37244 53829
rect 32306 53767 32307 53769
rect 32241 53766 32307 53767
rect 37243 53767 37244 53769
rect 37308 53767 37309 53831
rect 37243 53766 37309 53767
rect 39369 53831 39435 53832
rect 39369 53767 39370 53831
rect 39434 53829 39435 53831
rect 46005 53831 46071 53832
rect 46005 53829 46006 53831
rect 39434 53769 46006 53829
rect 39434 53767 39435 53769
rect 39369 53766 39435 53767
rect 46005 53767 46006 53769
rect 46070 53767 46071 53831
rect 46005 53766 46071 53767
rect 46497 53831 46563 53832
rect 46497 53767 46498 53831
rect 46562 53829 46563 53831
rect 54767 53831 54833 53832
rect 54767 53829 54768 53831
rect 46562 53769 54768 53829
rect 46562 53767 46563 53769
rect 46497 53766 46563 53767
rect 54767 53767 54768 53769
rect 54832 53767 54833 53831
rect 54767 53766 54833 53767
rect -11410 53703 -11344 53704
rect -11410 53639 -11409 53703
rect -11345 53701 -11344 53703
rect -7181 53703 -7115 53704
rect -7181 53701 -7180 53703
rect -11345 53641 -7180 53701
rect -11345 53639 -11344 53641
rect -11410 53638 -11344 53639
rect -7181 53639 -7180 53641
rect -7116 53701 -7115 53703
rect 165 53703 231 53704
rect 165 53701 166 53703
rect -7116 53641 166 53701
rect -7116 53639 -7115 53641
rect -7181 53638 -7115 53639
rect 165 53639 166 53641
rect 230 53639 231 53703
rect 165 53638 231 53639
rect 2195 53703 2261 53704
rect 2195 53639 2196 53703
rect 2260 53701 2261 53703
rect 3729 53703 3795 53704
rect 3729 53701 3730 53703
rect 2260 53641 3730 53701
rect 2260 53639 2261 53641
rect 2195 53638 2261 53639
rect 3729 53639 3730 53641
rect 3794 53639 3795 53703
rect 3729 53638 3795 53639
rect 6114 53703 6180 53704
rect 6114 53639 6115 53703
rect 6179 53701 6180 53703
rect 10343 53703 10409 53704
rect 10343 53701 10344 53703
rect 6179 53641 10344 53701
rect 6179 53639 6180 53641
rect 6114 53638 6180 53639
rect 10343 53639 10344 53641
rect 10408 53701 10409 53703
rect 14421 53703 14487 53704
rect 14421 53701 14422 53703
rect 10408 53641 14422 53701
rect 10408 53639 10409 53641
rect 10343 53638 10409 53639
rect 14421 53639 14422 53641
rect 14486 53639 14487 53703
rect 14421 53638 14487 53639
rect 14876 53703 14942 53704
rect 14876 53639 14877 53703
rect 14941 53701 14942 53703
rect 19105 53703 19171 53704
rect 19105 53701 19106 53703
rect 14941 53641 19106 53701
rect 14941 53639 14942 53641
rect 14876 53638 14942 53639
rect 19105 53639 19106 53641
rect 19170 53701 19171 53703
rect 21549 53703 21615 53704
rect 21549 53701 21550 53703
rect 19170 53641 21550 53701
rect 19170 53639 19171 53641
rect 19105 53638 19171 53639
rect 21549 53639 21550 53641
rect 21614 53639 21615 53703
rect 21549 53638 21615 53639
rect 23638 53703 23704 53704
rect 23638 53639 23639 53703
rect 23703 53701 23704 53703
rect 27867 53703 27933 53704
rect 27867 53701 27868 53703
rect 23703 53641 27868 53701
rect 23703 53639 23704 53641
rect 23638 53638 23704 53639
rect 27867 53639 27868 53641
rect 27932 53701 27933 53703
rect 28677 53703 28743 53704
rect 28677 53701 28678 53703
rect 27932 53641 28678 53701
rect 27932 53639 27933 53641
rect 27867 53638 27933 53639
rect 28677 53639 28678 53641
rect 28742 53639 28743 53703
rect 28677 53638 28743 53639
rect 32400 53703 32466 53704
rect 32400 53639 32401 53703
rect 32465 53701 32466 53703
rect 35805 53703 35871 53704
rect 35805 53701 35806 53703
rect 32465 53641 35806 53701
rect 32465 53639 32466 53641
rect 32400 53638 32466 53639
rect 35805 53639 35806 53641
rect 35870 53701 35871 53703
rect 36629 53703 36695 53704
rect 36629 53701 36630 53703
rect 35870 53641 36630 53701
rect 35870 53639 35871 53641
rect 35805 53638 35871 53639
rect 36629 53639 36630 53641
rect 36694 53639 36695 53703
rect 36629 53638 36695 53639
rect 41162 53703 41228 53704
rect 41162 53639 41163 53703
rect 41227 53701 41228 53703
rect 42933 53703 42999 53704
rect 42933 53701 42934 53703
rect 41227 53641 42934 53701
rect 41227 53639 41228 53641
rect 41162 53638 41228 53639
rect 42933 53639 42934 53641
rect 42998 53701 42999 53703
rect 45391 53703 45457 53704
rect 45391 53701 45392 53703
rect 42998 53641 45392 53701
rect 42998 53639 42999 53641
rect 42933 53638 42999 53639
rect 45391 53639 45392 53641
rect 45456 53639 45457 53703
rect 45391 53638 45457 53639
rect 49924 53703 49990 53704
rect 49924 53639 49925 53703
rect 49989 53701 49990 53703
rect 50061 53703 50127 53704
rect 50061 53701 50062 53703
rect 49989 53641 50062 53701
rect 49989 53639 49990 53641
rect 49924 53638 49990 53639
rect 50061 53639 50062 53641
rect 50126 53701 50127 53703
rect 54153 53703 54219 53704
rect 54153 53701 54154 53703
rect 50126 53641 54154 53701
rect 50126 53639 50127 53641
rect 50061 53638 50127 53639
rect 54153 53639 54154 53641
rect 54218 53639 54219 53703
rect 54153 53638 54219 53639
rect 36462 48035 36528 48036
rect 36462 47971 36463 48035
rect 36527 48033 36528 48035
rect 57128 48035 57194 48036
rect 57128 48033 57129 48035
rect 36527 47973 57129 48033
rect 36527 47971 36528 47973
rect 36462 47970 36528 47971
rect 57128 47971 57129 47973
rect 57193 47971 57194 48035
rect 57128 47970 57194 47971
rect 32518 47907 32584 47908
rect 32518 47843 32519 47907
rect 32583 47905 32584 47907
rect 48366 47907 48432 47908
rect 48366 47905 48367 47907
rect 32583 47845 48367 47905
rect 32583 47843 32584 47845
rect 32518 47842 32584 47843
rect 48366 47843 48367 47845
rect 48431 47843 48432 47907
rect 48366 47842 48432 47843
rect 28574 47779 28640 47780
rect 28574 47715 28575 47779
rect 28639 47777 28640 47779
rect 39604 47779 39670 47780
rect 39604 47777 39605 47779
rect 28639 47717 39605 47777
rect 28639 47715 28640 47717
rect 28574 47714 28640 47715
rect 39604 47715 39605 47717
rect 39669 47715 39670 47779
rect 39604 47714 39670 47715
rect 24630 47651 24696 47652
rect 24630 47587 24631 47651
rect 24695 47649 24696 47651
rect 30842 47651 30908 47652
rect 30842 47649 30843 47651
rect 24695 47589 30843 47649
rect 24695 47587 24696 47589
rect 24630 47586 24696 47587
rect 30842 47587 30843 47589
rect 30907 47587 30908 47651
rect 30842 47586 30908 47587
rect 20686 47523 20752 47524
rect 20686 47459 20687 47523
rect 20751 47521 20752 47523
rect 22080 47523 22146 47524
rect 22080 47521 22081 47523
rect 20751 47461 22081 47521
rect 20751 47459 20752 47461
rect 20686 47458 20752 47459
rect 22080 47459 22081 47461
rect 22145 47459 22146 47523
rect 22080 47458 22146 47459
rect 13318 47395 13384 47396
rect 13318 47331 13319 47395
rect 13383 47393 13384 47395
rect 16742 47395 16808 47396
rect 16742 47393 16743 47395
rect 13383 47333 16743 47393
rect 13383 47331 13384 47333
rect 13318 47330 13384 47331
rect 16742 47331 16743 47333
rect 16807 47331 16808 47395
rect 16742 47330 16808 47331
rect 4556 47267 4622 47268
rect 4556 47203 4557 47267
rect 4621 47265 4622 47267
rect 12798 47267 12864 47268
rect 12798 47265 12799 47267
rect 4621 47205 12799 47265
rect 4621 47203 4622 47205
rect 4556 47202 4622 47203
rect 12798 47203 12799 47205
rect 12863 47203 12864 47267
rect 12798 47202 12864 47203
rect -4206 47139 -4140 47140
rect -4206 47075 -4205 47139
rect -4141 47137 -4140 47139
rect 8854 47139 8920 47140
rect 8854 47137 8855 47139
rect -4141 47077 8855 47137
rect -4141 47075 -4140 47077
rect -4206 47074 -4140 47075
rect 8854 47075 8855 47077
rect 8919 47075 8920 47139
rect 8854 47074 8920 47075
rect 688 42540 44080 42600
rect 41585 26826 41651 26827
rect 41585 26762 41586 26826
rect 41650 26762 41651 26826
rect 41585 26761 41651 26762
rect 48679 26826 48745 26827
rect 48679 26762 48680 26826
rect 48744 26824 48745 26826
rect 52225 26826 52291 26827
rect 52225 26824 52226 26826
rect 48744 26764 52226 26824
rect 48744 26762 48745 26764
rect 48679 26761 48745 26762
rect 52225 26762 52226 26764
rect 52290 26762 52291 26826
rect 52225 26761 52291 26762
rect 41588 25576 41648 26761
rect 41272 25516 41648 25576
<< metal5 >>
rect 51500 20625 51820 20945
use And_Gate  And_Gate_0
timestamp 1757220954
transform 1 0 -10715 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_1
timestamp 1757220954
transform 1 0 -1953 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_2
timestamp 1757220954
transform 1 0 6809 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_3
timestamp 1757220954
transform 1 0 15571 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_4
timestamp 1757220954
transform 1 0 24333 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_5
timestamp 1757220954
transform 1 0 33095 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_6
timestamp 1757220954
transform 1 0 41857 0 1 51955
box -1558 -210 544 1618
use And_Gate  And_Gate_7
timestamp 1757220954
transform 1 0 50619 0 1 51955
box -1558 -210 544 1618
use CDAC_v3  CDAC_v3_0
timestamp 1757231656
transform 1 0 960 0 1 288
box -1004 -280 43852 46735
use Comparator  Comparator_0
timestamp 1756559655
transform -1 0 80195 0 1 12366
box 24473 -2307 30902 29735
use D_FlipFlop  D_FlipFlop_0
timestamp 1757226713
transform 1 0 48670 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_1
timestamp 1757226713
transform 1 0 39908 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1757226713
transform 1 0 31146 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1757226713
transform 1 0 22384 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1757226713
transform 1 0 4860 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1757226713
transform 1 0 13622 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1757226713
transform 1 0 -3902 0 1 49883
box 0 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1757226713
transform 1 0 -12664 0 1 49883
box 0 -1796 8762 1842
use Nand_Gate  Nand_Gate_0
timestamp 1757220954
transform -1 0 4506 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_1
timestamp 1757220954
transform -1 0 -4256 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_2
timestamp 1757220954
transform -1 0 13268 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_3
timestamp 1757220954
transform -1 0 30792 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_4
timestamp 1757220954
transform -1 0 39554 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_5
timestamp 1757220954
transform -1 0 48316 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_6
timestamp 1757220954
transform -1 0 22030 0 1 52275
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_7
timestamp 1757220954
transform -1 0 57078 0 1 52275
box 1906 -530 3264 1298
use Ring_Counter  Ring_Counter_0
timestamp 1757226903
transform 0 1 60854 -1 0 63603
box 606 -68805 9368 -8143
<< labels >>
flabel metal4 -4141 47077 8855 47137 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal4 4621 47205 12799 47265 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal4 13383 47333 16743 47393 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal4 20751 47461 22081 47521 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal4 24695 47589 30843 47649 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal4 28639 47717 39605 47777 0 FreeSans 160 0 0 0 Q5
port 8 nsew
flabel metal4 32583 47845 48367 47905 0 FreeSans 160 0 0 0 Q6
port 9 nsew
flabel metal4 36527 47973 57129 48033 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal4 688 42540 44080 42600 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal5 51500 20625 51820 20945 0 FreeSans 1120 0 0 0 Vin
port 13 nsew
flabel metal1 50226 10356 55345 10402 0 FreeSans 160 0 0 0 Vbias
port 11 nsew
flabel metal3 -6421 61680 47040 61740 0 FreeSans 160 0 0 0 EN
port 1 nsew
flabel metal3 19350 52906 19410 60683 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 57652 47014 57712 61677 0 FreeSans 160 90 0 0 VDD
port 12 nsew
<< end >>
