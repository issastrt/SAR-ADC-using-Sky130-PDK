** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-10-12_02-22-36/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0.000000u 0.242266 8.500000u 0.242266 8.500001u 0.230851 17.000000u 0.230851 17.000001u 0.215262 25.500000u
+ 0.215262 25.500001u 0.231873 34.000000u 0.231873 34.000001u 0.258920 42.500000u 0.258920 42.500001u 0.331710 51.000000u 0.331710
+ 51.000001u 0.359779 59.500000u 0.359779 59.500001u 0.354582 68.000000u 0.354582 68.000001u 0.328601 76.500000u 0.328601 76.500001u 0.295336
+ 85.000000u 0.295336 85.000001u 0.301555 93.500000u 0.301555 93.500001u 0.331710 102.000000u 0.331710 102.000001u 0.337971 110.500000u
+ 0.337971 110.500001u 0.373323 119.000000u 0.373323 119.000001u 0.382651 127.500000u 0.382651 127.500001u 0.377454 136.000000u 0.377454
+ 136.000001u 0.366040 144.500000u 0.366040 144.500001u 0.343167 153.000000u 0.343167 153.000001u 0.369149 161.500000u 0.369149 161.500001u
+ 0.398282 170.000000u 0.398282)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=-40
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 170u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-10-12_02-22-36/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
