magic
tech sky130A
magscale 1 2
timestamp 1757220954
<< metal1 >>
rect -1558 1572 544 1618
rect -1209 414 -1163 946
rect -595 414 -549 946
rect -372 642 195 688
rect 372 336 418 1033
rect -1558 -210 544 -164
use Inverter  Inverter_0
timestamp 1757220954
transform 1 0 -1566 0 1 676
box 1366 -886 2110 942
use Nand_Gate  Nand_Gate_0
timestamp 1757220954
transform 1 0 -3464 0 1 320
box 1906 -530 3264 1298
<< labels >>
flabel metal1 -1558 -210 544 -164 0 FreeSans 160 0 0 0 GND
port 0 nsew
flabel metal1 -1558 1572 544 1618 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 -1209 414 -1163 946 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 -595 414 -549 946 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal1 372 336 418 1033 0 FreeSans 160 90 0 0 Vout
port 4 nsew
<< end >>
