** sch_path: /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_20-48-13/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 0.557647058750 8.5u 0.557647058750 8.500001u 0.559411764625 17u 0.559411764625 17.000001u 0.561176470500 25.5u
+ 0.561176470500 25.500001u 0.562941176375 34u 0.562941176375 34.000001u 0.564705882250 42.5u 0.564705882250 42.500001u 0.566470588125 51u
+ 0.566470588125 51.000001u 0.568235294000 59.5u 0.568235294000 59.500001u 0.570000000000 68u 0.570000000000 68.000001u 0.571764705875 76.5u
+ 0.571764705875 76.500001u 0.573529411750 85u 0.573529411750 85.000001u 0.575294117625 93.5u 0.575294117625 93.500001u 0.577058823500 102u
+ 0.577058823500 102.000001u 0.578823529375 110.5u 0.578823529375 110.500001u 0.580588235250 119u 0.580588235250 119.000001u 0.582352941125 127.5u
+ 0.582352941125 127.500001u 0.584117647000 136u 0.584117647000 136.000001u 0.585882352875 144.5u 0.585882352875 144.500001u 0.587647058750 153u
+ 0.587647058750 153.000001u 0.589411764625 161.5u 0.589411764625 161.500001u 0.591176470500 170u 0.591176470500 170.000001u 0.592941176375 178.5u
+ 0.592941176375 178.500001u 0.594705882250 187u 0.594705882250 187.000001u 0.596470588125 195.5u 0.596470588125 195.500001u 0.598235294000 204u
+ 0.598235294000 204.000001u 0.600000000000 212.5u 0.600000000000 212.500001u 0.601764705875 221u 0.601764705875 221.000001u 0.603529411750 229.5u
+ 0.603529411750 229.500001u 0.605294117625 238u 0.605294117625 238.000001u 0.607058823500 246.5u 0.607058823500 246.500001u 0.608823529375 255u
+ 0.608823529375 255.000001u 0.610588235250 263.5u 0.610588235250 263.500001u 0.612352941125 272u 0.612352941125 272.000001u 0.614117647000 280.5u
+ 0.614117647000 280.500001u 0.615882352875 289u 0.615882352875 289.000001u 0.617647058750 297.5u 0.617647058750 297.500001u 0.619411764625 306u
+ 0.619411764625 306.000001u 0.621176470500 314.5u 0.621176470500 314.500001u 0.622941176375 323u 0.622941176375 323.000001u 0.624705882250 331.5u
+ 0.624705882250 331.500001u 0.626470588125 340u 0.626470588125 340.000001u 0.628235294000 348.5u 0.628235294000 348.500001u 0.630000000000 357u
+ 0.630000000000 357.000001u 0.631764705875 365.5u 0.631764705875 365.500001u 0.633529411750 374u 0.633529411750 374.000001u 0.635294117625 382.5u
+ 0.635294117625 382.500001u 0.637058823500 391u 0.637058823500 391.000001u 0.638823529375 399.5u 0.638823529375 399.500001u 0.640588235250 408u
+ 0.640588235250 408.000001u 0.642352941125 416.5u 0.642352941125 416.500001u 0.644117647000 425u 0.644117647000 425.000001u 0.645882352875 433.5u
+ 0.645882352875 433.500001u 0.647647058750 442u 0.647647058750 442.000001u 0.649411764625 450.5u 0.649411764625 450.500001u 0.651176470500 459u
+ 0.651176470500 459.000001u 0.652941176375 467.5u 0.652941176375 467.500001u 0.654705882250 476u 0.654705882250 476.000001u 0.656470588125 484.5u
+ 0.656470588125 484.500001u 0.658235294000 493u 0.658235294000 493.000001u 0.660000000000 501.5u 0.660000000000 501.500001u 0.661764705875 510u
+ 0.661764705875 510.000001u 0.663529411750 518.5u 0.663529411750 518.500001u 0.665294117625 527u 0.665294117625 527.000001u 0.667058823500 535.5u
+ 0.667058823500 535.500001u 0.668823529375 544u 0.668823529375 544.000001u 0.670588235250 552.5u 0.670588235250 552.500001u 0.672352941125 561u
+ 0.672352941125 561.000001u 0.674117647000 569.5u 0.674117647000 569.500001u 0.675882352875 578u 0.675882352875 578.000001u 0.677647058750 586.5u
+ 0.677647058750 586.500001u 0.679411764625 595u 0.679411764625 595.000001u 0.681176470500 603.5u 0.681176470500 603.500001u 0.682941176375 612u
+ 0.682941176375 612.000001u 0.684705882250 620.5u 0.684705882250 620.500001u 0.686470588125 629u 0.686470588125 629.000001u 0.688235294000 637.5u
+ 0.688235294000 637.500001u 0.690000000000 646u 0.690000000000 646.000001u 0.691764705875 654.5u 0.691764705875 654.500001u 0.693529411750 663u
+ 0.693529411750 663.000001u 0.695294117625 671.5u 0.695294117625 671.500001u 0.697058823500 680u 0.697058823500)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/samantha/cace/SAR-ADC-using-Sky130-PDK/netlist/schematic/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 680u uic
  wrdata /home/samantha/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-02_20-48-13/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
