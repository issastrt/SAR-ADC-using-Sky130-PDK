magic
tech sky130A
magscale 1 2
timestamp 1755761378
<< metal1 >>
rect 11040 36583 97170 36629
rect 19709 35780 19773 35786
rect 19709 35728 19715 35780
rect 19767 35728 19773 35780
rect 19709 35722 19773 35728
rect 22508 35780 22572 35786
rect 22508 35728 22514 35780
rect 22566 35728 22572 35780
rect 22508 35722 22572 35728
rect 30749 35780 30813 35786
rect 30749 35728 30755 35780
rect 30807 35728 30813 35780
rect 30749 35722 30813 35728
rect 33548 35780 33612 35786
rect 33548 35728 33554 35780
rect 33606 35728 33612 35780
rect 33548 35722 33612 35728
rect 41789 35780 41853 35786
rect 41789 35728 41795 35780
rect 41847 35728 41853 35780
rect 41789 35722 41853 35728
rect 44588 35780 44652 35786
rect 44588 35728 44594 35780
rect 44646 35728 44652 35780
rect 44588 35722 44652 35728
rect 52829 35780 52893 35786
rect 52829 35728 52835 35780
rect 52887 35728 52893 35780
rect 52829 35722 52893 35728
rect 55628 35780 55692 35786
rect 55628 35728 55634 35780
rect 55686 35728 55692 35780
rect 55628 35722 55692 35728
rect 63869 35780 63933 35786
rect 63869 35728 63875 35780
rect 63927 35728 63933 35780
rect 63869 35722 63933 35728
rect 66668 35780 66732 35786
rect 66668 35728 66674 35780
rect 66726 35728 66732 35780
rect 66668 35722 66732 35728
rect 74909 35780 74973 35786
rect 74909 35728 74915 35780
rect 74967 35728 74973 35780
rect 74909 35722 74973 35728
rect 77708 35780 77772 35786
rect 77708 35728 77714 35780
rect 77766 35728 77772 35780
rect 77708 35722 77772 35728
rect 85949 35780 86013 35786
rect 85949 35728 85955 35780
rect 86007 35728 86013 35780
rect 85949 35722 86013 35728
rect 88748 35780 88812 35786
rect 88748 35728 88754 35780
rect 88806 35728 88812 35780
rect 88748 35722 88812 35728
rect 87549 34850 87613 34856
rect 87549 34847 87555 34850
rect 11128 34801 87555 34847
rect 87549 34798 87555 34801
rect 87607 34847 87613 34850
rect 87607 34801 97170 34847
rect 87607 34798 87613 34801
rect 87549 34792 87613 34798
rect 96766 33294 96830 33300
rect 96766 33242 96772 33294
rect 96824 33242 96830 33294
rect 96766 33236 96830 33242
rect 86765 33068 86829 33074
rect 86765 33065 86771 33068
rect 11040 33019 86771 33065
rect 86765 33016 86771 33019
rect 86823 33065 86829 33068
rect 86823 33019 97170 33065
rect 86823 33016 86829 33019
rect 86765 33010 86829 33016
rect 86765 3613 86829 3619
rect 86765 3610 86771 3613
rect 88 3564 86771 3610
rect 86765 3561 86771 3564
rect 86823 3610 86829 3613
rect 86823 3564 97198 3610
rect 86823 3561 86829 3564
rect 86765 3555 86829 3561
rect 1656 3387 1720 3393
rect 1656 3335 1662 3387
rect 1714 3335 1720 3387
rect 1656 3329 1720 3335
rect 12696 3387 12760 3393
rect 12696 3335 12702 3387
rect 12754 3335 12760 3387
rect 12696 3329 12760 3335
rect 23736 3387 23800 3393
rect 23736 3335 23742 3387
rect 23794 3335 23800 3387
rect 23736 3329 23800 3335
rect 34776 3387 34840 3393
rect 34776 3335 34782 3387
rect 34834 3335 34840 3387
rect 34776 3329 34840 3335
rect 45816 3387 45880 3393
rect 45816 3335 45822 3387
rect 45874 3335 45880 3387
rect 45816 3329 45880 3335
rect 56856 3387 56920 3393
rect 56856 3335 56862 3387
rect 56914 3335 56920 3387
rect 56856 3329 56920 3335
rect 67896 3387 67960 3393
rect 67896 3335 67902 3387
rect 67954 3335 67960 3387
rect 67896 3329 67960 3335
rect 78936 3387 79000 3393
rect 78936 3335 78942 3387
rect 78994 3335 79000 3387
rect 78936 3329 79000 3335
rect 89976 3387 90040 3393
rect 89976 3335 89982 3387
rect 90034 3335 90040 3387
rect 89976 3329 90040 3335
rect 96766 3387 96830 3393
rect 96766 3335 96772 3387
rect 96824 3335 96830 3387
rect 96766 3329 96830 3335
rect 8446 2761 8510 2767
rect 8446 2709 8452 2761
rect 8504 2709 8510 2761
rect 8446 2703 8510 2709
rect 11245 2761 11309 2767
rect 11245 2709 11251 2761
rect 11303 2709 11309 2761
rect 11245 2703 11309 2709
rect 19486 2761 19550 2767
rect 19486 2709 19492 2761
rect 19544 2709 19550 2761
rect 19486 2703 19550 2709
rect 22285 2761 22349 2767
rect 22285 2709 22291 2761
rect 22343 2709 22349 2761
rect 22285 2703 22349 2709
rect 30526 2761 30590 2767
rect 30526 2709 30532 2761
rect 30584 2709 30590 2761
rect 30526 2703 30590 2709
rect 33325 2761 33389 2767
rect 33325 2709 33331 2761
rect 33383 2709 33389 2761
rect 33325 2703 33389 2709
rect 41566 2761 41630 2767
rect 41566 2709 41572 2761
rect 41624 2709 41630 2761
rect 41566 2703 41630 2709
rect 44365 2761 44429 2767
rect 44365 2709 44371 2761
rect 44423 2709 44429 2761
rect 44365 2703 44429 2709
rect 52606 2761 52670 2767
rect 52606 2709 52612 2761
rect 52664 2709 52670 2761
rect 52606 2703 52670 2709
rect 55405 2761 55469 2767
rect 55405 2709 55411 2761
rect 55463 2709 55469 2761
rect 55405 2703 55469 2709
rect 63646 2761 63710 2767
rect 63646 2709 63652 2761
rect 63704 2709 63710 2761
rect 63646 2703 63710 2709
rect 66445 2761 66509 2767
rect 66445 2709 66451 2761
rect 66503 2709 66509 2761
rect 66445 2703 66509 2709
rect 74686 2761 74750 2767
rect 74686 2709 74692 2761
rect 74744 2709 74750 2761
rect 74686 2703 74750 2709
rect 77485 2761 77549 2767
rect 77485 2709 77491 2761
rect 77543 2709 77549 2761
rect 77485 2703 77549 2709
rect 85726 2761 85790 2767
rect 85726 2709 85732 2761
rect 85784 2709 85790 2761
rect 85726 2703 85790 2709
rect 88525 2761 88589 2767
rect 88525 2709 88531 2761
rect 88583 2709 88589 2761
rect 88525 2703 88589 2709
rect 5730 1831 5794 1837
rect 5730 1828 5736 1831
rect 88 1782 5736 1828
rect 5730 1779 5736 1782
rect 5788 1828 5794 1831
rect 16770 1831 16834 1837
rect 16770 1828 16776 1831
rect 5788 1782 16776 1828
rect 5788 1779 5794 1782
rect 5730 1773 5794 1779
rect 16770 1779 16776 1782
rect 16828 1828 16834 1831
rect 27810 1831 27874 1837
rect 27810 1828 27816 1831
rect 16828 1782 27816 1828
rect 16828 1779 16834 1782
rect 16770 1773 16834 1779
rect 27810 1779 27816 1782
rect 27868 1828 27874 1831
rect 38850 1831 38914 1837
rect 38850 1828 38856 1831
rect 27868 1782 38856 1828
rect 27868 1779 27874 1782
rect 27810 1773 27874 1779
rect 38850 1779 38856 1782
rect 38908 1828 38914 1831
rect 49890 1831 49954 1837
rect 49890 1828 49896 1831
rect 38908 1782 49896 1828
rect 38908 1779 38914 1782
rect 38850 1773 38914 1779
rect 49890 1779 49896 1782
rect 49948 1828 49954 1831
rect 60930 1831 60994 1837
rect 60930 1828 60936 1831
rect 49948 1782 60936 1828
rect 49948 1779 49954 1782
rect 49890 1773 49954 1779
rect 60930 1779 60936 1782
rect 60988 1828 60994 1831
rect 71970 1831 72034 1837
rect 71970 1828 71976 1831
rect 60988 1782 71976 1828
rect 60988 1779 60994 1782
rect 60930 1773 60994 1779
rect 71970 1779 71976 1782
rect 72028 1828 72034 1831
rect 83010 1831 83074 1837
rect 83010 1828 83016 1831
rect 72028 1782 83016 1828
rect 72028 1779 72034 1782
rect 71970 1773 72034 1779
rect 83010 1779 83016 1782
rect 83068 1828 83074 1831
rect 87549 1831 87613 1837
rect 87549 1828 87555 1831
rect 83068 1782 87555 1828
rect 83068 1779 83074 1782
rect 83010 1773 83074 1779
rect 87549 1779 87555 1782
rect 87607 1828 87613 1831
rect 94050 1831 94114 1837
rect 94050 1828 94056 1831
rect 87607 1782 94056 1828
rect 87607 1779 87613 1782
rect 87549 1773 87613 1779
rect 94050 1779 94056 1782
rect 94108 1828 94114 1831
rect 94108 1782 97170 1828
rect 94108 1779 94114 1782
rect 94050 1773 94114 1779
rect 5730 1575 5794 1581
rect 5730 1523 5736 1575
rect 5788 1523 5794 1575
rect 5730 1517 5794 1523
rect 16770 1575 16834 1581
rect 16770 1523 16776 1575
rect 16828 1523 16834 1575
rect 16770 1517 16834 1523
rect 27810 1575 27874 1581
rect 27810 1523 27816 1575
rect 27868 1523 27874 1575
rect 27810 1517 27874 1523
rect 38850 1575 38914 1581
rect 38850 1523 38856 1575
rect 38908 1523 38914 1575
rect 38850 1517 38914 1523
rect 49890 1575 49954 1581
rect 49890 1523 49896 1575
rect 49948 1523 49954 1575
rect 49890 1517 49954 1523
rect 60930 1575 60994 1581
rect 60930 1523 60936 1575
rect 60988 1523 60994 1575
rect 60930 1517 60994 1523
rect 71970 1575 72034 1581
rect 71970 1523 71976 1575
rect 72028 1523 72034 1575
rect 71970 1517 72034 1523
rect 83010 1575 83074 1581
rect 83010 1523 83016 1575
rect 83068 1523 83074 1575
rect 83010 1517 83074 1523
rect 94050 1575 94114 1581
rect 94050 1523 94056 1575
rect 94108 1523 94114 1575
rect 94050 1517 94114 1523
rect 88 0 97198 46
<< via1 >>
rect 19715 35728 19767 35780
rect 22514 35728 22566 35780
rect 30755 35728 30807 35780
rect 33554 35728 33606 35780
rect 41795 35728 41847 35780
rect 44594 35728 44646 35780
rect 52835 35728 52887 35780
rect 55634 35728 55686 35780
rect 63875 35728 63927 35780
rect 66674 35728 66726 35780
rect 74915 35728 74967 35780
rect 77714 35728 77766 35780
rect 85955 35728 86007 35780
rect 88754 35728 88806 35780
rect 87555 34798 87607 34850
rect 96772 33242 96824 33294
rect 86771 33016 86823 33068
rect 86771 3561 86823 3613
rect 1662 3335 1714 3387
rect 12702 3335 12754 3387
rect 23742 3335 23794 3387
rect 34782 3335 34834 3387
rect 45822 3335 45874 3387
rect 56862 3335 56914 3387
rect 67902 3335 67954 3387
rect 78942 3335 78994 3387
rect 89982 3335 90034 3387
rect 96772 3335 96824 3387
rect 8452 2709 8504 2761
rect 11251 2709 11303 2761
rect 19492 2709 19544 2761
rect 22291 2709 22343 2761
rect 30532 2709 30584 2761
rect 33331 2709 33383 2761
rect 41572 2709 41624 2761
rect 44371 2709 44423 2761
rect 52612 2709 52664 2761
rect 55411 2709 55463 2761
rect 63652 2709 63704 2761
rect 66451 2709 66503 2761
rect 74692 2709 74744 2761
rect 77491 2709 77543 2761
rect 85732 2709 85784 2761
rect 88531 2709 88583 2761
rect 5736 1779 5788 1831
rect 16776 1779 16828 1831
rect 27816 1779 27868 1831
rect 38856 1779 38908 1831
rect 49896 1779 49948 1831
rect 60936 1779 60988 1831
rect 71976 1779 72028 1831
rect 83016 1779 83068 1831
rect 87555 1779 87607 1831
rect 94056 1779 94108 1831
rect 5736 1523 5788 1575
rect 16776 1523 16828 1575
rect 27816 1523 27868 1575
rect 38856 1523 38908 1575
rect 49896 1523 49948 1575
rect 60936 1523 60988 1575
rect 71976 1523 72028 1575
rect 83016 1523 83068 1575
rect 94056 1523 94108 1575
<< metal2 >>
rect 322 35782 396 35791
rect 322 35726 331 35782
rect 387 35777 396 35782
rect 19709 35780 19773 35786
rect 387 35731 11523 35777
rect 387 35726 396 35731
rect 322 35717 396 35726
rect 19709 35728 19715 35780
rect 19767 35777 19773 35780
rect 22508 35780 22572 35786
rect 22508 35777 22514 35780
rect 19767 35731 22514 35777
rect 19767 35728 19773 35731
rect 19709 35722 19773 35728
rect 22508 35728 22514 35731
rect 22566 35728 22572 35780
rect 22508 35722 22572 35728
rect 30749 35780 30813 35786
rect 30749 35728 30755 35780
rect 30807 35777 30813 35780
rect 33548 35780 33612 35786
rect 33548 35777 33554 35780
rect 30807 35731 33554 35777
rect 30807 35728 30813 35731
rect 30749 35722 30813 35728
rect 33548 35728 33554 35731
rect 33606 35728 33612 35780
rect 33548 35722 33612 35728
rect 41789 35780 41853 35786
rect 41789 35728 41795 35780
rect 41847 35777 41853 35780
rect 44588 35780 44652 35786
rect 44588 35777 44594 35780
rect 41847 35731 44594 35777
rect 41847 35728 41853 35731
rect 41789 35722 41853 35728
rect 44588 35728 44594 35731
rect 44646 35728 44652 35780
rect 44588 35722 44652 35728
rect 52829 35780 52893 35786
rect 52829 35728 52835 35780
rect 52887 35777 52893 35780
rect 55628 35780 55692 35786
rect 55628 35777 55634 35780
rect 52887 35731 55634 35777
rect 52887 35728 52893 35731
rect 52829 35722 52893 35728
rect 55628 35728 55634 35731
rect 55686 35728 55692 35780
rect 55628 35722 55692 35728
rect 63869 35780 63933 35786
rect 63869 35728 63875 35780
rect 63927 35777 63933 35780
rect 66668 35780 66732 35786
rect 66668 35777 66674 35780
rect 63927 35731 66674 35777
rect 63927 35728 63933 35731
rect 63869 35722 63933 35728
rect 66668 35728 66674 35731
rect 66726 35728 66732 35780
rect 66668 35722 66732 35728
rect 74909 35780 74973 35786
rect 74909 35728 74915 35780
rect 74967 35777 74973 35780
rect 77708 35780 77772 35786
rect 77708 35777 77714 35780
rect 74967 35731 77714 35777
rect 74967 35728 74973 35731
rect 74909 35722 74973 35728
rect 77708 35728 77714 35731
rect 77766 35728 77772 35780
rect 77708 35722 77772 35728
rect 85949 35780 86013 35786
rect 85949 35728 85955 35780
rect 86007 35777 86013 35780
rect 88748 35780 88812 35786
rect 88748 35777 88754 35780
rect 86007 35731 88754 35777
rect 86007 35728 86013 35731
rect 85949 35722 86013 35728
rect 88748 35728 88754 35731
rect 88806 35728 88812 35780
rect 88748 35722 88812 35728
rect 16765 35662 16839 35671
rect 16765 35606 16774 35662
rect 16830 35606 16839 35662
rect 16765 35597 16839 35606
rect 23731 35662 23805 35671
rect 23731 35606 23740 35662
rect 23796 35606 23805 35662
rect 23731 35597 23805 35606
rect 34771 35662 34845 35671
rect 34771 35606 34780 35662
rect 34836 35606 34845 35662
rect 34771 35597 34845 35606
rect 45811 35662 45885 35671
rect 45811 35606 45820 35662
rect 45876 35606 45885 35662
rect 45811 35597 45885 35606
rect 56851 35662 56925 35671
rect 56851 35606 56860 35662
rect 56916 35606 56925 35662
rect 56851 35597 56925 35606
rect 67891 35662 67965 35671
rect 67891 35606 67900 35662
rect 67956 35606 67965 35662
rect 67891 35597 67965 35606
rect 78931 35662 79005 35671
rect 78931 35606 78940 35662
rect 78996 35606 79005 35662
rect 78931 35597 79005 35606
rect 89971 35662 90045 35671
rect 89971 35606 89980 35662
rect 90036 35606 90045 35662
rect 89971 35597 90045 35606
rect 87544 34852 87618 34861
rect 87544 34796 87553 34852
rect 87609 34796 87618 34852
rect 87544 34787 87618 34796
rect 12691 34042 12765 34051
rect 12691 33986 12700 34042
rect 12756 33986 12765 34042
rect 12691 33977 12765 33986
rect 27805 34042 27879 34051
rect 27805 33986 27814 34042
rect 27870 33986 27879 34042
rect 27805 33977 27879 33986
rect 38845 34042 38919 34051
rect 38845 33986 38854 34042
rect 38910 33986 38919 34042
rect 38845 33977 38919 33986
rect 49885 34042 49959 34051
rect 49885 33986 49894 34042
rect 49950 33986 49959 34042
rect 49885 33977 49959 33986
rect 60925 34042 60999 34051
rect 60925 33986 60934 34042
rect 60990 33986 60999 34042
rect 60925 33977 60999 33986
rect 71965 34042 72039 34051
rect 71965 33986 71974 34042
rect 72030 33986 72039 34042
rect 71965 33977 72039 33986
rect 83005 34042 83079 34051
rect 83005 33986 83014 34042
rect 83070 33986 83079 34042
rect 83005 33977 83079 33986
rect 94045 34042 94119 34051
rect 94045 33986 94054 34042
rect 94110 33986 94119 34042
rect 94045 33977 94119 33986
rect 96761 33296 96835 33305
rect 96761 33240 96770 33296
rect 96826 33240 96835 33296
rect 96761 33231 96835 33240
rect 86760 33070 86834 33079
rect 86760 33014 86769 33070
rect 86825 33014 86834 33070
rect 86760 33005 86834 33014
rect 16765 32978 16839 32987
rect 16765 32922 16774 32978
rect 16830 32973 16839 32978
rect 27805 32978 27879 32987
rect 27805 32973 27814 32978
rect 16830 32927 27814 32973
rect 16830 32922 16839 32927
rect 16765 32913 16839 32922
rect 27805 32922 27814 32927
rect 27870 32973 27879 32978
rect 38845 32978 38919 32987
rect 38845 32973 38854 32978
rect 27870 32927 38854 32973
rect 27870 32922 27879 32927
rect 27805 32913 27879 32922
rect 38845 32922 38854 32927
rect 38910 32973 38919 32978
rect 49885 32978 49959 32987
rect 49885 32973 49894 32978
rect 38910 32927 49894 32973
rect 38910 32922 38919 32927
rect 38845 32913 38919 32922
rect 49885 32922 49894 32927
rect 49950 32973 49959 32978
rect 60925 32978 60999 32987
rect 60925 32973 60934 32978
rect 49950 32927 60934 32973
rect 49950 32922 49959 32927
rect 49885 32913 49959 32922
rect 60925 32922 60934 32927
rect 60990 32973 60999 32978
rect 71965 32978 72039 32987
rect 71965 32973 71974 32978
rect 60990 32927 71974 32973
rect 60990 32922 60999 32927
rect 60925 32913 60999 32922
rect 71965 32922 71974 32927
rect 72030 32973 72039 32978
rect 83005 32978 83079 32987
rect 83005 32973 83014 32978
rect 72030 32927 83014 32973
rect 72030 32922 72039 32927
rect 71965 32913 72039 32922
rect 83005 32922 83014 32927
rect 83070 32973 83079 32978
rect 94045 32978 94119 32987
rect 94045 32973 94054 32978
rect 83070 32927 94054 32973
rect 83070 32922 83079 32927
rect 83005 32913 83079 32922
rect 94045 32922 94054 32927
rect 94110 32922 94119 32978
rect 94045 32913 94119 32922
rect 12691 32886 12765 32895
rect 12691 32830 12700 32886
rect 12756 32881 12765 32886
rect 23731 32886 23805 32895
rect 23731 32881 23740 32886
rect 12756 32835 23740 32881
rect 12756 32830 12765 32835
rect 12691 32821 12765 32830
rect 23731 32830 23740 32835
rect 23796 32881 23805 32886
rect 34771 32886 34845 32895
rect 34771 32881 34780 32886
rect 23796 32835 34780 32881
rect 23796 32830 23805 32835
rect 23731 32821 23805 32830
rect 34771 32830 34780 32835
rect 34836 32881 34845 32886
rect 45811 32886 45885 32895
rect 45811 32881 45820 32886
rect 34836 32835 45820 32881
rect 34836 32830 34845 32835
rect 34771 32821 34845 32830
rect 45811 32830 45820 32835
rect 45876 32881 45885 32886
rect 56851 32886 56925 32895
rect 56851 32881 56860 32886
rect 45876 32835 56860 32881
rect 45876 32830 45885 32835
rect 45811 32821 45885 32830
rect 56851 32830 56860 32835
rect 56916 32881 56925 32886
rect 67891 32886 67965 32895
rect 67891 32881 67900 32886
rect 56916 32835 67900 32881
rect 56916 32830 56925 32835
rect 56851 32821 56925 32830
rect 67891 32830 67900 32835
rect 67956 32881 67965 32886
rect 78931 32886 79005 32895
rect 78931 32881 78940 32886
rect 67956 32835 78940 32881
rect 67956 32830 67965 32835
rect 67891 32821 67965 32830
rect 78931 32830 78940 32835
rect 78996 32881 79005 32886
rect 89971 32886 90045 32895
rect 89971 32881 89980 32886
rect 78996 32835 89980 32881
rect 78996 32830 79005 32835
rect 78931 32821 79005 32830
rect 89971 32830 89980 32835
rect 90036 32830 90045 32886
rect 89971 32821 90045 32830
rect 1651 3799 1725 3808
rect 1651 3743 1660 3799
rect 1716 3794 1725 3799
rect 12691 3799 12765 3808
rect 12691 3794 12700 3799
rect 1716 3748 12700 3794
rect 1716 3743 1725 3748
rect 1651 3734 1725 3743
rect 12691 3743 12700 3748
rect 12756 3794 12765 3799
rect 23731 3799 23805 3808
rect 23731 3794 23740 3799
rect 12756 3748 23740 3794
rect 12756 3743 12765 3748
rect 12691 3734 12765 3743
rect 23731 3743 23740 3748
rect 23796 3794 23805 3799
rect 34771 3799 34845 3808
rect 34771 3794 34780 3799
rect 23796 3748 34780 3794
rect 23796 3743 23805 3748
rect 23731 3734 23805 3743
rect 34771 3743 34780 3748
rect 34836 3794 34845 3799
rect 45811 3799 45885 3808
rect 45811 3794 45820 3799
rect 34836 3748 45820 3794
rect 34836 3743 34845 3748
rect 34771 3734 34845 3743
rect 45811 3743 45820 3748
rect 45876 3794 45885 3799
rect 56851 3799 56925 3808
rect 56851 3794 56860 3799
rect 45876 3748 56860 3794
rect 45876 3743 45885 3748
rect 45811 3734 45885 3743
rect 56851 3743 56860 3748
rect 56916 3794 56925 3799
rect 67891 3799 67965 3808
rect 67891 3794 67900 3799
rect 56916 3748 67900 3794
rect 56916 3743 56925 3748
rect 56851 3734 56925 3743
rect 67891 3743 67900 3748
rect 67956 3794 67965 3799
rect 78931 3799 79005 3808
rect 78931 3794 78940 3799
rect 67956 3748 78940 3794
rect 67956 3743 67965 3748
rect 67891 3734 67965 3743
rect 78931 3743 78940 3748
rect 78996 3794 79005 3799
rect 89971 3799 90045 3808
rect 89971 3794 89980 3799
rect 78996 3748 89980 3794
rect 78996 3743 79005 3748
rect 78931 3734 79005 3743
rect 89971 3743 89980 3748
rect 90036 3743 90045 3799
rect 89971 3734 90045 3743
rect 5725 3707 5799 3716
rect 5725 3651 5734 3707
rect 5790 3702 5799 3707
rect 16765 3707 16839 3716
rect 16765 3702 16774 3707
rect 5790 3656 16774 3702
rect 5790 3651 5799 3656
rect 5725 3642 5799 3651
rect 16765 3651 16774 3656
rect 16830 3702 16839 3707
rect 27805 3707 27879 3716
rect 27805 3702 27814 3707
rect 16830 3656 27814 3702
rect 16830 3651 16839 3656
rect 16765 3642 16839 3651
rect 27805 3651 27814 3656
rect 27870 3702 27879 3707
rect 38845 3707 38919 3716
rect 38845 3702 38854 3707
rect 27870 3656 38854 3702
rect 27870 3651 27879 3656
rect 27805 3642 27879 3651
rect 38845 3651 38854 3656
rect 38910 3702 38919 3707
rect 49885 3707 49959 3716
rect 49885 3702 49894 3707
rect 38910 3656 49894 3702
rect 38910 3651 38919 3656
rect 38845 3642 38919 3651
rect 49885 3651 49894 3656
rect 49950 3702 49959 3707
rect 60925 3707 60999 3716
rect 60925 3702 60934 3707
rect 49950 3656 60934 3702
rect 49950 3651 49959 3656
rect 49885 3642 49959 3651
rect 60925 3651 60934 3656
rect 60990 3702 60999 3707
rect 71965 3707 72039 3716
rect 71965 3702 71974 3707
rect 60990 3656 71974 3702
rect 60990 3651 60999 3656
rect 60925 3642 60999 3651
rect 71965 3651 71974 3656
rect 72030 3702 72039 3707
rect 83005 3707 83079 3716
rect 83005 3702 83014 3707
rect 72030 3656 83014 3702
rect 72030 3651 72039 3656
rect 71965 3642 72039 3651
rect 83005 3651 83014 3656
rect 83070 3702 83079 3707
rect 94045 3707 94119 3716
rect 94045 3702 94054 3707
rect 83070 3656 94054 3702
rect 83070 3651 83079 3656
rect 83005 3642 83079 3651
rect 94045 3651 94054 3656
rect 94110 3651 94119 3707
rect 94045 3642 94119 3651
rect 86760 3615 86834 3624
rect 86760 3559 86769 3615
rect 86825 3559 86834 3615
rect 86760 3550 86834 3559
rect 1651 3389 1725 3398
rect 1651 3333 1660 3389
rect 1716 3333 1725 3389
rect 1651 3324 1725 3333
rect 12691 3389 12765 3398
rect 12691 3333 12700 3389
rect 12756 3333 12765 3389
rect 12691 3324 12765 3333
rect 23731 3389 23805 3398
rect 23731 3333 23740 3389
rect 23796 3333 23805 3389
rect 23731 3324 23805 3333
rect 34771 3389 34845 3398
rect 34771 3333 34780 3389
rect 34836 3333 34845 3389
rect 34771 3324 34845 3333
rect 45811 3389 45885 3398
rect 45811 3333 45820 3389
rect 45876 3333 45885 3389
rect 45811 3324 45885 3333
rect 56851 3389 56925 3398
rect 56851 3333 56860 3389
rect 56916 3333 56925 3389
rect 56851 3324 56925 3333
rect 67891 3389 67965 3398
rect 67891 3333 67900 3389
rect 67956 3333 67965 3389
rect 67891 3324 67965 3333
rect 78931 3389 79005 3398
rect 78931 3333 78940 3389
rect 78996 3333 79005 3389
rect 78931 3324 79005 3333
rect 89971 3389 90045 3398
rect 89971 3333 89980 3389
rect 90036 3333 90045 3389
rect 89971 3324 90045 3333
rect 96761 3389 96835 3398
rect 96761 3333 96770 3389
rect 96826 3333 96835 3389
rect 96761 3324 96835 3333
rect 8446 2761 8510 2767
rect 8446 2709 8452 2761
rect 8504 2758 8510 2761
rect 11245 2761 11309 2767
rect 11245 2758 11251 2761
rect 8504 2712 11251 2758
rect 8504 2709 8510 2712
rect 8446 2703 8510 2709
rect 11245 2709 11251 2712
rect 11303 2709 11309 2761
rect 11245 2703 11309 2709
rect 19486 2761 19550 2767
rect 19486 2709 19492 2761
rect 19544 2758 19550 2761
rect 22285 2761 22349 2767
rect 22285 2758 22291 2761
rect 19544 2712 22291 2758
rect 19544 2709 19550 2712
rect 19486 2703 19550 2709
rect 22285 2709 22291 2712
rect 22343 2709 22349 2761
rect 22285 2703 22349 2709
rect 30526 2761 30590 2767
rect 30526 2709 30532 2761
rect 30584 2758 30590 2761
rect 33325 2761 33389 2767
rect 33325 2758 33331 2761
rect 30584 2712 33331 2758
rect 30584 2709 30590 2712
rect 30526 2703 30590 2709
rect 33325 2709 33331 2712
rect 33383 2709 33389 2761
rect 33325 2703 33389 2709
rect 41566 2761 41630 2767
rect 41566 2709 41572 2761
rect 41624 2758 41630 2761
rect 44365 2761 44429 2767
rect 44365 2758 44371 2761
rect 41624 2712 44371 2758
rect 41624 2709 41630 2712
rect 41566 2703 41630 2709
rect 44365 2709 44371 2712
rect 44423 2709 44429 2761
rect 44365 2703 44429 2709
rect 52606 2761 52670 2767
rect 52606 2709 52612 2761
rect 52664 2758 52670 2761
rect 55405 2761 55469 2767
rect 55405 2758 55411 2761
rect 52664 2712 55411 2758
rect 52664 2709 52670 2712
rect 52606 2703 52670 2709
rect 55405 2709 55411 2712
rect 55463 2709 55469 2761
rect 55405 2703 55469 2709
rect 63646 2761 63710 2767
rect 63646 2709 63652 2761
rect 63704 2758 63710 2761
rect 66445 2761 66509 2767
rect 66445 2758 66451 2761
rect 63704 2712 66451 2758
rect 63704 2709 63710 2712
rect 63646 2703 63710 2709
rect 66445 2709 66451 2712
rect 66503 2709 66509 2761
rect 66445 2703 66509 2709
rect 74686 2761 74750 2767
rect 74686 2709 74692 2761
rect 74744 2758 74750 2761
rect 77485 2761 77549 2767
rect 77485 2758 77491 2761
rect 74744 2712 77491 2758
rect 74744 2709 74750 2712
rect 74686 2703 74750 2709
rect 77485 2709 77491 2712
rect 77543 2709 77549 2761
rect 77485 2703 77549 2709
rect 85726 2761 85790 2767
rect 85726 2709 85732 2761
rect 85784 2758 85790 2761
rect 88525 2761 88589 2767
rect 88525 2758 88531 2761
rect 85784 2712 88531 2758
rect 85784 2709 85790 2712
rect 85726 2703 85790 2709
rect 88525 2709 88531 2712
rect 88583 2709 88589 2761
rect 88525 2703 88589 2709
rect 5725 1833 5799 1842
rect 5725 1777 5734 1833
rect 5790 1777 5799 1833
rect 5725 1768 5799 1777
rect 16765 1833 16839 1842
rect 16765 1777 16774 1833
rect 16830 1777 16839 1833
rect 16765 1768 16839 1777
rect 27805 1833 27879 1842
rect 27805 1777 27814 1833
rect 27870 1777 27879 1833
rect 27805 1768 27879 1777
rect 38845 1833 38919 1842
rect 38845 1777 38854 1833
rect 38910 1777 38919 1833
rect 38845 1768 38919 1777
rect 49885 1833 49959 1842
rect 49885 1777 49894 1833
rect 49950 1777 49959 1833
rect 49885 1768 49959 1777
rect 60925 1833 60999 1842
rect 60925 1777 60934 1833
rect 60990 1777 60999 1833
rect 60925 1768 60999 1777
rect 71965 1833 72039 1842
rect 71965 1777 71974 1833
rect 72030 1777 72039 1833
rect 71965 1768 72039 1777
rect 83005 1833 83079 1842
rect 83005 1777 83014 1833
rect 83070 1777 83079 1833
rect 83005 1768 83079 1777
rect 87544 1833 87618 1842
rect 87544 1777 87553 1833
rect 87609 1777 87618 1833
rect 87544 1768 87618 1777
rect 94045 1833 94119 1842
rect 94045 1777 94054 1833
rect 94110 1777 94119 1833
rect 94045 1768 94119 1777
rect 5725 1577 5799 1586
rect 5725 1521 5734 1577
rect 5790 1521 5799 1577
rect 5725 1512 5799 1521
rect 16765 1577 16839 1586
rect 16765 1521 16774 1577
rect 16830 1521 16839 1577
rect 16765 1512 16839 1521
rect 27805 1577 27879 1586
rect 27805 1521 27814 1577
rect 27870 1521 27879 1577
rect 27805 1512 27879 1521
rect 38845 1577 38919 1586
rect 38845 1521 38854 1577
rect 38910 1521 38919 1577
rect 38845 1512 38919 1521
rect 49885 1577 49959 1586
rect 49885 1521 49894 1577
rect 49950 1521 49959 1577
rect 49885 1512 49959 1521
rect 60925 1577 60999 1586
rect 60925 1521 60934 1577
rect 60990 1521 60999 1577
rect 60925 1512 60999 1521
rect 71965 1577 72039 1586
rect 71965 1521 71974 1577
rect 72030 1521 72039 1577
rect 71965 1512 72039 1521
rect 83005 1577 83079 1586
rect 83005 1521 83014 1577
rect 83070 1521 83079 1577
rect 83005 1512 83079 1521
rect 94045 1577 94119 1586
rect 94045 1521 94054 1577
rect 94110 1521 94119 1577
rect 94045 1512 94119 1521
<< via2 >>
rect 331 35726 387 35782
rect 16774 35606 16830 35662
rect 23740 35606 23796 35662
rect 34780 35606 34836 35662
rect 45820 35606 45876 35662
rect 56860 35606 56916 35662
rect 67900 35606 67956 35662
rect 78940 35606 78996 35662
rect 89980 35606 90036 35662
rect 87553 34850 87609 34852
rect 87553 34798 87555 34850
rect 87555 34798 87607 34850
rect 87607 34798 87609 34850
rect 87553 34796 87609 34798
rect 12700 33986 12756 34042
rect 27814 33986 27870 34042
rect 38854 33986 38910 34042
rect 49894 33986 49950 34042
rect 60934 33986 60990 34042
rect 71974 33986 72030 34042
rect 83014 33986 83070 34042
rect 94054 33986 94110 34042
rect 96770 33294 96826 33296
rect 96770 33242 96772 33294
rect 96772 33242 96824 33294
rect 96824 33242 96826 33294
rect 96770 33240 96826 33242
rect 86769 33068 86825 33070
rect 86769 33016 86771 33068
rect 86771 33016 86823 33068
rect 86823 33016 86825 33068
rect 86769 33014 86825 33016
rect 16774 32922 16830 32978
rect 27814 32922 27870 32978
rect 38854 32922 38910 32978
rect 49894 32922 49950 32978
rect 60934 32922 60990 32978
rect 71974 32922 72030 32978
rect 83014 32922 83070 32978
rect 94054 32922 94110 32978
rect 12700 32830 12756 32886
rect 23740 32830 23796 32886
rect 34780 32830 34836 32886
rect 45820 32830 45876 32886
rect 56860 32830 56916 32886
rect 67900 32830 67956 32886
rect 78940 32830 78996 32886
rect 89980 32830 90036 32886
rect 1660 3743 1716 3799
rect 12700 3743 12756 3799
rect 23740 3743 23796 3799
rect 34780 3743 34836 3799
rect 45820 3743 45876 3799
rect 56860 3743 56916 3799
rect 67900 3743 67956 3799
rect 78940 3743 78996 3799
rect 89980 3743 90036 3799
rect 5734 3651 5790 3707
rect 16774 3651 16830 3707
rect 27814 3651 27870 3707
rect 38854 3651 38910 3707
rect 49894 3651 49950 3707
rect 60934 3651 60990 3707
rect 71974 3651 72030 3707
rect 83014 3651 83070 3707
rect 94054 3651 94110 3707
rect 86769 3613 86825 3615
rect 86769 3561 86771 3613
rect 86771 3561 86823 3613
rect 86823 3561 86825 3613
rect 86769 3559 86825 3561
rect 1660 3387 1716 3389
rect 1660 3335 1662 3387
rect 1662 3335 1714 3387
rect 1714 3335 1716 3387
rect 1660 3333 1716 3335
rect 12700 3387 12756 3389
rect 12700 3335 12702 3387
rect 12702 3335 12754 3387
rect 12754 3335 12756 3387
rect 12700 3333 12756 3335
rect 23740 3387 23796 3389
rect 23740 3335 23742 3387
rect 23742 3335 23794 3387
rect 23794 3335 23796 3387
rect 23740 3333 23796 3335
rect 34780 3387 34836 3389
rect 34780 3335 34782 3387
rect 34782 3335 34834 3387
rect 34834 3335 34836 3387
rect 34780 3333 34836 3335
rect 45820 3387 45876 3389
rect 45820 3335 45822 3387
rect 45822 3335 45874 3387
rect 45874 3335 45876 3387
rect 45820 3333 45876 3335
rect 56860 3387 56916 3389
rect 56860 3335 56862 3387
rect 56862 3335 56914 3387
rect 56914 3335 56916 3387
rect 56860 3333 56916 3335
rect 67900 3387 67956 3389
rect 67900 3335 67902 3387
rect 67902 3335 67954 3387
rect 67954 3335 67956 3387
rect 67900 3333 67956 3335
rect 78940 3387 78996 3389
rect 78940 3335 78942 3387
rect 78942 3335 78994 3387
rect 78994 3335 78996 3387
rect 78940 3333 78996 3335
rect 89980 3387 90036 3389
rect 89980 3335 89982 3387
rect 89982 3335 90034 3387
rect 90034 3335 90036 3387
rect 89980 3333 90036 3335
rect 96770 3387 96826 3389
rect 96770 3335 96772 3387
rect 96772 3335 96824 3387
rect 96824 3335 96826 3387
rect 96770 3333 96826 3335
rect 5734 1831 5790 1833
rect 5734 1779 5736 1831
rect 5736 1779 5788 1831
rect 5788 1779 5790 1831
rect 5734 1777 5790 1779
rect 16774 1831 16830 1833
rect 16774 1779 16776 1831
rect 16776 1779 16828 1831
rect 16828 1779 16830 1831
rect 16774 1777 16830 1779
rect 27814 1831 27870 1833
rect 27814 1779 27816 1831
rect 27816 1779 27868 1831
rect 27868 1779 27870 1831
rect 27814 1777 27870 1779
rect 38854 1831 38910 1833
rect 38854 1779 38856 1831
rect 38856 1779 38908 1831
rect 38908 1779 38910 1831
rect 38854 1777 38910 1779
rect 49894 1831 49950 1833
rect 49894 1779 49896 1831
rect 49896 1779 49948 1831
rect 49948 1779 49950 1831
rect 49894 1777 49950 1779
rect 60934 1831 60990 1833
rect 60934 1779 60936 1831
rect 60936 1779 60988 1831
rect 60988 1779 60990 1831
rect 60934 1777 60990 1779
rect 71974 1831 72030 1833
rect 71974 1779 71976 1831
rect 71976 1779 72028 1831
rect 72028 1779 72030 1831
rect 71974 1777 72030 1779
rect 83014 1831 83070 1833
rect 83014 1779 83016 1831
rect 83016 1779 83068 1831
rect 83068 1779 83070 1831
rect 83014 1777 83070 1779
rect 87553 1831 87609 1833
rect 87553 1779 87555 1831
rect 87555 1779 87607 1831
rect 87607 1779 87609 1831
rect 87553 1777 87609 1779
rect 94054 1831 94110 1833
rect 94054 1779 94056 1831
rect 94056 1779 94108 1831
rect 94108 1779 94110 1831
rect 94054 1777 94110 1779
rect 5734 1575 5790 1577
rect 5734 1523 5736 1575
rect 5736 1523 5788 1575
rect 5788 1523 5790 1575
rect 5734 1521 5790 1523
rect 16774 1575 16830 1577
rect 16774 1523 16776 1575
rect 16776 1523 16828 1575
rect 16828 1523 16830 1575
rect 16774 1521 16830 1523
rect 27814 1575 27870 1577
rect 27814 1523 27816 1575
rect 27816 1523 27868 1575
rect 27868 1523 27870 1575
rect 27814 1521 27870 1523
rect 38854 1575 38910 1577
rect 38854 1523 38856 1575
rect 38856 1523 38908 1575
rect 38908 1523 38910 1575
rect 38854 1521 38910 1523
rect 49894 1575 49950 1577
rect 49894 1523 49896 1575
rect 49896 1523 49948 1575
rect 49948 1523 49950 1575
rect 49894 1521 49950 1523
rect 60934 1575 60990 1577
rect 60934 1523 60936 1575
rect 60936 1523 60988 1575
rect 60988 1523 60990 1575
rect 60934 1521 60990 1523
rect 71974 1575 72030 1577
rect 71974 1523 71976 1575
rect 71976 1523 72028 1575
rect 72028 1523 72030 1575
rect 71974 1521 72030 1523
rect 83014 1575 83070 1577
rect 83014 1523 83016 1575
rect 83016 1523 83068 1575
rect 83068 1523 83070 1575
rect 83014 1521 83070 1523
rect 94054 1575 94110 1577
rect 94054 1523 94056 1575
rect 94056 1523 94108 1575
rect 94108 1523 94110 1575
rect 94054 1521 94110 1523
<< metal3 >>
rect 326 35782 392 35787
rect 326 35726 331 35782
rect 387 35726 392 35782
rect 326 35721 392 35726
rect 329 1577 389 35721
rect 16769 35662 16835 35667
rect 16769 35606 16774 35662
rect 16830 35606 16835 35662
rect 16769 35601 16835 35606
rect 23735 35662 23801 35667
rect 23735 35606 23740 35662
rect 23796 35606 23801 35662
rect 23735 35601 23801 35606
rect 34775 35662 34841 35667
rect 34775 35606 34780 35662
rect 34836 35606 34841 35662
rect 34775 35601 34841 35606
rect 45815 35662 45881 35667
rect 45815 35606 45820 35662
rect 45876 35606 45881 35662
rect 45815 35601 45881 35606
rect 56855 35662 56921 35667
rect 56855 35606 56860 35662
rect 56916 35606 56921 35662
rect 56855 35601 56921 35606
rect 67895 35662 67961 35667
rect 67895 35606 67900 35662
rect 67956 35606 67961 35662
rect 67895 35601 67961 35606
rect 78935 35662 79001 35667
rect 78935 35606 78940 35662
rect 78996 35606 79001 35662
rect 78935 35601 79001 35606
rect 89975 35662 90041 35667
rect 89975 35606 89980 35662
rect 90036 35606 90041 35662
rect 89975 35601 90041 35606
rect 13434 34856 13510 34862
rect 13434 34792 13440 34856
rect 13504 34792 13510 34856
rect 13434 34786 13510 34792
rect 12695 34042 12761 34047
rect 12695 33986 12700 34042
rect 12756 33986 12761 34042
rect 12695 33981 12761 33986
rect 12698 32891 12758 33981
rect 16772 32983 16832 35601
rect 16769 32978 16835 32983
rect 16769 32922 16774 32978
rect 16830 32922 16835 32978
rect 16769 32917 16835 32922
rect 12695 32886 12761 32891
rect 12695 32830 12700 32886
rect 12756 32830 12761 32886
rect 12695 32825 12761 32830
rect 12698 3804 12758 32825
rect 1655 3799 1721 3804
rect 1655 3743 1660 3799
rect 1716 3743 1721 3799
rect 1655 3738 1721 3743
rect 12695 3799 12761 3804
rect 12695 3743 12700 3799
rect 12756 3743 12761 3799
rect 12695 3738 12761 3743
rect 1658 3394 1718 3738
rect 5729 3707 5795 3712
rect 5729 3651 5734 3707
rect 5790 3651 5795 3707
rect 5729 3646 5795 3651
rect 1655 3389 1721 3394
rect 1655 3333 1660 3389
rect 1716 3333 1721 3389
rect 1655 3328 1721 3333
rect 5732 1838 5792 3646
rect 12698 3394 12758 3738
rect 16772 3712 16832 32917
rect 23738 32891 23798 35601
rect 24474 34856 24550 34862
rect 24474 34792 24480 34856
rect 24544 34792 24550 34856
rect 24474 34786 24550 34792
rect 27809 34042 27875 34047
rect 27809 33986 27814 34042
rect 27870 33986 27875 34042
rect 27809 33981 27875 33986
rect 27812 32983 27872 33981
rect 27809 32978 27875 32983
rect 27809 32922 27814 32978
rect 27870 32922 27875 32978
rect 27809 32917 27875 32922
rect 23735 32886 23801 32891
rect 23735 32830 23740 32886
rect 23796 32830 23801 32886
rect 23735 32825 23801 32830
rect 23738 3804 23798 32825
rect 23735 3799 23801 3804
rect 23735 3743 23740 3799
rect 23796 3743 23801 3799
rect 23735 3738 23801 3743
rect 16769 3707 16835 3712
rect 16769 3651 16774 3707
rect 16830 3651 16835 3707
rect 16769 3646 16835 3651
rect 12695 3389 12761 3394
rect 12695 3333 12700 3389
rect 12756 3333 12761 3389
rect 12695 3328 12761 3333
rect 5729 1833 5795 1838
rect 5729 1777 5734 1833
rect 5790 1777 5795 1833
rect 5729 1772 5795 1777
rect 6468 1837 6544 1843
rect 16772 1838 16832 3646
rect 23738 3394 23798 3738
rect 27812 3712 27872 32917
rect 34778 32891 34838 35601
rect 35514 34856 35590 34862
rect 35514 34792 35520 34856
rect 35584 34792 35590 34856
rect 35514 34786 35590 34792
rect 38849 34042 38915 34047
rect 38849 33986 38854 34042
rect 38910 33986 38915 34042
rect 38849 33981 38915 33986
rect 38852 32983 38912 33981
rect 38849 32978 38915 32983
rect 38849 32922 38854 32978
rect 38910 32922 38915 32978
rect 38849 32917 38915 32922
rect 34775 32886 34841 32891
rect 34775 32830 34780 32886
rect 34836 32830 34841 32886
rect 34775 32825 34841 32830
rect 34778 3804 34838 32825
rect 34775 3799 34841 3804
rect 34775 3743 34780 3799
rect 34836 3743 34841 3799
rect 34775 3738 34841 3743
rect 27809 3707 27875 3712
rect 27809 3651 27814 3707
rect 27870 3651 27875 3707
rect 27809 3646 27875 3651
rect 23735 3389 23801 3394
rect 23735 3333 23740 3389
rect 23796 3333 23801 3389
rect 23735 3328 23801 3333
rect 6468 1773 6474 1837
rect 6538 1773 6544 1837
rect 5732 1582 5792 1772
rect 6468 1767 6544 1773
rect 16769 1833 16835 1838
rect 16769 1777 16774 1833
rect 16830 1777 16835 1833
rect 16769 1772 16835 1777
rect 17508 1837 17584 1843
rect 27812 1838 27872 3646
rect 34778 3394 34838 3738
rect 38852 3712 38912 32917
rect 45818 32891 45878 35601
rect 46554 34856 46630 34862
rect 46554 34792 46560 34856
rect 46624 34792 46630 34856
rect 46554 34786 46630 34792
rect 49889 34042 49955 34047
rect 49889 33986 49894 34042
rect 49950 33986 49955 34042
rect 49889 33981 49955 33986
rect 49892 32983 49952 33981
rect 49889 32978 49955 32983
rect 49889 32922 49894 32978
rect 49950 32922 49955 32978
rect 49889 32917 49955 32922
rect 45815 32886 45881 32891
rect 45815 32830 45820 32886
rect 45876 32830 45881 32886
rect 45815 32825 45881 32830
rect 45818 3804 45878 32825
rect 45815 3799 45881 3804
rect 45815 3743 45820 3799
rect 45876 3743 45881 3799
rect 45815 3738 45881 3743
rect 38849 3707 38915 3712
rect 38849 3651 38854 3707
rect 38910 3651 38915 3707
rect 38849 3646 38915 3651
rect 34775 3389 34841 3394
rect 34775 3333 34780 3389
rect 34836 3333 34841 3389
rect 34775 3328 34841 3333
rect 17508 1773 17514 1837
rect 17578 1773 17584 1837
rect 16772 1582 16832 1772
rect 17508 1767 17584 1773
rect 27809 1833 27875 1838
rect 27809 1777 27814 1833
rect 27870 1777 27875 1833
rect 27809 1772 27875 1777
rect 28548 1837 28624 1843
rect 38852 1838 38912 3646
rect 45818 3394 45878 3738
rect 49892 3712 49952 32917
rect 56858 32891 56918 35601
rect 57594 34856 57670 34862
rect 57594 34792 57600 34856
rect 57664 34792 57670 34856
rect 57594 34786 57670 34792
rect 60929 34042 60995 34047
rect 60929 33986 60934 34042
rect 60990 33986 60995 34042
rect 60929 33981 60995 33986
rect 60932 32983 60992 33981
rect 60929 32978 60995 32983
rect 60929 32922 60934 32978
rect 60990 32922 60995 32978
rect 60929 32917 60995 32922
rect 56855 32886 56921 32891
rect 56855 32830 56860 32886
rect 56916 32830 56921 32886
rect 56855 32825 56921 32830
rect 56858 3804 56918 32825
rect 56855 3799 56921 3804
rect 56855 3743 56860 3799
rect 56916 3743 56921 3799
rect 56855 3738 56921 3743
rect 49889 3707 49955 3712
rect 49889 3651 49894 3707
rect 49950 3651 49955 3707
rect 49889 3646 49955 3651
rect 45815 3389 45881 3394
rect 45815 3333 45820 3389
rect 45876 3333 45881 3389
rect 45815 3328 45881 3333
rect 28548 1773 28554 1837
rect 28618 1773 28624 1837
rect 27812 1582 27872 1772
rect 28548 1767 28624 1773
rect 38849 1833 38915 1838
rect 38849 1777 38854 1833
rect 38910 1777 38915 1833
rect 38849 1772 38915 1777
rect 39588 1837 39664 1843
rect 49892 1838 49952 3646
rect 56858 3394 56918 3738
rect 60932 3712 60992 32917
rect 67898 32891 67958 35601
rect 68634 34856 68710 34862
rect 68634 34792 68640 34856
rect 68704 34792 68710 34856
rect 68634 34786 68710 34792
rect 71969 34042 72035 34047
rect 71969 33986 71974 34042
rect 72030 33986 72035 34042
rect 71969 33981 72035 33986
rect 71972 32983 72032 33981
rect 71969 32978 72035 32983
rect 71969 32922 71974 32978
rect 72030 32922 72035 32978
rect 71969 32917 72035 32922
rect 67895 32886 67961 32891
rect 67895 32830 67900 32886
rect 67956 32830 67961 32886
rect 67895 32825 67961 32830
rect 67898 3804 67958 32825
rect 67895 3799 67961 3804
rect 67895 3743 67900 3799
rect 67956 3743 67961 3799
rect 67895 3738 67961 3743
rect 60929 3707 60995 3712
rect 60929 3651 60934 3707
rect 60990 3651 60995 3707
rect 60929 3646 60995 3651
rect 56855 3389 56921 3394
rect 56855 3333 56860 3389
rect 56916 3333 56921 3389
rect 56855 3328 56921 3333
rect 39588 1773 39594 1837
rect 39658 1773 39664 1837
rect 38852 1582 38912 1772
rect 39588 1767 39664 1773
rect 49889 1833 49955 1838
rect 49889 1777 49894 1833
rect 49950 1777 49955 1833
rect 49889 1772 49955 1777
rect 50628 1837 50704 1843
rect 60932 1838 60992 3646
rect 67898 3394 67958 3738
rect 71972 3712 72032 32917
rect 78938 32891 78998 35601
rect 79674 34856 79750 34862
rect 79674 34792 79680 34856
rect 79744 34792 79750 34856
rect 79674 34786 79750 34792
rect 87124 34856 87200 34862
rect 87124 34792 87130 34856
rect 87194 34792 87200 34856
rect 87124 34786 87200 34792
rect 87548 34852 87614 34857
rect 87548 34796 87553 34852
rect 87609 34796 87614 34852
rect 87548 34791 87614 34796
rect 83009 34042 83075 34047
rect 83009 33986 83014 34042
rect 83070 33986 83075 34042
rect 83009 33981 83075 33986
rect 83012 32983 83072 33981
rect 86764 33070 86830 33075
rect 86764 33014 86769 33070
rect 86825 33014 86830 33070
rect 86764 33009 86830 33014
rect 83009 32978 83075 32983
rect 83009 32922 83014 32978
rect 83070 32922 83075 32978
rect 83009 32917 83075 32922
rect 78935 32886 79001 32891
rect 78935 32830 78940 32886
rect 78996 32830 79001 32886
rect 78935 32825 79001 32830
rect 78938 3804 78998 32825
rect 78935 3799 79001 3804
rect 78935 3743 78940 3799
rect 78996 3743 79001 3799
rect 78935 3738 79001 3743
rect 71969 3707 72035 3712
rect 71969 3651 71974 3707
rect 72030 3651 72035 3707
rect 71969 3646 72035 3651
rect 67895 3389 67961 3394
rect 67895 3333 67900 3389
rect 67956 3333 67961 3389
rect 67895 3328 67961 3333
rect 50628 1773 50634 1837
rect 50698 1773 50704 1837
rect 49892 1582 49952 1772
rect 50628 1767 50704 1773
rect 60929 1833 60995 1838
rect 60929 1777 60934 1833
rect 60990 1777 60995 1833
rect 60929 1772 60995 1777
rect 61668 1837 61744 1843
rect 71972 1838 72032 3646
rect 78938 3394 78998 3738
rect 83012 3712 83072 32917
rect 83009 3707 83075 3712
rect 83009 3651 83014 3707
rect 83070 3651 83075 3707
rect 83009 3646 83075 3651
rect 78935 3389 79001 3394
rect 78935 3333 78940 3389
rect 78996 3333 79001 3389
rect 78935 3328 79001 3333
rect 61668 1773 61674 1837
rect 61738 1773 61744 1837
rect 60932 1582 60992 1772
rect 61668 1767 61744 1773
rect 71969 1833 72035 1838
rect 71969 1777 71974 1833
rect 72030 1777 72035 1833
rect 71969 1772 72035 1777
rect 72708 1837 72784 1843
rect 83012 1838 83072 3646
rect 86767 3620 86827 33009
rect 86764 3615 86830 3620
rect 86764 3559 86769 3615
rect 86825 3559 86830 3615
rect 86764 3554 86830 3559
rect 87132 1843 87192 34786
rect 72708 1773 72714 1837
rect 72778 1773 72784 1837
rect 71972 1582 72032 1772
rect 72708 1767 72784 1773
rect 83009 1833 83075 1838
rect 83009 1777 83014 1833
rect 83070 1777 83075 1833
rect 83009 1772 83075 1777
rect 83748 1837 83824 1843
rect 83748 1773 83754 1837
rect 83818 1773 83824 1837
rect 83012 1582 83072 1772
rect 83748 1767 83824 1773
rect 87124 1837 87200 1843
rect 87551 1838 87611 34791
rect 89978 32891 90038 35601
rect 90714 34856 90790 34862
rect 90714 34792 90720 34856
rect 90784 34792 90790 34856
rect 90714 34786 90790 34792
rect 94049 34042 94115 34047
rect 94049 33986 94054 34042
rect 94110 33986 94115 34042
rect 94049 33981 94115 33986
rect 94052 32983 94112 33981
rect 96765 33296 96831 33301
rect 96765 33240 96770 33296
rect 96826 33240 96831 33296
rect 96765 33235 96831 33240
rect 94049 32978 94115 32983
rect 94049 32922 94054 32978
rect 94110 32922 94115 32978
rect 94049 32917 94115 32922
rect 89975 32886 90041 32891
rect 89975 32830 89980 32886
rect 90036 32830 90041 32886
rect 89975 32825 90041 32830
rect 89978 3804 90038 32825
rect 89975 3799 90041 3804
rect 89975 3743 89980 3799
rect 90036 3743 90041 3799
rect 89975 3738 90041 3743
rect 89978 3394 90038 3738
rect 94052 3712 94112 32917
rect 94049 3707 94115 3712
rect 94049 3651 94054 3707
rect 94110 3651 94115 3707
rect 94049 3646 94115 3651
rect 89975 3389 90041 3394
rect 89975 3333 89980 3389
rect 90036 3333 90041 3389
rect 89975 3328 90041 3333
rect 94052 1838 94112 3646
rect 96768 3394 96828 33235
rect 96765 3389 96831 3394
rect 96765 3333 96770 3389
rect 96826 3333 96831 3389
rect 96765 3328 96831 3333
rect 87124 1773 87130 1837
rect 87194 1773 87200 1837
rect 87124 1767 87200 1773
rect 87548 1833 87614 1838
rect 87548 1777 87553 1833
rect 87609 1777 87614 1833
rect 87548 1772 87614 1777
rect 94049 1833 94115 1838
rect 94049 1777 94054 1833
rect 94110 1777 94115 1833
rect 94049 1772 94115 1777
rect 94788 1837 94864 1843
rect 94788 1773 94794 1837
rect 94858 1773 94864 1837
rect 94052 1582 94112 1772
rect 94788 1767 94864 1773
rect 5729 1577 5795 1582
rect 5729 1521 5734 1577
rect 5790 1521 5795 1577
rect 5729 1516 5795 1521
rect 16769 1577 16835 1582
rect 16769 1521 16774 1577
rect 16830 1521 16835 1577
rect 16769 1516 16835 1521
rect 27809 1577 27875 1582
rect 27809 1521 27814 1577
rect 27870 1521 27875 1577
rect 27809 1516 27875 1521
rect 38849 1577 38915 1582
rect 38849 1521 38854 1577
rect 38910 1521 38915 1577
rect 38849 1516 38915 1521
rect 49889 1577 49955 1582
rect 49889 1521 49894 1577
rect 49950 1521 49955 1577
rect 49889 1516 49955 1521
rect 60929 1577 60995 1582
rect 60929 1521 60934 1577
rect 60990 1521 60995 1577
rect 60929 1516 60995 1521
rect 71969 1577 72035 1582
rect 71969 1521 71974 1577
rect 72030 1521 72035 1577
rect 71969 1516 72035 1521
rect 83009 1577 83075 1582
rect 83009 1521 83014 1577
rect 83070 1521 83075 1577
rect 83009 1516 83075 1521
rect 94049 1577 94115 1582
rect 94049 1521 94054 1577
rect 94110 1521 94115 1577
rect 94049 1516 94115 1521
rect 97205 51 97265 3559
<< via3 >>
rect 13440 34792 13504 34856
rect 24480 34792 24544 34856
rect 35520 34792 35584 34856
rect 6474 1773 6538 1837
rect 46560 34792 46624 34856
rect 17514 1773 17578 1837
rect 57600 34792 57664 34856
rect 28554 1773 28618 1837
rect 68640 34792 68704 34856
rect 39594 1773 39658 1837
rect 79680 34792 79744 34856
rect 87130 34792 87194 34856
rect 50634 1773 50698 1837
rect 61674 1773 61738 1837
rect 72714 1773 72778 1837
rect 83754 1773 83818 1837
rect 90720 34792 90784 34856
rect 87130 1773 87194 1837
rect 94794 1773 94858 1837
<< metal4 >>
rect 13439 34856 13505 34857
rect 13439 34792 13440 34856
rect 13504 34854 13505 34856
rect 24479 34856 24545 34857
rect 24479 34854 24480 34856
rect 13504 34794 24480 34854
rect 13504 34792 13505 34794
rect 13439 34791 13505 34792
rect 24479 34792 24480 34794
rect 24544 34854 24545 34856
rect 35519 34856 35585 34857
rect 35519 34854 35520 34856
rect 24544 34794 35520 34854
rect 24544 34792 24545 34794
rect 24479 34791 24545 34792
rect 35519 34792 35520 34794
rect 35584 34854 35585 34856
rect 46559 34856 46625 34857
rect 46559 34854 46560 34856
rect 35584 34794 46560 34854
rect 35584 34792 35585 34794
rect 35519 34791 35585 34792
rect 46559 34792 46560 34794
rect 46624 34854 46625 34856
rect 57599 34856 57665 34857
rect 57599 34854 57600 34856
rect 46624 34794 57600 34854
rect 46624 34792 46625 34794
rect 46559 34791 46625 34792
rect 57599 34792 57600 34794
rect 57664 34854 57665 34856
rect 68639 34856 68705 34857
rect 68639 34854 68640 34856
rect 57664 34794 68640 34854
rect 57664 34792 57665 34794
rect 57599 34791 57665 34792
rect 68639 34792 68640 34794
rect 68704 34854 68705 34856
rect 79679 34856 79745 34857
rect 79679 34854 79680 34856
rect 68704 34794 79680 34854
rect 68704 34792 68705 34794
rect 68639 34791 68705 34792
rect 79679 34792 79680 34794
rect 79744 34854 79745 34856
rect 87129 34856 87195 34857
rect 87129 34854 87130 34856
rect 79744 34794 87130 34854
rect 79744 34792 79745 34794
rect 79679 34791 79745 34792
rect 87129 34792 87130 34794
rect 87194 34854 87195 34856
rect 90719 34856 90785 34857
rect 90719 34854 90720 34856
rect 87194 34794 90720 34854
rect 87194 34792 87195 34794
rect 87129 34791 87195 34792
rect 90719 34792 90720 34794
rect 90784 34792 90785 34856
rect 90719 34791 90785 34792
rect 6473 1837 6539 1838
rect 6473 1773 6474 1837
rect 6538 1835 6539 1837
rect 17513 1837 17579 1838
rect 17513 1835 17514 1837
rect 6538 1775 17514 1835
rect 6538 1773 6539 1775
rect 6473 1772 6539 1773
rect 17513 1773 17514 1775
rect 17578 1835 17579 1837
rect 28553 1837 28619 1838
rect 28553 1835 28554 1837
rect 17578 1775 28554 1835
rect 17578 1773 17579 1775
rect 17513 1772 17579 1773
rect 28553 1773 28554 1775
rect 28618 1835 28619 1837
rect 39593 1837 39659 1838
rect 39593 1835 39594 1837
rect 28618 1775 39594 1835
rect 28618 1773 28619 1775
rect 28553 1772 28619 1773
rect 39593 1773 39594 1775
rect 39658 1835 39659 1837
rect 50633 1837 50699 1838
rect 50633 1835 50634 1837
rect 39658 1775 50634 1835
rect 39658 1773 39659 1775
rect 39593 1772 39659 1773
rect 50633 1773 50634 1775
rect 50698 1835 50699 1837
rect 61673 1837 61739 1838
rect 61673 1835 61674 1837
rect 50698 1775 61674 1835
rect 50698 1773 50699 1775
rect 50633 1772 50699 1773
rect 61673 1773 61674 1775
rect 61738 1835 61739 1837
rect 72713 1837 72779 1838
rect 72713 1835 72714 1837
rect 61738 1775 72714 1835
rect 61738 1773 61739 1775
rect 61673 1772 61739 1773
rect 72713 1773 72714 1775
rect 72778 1835 72779 1837
rect 83753 1837 83819 1838
rect 83753 1835 83754 1837
rect 72778 1775 83754 1835
rect 72778 1773 72779 1775
rect 72713 1772 72779 1773
rect 83753 1773 83754 1775
rect 83818 1835 83819 1837
rect 87129 1837 87195 1838
rect 87129 1835 87130 1837
rect 83818 1775 87130 1835
rect 83818 1773 83819 1775
rect 83753 1772 83819 1773
rect 87129 1773 87130 1775
rect 87194 1835 87195 1837
rect 94793 1837 94859 1838
rect 94793 1835 94794 1837
rect 87194 1775 94794 1835
rect 87194 1773 87195 1775
rect 87129 1772 87195 1773
rect 94793 1773 94794 1775
rect 94858 1773 94859 1837
rect 94793 1772 94859 1773
use D_FlipFlop  D_FlipFlop_1
timestamp 1755760262
transform 1 0 22168 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1755760262
transform 1 0 33208 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1755760262
transform 1 0 44248 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1755760262
transform 1 0 55288 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1755760262
transform 1 0 66328 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1755760262
transform 1 0 88408 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1755760262
transform 1 0 77368 0 1 34801
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_8
timestamp 1755760262
transform -1 0 19890 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_9
timestamp 1755760262
transform -1 0 86130 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_10
timestamp 1755760262
transform -1 0 97170 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_11
timestamp 1755760262
transform -1 0 75090 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_12
timestamp 1755760262
transform -1 0 64050 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_13
timestamp 1755760262
transform -1 0 53010 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_14
timestamp 1755760262
transform -1 0 41970 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_15
timestamp 1755760262
transform -1 0 30930 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_16
timestamp 1755760262
transform -1 0 8850 0 1 1782
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_17
timestamp 1755760262
transform 1 0 11128 0 1 34801
box -102 -1796 8762 1842
<< labels >>
flabel metal2 19767 35731 22514 35777 0 FreeSans 160 0 0 0 Q0
port 0 nsew
flabel metal2 30807 35731 33554 35777 0 FreeSans 160 0 0 0 Q1
port 1 nsew
flabel metal2 41847 35731 44594 35777 0 FreeSans 160 0 0 0 Q2
port 2 nsew
flabel metal2 52887 35731 55634 35777 0 FreeSans 160 0 0 0 Q3
port 3 nsew
flabel metal2 63927 35731 66674 35777 0 FreeSans 160 0 0 0 Q4
port 4 nsew
flabel metal2 74967 35731 77714 35777 0 FreeSans 160 0 0 0 Q5
port 5 nsew
flabel metal2 86007 35731 88754 35777 0 FreeSans 160 0 0 0 Q6
port 6 nsew
flabel metal3 96768 3389 96828 33240 0 FreeSans 160 0 0 0 Q7
port 7 nsew
flabel metal2 85784 2712 88531 2758 0 FreeSans 160 0 0 0 Q8
port 8 nsew
flabel metal2 74744 2712 77491 2758 0 FreeSans 160 0 0 0 Q9
port 9 nsew
flabel metal2 63704 2712 66451 2758 0 FreeSans 160 0 0 0 Q10
port 10 nsew
flabel metal2 52664 2712 55411 2758 0 FreeSans 160 0 0 0 Q11
port 11 nsew
flabel metal2 41624 2712 44371 2758 0 FreeSans 160 0 0 0 Q12
port 12 nsew
flabel metal2 30590 2712 33331 2758 0 FreeSans 160 0 0 0 Q13
port 13 nsew
flabel metal2 19544 2712 22291 2758 0 FreeSans 160 0 0 0 Q14
port 14 nsew
flabel metal2 8504 2712 11251 2758 0 FreeSans 160 0 0 0 Q15
port 15 nsew
flabel metal2 78996 3748 89980 3794 0 FreeSans 160 0 0 0 EN
port 16 nsew
flabel metal2 83070 3656 94054 3702 0 FreeSans 160 0 0 0 VDD
port 17 nsew
flabel metal3 97205 51 97265 3559 0 FreeSans 160 90 0 0 GND
port 20 nsew
flabel metal4 83818 1775 87130 1835 0 FreeSans 160 0 0 0 CLK
port 21 nsew
<< end >>
