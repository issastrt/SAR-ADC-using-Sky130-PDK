magic
tech sky130A
magscale 1 2
timestamp 1754907470
<< metal1 >>
rect 518 -68791 564 -8157
rect 9410 -9940 9456 -8157
rect 2304 -11944 2368 -11938
rect 2304 -11996 2310 -11944
rect 2362 -11996 2368 -11944
rect 2304 -12002 2368 -11996
rect 2304 -15508 2368 -15502
rect 2304 -15560 2310 -15508
rect 2362 -15560 2368 -15508
rect 2304 -15566 2368 -15560
rect 2304 -19072 2368 -19066
rect 2304 -19124 2310 -19072
rect 2362 -19124 2368 -19072
rect 2304 -19130 2368 -19124
rect 2304 -22636 2368 -22630
rect 2304 -22688 2310 -22636
rect 2362 -22688 2368 -22636
rect 2304 -22694 2368 -22688
rect 2304 -26200 2368 -26194
rect 2304 -26252 2310 -26200
rect 2362 -26252 2368 -26200
rect 2304 -26258 2368 -26252
rect 2304 -29764 2368 -29758
rect 2304 -29816 2310 -29764
rect 2362 -29816 2368 -29764
rect 2304 -29822 2368 -29816
rect 2304 -33328 2368 -33322
rect 2304 -33380 2310 -33328
rect 2362 -33380 2368 -33328
rect 2304 -33386 2368 -33380
rect 2304 -36892 2368 -36886
rect 2304 -36944 2310 -36892
rect 2362 -36944 2368 -36892
rect 2304 -36950 2368 -36944
rect 2304 -40456 2368 -40450
rect 2304 -40508 2310 -40456
rect 2362 -40508 2368 -40456
rect 2304 -40514 2368 -40508
rect 2304 -44020 2368 -44014
rect 2304 -44072 2310 -44020
rect 2362 -44072 2368 -44020
rect 2304 -44078 2368 -44072
rect 2304 -47584 2368 -47578
rect 2304 -47636 2310 -47584
rect 2362 -47636 2368 -47584
rect 2304 -47642 2368 -47636
rect 2304 -51148 2368 -51142
rect 2304 -51200 2310 -51148
rect 2362 -51200 2368 -51148
rect 2304 -51206 2368 -51200
rect 2304 -54712 2368 -54706
rect 2304 -54764 2310 -54712
rect 2362 -54764 2368 -54712
rect 2304 -54770 2368 -54764
rect 2304 -58276 2368 -58270
rect 2304 -58328 2310 -58276
rect 2362 -58328 2368 -58276
rect 2304 -58334 2368 -58328
rect 2304 -61840 2368 -61834
rect 2304 -61892 2310 -61840
rect 2362 -61892 2368 -61840
rect 2304 -61898 2368 -61892
rect 2304 -65404 2368 -65398
rect 2304 -65456 2310 -65404
rect 2362 -65456 2368 -65404
rect 2304 -65462 2368 -65456
rect 1699 -67009 1745 -66707
rect 9410 -67009 9456 -11767
<< via1 >>
rect 2310 -11996 2362 -11944
rect 2310 -15560 2362 -15508
rect 2310 -19124 2362 -19072
rect 2310 -22688 2362 -22636
rect 2310 -26252 2362 -26200
rect 2310 -29816 2362 -29764
rect 2310 -33380 2362 -33328
rect 2310 -36944 2362 -36892
rect 2310 -40508 2362 -40456
rect 2310 -44072 2362 -44020
rect 2310 -47636 2362 -47584
rect 2310 -51200 2362 -51148
rect 2310 -54764 2362 -54712
rect 2310 -58328 2362 -58276
rect 2310 -61892 2362 -61840
rect 2310 -65456 2362 -65404
<< metal2 >>
rect 2299 -9004 2373 -8995
rect 2299 -9060 2308 -9004
rect 2364 -9060 2373 -9004
rect 2299 -9069 2373 -9060
rect 1721 -10190 1795 -10181
rect 1721 -10246 1730 -10190
rect 1786 -10246 1795 -10190
rect 1721 -10255 1795 -10246
rect 2304 -11944 2368 -11938
rect 2304 -11996 2310 -11944
rect 2362 -11947 2368 -11944
rect 9060 -11942 9134 -11933
rect 9060 -11947 9069 -11942
rect 2362 -11993 9069 -11947
rect 2362 -11996 2368 -11993
rect 2304 -12002 2368 -11996
rect 9060 -11998 9069 -11993
rect 9125 -11998 9134 -11942
rect 9060 -12007 9134 -11998
rect 2005 -12688 2079 -12679
rect 2005 -12744 2014 -12688
rect 2070 -12744 2079 -12688
rect 2005 -12753 2079 -12744
rect 1721 -13242 1795 -13233
rect 1721 -13298 1730 -13242
rect 1786 -13298 1795 -13242
rect 1721 -13307 1795 -13298
rect 2304 -15508 2368 -15502
rect 2304 -15560 2310 -15508
rect 2362 -15511 2368 -15508
rect 9060 -15506 9134 -15497
rect 9060 -15511 9069 -15506
rect 2362 -15557 9069 -15511
rect 2362 -15560 2368 -15557
rect 2304 -15566 2368 -15560
rect 9060 -15562 9069 -15557
rect 9125 -15562 9134 -15506
rect 9060 -15571 9134 -15562
rect 2304 -19072 2368 -19066
rect 2304 -19124 2310 -19072
rect 2362 -19075 2368 -19072
rect 9060 -19070 9134 -19061
rect 9060 -19075 9069 -19070
rect 2362 -19121 9069 -19075
rect 2362 -19124 2368 -19121
rect 2304 -19130 2368 -19124
rect 9060 -19126 9069 -19121
rect 9125 -19126 9134 -19070
rect 9060 -19135 9134 -19126
rect 2304 -22636 2368 -22630
rect 2304 -22688 2310 -22636
rect 2362 -22639 2368 -22636
rect 9060 -22634 9134 -22625
rect 9060 -22639 9069 -22634
rect 2362 -22685 9069 -22639
rect 2362 -22688 2368 -22685
rect 2304 -22694 2368 -22688
rect 9060 -22690 9069 -22685
rect 9125 -22690 9134 -22634
rect 9060 -22699 9134 -22690
rect 2304 -26200 2368 -26194
rect 2304 -26252 2310 -26200
rect 2362 -26203 2368 -26200
rect 9060 -26198 9134 -26189
rect 9060 -26203 9069 -26198
rect 2362 -26249 9069 -26203
rect 2362 -26252 2368 -26249
rect 2304 -26258 2368 -26252
rect 9060 -26254 9069 -26249
rect 9125 -26254 9134 -26198
rect 9060 -26263 9134 -26254
rect 2304 -29764 2368 -29758
rect 2304 -29816 2310 -29764
rect 2362 -29767 2368 -29764
rect 9060 -29762 9134 -29753
rect 9060 -29767 9069 -29762
rect 2362 -29813 9069 -29767
rect 2362 -29816 2368 -29813
rect 2304 -29822 2368 -29816
rect 9060 -29818 9069 -29813
rect 9125 -29818 9134 -29762
rect 9060 -29827 9134 -29818
rect 2304 -33328 2368 -33322
rect 2304 -33380 2310 -33328
rect 2362 -33331 2368 -33328
rect 9060 -33326 9134 -33317
rect 9060 -33331 9069 -33326
rect 2362 -33377 9069 -33331
rect 2362 -33380 2368 -33377
rect 2304 -33386 2368 -33380
rect 9060 -33382 9069 -33377
rect 9125 -33382 9134 -33326
rect 9060 -33391 9134 -33382
rect 2304 -36892 2368 -36886
rect 2304 -36944 2310 -36892
rect 2362 -36895 2368 -36892
rect 9060 -36890 9134 -36881
rect 9060 -36895 9069 -36890
rect 2362 -36941 9069 -36895
rect 2362 -36944 2368 -36941
rect 2304 -36950 2368 -36944
rect 9060 -36946 9069 -36941
rect 9125 -36946 9134 -36890
rect 9060 -36955 9134 -36946
rect 2304 -40456 2368 -40450
rect 2304 -40508 2310 -40456
rect 2362 -40459 2368 -40456
rect 9060 -40454 9134 -40445
rect 9060 -40459 9069 -40454
rect 2362 -40505 9069 -40459
rect 2362 -40508 2368 -40505
rect 2304 -40514 2368 -40508
rect 9060 -40510 9069 -40505
rect 9125 -40510 9134 -40454
rect 9060 -40519 9134 -40510
rect 2304 -44020 2368 -44014
rect 2304 -44072 2310 -44020
rect 2362 -44023 2368 -44020
rect 9060 -44018 9134 -44009
rect 9060 -44023 9069 -44018
rect 2362 -44069 9069 -44023
rect 2362 -44072 2368 -44069
rect 2304 -44078 2368 -44072
rect 9060 -44074 9069 -44069
rect 9125 -44074 9134 -44018
rect 9060 -44083 9134 -44074
rect 2304 -47584 2368 -47578
rect 2304 -47636 2310 -47584
rect 2362 -47587 2368 -47584
rect 9060 -47582 9134 -47573
rect 9060 -47587 9069 -47582
rect 2362 -47633 9069 -47587
rect 2362 -47636 2368 -47633
rect 2304 -47642 2368 -47636
rect 9060 -47638 9069 -47633
rect 9125 -47638 9134 -47582
rect 9060 -47647 9134 -47638
rect 2304 -51148 2368 -51142
rect 2304 -51200 2310 -51148
rect 2362 -51151 2368 -51148
rect 9060 -51146 9134 -51137
rect 9060 -51151 9069 -51146
rect 2362 -51197 9069 -51151
rect 2362 -51200 2368 -51197
rect 2304 -51206 2368 -51200
rect 9060 -51202 9069 -51197
rect 9125 -51202 9134 -51146
rect 9060 -51211 9134 -51202
rect 2304 -54712 2368 -54706
rect 2304 -54764 2310 -54712
rect 2362 -54715 2368 -54712
rect 9060 -54710 9134 -54701
rect 9060 -54715 9069 -54710
rect 2362 -54761 9069 -54715
rect 2362 -54764 2368 -54761
rect 2304 -54770 2368 -54764
rect 9060 -54766 9069 -54761
rect 9125 -54766 9134 -54710
rect 9060 -54775 9134 -54766
rect 2304 -58276 2368 -58270
rect 2304 -58328 2310 -58276
rect 2362 -58279 2368 -58276
rect 9060 -58274 9134 -58265
rect 9060 -58279 9069 -58274
rect 2362 -58325 9069 -58279
rect 2362 -58328 2368 -58325
rect 2304 -58334 2368 -58328
rect 9060 -58330 9069 -58325
rect 9125 -58330 9134 -58274
rect 9060 -58339 9134 -58330
rect 2304 -61840 2368 -61834
rect 2304 -61892 2310 -61840
rect 2362 -61843 2368 -61840
rect 9060 -61838 9134 -61829
rect 9060 -61843 9069 -61838
rect 2362 -61889 9069 -61843
rect 2362 -61892 2368 -61889
rect 2304 -61898 2368 -61892
rect 9060 -61894 9069 -61889
rect 9125 -61894 9134 -61838
rect 9060 -61903 9134 -61894
rect 2304 -65404 2368 -65398
rect 2304 -65456 2310 -65404
rect 2362 -65407 2368 -65404
rect 9060 -65402 9134 -65393
rect 9060 -65407 9069 -65402
rect 2362 -65453 9069 -65407
rect 2362 -65456 2368 -65453
rect 2304 -65462 2368 -65456
rect 9060 -65458 9069 -65453
rect 9125 -65458 9134 -65402
rect 9060 -65467 9134 -65458
rect 2299 -66958 2373 -66949
rect 2299 -67014 2308 -66958
rect 2364 -66963 2373 -66958
rect 9060 -66958 9134 -66949
rect 9060 -66963 9069 -66958
rect 2364 -67009 9069 -66963
rect 2364 -67014 2373 -67009
rect 2299 -67023 2373 -67014
rect 9060 -67014 9069 -67009
rect 9125 -67014 9134 -66958
rect 9060 -67023 9134 -67014
<< via2 >>
rect 2308 -9060 2364 -9004
rect 1730 -10246 1786 -10190
rect 9069 -11998 9125 -11942
rect 2014 -12744 2070 -12688
rect 1730 -13298 1786 -13242
rect 9069 -15562 9125 -15506
rect 9069 -19126 9125 -19070
rect 9069 -22690 9125 -22634
rect 9069 -26254 9125 -26198
rect 9069 -29818 9125 -29762
rect 9069 -33382 9125 -33326
rect 9069 -36946 9125 -36890
rect 9069 -40510 9125 -40454
rect 9069 -44074 9125 -44018
rect 9069 -47638 9125 -47582
rect 9069 -51202 9125 -51146
rect 9069 -54766 9125 -54710
rect 9069 -58330 9125 -58274
rect 9069 -61894 9125 -61838
rect 9069 -65458 9125 -65402
rect 2308 -67014 2364 -66958
rect 9069 -67014 9125 -66958
<< metal3 >>
rect 2303 -9004 2369 -8999
rect 2303 -9060 2308 -9004
rect 2364 -9060 2369 -9004
rect 2303 -9065 2369 -9060
rect 1725 -10190 1791 -10185
rect 1725 -10246 1730 -10190
rect 1786 -10246 1791 -10190
rect 1725 -10251 1791 -10246
rect 1728 -13237 1788 -10251
rect 2012 -12683 2072 -10742
rect 1725 -13242 1791 -13237
rect 1725 -13298 1730 -13242
rect 1786 -13298 1791 -13242
rect 1725 -13303 1791 -13298
rect 1863 -67272 1923 -12686
rect 2009 -12688 2075 -12683
rect 2009 -12744 2014 -12688
rect 2070 -12744 2075 -12688
rect 2009 -12749 2075 -12744
rect 2012 -67826 2072 -13240
rect 2306 -66953 2366 -9065
rect 2303 -66958 2369 -66953
rect 2303 -67014 2308 -66958
rect 2364 -67014 2369 -66958
rect 2303 -67019 2369 -67014
rect 2920 -67272 2980 -9676
rect 9067 -11937 9127 -9580
rect 9064 -11942 9130 -11937
rect 9064 -11998 9069 -11942
rect 9125 -11998 9130 -11942
rect 9064 -12003 9130 -11998
rect 9067 -15501 9127 -13144
rect 9064 -15506 9130 -15501
rect 9064 -15562 9069 -15506
rect 9125 -15562 9130 -15506
rect 9064 -15567 9130 -15562
rect 9067 -19065 9127 -16708
rect 9064 -19070 9130 -19065
rect 9064 -19126 9069 -19070
rect 9125 -19126 9130 -19070
rect 9064 -19131 9130 -19126
rect 9067 -22629 9127 -20272
rect 9064 -22634 9130 -22629
rect 9064 -22690 9069 -22634
rect 9125 -22690 9130 -22634
rect 9064 -22695 9130 -22690
rect 9067 -26193 9127 -23836
rect 9064 -26198 9130 -26193
rect 9064 -26254 9069 -26198
rect 9125 -26254 9130 -26198
rect 9064 -26259 9130 -26254
rect 9067 -29757 9127 -27400
rect 9064 -29762 9130 -29757
rect 9064 -29818 9069 -29762
rect 9125 -29818 9130 -29762
rect 9064 -29823 9130 -29818
rect 9067 -33321 9127 -30964
rect 9064 -33326 9130 -33321
rect 9064 -33382 9069 -33326
rect 9125 -33382 9130 -33326
rect 9064 -33387 9130 -33382
rect 9067 -36885 9127 -34528
rect 9064 -36890 9130 -36885
rect 9064 -36946 9069 -36890
rect 9125 -36946 9130 -36890
rect 9064 -36951 9130 -36946
rect 9067 -40449 9127 -38092
rect 9064 -40454 9130 -40449
rect 9064 -40510 9069 -40454
rect 9125 -40510 9130 -40454
rect 9064 -40515 9130 -40510
rect 9067 -44013 9127 -41656
rect 9064 -44018 9130 -44013
rect 9064 -44074 9069 -44018
rect 9125 -44074 9130 -44018
rect 9064 -44079 9130 -44074
rect 9067 -47577 9127 -45220
rect 9064 -47582 9130 -47577
rect 9064 -47638 9069 -47582
rect 9125 -47638 9130 -47582
rect 9064 -47643 9130 -47638
rect 9067 -51141 9127 -48784
rect 9064 -51146 9130 -51141
rect 9064 -51202 9069 -51146
rect 9125 -51202 9130 -51146
rect 9064 -51207 9130 -51202
rect 9067 -54705 9127 -52348
rect 9064 -54710 9130 -54705
rect 9064 -54766 9069 -54710
rect 9125 -54766 9130 -54710
rect 9064 -54771 9130 -54766
rect 9067 -58269 9127 -55912
rect 9064 -58274 9130 -58269
rect 9064 -58330 9069 -58274
rect 9125 -58330 9130 -58274
rect 9064 -58335 9130 -58330
rect 9067 -61833 9127 -59476
rect 9064 -61838 9130 -61833
rect 9064 -61894 9069 -61838
rect 9125 -61894 9130 -61838
rect 9064 -61899 9130 -61894
rect 9067 -65397 9127 -63040
rect 9064 -65402 9130 -65397
rect 9064 -65458 9069 -65402
rect 9125 -65458 9130 -65402
rect 9064 -65463 9130 -65458
rect 9064 -66958 9130 -66953
rect 9064 -67014 9069 -66958
rect 9125 -67014 9130 -66958
rect 9064 -67019 9130 -67014
use D_FlipFlop  D_FlipFlop_0
timestamp 1754907470
transform 1 0 606 0 1 -9985
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_1
timestamp 1754907470
transform 1 0 606 0 1 -13549
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_2
timestamp 1754907470
transform 1 0 606 0 1 -17113
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_3
timestamp 1754907470
transform 1 0 606 0 1 -20677
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_4
timestamp 1754907470
transform 1 0 606 0 1 -24241
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_5
timestamp 1754907470
transform 1 0 606 0 1 -27805
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_6
timestamp 1754907470
transform 1 0 606 0 1 -31369
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_7
timestamp 1754907470
transform 1 0 606 0 1 -34933
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_8
timestamp 1754907470
transform 1 0 606 0 1 -38497
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_9
timestamp 1754907470
transform 1 0 606 0 1 -42061
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_10
timestamp 1754907470
transform 1 0 606 0 1 -45625
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_11
timestamp 1754907470
transform 1 0 606 0 1 -49189
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_12
timestamp 1754907470
transform 1 0 606 0 1 -52753
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_13
timestamp 1754907470
transform 1 0 606 0 1 -56317
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_14
timestamp 1754907470
transform 1 0 606 0 1 -59881
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_15
timestamp 1754907470
transform 1 0 606 0 1 -63445
box -88 -1782 8850 1828
use D_FlipFlop  D_FlipFlop_16
timestamp 1754907470
transform 1 0 606 0 1 -67009
box -88 -1782 8850 1828
<< labels >>
flabel metal3 2012 -67826 2072 -13240 0 FreeSans 160 90 0 0 VDD
port 19 nsew
flabel metal3 2920 -67272 2980 -9676 0 FreeSans 160 90 0 0 CLK
port 0 nsew
flabel metal3 1863 -67272 1923 -12686 0 FreeSans 160 90 0 0 EN
port 1 nsew
flabel metal3 9067 -11942 9127 -9580 0 FreeSans 160 0 0 0 Q0
port 3 nsew
flabel metal3 9067 -15506 9127 -13144 0 FreeSans 160 0 0 0 Q1
port 4 nsew
flabel metal3 9067 -19070 9127 -16708 0 FreeSans 160 0 0 0 Q2
port 5 nsew
flabel metal3 9067 -22634 9127 -20272 0 FreeSans 160 0 0 0 Q3
port 6 nsew
flabel metal3 9067 -26198 9127 -23836 0 FreeSans 160 0 0 0 Q4
port 7 nsew
flabel metal3 9067 -29762 9127 -27400 0 FreeSans 160 0 0 0 Q5
port 8 nsew
flabel metal3 9067 -33326 9127 -30964 0 FreeSans 160 0 0 0 Q6
port 9 nsew
flabel metal3 9067 -36890 9127 -34528 0 FreeSans 160 0 0 0 Q7
port 10 nsew
flabel metal3 9067 -40454 9127 -38092 0 FreeSans 160 0 0 0 Q8
port 11 nsew
flabel metal3 9067 -44018 9127 -41656 0 FreeSans 160 0 0 0 Q9
port 12 nsew
flabel metal3 9067 -47582 9127 -45220 0 FreeSans 160 0 0 0 Q10
port 13 nsew
flabel metal3 9067 -51146 9127 -48784 0 FreeSans 160 0 0 0 Q11
port 14 nsew
flabel metal3 9067 -54710 9127 -52348 0 FreeSans 160 0 0 0 Q12
port 15 nsew
flabel metal3 9067 -58274 9127 -55912 0 FreeSans 160 0 0 0 Q13
port 16 nsew
flabel metal3 9067 -61838 9127 -59476 0 FreeSans 160 0 0 0 Q14
port 17 nsew
flabel metal3 9067 -65402 9127 -63040 0 FreeSans 160 0 0 0 Q15
port 18 nsew
flabel metal1 518 -68791 564 -8157 0 FreeSans 160 90 0 0 GND
port 2 nsew
<< end >>
