** sch_path: /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-10_01-59-54/parameters/DNL/run_0/sar_output_dnl.sch
**.subckt sar_output_dnl
VVDD VDD GND DC 1.8
VVGND VGND GND DC 0
VVbias Vbias GND DC -0.9
VVin Vin GND PWL(0u 1.2 8.5u 1.2 8.500001u 1.201764705875 17.0u 1.201764705875 17.000001u 1.20352941175 25.5u 1.20352941175
+ 25.500001u 1.205294117625 34.0u 1.205294117625 34.000001u 1.2070588235 42.5u 1.2070588235 42.500001u 1.208823529375 51.0u 1.208823529375
+ 51.000001u 1.21058823525 59.5u 1.21058823525 59.500001u 1.212352941125 68.0u 1.212352941125 68.000001u 1.214117647 76.5u 1.214117647
+ 76.500001u 1.215882352875 85.0u 1.215882352875 85.000001u 1.21764705875 93.5u 1.21764705875 93.500001u 1.219411764625 102.0u 1.219411764625
+ 102.000001u 1.2211764705 110.5u 1.2211764705 110.500001u 1.222941176375 119.0u 1.222941176375 119.000001u 1.22470588225 127.5u 1.22470588225
+ 127.500001u 1.226470588125 136.0u 1.226470588125 136.000001u 1.228235294 144.5u 1.228235294 144.500001u 1.23 153.0u 1.23 153.000001u
+ 1.231764705875 161.5u 1.231764705875 161.500001u 1.23352941175 170.0u 1.23352941175 170.000001u 1.235294117625 178.5u 1.235294117625)
R1 net1 GND 0.01 m=1
Rout GND Q7 100000000.0 m=1
Rout1 GND Q6 100000000.0 m=1
Rout2 GND Q5 100000000.0 m=1
Rout3 GND Q4 100000000.0 m=1
Rout4 GND Q3 100000000.0 m=1
Rout5 GND Q2 100000000.0 m=1
Rout6 GND Q1 100000000.0 m=1
Rout7 GND Q0 100000000.0 m=1
x1 VDD Vin Q0 Vbias EN Q1 CLK Q2 Q3 Q4 Q5 Q6 Q7 VGND SAR-ADC-using-Sky130-PDK
VEN EN net1 PULSE(1.8 0 0 100ps 100ps 0.25u 0)
VCLK CLK GND PULSE(1.8 0 0 100p 100p 0.25u 0.5u)
**** begin user architecture code

* CACE gensim simulation file sar_output_dnl_0
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the current through the DAC.  Include both current through vdd and VREFH

.include /home/ece/cace/SAR-ADC-using-Sky130-PDK/netlist/rcx/SAR-ADC-using-Sky130-PDK.spice
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

.option TEMP=27
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1




.control
set wr_singlescale

  tran 0.5u 178.5u uic
  wrdata /home/ece/cace/SAR-ADC-using-Sky130-PDK/runs/RUN_2025-09-10_01-59-54/parameters/DNL/run_0/sar_output_dnl_0.data V(Vin) V(Q7) V(Q6) V(Q5) V(Q4) V(Q3) V(Q2) V(Q1) V(Q0)

end

quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
