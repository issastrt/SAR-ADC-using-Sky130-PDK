magic
tech sky130A
magscale 1 2
timestamp 1757097579
use CDAC  CDAC_0
timestamp 1757096721
transform 1 0 39078 0 1 6805
box -39092 -6796 55448 26024
use Comparator  Comparator_0
timestamp 1756559655
transform 1 0 71592 0 1 -4769
box 24473 -2307 30902 29735
use D_FlipFlop  D_FlipFlop_0
timestamp 1757097579
transform 1 0 60852 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_1
timestamp 1757097579
transform 1 0 52090 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_2
timestamp 1757097579
transform 1 0 43328 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_3
timestamp 1757097579
transform 1 0 34566 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_4
timestamp 1757097579
transform 1 0 17042 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_5
timestamp 1757097579
transform 1 0 25804 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_6
timestamp 1757097579
transform 1 0 8280 0 1 -5691
box 0 -1782 8762 1828
use D_FlipFlop  D_FlipFlop_7
timestamp 1757097579
transform 1 0 -482 0 1 -5691
box 0 -1782 8762 1828
<< end >>
