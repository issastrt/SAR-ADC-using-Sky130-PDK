magic
tech sky130A
magscale 1 2
timestamp 1761301090
<< nwell >>
rect 1296 -684 1338 198
rect 1961 -503 1989 -3
rect 2072 -234 2460 -66
rect 3226 -684 3268 198
<< pwell >>
rect 3135 -834 3205 -764
rect 1438 -1072 1518 -992
rect 2432 -1280 2512 -1200
<< mvpsubdiff >>
rect 1344 -816 1404 -782
rect 3160 -816 3220 -782
rect 1344 -842 1378 -816
rect 1344 -1456 1378 -1430
rect 3186 -842 3220 -816
rect 3186 -1456 3220 -1430
rect 1344 -1490 1404 -1456
rect 3160 -1490 3220 -1456
<< mvpsubdiffcont >>
rect 1404 -816 3160 -782
rect 1344 -1430 1378 -842
rect 3186 -1430 3220 -842
rect 1404 -1490 3160 -1456
<< locali >>
rect 1512 238 1824 244
rect 1512 204 1518 238
rect 1818 204 1824 238
rect 1512 86 1824 204
rect 2126 238 2438 244
rect 2126 204 2132 238
rect 2432 204 2438 238
rect 2126 86 2438 204
rect 2740 238 3052 244
rect 2740 204 2746 238
rect 3046 204 3052 238
rect 2740 86 3052 204
rect 1344 -816 1404 -782
rect 3160 -816 3220 -782
rect 1344 -842 1378 -816
rect 1344 -1456 1378 -1430
rect 3186 -842 3220 -816
rect 3186 -1456 3220 -1430
rect 1344 -1490 1404 -1456
rect 3160 -1490 3220 -1456
rect 1440 -1544 1896 -1490
rect 1440 -1578 1446 -1544
rect 1890 -1578 1896 -1544
rect 1440 -1584 1896 -1578
rect 2054 -1544 2510 -1490
rect 2054 -1578 2060 -1544
rect 2504 -1578 2510 -1544
rect 2054 -1584 2510 -1578
rect 2668 -1544 3124 -1490
rect 2668 -1578 2674 -1544
rect 3118 -1578 3124 -1544
rect 2668 -1584 3124 -1578
<< viali >>
rect 1518 204 1818 238
rect 2132 204 2432 238
rect 2746 204 3046 238
rect 1446 -1578 1890 -1544
rect 2060 -1578 2504 -1544
rect 2674 -1578 3118 -1544
<< metal1 >>
rect 1296 238 3268 261
rect 1296 204 1518 238
rect 1818 204 2132 238
rect 2432 204 2746 238
rect 3046 204 3268 238
rect 1296 181 3268 204
rect 1596 -58 1740 22
rect 2210 -58 2354 22
rect 2654 -99 2734 181
rect 2824 -58 2968 22
rect 1510 -321 1590 -99
rect 1510 -373 1524 -321
rect 1576 -373 1590 -321
rect 1510 -387 1590 -373
rect 1746 -307 1826 -99
rect 2160 -107 2204 -99
rect 2124 -307 2204 -107
rect 1746 -387 2204 -307
rect 2360 -113 2440 -99
rect 2360 -165 2374 -113
rect 2426 -165 2440 -113
rect 2360 -387 2440 -165
rect 2654 -179 2818 -99
rect 2738 -387 2818 -179
rect 2974 -307 3054 -99
rect 2974 -387 3210 -307
rect 1596 -508 1740 -428
rect 1628 -773 1708 -508
rect 1628 -825 1642 -773
rect 1694 -825 1708 -773
rect 1628 -880 1708 -825
rect 1524 -960 1812 -880
rect 1935 -992 2015 -387
rect 2210 -508 2354 -428
rect 2824 -508 2968 -428
rect 2242 -549 2322 -508
rect 2856 -549 2936 -508
rect 2242 -629 2936 -549
rect 2242 -880 2322 -629
rect 2856 -880 2936 -629
rect 3130 -773 3210 -387
rect 3130 -825 3144 -773
rect 3196 -825 3210 -773
rect 2138 -960 2426 -880
rect 2752 -960 3040 -880
rect 3130 -992 3210 -825
rect 1438 -1006 1518 -992
rect 1438 -1058 1452 -1006
rect 1504 -1058 1518 -1006
rect 1438 -1280 1518 -1058
rect 1818 -1038 2132 -992
rect 1818 -1280 1898 -1038
rect 2052 -1280 2132 -1038
rect 2432 -1214 2512 -992
rect 2666 -1200 2746 -992
rect 2432 -1266 2446 -1214
rect 2498 -1266 2512 -1214
rect 2432 -1280 2512 -1266
rect 2582 -1280 2746 -1200
rect 3046 -1072 3210 -992
rect 3046 -1280 3126 -1072
rect 1524 -1392 1812 -1312
rect 2138 -1392 2426 -1312
rect 2582 -1521 2662 -1280
rect 2752 -1392 3040 -1312
rect 1296 -1544 3268 -1521
rect 1296 -1578 1446 -1544
rect 1890 -1578 2060 -1544
rect 2504 -1578 2674 -1544
rect 3118 -1578 3268 -1544
rect 1296 -1601 3268 -1578
<< via1 >>
rect 1524 -373 1576 -321
rect 2374 -165 2426 -113
rect 1642 -825 1694 -773
rect 3144 -825 3196 -773
rect 1452 -1058 1504 -1006
rect 2446 -1266 2498 -1214
<< metal2 >>
rect 2052 -111 2440 -99
rect 2052 -167 2064 -111
rect 2120 -113 2440 -111
rect 2120 -165 2374 -113
rect 2426 -165 2440 -113
rect 2120 -167 2440 -165
rect 2052 -179 2440 -167
rect 1510 -319 1898 -307
rect 1510 -321 1830 -319
rect 1510 -373 1524 -321
rect 1576 -373 1830 -321
rect 1510 -375 1830 -373
rect 1886 -375 1898 -319
rect 1510 -387 1898 -375
rect 1628 -773 3210 -759
rect 1628 -825 1642 -773
rect 1694 -825 3144 -773
rect 3196 -825 3210 -773
rect 1628 -839 3210 -825
rect 1438 -1004 2132 -992
rect 1438 -1006 2064 -1004
rect 1438 -1058 1452 -1006
rect 1504 -1058 2064 -1006
rect 1438 -1060 2064 -1058
rect 2120 -1060 2132 -1004
rect 1438 -1072 2132 -1060
rect 1818 -1212 2512 -1200
rect 1818 -1268 1830 -1212
rect 1886 -1214 2512 -1212
rect 1886 -1266 2446 -1214
rect 2498 -1266 2512 -1214
rect 1886 -1268 2512 -1266
rect 1818 -1280 2512 -1268
<< via2 >>
rect 2064 -167 2120 -111
rect 1830 -375 1886 -319
rect 2064 -1060 2120 -1004
rect 1830 -1268 1886 -1212
<< metal3 >>
rect 2059 -111 2125 -106
rect 2059 -167 2064 -111
rect 2120 -167 2125 -111
rect 2059 -172 2125 -167
rect 1825 -319 1891 -314
rect 1825 -375 1830 -319
rect 1886 -375 1891 -319
rect 1825 -380 1891 -375
rect 1828 -1207 1888 -380
rect 2062 -999 2122 -172
rect 2059 -1004 2125 -999
rect 2059 -1060 2064 -1004
rect 2120 -1060 2125 -1004
rect 2059 -1065 2125 -1060
rect 1825 -1212 1891 -1207
rect 1825 -1268 1830 -1212
rect 1886 -1268 1891 -1212
rect 1825 -1273 1891 -1268
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM1
timestamp 1757220954
transform 1 0 1668 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM2
timestamp 1757220954
transform 1 0 2282 0 1 -1136
box -372 -402 372 402
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM3
timestamp 1757220954
transform 1 0 2282 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM4
timestamp 1757220954
transform 1 0 1668 0 1 -1136
box -372 -402 372 402
use sky130_fd_pr__pfet_g5v0d10v5_CY7YBN  XM5
timestamp 1757220954
transform 1 0 2896 0 1 -243
box -330 -441 330 441
use sky130_fd_pr__nfet_g5v0d10v5_3Y2F6P  XM6
timestamp 1757220954
transform 1 0 2896 0 1 -1136
box -372 -402 372 402
<< labels >>
flabel metal1 1296 -1584 3268 -1538 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal1 1296 198 3268 244 0 FreeSans 160 0 0 0 VDD
port 3 nsew
flabel metal1 2259 -612 2919 -566 0 FreeSans 160 0 0 0 Vref
port 4 nsew
flabel metal1 1952 -1038 1998 -341 0 FreeSans 160 0 0 0 Z
port 5 nsew
flabel metal3 1828 -1212 1888 -375 0 FreeSans 160 0 0 0 B
port 1 nsew
flabel metal3 2062 -1004 2122 -167 0 FreeSans 160 0 0 0 A
port 0 nsew
<< end >>
