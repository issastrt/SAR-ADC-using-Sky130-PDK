magic
tech sky130A
magscale 1 2
timestamp 1756559655
<< dnwell >>
rect 24583 14110 26613 29565
rect 24583 -1560 30792 14110
rect 24560 -2160 30792 -1560
rect 24583 -2191 30792 -2160
rect 24583 -2197 26613 -2191
<< nwell >>
rect 24473 29359 26723 29675
rect 24473 -1985 24795 29359
rect 26407 14220 26723 29359
rect 28818 18606 29237 29200
rect 29235 16606 29951 18606
rect 26407 13904 30902 14220
rect 30586 -1985 30902 13904
rect 24473 -2307 30902 -1985
<< pwell >>
rect 24850 12337 26328 29265
rect 24850 617 28850 12337
rect 24850 -1964 29969 617
rect 27899 -1985 27965 -1964
rect 28952 -1985 29018 -1964
<< mvnsubdiff >>
rect 24540 29588 26656 29608
rect 24540 29554 24634 29588
rect 26576 29554 26656 29588
rect 24540 29534 26656 29554
rect 24540 29528 24620 29534
rect 24540 -2146 24560 29528
rect 24600 -2146 24620 29528
rect 26582 29528 26656 29534
rect 26582 14157 26602 29528
rect 26636 14157 26656 29528
rect 26582 14153 26656 14157
rect 26582 14133 30835 14153
rect 26582 14099 26672 14133
rect 30755 14099 30835 14133
rect 26582 14079 30835 14099
rect 24540 -2160 24620 -2146
rect 30761 14073 30835 14079
rect 30761 -2154 30781 14073
rect 30815 -2154 30835 14073
rect 30761 -2160 30835 -2154
rect 24540 -2180 30835 -2160
rect 24540 -2220 24620 -2180
rect 30755 -2220 30835 -2180
rect 24540 -2240 30835 -2220
<< mvnsubdiffcont >>
rect 24634 29554 26576 29588
rect 24560 -2146 24600 29528
rect 26602 14157 26636 29528
rect 26672 14099 30755 14133
rect 30781 -2154 30815 14073
rect 24620 -2220 30755 -2180
<< locali >>
rect 24634 29715 26576 29721
rect 24634 29681 24640 29715
rect 26570 29681 26576 29715
rect 24634 29588 26576 29681
rect 24560 29554 24634 29588
rect 26576 29554 26636 29588
rect 24560 29528 24600 29554
rect 26602 29528 26636 29554
rect 27657 29240 28743 29246
rect 27657 29206 27663 29240
rect 28737 29206 28743 29240
rect 27657 29088 28743 29206
rect 29313 29240 29873 29246
rect 29313 29206 29319 29240
rect 29867 29206 29873 29240
rect 29313 29088 29873 29206
rect 26602 14133 26636 14157
rect 26602 14099 26672 14133
rect 30755 14099 30815 14133
rect 30781 14073 30815 14099
rect 24982 -1970 26196 -1829
rect 24982 -2004 24988 -1970
rect 26190 -2004 26196 -1970
rect 24982 -2010 26196 -2004
rect 27426 -1970 28438 -1817
rect 27426 -2004 27432 -1970
rect 28432 -2004 28438 -1970
rect 27426 -2010 28438 -2004
rect 29457 -1970 29825 -1817
rect 29457 -2004 29463 -1970
rect 29819 -2004 29825 -1970
rect 29457 -2010 29825 -2004
rect 24560 -2180 24600 -2146
rect 30781 -2180 30815 -2154
rect 24560 -2220 24620 -2180
rect 30755 -2220 30815 -2180
<< viali >>
rect 24640 29681 26570 29715
rect 27663 29206 28737 29240
rect 29319 29206 29867 29240
rect 24988 -2004 26190 -1970
rect 27432 -2004 28432 -1970
rect 29463 -2004 29819 -1970
<< metal1 >>
rect 26721 29724 26785 29730
rect 26721 29721 26727 29724
rect 24473 29715 26727 29721
rect 24473 29681 24640 29715
rect 26570 29681 26727 29715
rect 24473 29675 26727 29681
rect 25016 28832 26162 29675
rect 26721 29672 26727 29675
rect 26779 29672 26785 29724
rect 26721 29666 26785 29672
rect 26721 29249 26785 29255
rect 26721 29197 26727 29249
rect 26779 29246 26785 29249
rect 26779 29240 29951 29246
rect 26779 29206 27663 29240
rect 28737 29206 29319 29240
rect 29867 29206 29951 29240
rect 26779 29200 29951 29206
rect 26779 29197 26785 29200
rect 26721 29191 26785 29197
rect 28177 28903 28223 29200
rect 29391 28903 29437 29200
rect 28089 28857 28311 28903
rect 29391 28857 29441 28903
rect 26057 28818 26103 28832
rect 28603 18952 28682 18958
rect 28603 18949 28624 18952
rect 27785 18871 27831 18923
rect 28569 18903 28624 18949
rect 28618 18900 28624 18903
rect 28676 18900 28682 18952
rect 28618 18894 28682 18900
rect 27718 18865 27831 18871
rect 27718 18813 27724 18865
rect 27776 18862 27831 18865
rect 27776 18816 28559 18862
rect 27776 18813 27782 18816
rect 27718 18807 27782 18813
rect 29690 16957 29754 16963
rect 29690 16905 29696 16957
rect 29748 16905 29754 16957
rect 29690 16899 29754 16905
rect 29561 16865 29625 16871
rect 29561 16813 29567 16865
rect 29619 16813 29625 16865
rect 29561 16807 29625 16813
rect 27905 12160 27969 12166
rect 27905 12108 27911 12160
rect 27963 12108 27969 12160
rect 27905 12102 27969 12108
rect 27718 12061 27782 12067
rect 27718 12009 27724 12061
rect 27776 12009 27782 12061
rect 27718 12003 27782 12009
rect 28618 12062 28682 12068
rect 28618 12010 28624 12062
rect 28676 12010 28682 12062
rect 28618 12004 28682 12010
rect 27975 9133 28039 9139
rect 27975 9081 27981 9133
rect 28033 9081 28039 9133
rect 27975 9075 28039 9081
rect 28361 9133 28425 9139
rect 28361 9081 28367 9133
rect 28419 9081 28425 9133
rect 28361 9075 28425 9081
rect 28503 9032 28567 9038
rect 28503 8980 28509 9032
rect 28561 8980 28567 9032
rect 28503 8974 28567 8980
rect 28093 2275 28157 2281
rect 28093 2223 28099 2275
rect 28151 2223 28157 2275
rect 28093 2217 28157 2223
rect 29738 292 29802 298
rect 29738 240 29744 292
rect 29796 240 29802 292
rect 29738 234 29802 240
rect 27460 -1581 27506 -1564
rect 25981 -1587 26045 -1581
rect 25981 -1639 25987 -1587
rect 26039 -1639 26045 -1587
rect 25981 -1645 26045 -1639
rect 27451 -1587 27515 -1581
rect 27451 -1639 27457 -1587
rect 27509 -1639 27515 -1587
rect 27451 -1645 27515 -1639
rect 27709 -1587 27773 -1581
rect 27709 -1639 27715 -1587
rect 27767 -1639 27773 -1587
rect 27709 -1645 27773 -1639
rect 28351 -1587 28415 -1581
rect 28351 -1639 28357 -1587
rect 28409 -1639 28415 -1587
rect 28351 -1645 28415 -1639
rect 29480 -1587 29544 -1581
rect 29480 -1639 29486 -1587
rect 29538 -1639 29544 -1587
rect 29480 -1645 29544 -1639
rect 27460 -1673 27506 -1645
rect 27460 -1719 29737 -1673
rect 27900 -1961 27964 -1955
rect 27900 -1964 27906 -1961
rect 24850 -1970 27906 -1964
rect 27958 -1964 27964 -1961
rect 28953 -1961 29017 -1955
rect 28953 -1964 28959 -1961
rect 27958 -1970 28959 -1964
rect 24850 -2004 24988 -1970
rect 26190 -2004 27432 -1970
rect 28432 -2004 28959 -1970
rect 24850 -2010 27906 -2004
rect 27900 -2013 27906 -2010
rect 27958 -2010 28959 -2004
rect 27958 -2013 27964 -2010
rect 27900 -2019 27964 -2013
rect 28953 -2013 28959 -2010
rect 29011 -1964 29017 -1961
rect 29011 -1970 29969 -1964
rect 29011 -2004 29463 -1970
rect 29819 -2004 29969 -1970
rect 29011 -2010 29969 -2004
rect 29011 -2013 29017 -2010
rect 28953 -2019 29017 -2013
<< via1 >>
rect 26727 29672 26779 29724
rect 26727 29197 26779 29249
rect 28624 18900 28676 18952
rect 27724 18813 27776 18865
rect 29696 16905 29748 16957
rect 29567 16813 29619 16865
rect 27911 12108 27963 12160
rect 27724 12009 27776 12061
rect 28624 12010 28676 12062
rect 27981 9081 28033 9133
rect 28367 9081 28419 9133
rect 28509 8980 28561 9032
rect 28099 2223 28151 2275
rect 29744 240 29796 292
rect 25987 -1639 26039 -1587
rect 27457 -1639 27509 -1587
rect 27715 -1639 27767 -1587
rect 28357 -1639 28409 -1587
rect 29486 -1639 29538 -1587
rect 27906 -1970 27958 -1961
rect 27906 -2004 27958 -1970
rect 27906 -2013 27958 -2004
rect 28959 -2013 29011 -1961
<< metal2 >>
rect 26716 29726 26790 29735
rect 26716 29670 26725 29726
rect 26781 29670 26790 29726
rect 26716 29661 26790 29670
rect 26716 29251 26790 29260
rect 26716 29195 26725 29251
rect 26781 29195 26790 29251
rect 26716 29186 26790 29195
rect 28613 18954 28687 18963
rect 28613 18898 28622 18954
rect 28678 18898 28687 18954
rect 28613 18889 28687 18898
rect 27713 18867 27787 18876
rect 27713 18811 27722 18867
rect 27778 18811 27787 18867
rect 27713 18802 27787 18811
rect 29690 16957 29754 16963
rect 29690 16905 29696 16957
rect 29748 16954 29754 16957
rect 30164 16959 30238 16968
rect 30164 16954 30173 16959
rect 29748 16908 30173 16954
rect 29748 16905 29754 16908
rect 29690 16899 29754 16905
rect 30164 16903 30173 16908
rect 30229 16903 30238 16959
rect 30164 16894 30238 16903
rect 28613 16867 28687 16876
rect 28613 16811 28622 16867
rect 28678 16862 28687 16867
rect 29556 16867 29630 16876
rect 29556 16862 29565 16867
rect 28678 16816 29565 16862
rect 28678 16811 28687 16816
rect 28613 16802 28687 16811
rect 29556 16811 29565 16816
rect 29621 16811 29630 16867
rect 29556 16802 29630 16811
rect 27900 12162 27974 12171
rect 27900 12106 27909 12162
rect 27965 12106 27974 12162
rect 27900 12097 27974 12106
rect 27713 12063 27787 12072
rect 27713 12007 27722 12063
rect 27778 12007 27787 12063
rect 27713 11998 27787 12007
rect 28613 12064 28687 12073
rect 28613 12008 28622 12064
rect 28678 12008 28687 12064
rect 28613 11999 28687 12008
rect 27975 9133 28039 9139
rect 27975 9081 27981 9133
rect 28033 9130 28039 9133
rect 28163 9135 28237 9144
rect 28163 9130 28172 9135
rect 28033 9084 28172 9130
rect 28033 9081 28039 9084
rect 27975 9075 28039 9081
rect 28163 9079 28172 9084
rect 28228 9130 28237 9135
rect 28361 9133 28425 9139
rect 28361 9130 28367 9133
rect 28228 9084 28367 9130
rect 28228 9079 28237 9084
rect 28163 9070 28237 9079
rect 28361 9081 28367 9084
rect 28419 9081 28425 9133
rect 28361 9075 28425 9081
rect 28498 9034 28572 9043
rect 28498 8978 28507 9034
rect 28563 8978 28572 9034
rect 28498 8969 28572 8978
rect 28088 2277 28162 2286
rect 28088 2221 28097 2277
rect 28153 2221 28162 2277
rect 28088 2212 28162 2221
rect 29738 292 29802 298
rect 29738 240 29744 292
rect 29796 289 29802 292
rect 30164 294 30238 303
rect 30164 289 30173 294
rect 29796 243 30173 289
rect 29796 240 29802 243
rect 29738 234 29802 240
rect 30164 238 30173 243
rect 30229 238 30238 294
rect 30164 229 30238 238
rect 25981 -1587 26045 -1581
rect 25981 -1639 25987 -1587
rect 26039 -1590 26045 -1587
rect 27451 -1587 27515 -1581
rect 27451 -1590 27457 -1587
rect 26039 -1636 27457 -1590
rect 26039 -1639 26045 -1636
rect 25981 -1645 26045 -1639
rect 27451 -1639 27457 -1636
rect 27509 -1639 27515 -1587
rect 27451 -1645 27515 -1639
rect 27709 -1587 27773 -1581
rect 27709 -1639 27715 -1587
rect 27767 -1590 27773 -1587
rect 27895 -1585 27969 -1576
rect 27895 -1590 27904 -1585
rect 27767 -1636 27904 -1590
rect 27767 -1639 27773 -1636
rect 27709 -1645 27773 -1639
rect 27895 -1641 27904 -1636
rect 27960 -1590 27969 -1585
rect 28351 -1587 28415 -1581
rect 28351 -1590 28357 -1587
rect 27960 -1636 28357 -1590
rect 27960 -1641 27969 -1636
rect 27895 -1650 27969 -1641
rect 28351 -1639 28357 -1636
rect 28409 -1590 28415 -1587
rect 28948 -1585 29022 -1576
rect 28948 -1590 28957 -1585
rect 28409 -1636 28957 -1590
rect 28409 -1639 28415 -1636
rect 28351 -1645 28415 -1639
rect 28948 -1641 28957 -1636
rect 29013 -1590 29022 -1585
rect 29480 -1587 29544 -1581
rect 29480 -1590 29486 -1587
rect 29013 -1636 29486 -1590
rect 29013 -1641 29022 -1636
rect 28948 -1650 29022 -1641
rect 29480 -1639 29486 -1636
rect 29538 -1639 29544 -1587
rect 29480 -1645 29544 -1639
rect 27895 -1959 27969 -1950
rect 27895 -2015 27904 -1959
rect 27960 -2015 27969 -1959
rect 27895 -2024 27969 -2015
rect 28948 -1959 29022 -1950
rect 28948 -2015 28957 -1959
rect 29013 -2015 29022 -1959
rect 28948 -2024 29022 -2015
<< via2 >>
rect 26725 29724 26781 29726
rect 26725 29672 26727 29724
rect 26727 29672 26779 29724
rect 26779 29672 26781 29724
rect 26725 29670 26781 29672
rect 26725 29249 26781 29251
rect 26725 29197 26727 29249
rect 26727 29197 26779 29249
rect 26779 29197 26781 29249
rect 26725 29195 26781 29197
rect 28622 18952 28678 18954
rect 28622 18900 28624 18952
rect 28624 18900 28676 18952
rect 28676 18900 28678 18952
rect 28622 18898 28678 18900
rect 27722 18865 27778 18867
rect 27722 18813 27724 18865
rect 27724 18813 27776 18865
rect 27776 18813 27778 18865
rect 27722 18811 27778 18813
rect 30173 16903 30229 16959
rect 28622 16811 28678 16867
rect 29565 16865 29621 16867
rect 29565 16813 29567 16865
rect 29567 16813 29619 16865
rect 29619 16813 29621 16865
rect 29565 16811 29621 16813
rect 27909 12160 27965 12162
rect 27909 12108 27911 12160
rect 27911 12108 27963 12160
rect 27963 12108 27965 12160
rect 27909 12106 27965 12108
rect 27722 12061 27778 12063
rect 27722 12009 27724 12061
rect 27724 12009 27776 12061
rect 27776 12009 27778 12061
rect 27722 12007 27778 12009
rect 28622 12062 28678 12064
rect 28622 12010 28624 12062
rect 28624 12010 28676 12062
rect 28676 12010 28678 12062
rect 28622 12008 28678 12010
rect 28172 9079 28228 9135
rect 28507 9032 28563 9034
rect 28507 8980 28509 9032
rect 28509 8980 28561 9032
rect 28561 8980 28563 9032
rect 28507 8978 28563 8980
rect 28097 2275 28153 2277
rect 28097 2223 28099 2275
rect 28099 2223 28151 2275
rect 28151 2223 28153 2275
rect 28097 2221 28153 2223
rect 30173 238 30229 294
rect 27904 -1641 27960 -1585
rect 28957 -1641 29013 -1585
rect 27904 -1961 27960 -1959
rect 27904 -2013 27906 -1961
rect 27906 -2013 27958 -1961
rect 27958 -2013 27960 -1961
rect 27904 -2015 27960 -2013
rect 28957 -1961 29013 -1959
rect 28957 -2013 28959 -1961
rect 28959 -2013 29011 -1961
rect 29011 -2013 29013 -1961
rect 28957 -2015 29013 -2013
<< metal3 >>
rect 26720 29726 26786 29731
rect 26720 29670 26725 29726
rect 26781 29670 26786 29726
rect 26720 29665 26786 29670
rect 26723 29256 26783 29665
rect 26720 29251 26786 29256
rect 26720 29195 26725 29251
rect 26781 29195 26786 29251
rect 26720 29190 26786 29195
rect 28617 18954 28683 18959
rect 28617 18898 28622 18954
rect 28678 18898 28683 18954
rect 28617 18893 28683 18898
rect 27717 18867 27783 18872
rect 27717 18811 27722 18867
rect 27778 18811 27783 18867
rect 27717 18806 27783 18811
rect 27720 12068 27780 18806
rect 28620 16872 28680 18893
rect 30168 16959 30234 16964
rect 30168 16903 30173 16959
rect 30229 16903 30234 16959
rect 30168 16898 30234 16903
rect 28617 16867 28683 16872
rect 28617 16811 28622 16867
rect 28678 16811 28683 16867
rect 28617 16806 28683 16811
rect 29560 16867 29626 16872
rect 29560 16811 29565 16867
rect 29621 16811 29626 16867
rect 29560 16806 29626 16811
rect 27899 12475 27975 12481
rect 27899 12411 27905 12475
rect 27969 12411 27975 12475
rect 27899 12405 27975 12411
rect 27907 12167 27967 12405
rect 27904 12162 27970 12167
rect 27904 12106 27909 12162
rect 27965 12106 27970 12162
rect 27904 12101 27970 12106
rect 28620 12069 28680 16806
rect 29563 13429 29623 16806
rect 29555 13423 29631 13429
rect 29555 13359 29561 13423
rect 29625 13359 29631 13423
rect 29555 13353 29631 13359
rect 27717 12063 27783 12068
rect 27717 12007 27722 12063
rect 27778 12007 27783 12063
rect 27717 12002 27783 12007
rect 28617 12064 28683 12069
rect 28617 12008 28622 12064
rect 28678 12008 28683 12064
rect 28617 12003 28683 12008
rect 30171 11311 30231 16898
rect 30163 11305 30239 11311
rect 30163 11241 30169 11305
rect 30233 11241 30239 11305
rect 30163 11235 30239 11241
rect 28167 9135 28233 9140
rect 28167 9079 28172 9135
rect 28228 9079 28233 9135
rect 28167 9074 28233 9079
rect 28170 2466 28230 9074
rect 28502 9034 28568 9039
rect 28502 8978 28507 9034
rect 28563 8978 28568 9034
rect 28502 8973 28568 8978
rect 28505 8735 28565 8973
rect 28497 8729 28573 8735
rect 28497 8665 28503 8729
rect 28567 8665 28573 8729
rect 28497 8659 28573 8665
rect 28947 5357 29023 5363
rect 28947 5293 28953 5357
rect 29017 5293 29023 5357
rect 28947 5287 29023 5293
rect 28096 2406 28230 2466
rect 28096 2282 28156 2406
rect 28092 2277 28158 2282
rect 28092 2221 28097 2277
rect 28153 2221 28158 2277
rect 28092 2216 28158 2221
rect 28955 -1580 29015 5287
rect 30171 299 30231 11235
rect 30168 294 30234 299
rect 30168 238 30173 294
rect 30229 238 30234 294
rect 30168 233 30234 238
rect 27899 -1585 27965 -1580
rect 27899 -1641 27904 -1585
rect 27960 -1641 27965 -1585
rect 27899 -1646 27965 -1641
rect 28952 -1585 29018 -1580
rect 28952 -1641 28957 -1585
rect 29013 -1641 29018 -1585
rect 28952 -1646 29018 -1641
rect 27902 -1954 27962 -1646
rect 28955 -1954 29015 -1646
rect 27899 -1959 27965 -1954
rect 27899 -2015 27904 -1959
rect 27960 -2015 27965 -1959
rect 27899 -2020 27965 -2015
rect 28952 -1959 29018 -1954
rect 28952 -2015 28957 -1959
rect 29013 -2015 29018 -1959
rect 28952 -2020 29018 -2015
<< via3 >>
rect 27905 12411 27969 12475
rect 29561 13359 29625 13423
rect 30169 11241 30233 11305
rect 28503 8665 28567 8729
rect 28953 5293 29017 5357
<< via4 >>
rect 29475 13423 29711 13509
rect 29475 13359 29561 13423
rect 29561 13359 29625 13423
rect 29625 13359 29711 13423
rect 29475 13273 29711 13359
rect 27819 12475 28055 12561
rect 27819 12411 27905 12475
rect 27905 12411 27969 12475
rect 27969 12411 28055 12475
rect 27819 12325 28055 12411
rect 30083 11305 30319 11391
rect 30083 11241 30169 11305
rect 30169 11241 30233 11305
rect 30233 11241 30319 11305
rect 30083 11155 30319 11241
rect 28417 8729 28653 8815
rect 28417 8665 28503 8729
rect 28503 8665 28567 8729
rect 28567 8665 28653 8729
rect 28417 8579 28653 8665
rect 28867 5357 29103 5443
rect 28867 5293 28953 5357
rect 28953 5293 29017 5357
rect 29017 5293 29103 5357
rect 28867 5207 29103 5293
<< metal5 >>
rect 29433 13509 29753 13533
rect 29433 13273 29475 13509
rect 29711 13273 29753 13509
rect 27777 12561 28097 12881
rect 27777 12325 27819 12561
rect 28055 12325 28097 12561
rect 27777 12301 28097 12325
rect 29433 12128 29753 13273
rect 29103 11391 30343 11433
rect 29103 11155 30083 11391
rect 30319 11155 30343 11391
rect 29103 11113 30343 11155
rect 28375 8815 28695 8839
rect 28375 8579 28417 8815
rect 28653 8579 28695 8815
rect 28375 8259 28695 8579
rect 29433 6180 29753 11113
rect 28835 5443 30165 5485
rect 28835 5207 28867 5443
rect 29103 5207 30165 5443
rect 28835 5165 30165 5207
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_0
timestamp 1756481424
transform 0 1 29593 -1 0 6071
box -884 -281 906 281
use sky130_fd_pr__cap_mim_m3_2_AZGBXE  sky130_fd_pr__cap_mim_m3_2_AZGBXE_1
timestamp 1756481424
transform 0 1 29593 -1 0 12019
box -884 -281 906 281
use sky130_fd_pr__nfet_g5v0d10v5_94KJBV  sky130_fd_pr__nfet_g5v0d10v5_94KJBV_0
timestamp 1756538730
transform 1 0 27878 0 1 10565
box -328 -1758 328 1758
use sky130_fd_pr__nfet_g5v0d10v5_94KJBV  sky130_fd_pr__nfet_g5v0d10v5_94KJBV_1
timestamp 1756538730
transform 1 0 28522 0 1 10565
box -328 -1758 328 1758
use sky130_fd_pr__nfet_g5v0d10v5_DTGLBV  sky130_fd_pr__nfet_g5v0d10v5_DTGLBV_1
timestamp 1756538730
transform 1 0 28254 0 1 359
box -328 -2258 328 2258
use sky130_fd_pr__nfet_g5v0d10v5_DTGLBV  sky130_fd_pr__nfet_g5v0d10v5_DTGLBV_2
timestamp 1756538730
transform 1 0 27610 0 1 359
box -328 -2258 328 2258
use sky130_fd_pr__res_xhigh_po_5p73_2WP2GG  sky130_fd_pr__res_xhigh_po_5p73_2WP2GG_0
timestamp 1756481424
transform 1 0 25589 0 1 13683
box -739 -15582 739 15582
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM3
timestamp 1756481424
transform 1 0 27937 0 1 23903
box -358 -5297 358 5297
use sky130_fd_pr__pfet_g5v0d10v5_U7VG7Q  XM4
timestamp 1756481424
transform 1 0 28463 0 1 23903
box -358 -5297 358 5297
use sky130_fd_pr__nfet_g5v0d10v5_Q3M7H8  XM6
timestamp 1756481424
transform 1 0 29641 0 1 -641
box -328 -1258 328 1258
use sky130_fd_pr__pfet_g5v0d10v5_UX3D7Q  XM9
timestamp 1756481424
transform 1 0 29593 0 1 22903
box -358 -6297 358 6297
<< labels >>
flabel metal5 27777 12561 28097 12881 0 FreeSans 800 0 0 0 Vinm
port 3 nsew
flabel metal5 29433 6180 29753 10857 0 FreeSans 800 0 0 0 Vout
port 5 nsew
flabel metal1 26723 29200 27663 29246 0 FreeSans 160 0 0 0 VDD
port 2 nsew
flabel metal1 25175 -2010 27906 -1964 0 FreeSans 160 0 0 0 VSS
port 6 nsew
flabel metal5 28375 8259 28695 8579 0 FreeSans 800 0 0 0 Vinp
port 4 nsew
<< end >>
