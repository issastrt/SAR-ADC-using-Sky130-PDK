magic
tech sky130A
magscale 1 2
timestamp 1756274891
<< nwell >>
rect 48421 48259 49779 49141
rect 70501 48259 71859 49141
rect 92581 48259 93939 49141
<< pwell >>
rect 77420 21858 77480 21904
<< metal1 >>
rect 60043 48518 60107 48524
rect 48770 48266 48816 48515
rect 60043 48466 60049 48518
rect 60101 48466 60107 48518
rect 82123 48518 82187 48524
rect 60043 48460 60107 48466
rect 49598 48432 49662 48438
rect 49598 48380 49604 48432
rect 49656 48380 49662 48432
rect 49598 48374 49662 48380
rect 59429 48432 59493 48438
rect 59429 48380 59435 48432
rect 59487 48380 59493 48432
rect 59429 48374 59493 48380
rect 70850 48266 70896 48515
rect 82123 48466 82129 48518
rect 82181 48466 82187 48518
rect 104203 48518 104267 48524
rect 82123 48460 82187 48466
rect 71678 48432 71742 48438
rect 71678 48380 71684 48432
rect 71736 48380 71742 48432
rect 71678 48374 71742 48380
rect 81509 48432 81573 48438
rect 81509 48380 81515 48432
rect 81567 48380 81573 48432
rect 81509 48374 81573 48380
rect 92930 48266 92976 48515
rect 104203 48466 104209 48518
rect 104261 48466 104267 48518
rect 104203 48460 104267 48466
rect 126283 48518 126347 48524
rect 126283 48466 126289 48518
rect 126341 48466 126347 48518
rect 126283 48460 126347 48466
rect 93758 48432 93822 48438
rect 93758 48380 93764 48432
rect 93816 48380 93822 48432
rect 93758 48374 93822 48380
rect 103589 48432 103653 48438
rect 103589 48380 103595 48432
rect 103647 48380 103653 48432
rect 103589 48374 103653 48380
rect 115838 48432 115902 48438
rect 115838 48380 115844 48432
rect 115896 48380 115902 48432
rect 115838 48374 115902 48380
rect 125669 48432 125733 48438
rect 125669 48380 125675 48432
rect 125727 48380 125733 48432
rect 125669 48374 125733 48380
rect 127250 48401 127314 48407
rect 127250 48349 127256 48401
rect 127308 48349 127314 48401
rect 127250 48343 127314 48349
rect 48761 48260 48825 48266
rect 48761 48208 48767 48260
rect 48819 48208 48825 48260
rect 48761 48202 48825 48208
rect 49375 48260 49439 48266
rect 49375 48208 49381 48260
rect 49433 48208 49439 48260
rect 49375 48202 49439 48208
rect 70841 48260 70905 48266
rect 70841 48208 70847 48260
rect 70899 48208 70905 48260
rect 70841 48202 70905 48208
rect 71455 48260 71519 48266
rect 71455 48208 71461 48260
rect 71513 48208 71519 48260
rect 71455 48202 71519 48208
rect 92921 48260 92985 48266
rect 92921 48208 92927 48260
rect 92979 48208 92985 48260
rect 92921 48202 92985 48208
rect 93535 48260 93599 48266
rect 93535 48208 93541 48260
rect 93593 48208 93599 48260
rect 93535 48202 93599 48208
rect 115001 48260 115065 48266
rect 115001 48208 115007 48260
rect 115059 48208 115065 48260
rect 115001 48202 115065 48208
rect 115615 48260 115679 48266
rect 115615 48208 115621 48260
rect 115673 48208 115679 48260
rect 115615 48202 115679 48208
rect 48770 47983 48816 48202
rect 70850 47983 70896 48202
rect 92930 47983 92976 48202
rect 61010 47961 61074 47967
rect 61010 47909 61016 47961
rect 61068 47909 61074 47961
rect 61010 47903 61074 47909
rect 77463 45581 77527 45587
rect 77463 45529 77469 45581
rect 77521 45529 77527 45581
rect 77463 45523 77527 45529
rect 77459 42450 77523 42456
rect 77459 42398 77465 42450
rect 77517 42398 77523 42450
rect 77459 42392 77523 42398
rect 77459 38878 77523 38884
rect 77459 38826 77465 38878
rect 77517 38826 77523 38878
rect 77459 38820 77523 38826
rect 77459 35322 77523 35328
rect 77459 35270 77465 35322
rect 77517 35270 77523 35322
rect 77459 35264 77523 35270
rect 77411 29035 77475 29041
rect 77411 28983 77417 29035
rect 77469 28983 77475 29035
rect 77411 28977 77475 28983
rect 77411 25471 77475 25477
rect 77411 25419 77417 25471
rect 77469 25419 77475 25471
rect 77411 25413 77475 25419
rect 77411 21902 77475 21908
rect 77411 21850 77417 21902
rect 77469 21850 77475 21902
rect 77411 21844 77475 21850
rect 77411 18957 77475 18963
rect 77411 18905 77417 18957
rect 77469 18905 77475 18957
rect 77411 18899 77475 18905
rect 49970 17917 50034 17923
rect 49970 17865 49976 17917
rect 50028 17865 50034 17917
rect 49970 17859 50034 17865
rect 72050 17917 72114 17923
rect 72050 17865 72056 17917
rect 72108 17865 72114 17917
rect 72050 17859 72114 17865
rect 94129 17917 94193 17923
rect 94129 17865 94135 17917
rect 94187 17865 94193 17917
rect 94129 17859 94193 17865
rect 116210 17917 116274 17923
rect 116210 17865 116216 17917
rect 116268 17865 116274 17917
rect 116210 17859 116274 17865
rect 38558 17744 38622 17750
rect 38558 17692 38564 17744
rect 38616 17692 38622 17744
rect 38558 17686 38622 17692
rect 49003 17744 49067 17750
rect 49003 17692 49009 17744
rect 49061 17692 49067 17744
rect 49003 17686 49067 17692
rect 60638 17744 60702 17750
rect 60638 17692 60644 17744
rect 60696 17692 60702 17744
rect 60638 17686 60702 17692
rect 71083 17744 71147 17750
rect 71083 17692 71089 17744
rect 71141 17692 71147 17744
rect 71083 17686 71147 17692
rect 82718 17744 82782 17750
rect 82718 17692 82724 17744
rect 82776 17692 82782 17744
rect 82718 17686 82782 17692
rect 93163 17744 93227 17750
rect 93163 17692 93169 17744
rect 93221 17692 93227 17744
rect 93163 17686 93227 17692
rect 104798 17744 104862 17750
rect 104798 17692 104804 17744
rect 104856 17692 104862 17744
rect 104798 17686 104862 17692
rect 115243 17744 115307 17750
rect 115243 17692 115249 17744
rect 115301 17692 115307 17744
rect 115243 17686 115307 17692
rect 37721 17572 37785 17578
rect 37721 17520 37727 17572
rect 37779 17520 37785 17572
rect 37721 17514 37785 17520
rect 38335 17572 38399 17578
rect 38335 17520 38341 17572
rect 38393 17520 38399 17572
rect 38335 17514 38399 17520
rect 59801 17572 59865 17578
rect 59801 17520 59807 17572
rect 59859 17520 59865 17572
rect 59801 17514 59865 17520
rect 60415 17572 60479 17578
rect 60415 17520 60421 17572
rect 60473 17520 60479 17572
rect 60415 17514 60479 17520
rect 81881 17572 81945 17578
rect 81881 17520 81887 17572
rect 81939 17520 81945 17572
rect 81881 17514 81945 17520
rect 82495 17572 82559 17578
rect 82495 17520 82501 17572
rect 82553 17520 82559 17572
rect 82495 17514 82559 17520
rect 103961 17572 104025 17578
rect 103961 17520 103967 17572
rect 104019 17520 104025 17572
rect 103961 17514 104025 17520
rect 104575 17572 104639 17578
rect 104575 17520 104581 17572
rect 104633 17520 104639 17572
rect 104575 17514 104639 17520
rect 48389 17344 48453 17350
rect 48389 17292 48395 17344
rect 48447 17292 48453 17344
rect 48389 17286 48453 17292
rect 70469 17344 70533 17350
rect 70469 17292 70475 17344
rect 70527 17292 70533 17344
rect 70469 17286 70533 17292
rect 92549 17344 92613 17350
rect 92549 17292 92555 17344
rect 92607 17292 92613 17344
rect 92549 17286 92613 17292
rect 114629 17344 114693 17350
rect 114629 17292 114635 17344
rect 114687 17292 114693 17344
rect 114629 17286 114693 17292
rect 135448 16601 140076 16647
<< via1 >>
rect 60049 48466 60101 48518
rect 49604 48380 49656 48432
rect 59435 48380 59487 48432
rect 82129 48466 82181 48518
rect 71684 48380 71736 48432
rect 81515 48380 81567 48432
rect 104209 48466 104261 48518
rect 126289 48466 126341 48518
rect 93764 48380 93816 48432
rect 103595 48380 103647 48432
rect 115844 48380 115896 48432
rect 125675 48380 125727 48432
rect 127256 48349 127308 48401
rect 48767 48208 48819 48260
rect 49381 48208 49433 48260
rect 70847 48208 70899 48260
rect 71461 48208 71513 48260
rect 92927 48208 92979 48260
rect 93541 48208 93593 48260
rect 115007 48208 115059 48260
rect 115621 48208 115673 48260
rect 61016 47909 61068 47961
rect 77469 45529 77521 45581
rect 77465 42398 77517 42450
rect 77465 38826 77517 38878
rect 77465 35270 77517 35322
rect 77417 28983 77469 29035
rect 77417 25419 77469 25471
rect 77417 21850 77469 21902
rect 77417 18905 77469 18957
rect 49976 17865 50028 17917
rect 72056 17865 72108 17917
rect 94135 17865 94187 17917
rect 116216 17865 116268 17917
rect 38564 17692 38616 17744
rect 49009 17692 49061 17744
rect 60644 17692 60696 17744
rect 71089 17692 71141 17744
rect 82724 17692 82776 17744
rect 93169 17692 93221 17744
rect 104804 17692 104856 17744
rect 115249 17692 115301 17744
rect 37727 17520 37779 17572
rect 38341 17520 38393 17572
rect 59807 17520 59859 17572
rect 60421 17520 60473 17572
rect 81887 17520 81939 17572
rect 82501 17520 82553 17572
rect 103967 17520 104019 17572
rect 104581 17520 104633 17572
rect 48395 17292 48447 17344
rect 70475 17292 70527 17344
rect 92555 17292 92607 17344
rect 114635 17292 114687 17344
<< metal2 >>
rect 48027 52317 48101 52326
rect 48027 52261 48036 52317
rect 48092 52261 48101 52317
rect 48027 52252 48101 52261
rect 59067 52317 59141 52326
rect 59067 52261 59076 52317
rect 59132 52261 59141 52317
rect 59067 52252 59141 52261
rect 70107 52317 70181 52326
rect 70107 52261 70116 52317
rect 70172 52261 70181 52317
rect 70107 52252 70181 52261
rect 81147 52317 81221 52326
rect 81147 52261 81156 52317
rect 81212 52261 81221 52317
rect 81147 52252 81221 52261
rect 92187 52317 92261 52326
rect 92187 52261 92196 52317
rect 92252 52261 92261 52317
rect 92187 52252 92261 52261
rect 103227 52317 103301 52326
rect 103227 52261 103236 52317
rect 103292 52261 103301 52317
rect 103227 52252 103301 52261
rect 114267 52317 114341 52326
rect 114267 52261 114276 52317
rect 114332 52261 114341 52317
rect 114267 52252 114341 52261
rect 60043 48518 60107 48524
rect 60043 48515 60049 48518
rect 60007 48469 60049 48515
rect 60043 48466 60049 48469
rect 60101 48515 60107 48518
rect 82123 48518 82187 48524
rect 82123 48515 82129 48518
rect 60101 48469 82129 48515
rect 60101 48466 60107 48469
rect 60043 48460 60107 48466
rect 82123 48466 82129 48469
rect 82181 48515 82187 48518
rect 104203 48518 104267 48524
rect 104203 48515 104209 48518
rect 82181 48469 104209 48515
rect 82181 48466 82187 48469
rect 82123 48460 82187 48466
rect 104203 48466 104209 48469
rect 104261 48515 104267 48518
rect 126283 48518 126347 48524
rect 126283 48515 126289 48518
rect 104261 48469 126289 48515
rect 104261 48466 104267 48469
rect 104203 48460 104267 48466
rect 126283 48466 126289 48469
rect 126341 48466 126347 48518
rect 126283 48460 126347 48466
rect 49598 48432 49662 48438
rect 49598 48380 49604 48432
rect 49656 48429 49662 48432
rect 59429 48432 59493 48438
rect 59429 48429 59435 48432
rect 49656 48383 59435 48429
rect 49656 48380 49662 48383
rect 49598 48374 49662 48380
rect 59429 48380 59435 48383
rect 59487 48380 59493 48432
rect 59429 48374 59493 48380
rect 71678 48432 71742 48438
rect 71678 48380 71684 48432
rect 71736 48429 71742 48432
rect 81509 48432 81573 48438
rect 81509 48429 81515 48432
rect 71736 48383 81515 48429
rect 71736 48380 71742 48383
rect 71678 48374 71742 48380
rect 81509 48380 81515 48383
rect 81567 48380 81573 48432
rect 81509 48374 81573 48380
rect 93758 48432 93822 48438
rect 93758 48380 93764 48432
rect 93816 48429 93822 48432
rect 103589 48432 103653 48438
rect 103589 48429 103595 48432
rect 93816 48383 103595 48429
rect 93816 48380 93822 48383
rect 93758 48374 93822 48380
rect 103589 48380 103595 48383
rect 103647 48380 103653 48432
rect 103589 48374 103653 48380
rect 115838 48432 115902 48438
rect 115838 48380 115844 48432
rect 115896 48429 115902 48432
rect 125669 48432 125733 48438
rect 125669 48429 125675 48432
rect 115896 48383 125675 48429
rect 115896 48380 115902 48383
rect 115838 48374 115902 48380
rect 125669 48380 125675 48383
rect 125727 48380 125733 48432
rect 125669 48374 125733 48380
rect 127245 48403 127319 48412
rect 127245 48347 127254 48403
rect 127310 48347 127319 48403
rect 127245 48338 127319 48347
rect 128604 48403 128678 48412
rect 128604 48347 128613 48403
rect 128669 48347 128678 48403
rect 128604 48338 128678 48347
rect 48027 48262 48101 48271
rect 48027 48206 48036 48262
rect 48092 48257 48101 48262
rect 48761 48260 48825 48266
rect 48761 48257 48767 48260
rect 48092 48211 48767 48257
rect 48092 48206 48101 48211
rect 48027 48197 48101 48206
rect 48761 48208 48767 48211
rect 48819 48208 48825 48260
rect 48761 48202 48825 48208
rect 49375 48260 49439 48266
rect 49375 48208 49381 48260
rect 49433 48257 49439 48260
rect 59067 48262 59141 48271
rect 59067 48257 59076 48262
rect 49433 48211 59076 48257
rect 49433 48208 49439 48211
rect 49375 48202 49439 48208
rect 59067 48206 59076 48211
rect 59132 48206 59141 48262
rect 59067 48197 59141 48206
rect 70107 48262 70181 48271
rect 70107 48206 70116 48262
rect 70172 48257 70181 48262
rect 70841 48260 70905 48266
rect 70841 48257 70847 48260
rect 70172 48211 70847 48257
rect 70172 48206 70181 48211
rect 70107 48197 70181 48206
rect 70841 48208 70847 48211
rect 70899 48208 70905 48260
rect 70841 48202 70905 48208
rect 71455 48260 71519 48266
rect 71455 48208 71461 48260
rect 71513 48257 71519 48260
rect 81147 48262 81221 48271
rect 81147 48257 81156 48262
rect 71513 48211 81156 48257
rect 71513 48208 71519 48211
rect 71455 48202 71519 48208
rect 81147 48206 81156 48211
rect 81212 48206 81221 48262
rect 81147 48197 81221 48206
rect 92187 48262 92261 48271
rect 92187 48206 92196 48262
rect 92252 48257 92261 48262
rect 92921 48260 92985 48266
rect 92921 48257 92927 48260
rect 92252 48211 92927 48257
rect 92252 48206 92261 48211
rect 92187 48197 92261 48206
rect 92921 48208 92927 48211
rect 92979 48208 92985 48260
rect 92921 48202 92985 48208
rect 93535 48260 93599 48266
rect 93535 48208 93541 48260
rect 93593 48257 93599 48260
rect 103227 48262 103301 48271
rect 103227 48257 103236 48262
rect 93593 48211 103236 48257
rect 93593 48208 93599 48211
rect 93535 48202 93599 48208
rect 103227 48206 103236 48211
rect 103292 48206 103301 48262
rect 103227 48197 103301 48206
rect 114267 48262 114341 48271
rect 114267 48206 114276 48262
rect 114332 48257 114341 48262
rect 115001 48260 115065 48266
rect 115001 48257 115007 48260
rect 114332 48211 115007 48257
rect 114332 48206 114341 48211
rect 114267 48197 114341 48206
rect 115001 48208 115007 48211
rect 115059 48208 115065 48260
rect 115001 48202 115065 48208
rect 115615 48260 115679 48266
rect 115615 48208 115621 48260
rect 115673 48257 115679 48260
rect 124832 48262 124906 48271
rect 124832 48257 124841 48262
rect 115673 48211 124841 48257
rect 115673 48208 115679 48211
rect 115615 48202 115679 48208
rect 124832 48206 124841 48211
rect 124897 48206 124906 48262
rect 124832 48197 124906 48206
rect 61005 47963 61079 47972
rect 61005 47907 61014 47963
rect 61070 47907 61079 47963
rect 61005 47898 61079 47907
rect 134008 46594 134082 46603
rect 134008 46589 134017 46594
rect 133446 46543 134017 46589
rect 134008 46538 134017 46543
rect 134073 46538 134082 46594
rect 134008 46529 134082 46538
rect 77463 45581 77527 45587
rect 77463 45529 77469 45581
rect 77521 45578 77527 45581
rect 125313 45583 125387 45592
rect 125313 45578 125322 45583
rect 77521 45532 125322 45578
rect 77521 45529 77527 45532
rect 77463 45523 77527 45529
rect 125313 45527 125322 45532
rect 125378 45527 125387 45583
rect 125313 45518 125387 45527
rect 134008 43030 134082 43039
rect 134008 43025 134017 43030
rect 133446 42979 134017 43025
rect 134008 42974 134017 42979
rect 134073 42974 134082 43030
rect 134008 42965 134082 42974
rect 77459 42450 77523 42456
rect 77459 42398 77465 42450
rect 77517 42447 77523 42450
rect 77517 42401 125327 42447
rect 77517 42398 77523 42401
rect 77459 42392 77523 42398
rect 134008 39466 134082 39475
rect 134008 39461 134017 39466
rect 133446 39415 134017 39461
rect 134008 39410 134017 39415
rect 134073 39410 134082 39466
rect 134008 39401 134082 39410
rect 77459 38878 77523 38884
rect 77459 38826 77465 38878
rect 77517 38875 77523 38878
rect 77517 38829 125376 38875
rect 77517 38826 77523 38829
rect 77459 38820 77523 38826
rect 134008 35902 134082 35911
rect 134008 35897 134017 35902
rect 133446 35851 134017 35897
rect 134008 35846 134017 35851
rect 134073 35846 134082 35902
rect 134008 35837 134082 35846
rect 77459 35322 77523 35328
rect 77459 35270 77465 35322
rect 77517 35319 77523 35322
rect 77517 35273 125328 35319
rect 77517 35270 77523 35273
rect 77459 35264 77523 35270
rect 134008 30222 134082 30231
rect 134008 30218 134017 30222
rect 133446 30172 134017 30218
rect 134008 30166 134017 30172
rect 134073 30166 134082 30222
rect 134008 30157 134082 30166
rect 77411 29035 77475 29041
rect 77411 28983 77417 29035
rect 77469 29032 77475 29035
rect 77469 28986 125387 29032
rect 77469 28983 77475 28986
rect 77411 28977 77475 28983
rect 134008 26659 134082 26668
rect 134008 26654 134017 26659
rect 133446 26608 134017 26654
rect 134008 26603 134017 26608
rect 134073 26603 134082 26659
rect 134008 26594 134082 26603
rect 77411 25471 77475 25477
rect 77411 25419 77417 25471
rect 77469 25468 77475 25471
rect 77469 25422 125387 25468
rect 77469 25419 77475 25422
rect 77411 25413 77475 25419
rect 134008 23095 134082 23104
rect 134008 23090 134017 23095
rect 133446 23044 134017 23090
rect 134008 23039 134017 23044
rect 134073 23039 134082 23095
rect 134008 23030 134082 23039
rect 77411 21904 77475 21908
rect 77411 21902 125387 21904
rect 77411 21850 77417 21902
rect 77469 21858 125387 21902
rect 77469 21850 77475 21858
rect 77411 21844 77475 21850
rect 134008 19531 134082 19540
rect 134008 19526 134017 19531
rect 133446 19480 134017 19526
rect 134008 19475 134017 19480
rect 134073 19475 134082 19531
rect 134008 19466 134082 19475
rect 77411 18957 77475 18963
rect 77411 18905 77417 18957
rect 77469 18948 77475 18957
rect 77469 18905 125332 18948
rect 77411 18902 125332 18905
rect 77411 18899 77475 18902
rect 49965 17919 50039 17928
rect 49965 17863 49974 17919
rect 50030 17863 50039 17919
rect 49965 17854 50039 17863
rect 72045 17919 72119 17928
rect 72045 17863 72054 17919
rect 72110 17863 72119 17919
rect 72045 17854 72119 17863
rect 94124 17919 94198 17928
rect 94124 17863 94133 17919
rect 94189 17863 94198 17919
rect 94124 17854 94198 17863
rect 116205 17919 116279 17928
rect 116205 17863 116214 17919
rect 116270 17863 116279 17919
rect 116205 17854 116279 17863
rect 38558 17744 38622 17750
rect 38558 17692 38564 17744
rect 38616 17741 38622 17744
rect 49003 17744 49067 17750
rect 49003 17741 49009 17744
rect 38616 17695 49009 17741
rect 38616 17692 38622 17695
rect 38558 17686 38622 17692
rect 49003 17692 49009 17695
rect 49061 17692 49067 17744
rect 49003 17686 49067 17692
rect 60638 17744 60702 17750
rect 60638 17692 60644 17744
rect 60696 17741 60702 17744
rect 71083 17744 71147 17750
rect 71083 17741 71089 17744
rect 60696 17695 71089 17741
rect 60696 17692 60702 17695
rect 60638 17686 60702 17692
rect 71083 17692 71089 17695
rect 71141 17692 71147 17744
rect 71083 17686 71147 17692
rect 82718 17744 82782 17750
rect 82718 17692 82724 17744
rect 82776 17741 82782 17744
rect 93163 17744 93227 17750
rect 93163 17741 93169 17744
rect 82776 17695 93169 17741
rect 82776 17692 82782 17695
rect 82718 17686 82782 17692
rect 93163 17692 93169 17695
rect 93221 17692 93227 17744
rect 93163 17686 93227 17692
rect 104798 17744 104862 17750
rect 104798 17692 104804 17744
rect 104856 17741 104862 17744
rect 115243 17744 115307 17750
rect 115243 17741 115249 17744
rect 104856 17695 115249 17741
rect 104856 17692 104862 17695
rect 104798 17686 104862 17692
rect 115243 17692 115249 17695
rect 115301 17692 115307 17744
rect 115243 17686 115307 17692
rect 37082 17574 37156 17583
rect 37082 17518 37091 17574
rect 37147 17569 37156 17574
rect 37721 17572 37785 17578
rect 37721 17569 37727 17572
rect 37147 17523 37727 17569
rect 37147 17518 37156 17523
rect 37082 17509 37156 17518
rect 37721 17520 37727 17523
rect 37779 17520 37785 17572
rect 37721 17514 37785 17520
rect 38335 17572 38399 17578
rect 38335 17520 38341 17572
rect 38393 17569 38399 17572
rect 48122 17574 48196 17583
rect 48122 17569 48131 17574
rect 38393 17523 48131 17569
rect 38393 17520 38399 17523
rect 38335 17514 38399 17520
rect 48122 17518 48131 17523
rect 48187 17518 48196 17574
rect 48122 17509 48196 17518
rect 59162 17574 59236 17583
rect 59162 17518 59171 17574
rect 59227 17569 59236 17574
rect 59801 17572 59865 17578
rect 59801 17569 59807 17572
rect 59227 17523 59807 17569
rect 59227 17518 59236 17523
rect 59162 17509 59236 17518
rect 59801 17520 59807 17523
rect 59859 17520 59865 17572
rect 59801 17514 59865 17520
rect 60415 17572 60479 17578
rect 60415 17520 60421 17572
rect 60473 17569 60479 17572
rect 70202 17574 70276 17583
rect 70202 17569 70211 17574
rect 60473 17523 70211 17569
rect 60473 17520 60479 17523
rect 60415 17514 60479 17520
rect 70202 17518 70211 17523
rect 70267 17518 70276 17574
rect 70202 17509 70276 17518
rect 81242 17574 81316 17583
rect 81242 17518 81251 17574
rect 81307 17569 81316 17574
rect 81881 17572 81945 17578
rect 81881 17569 81887 17572
rect 81307 17523 81887 17569
rect 81307 17518 81316 17523
rect 81242 17509 81316 17518
rect 81881 17520 81887 17523
rect 81939 17520 81945 17572
rect 81881 17514 81945 17520
rect 82495 17572 82559 17578
rect 82495 17520 82501 17572
rect 82553 17569 82559 17572
rect 92282 17574 92356 17583
rect 92282 17569 92291 17574
rect 82553 17523 92291 17569
rect 82553 17520 82559 17523
rect 82495 17514 82559 17520
rect 92282 17518 92291 17523
rect 92347 17518 92356 17574
rect 92282 17509 92356 17518
rect 103322 17574 103396 17583
rect 103322 17518 103331 17574
rect 103387 17569 103396 17574
rect 103961 17572 104025 17578
rect 103961 17569 103967 17572
rect 103387 17523 103967 17569
rect 103387 17518 103396 17523
rect 103322 17509 103396 17518
rect 103961 17520 103967 17523
rect 104019 17520 104025 17572
rect 103961 17514 104025 17520
rect 104575 17572 104639 17578
rect 104575 17520 104581 17572
rect 104633 17569 104639 17572
rect 114362 17574 114436 17583
rect 114362 17569 114371 17574
rect 104633 17523 114371 17569
rect 104633 17520 104639 17523
rect 104575 17514 104639 17520
rect 114362 17518 114371 17523
rect 114427 17518 114436 17574
rect 114362 17509 114436 17518
rect 48389 17344 48453 17350
rect 48389 17292 48395 17344
rect 48447 17341 48453 17344
rect 70469 17344 70533 17350
rect 70469 17341 70475 17344
rect 48447 17295 70475 17341
rect 48447 17292 48453 17295
rect 48389 17286 48453 17292
rect 70469 17292 70475 17295
rect 70527 17341 70533 17344
rect 92549 17344 92613 17350
rect 92549 17341 92555 17344
rect 70527 17295 92555 17341
rect 70527 17292 70533 17295
rect 70469 17286 70533 17292
rect 92549 17292 92555 17295
rect 92607 17341 92613 17344
rect 114629 17344 114693 17350
rect 114629 17341 114635 17344
rect 92607 17295 114635 17341
rect 92607 17292 92613 17295
rect 92549 17286 92613 17292
rect 114629 17292 114635 17295
rect 114687 17292 114693 17344
rect 114629 17286 114693 17292
rect 37082 15542 37156 15551
rect 37082 15486 37091 15542
rect 37147 15486 37156 15542
rect 37082 15477 37156 15486
rect 48121 15542 48196 15551
rect 48121 15486 48131 15542
rect 48187 15486 48196 15542
rect 48121 15477 48196 15486
rect 59162 15542 59236 15551
rect 59162 15486 59171 15542
rect 59227 15486 59236 15542
rect 59162 15477 59236 15486
rect 70202 15542 70276 15551
rect 70202 15486 70211 15542
rect 70267 15486 70276 15542
rect 70202 15477 70276 15486
rect 81242 15542 81316 15551
rect 81242 15486 81251 15542
rect 81307 15486 81316 15542
rect 81242 15477 81316 15486
rect 92282 15542 92356 15551
rect 92282 15486 92291 15542
rect 92347 15486 92356 15542
rect 92282 15477 92356 15486
rect 103322 15542 103396 15551
rect 103322 15486 103331 15542
rect 103387 15486 103396 15542
rect 103322 15477 103396 15486
rect 114362 15542 114436 15551
rect 114362 15486 114371 15542
rect 114427 15486 114436 15542
rect 114362 15477 114436 15486
<< via2 >>
rect 48036 52261 48092 52317
rect 59076 52261 59132 52317
rect 70116 52261 70172 52317
rect 81156 52261 81212 52317
rect 92196 52261 92252 52317
rect 103236 52261 103292 52317
rect 114276 52261 114332 52317
rect 127254 48401 127310 48403
rect 127254 48349 127256 48401
rect 127256 48349 127308 48401
rect 127308 48349 127310 48401
rect 127254 48347 127310 48349
rect 128613 48347 128669 48403
rect 48036 48206 48092 48262
rect 59076 48206 59132 48262
rect 70116 48206 70172 48262
rect 81156 48206 81212 48262
rect 92196 48206 92252 48262
rect 103236 48206 103292 48262
rect 114276 48206 114332 48262
rect 124841 48206 124897 48262
rect 61014 47961 61070 47963
rect 61014 47909 61016 47961
rect 61016 47909 61068 47961
rect 61068 47909 61070 47961
rect 61014 47907 61070 47909
rect 134017 46538 134073 46594
rect 125322 45527 125378 45583
rect 134017 42974 134073 43030
rect 134017 39410 134073 39466
rect 134017 35846 134073 35902
rect 134017 30166 134073 30222
rect 134017 26603 134073 26659
rect 134017 23039 134073 23095
rect 134017 19475 134073 19531
rect 49974 17917 50030 17919
rect 49974 17865 49976 17917
rect 49976 17865 50028 17917
rect 50028 17865 50030 17917
rect 49974 17863 50030 17865
rect 72054 17917 72110 17919
rect 72054 17865 72056 17917
rect 72056 17865 72108 17917
rect 72108 17865 72110 17917
rect 72054 17863 72110 17865
rect 94133 17917 94189 17919
rect 94133 17865 94135 17917
rect 94135 17865 94187 17917
rect 94187 17865 94189 17917
rect 94133 17863 94189 17865
rect 116214 17917 116270 17919
rect 116214 17865 116216 17917
rect 116216 17865 116268 17917
rect 116268 17865 116270 17917
rect 116214 17863 116270 17865
rect 37091 17518 37147 17574
rect 48131 17518 48187 17574
rect 59171 17518 59227 17574
rect 70211 17518 70267 17574
rect 81251 17518 81307 17574
rect 92291 17518 92347 17574
rect 103331 17518 103387 17574
rect 114371 17518 114427 17574
rect 37091 15486 37147 15542
rect 48131 15486 48187 15542
rect 59171 15486 59227 15542
rect 70211 15486 70267 15542
rect 81251 15486 81307 15542
rect 92291 15486 92347 15542
rect 103331 15486 103387 15542
rect 114371 15486 114427 15542
<< metal3 >>
rect 48031 52317 48097 52322
rect 48031 52261 48036 52317
rect 48092 52261 48097 52317
rect 48031 52256 48097 52261
rect 59071 52317 59137 52322
rect 59071 52261 59076 52317
rect 59132 52261 59137 52317
rect 59071 52256 59137 52261
rect 70111 52317 70177 52322
rect 70111 52261 70116 52317
rect 70172 52261 70177 52317
rect 70111 52256 70177 52261
rect 81151 52317 81217 52322
rect 81151 52261 81156 52317
rect 81212 52261 81217 52317
rect 81151 52256 81217 52261
rect 92191 52317 92257 52322
rect 92191 52261 92196 52317
rect 92252 52261 92257 52317
rect 92191 52256 92257 52261
rect 103231 52317 103297 52322
rect 103231 52261 103236 52317
rect 103292 52261 103297 52317
rect 103231 52256 103297 52261
rect 114271 52317 114337 52322
rect 114271 52261 114276 52317
rect 114332 52261 114337 52317
rect 114271 52256 114337 52261
rect 48034 48267 48094 52256
rect 59074 48267 59134 52256
rect 70114 48267 70174 52256
rect 81154 48267 81214 52256
rect 92194 48267 92254 52256
rect 103234 48267 103294 52256
rect 114274 48267 114334 52256
rect 127252 48413 127312 48466
rect 127244 48407 127320 48413
rect 127244 48343 127250 48407
rect 127314 48343 127320 48407
rect 127244 48337 127320 48343
rect 128603 48407 128679 48413
rect 128603 48343 128609 48407
rect 128673 48343 128679 48407
rect 128603 48337 128679 48343
rect 127252 48314 127312 48337
rect 48031 48262 48097 48267
rect 48031 48206 48036 48262
rect 48092 48206 48097 48262
rect 48031 48201 48097 48206
rect 59071 48262 59137 48267
rect 59071 48206 59076 48262
rect 59132 48206 59137 48262
rect 59071 48201 59137 48206
rect 70111 48262 70177 48267
rect 70111 48206 70116 48262
rect 70172 48206 70177 48262
rect 70111 48201 70177 48206
rect 81151 48262 81217 48267
rect 81151 48206 81156 48262
rect 81212 48206 81217 48262
rect 81151 48201 81217 48206
rect 92191 48262 92257 48267
rect 92191 48206 92196 48262
rect 92252 48206 92257 48262
rect 92191 48201 92257 48206
rect 103231 48262 103297 48267
rect 103231 48206 103236 48262
rect 103292 48206 103297 48262
rect 103231 48201 103297 48206
rect 114271 48262 114337 48267
rect 114271 48206 114276 48262
rect 114332 48206 114337 48262
rect 114271 48201 114337 48206
rect 124836 48262 124902 48267
rect 124836 48206 124841 48262
rect 124897 48206 124902 48262
rect 124836 48201 124902 48206
rect 48034 47786 48094 48201
rect 61012 47973 61072 48040
rect 61004 47967 61080 47973
rect 61004 47903 61010 47967
rect 61074 47903 61080 47967
rect 61004 47897 61080 47903
rect 61012 47854 61072 47897
rect 48026 47780 48102 47786
rect 48026 47716 48032 47780
rect 48096 47716 48102 47780
rect 48026 47710 48102 47716
rect 70114 43724 70174 48201
rect 70106 43718 70182 43724
rect 70106 43654 70112 43718
rect 70176 43654 70182 43718
rect 70106 43648 70182 43654
rect 83092 42167 83152 47958
rect 83084 42161 83160 42167
rect 83084 42097 83090 42161
rect 83154 42097 83160 42161
rect 83084 42091 83160 42097
rect 92194 38361 92254 48201
rect 105172 38516 105232 47960
rect 105164 38510 105240 38516
rect 105164 38446 105170 38510
rect 105234 38446 105240 38510
rect 105164 38440 105240 38446
rect 92186 38355 92262 38361
rect 92186 38291 92192 38355
rect 92256 38291 92262 38355
rect 92186 38285 92262 38291
rect 114274 34859 114334 48201
rect 125317 45583 125383 45588
rect 125317 45527 125322 45583
rect 125378 45527 125383 45583
rect 125317 45522 125383 45527
rect 128611 34982 128671 48337
rect 131459 47967 131535 47973
rect 131459 47903 131465 47967
rect 131529 47903 131535 47967
rect 131459 47897 131535 47903
rect 131467 45848 131527 47897
rect 132516 47780 132592 47786
rect 132516 47716 132522 47780
rect 132586 47716 132592 47780
rect 132516 47710 132592 47716
rect 132524 46357 132584 47710
rect 134012 46594 134078 46599
rect 134012 46538 134017 46594
rect 134073 46538 134078 46594
rect 134012 46533 134078 46538
rect 132516 43718 132592 43724
rect 132516 43654 132522 43718
rect 132586 43654 132592 43718
rect 132516 43648 132592 43654
rect 132524 42825 132584 43648
rect 134015 43035 134075 46533
rect 134012 43030 134078 43035
rect 134012 42974 134017 43030
rect 134073 42974 134078 43030
rect 134012 42969 134078 42974
rect 131459 42161 131535 42167
rect 131459 42097 131465 42161
rect 131529 42097 131535 42161
rect 131459 42091 131535 42097
rect 134015 39471 134075 42969
rect 134012 39466 134078 39471
rect 134012 39410 134017 39466
rect 134073 39410 134078 39466
rect 134012 39405 134078 39410
rect 131459 38510 131535 38516
rect 131459 38446 131465 38510
rect 131529 38446 131535 38510
rect 131459 38440 131535 38446
rect 132516 38355 132592 38361
rect 132516 38291 132522 38355
rect 132586 38291 132592 38355
rect 132516 38285 132592 38291
rect 134015 35907 134075 39405
rect 134012 35902 134078 35907
rect 134012 35846 134017 35902
rect 134073 35846 134078 35902
rect 134012 35841 134078 35846
rect 128603 34976 128679 34982
rect 128603 34912 128609 34976
rect 128673 34912 128679 34976
rect 128603 34906 128679 34912
rect 131459 34976 131535 34982
rect 131459 34912 131465 34976
rect 131529 34912 131535 34976
rect 131459 34906 131535 34912
rect 114266 34853 114342 34859
rect 114266 34789 114272 34853
rect 114336 34789 114342 34853
rect 114266 34783 114342 34789
rect 132516 34853 132592 34859
rect 132516 34789 132522 34853
rect 132586 34789 132592 34853
rect 132516 34783 132592 34789
rect 134015 30227 134075 35841
rect 137450 32768 137510 32848
rect 137442 32762 137518 32768
rect 137442 32698 137448 32762
rect 137512 32698 137518 32762
rect 137442 32692 137518 32698
rect 137450 32612 137510 32692
rect 134012 30222 134078 30227
rect 134012 30166 134017 30222
rect 134073 30166 134078 30222
rect 134012 30161 134078 30166
rect 114361 29637 114437 29643
rect 114361 29573 114367 29637
rect 114431 29573 114437 29637
rect 114361 29567 114437 29573
rect 132516 29637 132592 29643
rect 132516 29573 132522 29637
rect 132586 29573 132592 29637
rect 132516 29567 132592 29573
rect 94123 26088 94199 26094
rect 94123 26024 94129 26088
rect 94193 26024 94199 26088
rect 94123 26018 94199 26024
rect 92281 25898 92357 25904
rect 92281 25834 92287 25898
rect 92351 25834 92357 25898
rect 92281 25828 92357 25834
rect 70201 22509 70277 22515
rect 70201 22445 70207 22509
rect 70271 22445 70277 22509
rect 70201 22439 70277 22445
rect 49964 18605 50040 18611
rect 49964 18541 49970 18605
rect 50034 18541 50040 18605
rect 49964 18535 50040 18541
rect 48121 18349 48197 18355
rect 48121 18285 48127 18349
rect 48191 18285 48197 18349
rect 48121 18279 48197 18285
rect 48129 17579 48189 18279
rect 49972 17924 50032 18535
rect 49969 17919 50035 17924
rect 49969 17863 49974 17919
rect 50030 17863 50035 17919
rect 49969 17858 50035 17863
rect 70209 17579 70269 22439
rect 72044 22279 72120 22285
rect 72044 22215 72050 22279
rect 72114 22215 72120 22279
rect 72044 22209 72120 22215
rect 72052 17924 72112 22209
rect 72049 17919 72115 17924
rect 72049 17863 72054 17919
rect 72110 17863 72115 17919
rect 72049 17858 72115 17863
rect 92289 17579 92349 25828
rect 94131 17924 94191 26018
rect 94128 17919 94194 17924
rect 94128 17863 94133 17919
rect 94189 17863 94194 17919
rect 94128 17858 94194 17863
rect 114369 17579 114429 29567
rect 116204 29481 116280 29487
rect 116204 29417 116210 29481
rect 116274 29417 116280 29481
rect 116204 29411 116280 29417
rect 131459 29481 131535 29488
rect 131459 29417 131465 29481
rect 131529 29417 131535 29481
rect 131459 29411 131535 29417
rect 116212 17924 116272 29411
rect 134015 26664 134075 30161
rect 134012 26659 134078 26664
rect 134012 26603 134017 26659
rect 134073 26603 134078 26659
rect 134012 26598 134078 26603
rect 132516 26088 132592 26094
rect 132516 26024 132522 26088
rect 132586 26024 132592 26088
rect 132516 26018 132592 26024
rect 134015 23100 134075 26598
rect 134012 23095 134078 23100
rect 134012 23039 134017 23095
rect 134073 23039 134078 23095
rect 134012 23034 134078 23039
rect 132516 22509 132592 22515
rect 132516 22445 132522 22509
rect 132586 22445 132592 22509
rect 132516 22439 132592 22445
rect 131459 22279 131535 22285
rect 131459 22215 131465 22279
rect 131529 22215 131535 22279
rect 131459 22209 131535 22215
rect 134015 19536 134075 23034
rect 134012 19531 134078 19536
rect 134012 19475 134017 19531
rect 134073 19475 134078 19531
rect 134012 19470 134078 19475
rect 131459 18605 131535 18611
rect 131459 18541 131465 18605
rect 131529 18541 131535 18605
rect 131459 18535 131535 18541
rect 132516 18349 132592 18355
rect 132516 18285 132522 18349
rect 132586 18285 132592 18349
rect 132516 18279 132592 18285
rect 116209 17919 116275 17924
rect 116209 17863 116214 17919
rect 116270 17863 116275 17919
rect 116209 17858 116275 17863
rect 37086 17574 37152 17579
rect 37086 17518 37091 17574
rect 37147 17518 37152 17574
rect 37086 17513 37152 17518
rect 48126 17574 48192 17579
rect 48126 17518 48131 17574
rect 48187 17518 48192 17574
rect 48126 17513 48192 17518
rect 59166 17574 59232 17579
rect 59166 17518 59171 17574
rect 59227 17518 59232 17574
rect 59166 17513 59232 17518
rect 70206 17574 70272 17579
rect 70206 17518 70211 17574
rect 70267 17518 70272 17574
rect 70206 17513 70272 17518
rect 81246 17574 81312 17579
rect 81246 17518 81251 17574
rect 81307 17518 81312 17574
rect 81246 17513 81312 17518
rect 92286 17574 92352 17579
rect 92286 17518 92291 17574
rect 92347 17518 92352 17574
rect 92286 17513 92352 17518
rect 103326 17574 103392 17579
rect 103326 17518 103331 17574
rect 103387 17518 103392 17574
rect 103326 17513 103392 17518
rect 114366 17574 114432 17579
rect 114366 17518 114371 17574
rect 114427 17518 114432 17574
rect 114366 17513 114432 17518
rect 37089 15547 37149 17513
rect 48129 15547 48189 17513
rect 59169 15547 59229 17513
rect 70209 15547 70269 17513
rect 81249 15547 81309 17513
rect 92289 15547 92349 17513
rect 103329 15547 103389 17513
rect 114369 15547 114429 17513
rect 37086 15542 37152 15547
rect 37086 15486 37091 15542
rect 37147 15486 37152 15542
rect 37086 15481 37152 15486
rect 48126 15542 48192 15547
rect 48126 15486 48131 15542
rect 48187 15486 48192 15542
rect 48126 15481 48192 15486
rect 59166 15542 59232 15547
rect 59166 15486 59171 15542
rect 59227 15486 59232 15542
rect 59166 15481 59232 15486
rect 70206 15542 70272 15547
rect 70206 15486 70211 15542
rect 70267 15486 70272 15542
rect 70206 15481 70272 15486
rect 81246 15542 81312 15547
rect 81246 15486 81251 15542
rect 81307 15486 81312 15542
rect 81246 15481 81312 15486
rect 92286 15542 92352 15547
rect 92286 15486 92291 15542
rect 92347 15486 92352 15542
rect 92286 15481 92352 15486
rect 103326 15542 103392 15547
rect 103326 15486 103331 15542
rect 103387 15486 103392 15542
rect 103326 15481 103392 15486
rect 114366 15542 114432 15547
rect 114366 15486 114371 15542
rect 114427 15486 114432 15542
rect 114366 15481 114432 15486
<< via3 >>
rect 127250 48403 127314 48407
rect 127250 48347 127254 48403
rect 127254 48347 127310 48403
rect 127310 48347 127314 48403
rect 127250 48343 127314 48347
rect 128609 48403 128673 48407
rect 128609 48347 128613 48403
rect 128613 48347 128669 48403
rect 128669 48347 128673 48403
rect 128609 48343 128673 48347
rect 61010 47963 61074 47967
rect 61010 47907 61014 47963
rect 61014 47907 61070 47963
rect 61070 47907 61074 47963
rect 61010 47903 61074 47907
rect 48032 47716 48096 47780
rect 70112 43654 70176 43718
rect 83090 42097 83154 42161
rect 105170 38446 105234 38510
rect 92192 38291 92256 38355
rect 131465 47903 131529 47967
rect 132522 47716 132586 47780
rect 132522 43654 132586 43718
rect 131465 42097 131529 42161
rect 131465 38446 131529 38510
rect 132522 38291 132586 38355
rect 128609 34912 128673 34976
rect 131465 34912 131529 34976
rect 114272 34789 114336 34853
rect 132522 34789 132586 34853
rect 137448 32698 137512 32762
rect 114367 29573 114431 29637
rect 132522 29573 132586 29637
rect 94129 26024 94193 26088
rect 92287 25834 92351 25898
rect 70207 22445 70271 22509
rect 49970 18541 50034 18605
rect 48127 18285 48191 18349
rect 72050 22215 72114 22279
rect 116210 29417 116274 29481
rect 131465 29417 131529 29481
rect 132522 26024 132586 26088
rect 132522 22445 132586 22509
rect 131465 22215 131529 22279
rect 131465 18541 131529 18605
rect 132522 18285 132586 18349
<< metal4 >>
rect 127249 48407 127315 48408
rect 127249 48343 127250 48407
rect 127314 48405 127315 48407
rect 128608 48407 128674 48408
rect 128608 48405 128609 48407
rect 127314 48345 128609 48405
rect 127314 48343 127315 48345
rect 127249 48342 127315 48343
rect 128608 48343 128609 48345
rect 128673 48343 128674 48407
rect 128608 48342 128674 48343
rect 61009 47967 61075 47968
rect 61009 47903 61010 47967
rect 61074 47965 61075 47967
rect 131464 47967 131530 47968
rect 131464 47965 131465 47967
rect 61074 47905 131465 47965
rect 61074 47903 61075 47905
rect 61009 47902 61075 47903
rect 131464 47903 131465 47905
rect 131529 47903 131530 47967
rect 131464 47902 131530 47903
rect 48031 47780 48097 47781
rect 48031 47716 48032 47780
rect 48096 47778 48097 47780
rect 132521 47780 132587 47781
rect 132521 47778 132522 47780
rect 48096 47718 132522 47778
rect 48096 47716 48097 47718
rect 48031 47715 48097 47716
rect 132521 47716 132522 47718
rect 132586 47716 132587 47780
rect 132521 47715 132587 47716
rect 70111 43718 70177 43719
rect 70111 43654 70112 43718
rect 70176 43716 70177 43718
rect 132521 43718 132587 43719
rect 132521 43716 132522 43718
rect 70176 43656 132522 43716
rect 70176 43654 70177 43656
rect 70111 43653 70177 43654
rect 132521 43654 132522 43656
rect 132586 43654 132587 43718
rect 132521 43653 132587 43654
rect 83089 42161 83155 42162
rect 83089 42097 83090 42161
rect 83154 42159 83155 42161
rect 131464 42161 131530 42162
rect 131464 42159 131465 42161
rect 83154 42099 131465 42159
rect 83154 42097 83155 42099
rect 83089 42096 83155 42097
rect 131464 42097 131465 42099
rect 131529 42097 131530 42161
rect 131464 42096 131530 42097
rect 105169 38510 105235 38511
rect 105169 38446 105170 38510
rect 105234 38508 105235 38510
rect 131464 38510 131530 38511
rect 131464 38508 131465 38510
rect 105234 38448 131465 38508
rect 105234 38446 105235 38448
rect 105169 38445 105235 38446
rect 131464 38446 131465 38448
rect 131529 38446 131530 38510
rect 131464 38445 131530 38446
rect 92191 38355 92257 38356
rect 92191 38291 92192 38355
rect 92256 38353 92257 38355
rect 132521 38355 132587 38356
rect 132521 38353 132522 38355
rect 92256 38293 132522 38353
rect 92256 38291 92257 38293
rect 92191 38290 92257 38291
rect 132521 38291 132522 38293
rect 132586 38291 132587 38355
rect 132521 38290 132587 38291
rect 128608 34976 128674 34977
rect 128608 34912 128609 34976
rect 128673 34974 128674 34976
rect 131464 34976 131530 34977
rect 131464 34974 131465 34976
rect 128673 34914 131465 34974
rect 128673 34912 128674 34914
rect 128608 34911 128674 34912
rect 131464 34912 131465 34914
rect 131529 34912 131530 34976
rect 131464 34911 131530 34912
rect 114266 34853 114342 34859
rect 114266 34789 114272 34853
rect 114336 34851 114342 34853
rect 132521 34853 132587 34854
rect 132521 34851 132522 34853
rect 114336 34791 132522 34851
rect 114336 34789 114342 34791
rect 114266 34783 114342 34789
rect 132521 34789 132522 34791
rect 132586 34789 132587 34853
rect 132521 34788 132587 34789
rect 121458 32700 137362 32760
rect 114366 29637 114432 29638
rect 114366 29573 114367 29637
rect 114431 29635 114432 29637
rect 132521 29637 132587 29638
rect 132521 29635 132522 29637
rect 114431 29575 132522 29635
rect 114431 29573 114432 29575
rect 114366 29572 114432 29573
rect 132521 29573 132522 29575
rect 132586 29573 132587 29637
rect 132521 29572 132587 29573
rect 116209 29481 116275 29482
rect 116209 29417 116210 29481
rect 116274 29479 116275 29481
rect 131464 29481 131530 29482
rect 131464 29479 131465 29481
rect 116274 29419 131465 29479
rect 116274 29417 116275 29419
rect 116209 29416 116275 29417
rect 131464 29417 131465 29419
rect 131529 29417 131530 29481
rect 131464 29416 131530 29417
rect 94128 26088 94194 26089
rect 94128 26024 94129 26088
rect 94193 26086 94194 26088
rect 132521 26088 132587 26089
rect 132521 26086 132522 26088
rect 94193 26026 132522 26086
rect 94193 26024 94194 26026
rect 94128 26023 94194 26024
rect 132521 26024 132522 26026
rect 132586 26024 132587 26088
rect 132521 26023 132587 26024
rect 92286 25898 92352 25899
rect 92286 25834 92287 25898
rect 92351 25896 92352 25898
rect 92351 25836 132432 25896
rect 92351 25834 92352 25836
rect 92286 25833 92352 25834
rect 70206 22509 70272 22510
rect 70206 22445 70207 22509
rect 70271 22507 70272 22509
rect 132521 22509 132587 22510
rect 132521 22507 132522 22509
rect 70271 22447 132522 22507
rect 70271 22445 70272 22447
rect 70206 22444 70272 22445
rect 132521 22445 132522 22447
rect 132586 22445 132587 22509
rect 132521 22444 132587 22445
rect 72049 22279 72115 22280
rect 72049 22215 72050 22279
rect 72114 22277 72115 22279
rect 131464 22279 131530 22280
rect 131464 22277 131465 22279
rect 72114 22217 131465 22277
rect 72114 22215 72115 22217
rect 72049 22214 72115 22215
rect 131464 22215 131465 22217
rect 131529 22215 131530 22279
rect 132609 22217 134302 22277
rect 131464 22214 131530 22215
rect 49969 18605 50035 18606
rect 49969 18541 49970 18605
rect 50034 18603 50035 18605
rect 131464 18605 131530 18606
rect 131464 18603 131465 18605
rect 50034 18543 131465 18603
rect 50034 18541 50035 18543
rect 49969 18540 50035 18541
rect 131464 18541 131465 18543
rect 131529 18541 131530 18605
rect 131464 18540 131530 18541
rect 48126 18349 48192 18350
rect 48126 18285 48127 18349
rect 48191 18347 48192 18349
rect 132521 18349 132587 18350
rect 132521 18347 132522 18349
rect 48191 18287 132522 18347
rect 48191 18285 48192 18287
rect 48126 18284 48192 18285
rect 132521 18285 132522 18287
rect 132586 18285 132587 18349
rect 132521 18284 132587 18285
<< via4 >>
rect 137362 32762 137598 32848
rect 137362 32698 137448 32762
rect 137448 32698 137512 32762
rect 137512 32698 137598 32762
rect 137362 32612 137598 32698
rect 121458 30826 121694 31062
<< metal5 >>
rect 137320 32848 137640 32872
rect 137320 32612 137362 32848
rect 137598 32612 137640 32848
rect 137320 31172 137640 32612
rect 136794 26888 137114 27468
use And_Gate  And_Gate_0
timestamp 1756271862
transform 1 0 71687 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_1
timestamp 1756271862
transform 1 0 49607 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_2
timestamp 1756271862
transform 1 0 93767 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_3
timestamp 1756271862
transform 1 0 115847 0 1 16881
box -1558 -210 544 1618
use And_Gate  And_Gate_4
timestamp 1756271862
transform 1 0 82727 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_5
timestamp 1756271862
transform 1 0 60647 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_6
timestamp 1756271862
transform 1 0 104807 0 1 47569
box -1558 -210 544 1618
use And_Gate  And_Gate_7
timestamp 1756271862
transform 1 0 126887 0 1 47710
box -1558 -210 544 1618
use CDAC8  CDAC8_0
timestamp 1756271862
transform 1 0 68478 0 1 21136
box -39092 -2552 55448 26024
use comparator  comparator_0
timestamp 1755326863
transform -1 0 165417 0 1 18611
box 25341 -2024 30343 29246
use D_FlipFlop  D_FlipFlop_0
timestamp 1756271862
transform -1 0 133841 0 1 45613
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_1
timestamp 1756271862
transform -1 0 133841 0 1 34921
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_2
timestamp 1756271862
transform -1 0 133841 0 1 38485
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_3
timestamp 1756271862
transform -1 0 133841 0 1 42049
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_4
timestamp 1756271862
transform -1 0 133841 0 1 29242
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_5
timestamp 1756271862
transform -1 0 133841 0 1 25678
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_6
timestamp 1756271862
transform -1 0 133841 0 1 22114
box -102 -1796 8762 1842
use D_FlipFlop  D_FlipFlop_7
timestamp 1756271862
transform -1 0 133841 0 1 18550
box -102 -1796 8762 1842
use Nand_Gate  Nand_Gate_0
timestamp 1756271862
transform 1 0 68595 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_1
timestamp 1756271862
transform 1 0 101715 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_2
timestamp 1756271862
transform 1 0 90675 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_3
timestamp 1756271862
transform 1 0 46515 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_4
timestamp 1756271862
transform 1 0 35475 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_5
timestamp 1756271862
transform 1 0 112755 0 1 47889
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_6
timestamp 1756271862
transform 1 0 79635 0 1 17201
box 1906 -530 3264 1298
use Nand_Gate  Nand_Gate_7
timestamp 1756271862
transform 1 0 57555 0 1 17201
box 1906 -530 3264 1298
use RingCounter  RingCounter_0
timestamp 1756271862
transform 1 0 28071 0 1 12779
box -2592 -14 99850 40399
<< labels >>
flabel metal2 77469 18902 125332 18948 0 FreeSans 160 0 0 0 Q0
port 0 nsew
flabel metal2 77469 21858 125387 21904 0 FreeSans 160 0 0 0 Q1
port 1 nsew
flabel metal2 77469 25422 125387 25468 0 FreeSans 160 0 0 0 Q2
port 2 nsew
flabel metal2 77469 28986 125387 29032 0 FreeSans 160 0 0 0 Q3
port 3 nsew
flabel metal2 77517 35273 125328 35319 0 FreeSans 160 0 0 0 Q4
port 4 nsew
flabel metal2 77517 38829 125376 38875 0 FreeSans 160 0 0 0 Q5
port 5 nsew
flabel metal2 77517 42401 125327 42447 0 FreeSans 160 0 0 0 Q6
port 6 nsew
flabel metal2 77521 45532 125322 45578 0 FreeSans 160 0 0 0 Q7
port 7 nsew
flabel metal5 136794 26888 137114 27468 0 FreeSans 800 0 0 0 Vin
port 8 nsew
flabel metal1 135448 16601 140076 16647 0 FreeSans 160 0 0 0 Vbias
port 9 nsew
flabel metal1 92930 47983 92976 48515 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 70850 47983 70896 48515 0 FreeSans 160 0 0 0 A
port 2 nsew
flabel metal1 48770 47983 48816 48515 0 FreeSans 160 0 0 0 A
port 2 nsew
<< end >>
